VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_signal_buffering_alt
  CLASS BLOCK ;
  FOREIGN gpio_signal_buffering_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN mgmt_io_in_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 3540.800 3384.860 3542.390 ;
      LAYER mcon ;
        RECT 3384.690 3541.300 3384.860 3542.390 ;
      LAYER met1 ;
        RECT 3381.760 3542.085 3381.900 3575.605 ;
        RECT 3381.760 3541.765 3382.020 3542.085 ;
        RECT 3384.640 3541.240 3384.900 3542.450 ;
      LAYER via ;
        RECT 3381.760 3541.795 3382.020 3542.055 ;
        RECT 3384.640 3541.300 3384.900 3542.390 ;
      LAYER met2 ;
        RECT 3381.730 3541.935 3382.050 3542.055 ;
        RECT 3384.610 3541.935 3384.930 3542.390 ;
        RECT 3381.310 3541.795 3384.930 3541.935 ;
        RECT 3384.610 3541.300 3384.930 3541.795 ;
    END
  END mgmt_io_in_unbuf[13]
  PIN mgmt_io_out_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 3540.895 3388.770 3541.065 ;
        RECT 3387.410 3540.810 3388.290 3540.895 ;
        RECT 3387.410 3540.225 3387.580 3540.810 ;
        RECT 3386.560 3540.055 3387.580 3540.225 ;
        RECT 3387.410 3539.385 3387.580 3540.055 ;
        RECT 3386.560 3539.215 3387.580 3539.385 ;
        RECT 3387.410 3538.545 3387.580 3539.215 ;
        RECT 3386.560 3538.375 3387.580 3538.545 ;
        RECT 3388.120 3540.225 3388.290 3540.810 ;
        RECT 3388.120 3540.055 3388.770 3540.225 ;
        RECT 3388.120 3539.385 3388.290 3540.055 ;
        RECT 3388.120 3539.215 3388.770 3539.385 ;
        RECT 3388.120 3538.545 3388.290 3539.215 ;
        RECT 3388.120 3538.375 3388.770 3538.545 ;
      LAYER met1 ;
        RECT 3381.480 3541.115 3381.620 3574.605 ;
        RECT 3381.480 3540.795 3381.740 3541.115 ;
        RECT 3387.350 3540.760 3388.320 3541.020 ;
      LAYER via ;
        RECT 3381.480 3540.825 3381.740 3541.085 ;
        RECT 3387.410 3540.760 3388.260 3541.020 ;
      LAYER met2 ;
        RECT 3381.450 3540.965 3381.770 3541.085 ;
        RECT 3387.410 3540.965 3388.260 3541.050 ;
        RECT 3381.310 3540.825 3388.260 3540.965 ;
        RECT 3387.410 3540.730 3388.260 3540.825 ;
    END
  END mgmt_io_out_buf[13]
  PIN mgmt_io_in_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2230.700 3384.860 2232.290 ;
      LAYER mcon ;
        RECT 3384.690 2231.200 3384.860 2232.290 ;
      LAYER met1 ;
        RECT 3381.200 2231.985 3381.340 2281.275 ;
        RECT 3381.200 2231.665 3381.460 2231.985 ;
        RECT 3384.640 2231.140 3384.900 2232.350 ;
      LAYER via ;
        RECT 3381.200 2231.695 3381.460 2231.955 ;
        RECT 3384.640 2231.200 3384.900 2232.290 ;
      LAYER met2 ;
        RECT 3381.170 2231.835 3381.490 2231.955 ;
        RECT 3384.610 2231.835 3384.930 2232.290 ;
        RECT 3377.950 2231.695 3384.930 2231.835 ;
        RECT 3384.610 2231.200 3384.930 2231.695 ;
    END
  END mgmt_io_in_unbuf[12]
  PIN mgmt_io_in_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2224.720 3384.860 2226.310 ;
      LAYER mcon ;
        RECT 3384.690 2225.220 3384.860 2226.310 ;
      LAYER met1 ;
        RECT 3380.640 2226.005 3380.780 2279.275 ;
        RECT 3380.640 2225.685 3380.900 2226.005 ;
        RECT 3384.640 2225.160 3384.900 2226.370 ;
      LAYER via ;
        RECT 3380.640 2225.715 3380.900 2225.975 ;
        RECT 3384.640 2225.220 3384.900 2226.310 ;
      LAYER met2 ;
        RECT 3380.610 2225.855 3380.930 2225.975 ;
        RECT 3384.610 2225.855 3384.930 2226.310 ;
        RECT 3377.950 2225.715 3384.930 2225.855 ;
        RECT 3384.610 2225.220 3384.930 2225.715 ;
    END
  END mgmt_io_in_unbuf[11]
  PIN mgmt_io_in_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2218.740 3384.860 2220.330 ;
      LAYER mcon ;
        RECT 3384.690 2219.240 3384.860 2220.330 ;
      LAYER met1 ;
        RECT 3380.080 2220.025 3380.220 2277.275 ;
        RECT 3380.080 2219.705 3380.340 2220.025 ;
        RECT 3384.640 2219.180 3384.900 2220.390 ;
      LAYER via ;
        RECT 3380.080 2219.735 3380.340 2219.995 ;
        RECT 3384.640 2219.240 3384.900 2220.330 ;
      LAYER met2 ;
        RECT 3380.050 2219.875 3380.370 2219.995 ;
        RECT 3384.610 2219.875 3384.930 2220.330 ;
        RECT 3377.950 2219.735 3384.930 2219.875 ;
        RECT 3384.610 2219.240 3384.930 2219.735 ;
    END
  END mgmt_io_in_unbuf[10]
  PIN mgmt_io_in_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2212.760 3384.860 2214.350 ;
      LAYER mcon ;
        RECT 3384.690 2213.260 3384.860 2214.350 ;
      LAYER met1 ;
        RECT 3379.520 2214.045 3379.660 2275.275 ;
        RECT 3379.520 2213.725 3379.780 2214.045 ;
        RECT 3384.640 2213.200 3384.900 2214.410 ;
      LAYER via ;
        RECT 3379.520 2213.755 3379.780 2214.015 ;
        RECT 3384.640 2213.260 3384.900 2214.350 ;
      LAYER met2 ;
        RECT 3379.490 2213.895 3379.810 2214.015 ;
        RECT 3384.610 2213.895 3384.930 2214.350 ;
        RECT 3377.950 2213.755 3384.930 2213.895 ;
        RECT 3384.610 2213.260 3384.930 2213.755 ;
    END
  END mgmt_io_in_unbuf[9]
  PIN mgmt_io_in_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2206.780 3384.860 2208.370 ;
      LAYER mcon ;
        RECT 3384.690 2207.280 3384.860 2208.370 ;
      LAYER met1 ;
        RECT 3378.960 2208.065 3379.100 2273.275 ;
        RECT 3378.960 2207.745 3379.220 2208.065 ;
        RECT 3384.640 2207.220 3384.900 2208.430 ;
      LAYER via ;
        RECT 3378.960 2207.775 3379.220 2208.035 ;
        RECT 3384.640 2207.280 3384.900 2208.370 ;
      LAYER met2 ;
        RECT 3378.930 2207.915 3379.250 2208.035 ;
        RECT 3384.610 2207.915 3384.930 2208.370 ;
        RECT 3377.950 2207.775 3384.930 2207.915 ;
        RECT 3384.610 2207.280 3384.930 2207.775 ;
    END
  END mgmt_io_in_unbuf[8]
  PIN mgmt_io_in_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2200.800 3384.860 2202.390 ;
      LAYER mcon ;
        RECT 3384.690 2201.300 3384.860 2202.390 ;
      LAYER met1 ;
        RECT 3378.400 2202.085 3378.540 2271.275 ;
        RECT 3378.400 2201.765 3378.660 2202.085 ;
        RECT 3384.640 2201.240 3384.900 2202.450 ;
      LAYER via ;
        RECT 3378.400 2201.795 3378.660 2202.055 ;
        RECT 3384.640 2201.300 3384.900 2202.390 ;
      LAYER met2 ;
        RECT 3378.370 2201.935 3378.690 2202.055 ;
        RECT 3384.610 2201.935 3384.930 2202.390 ;
        RECT 3377.950 2201.795 3384.930 2201.935 ;
        RECT 3384.610 2201.300 3384.930 2201.795 ;
    END
  END mgmt_io_in_unbuf[7]
  PIN mgmt_io_out_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2200.895 3388.770 2201.065 ;
        RECT 3387.410 2200.810 3388.290 2200.895 ;
        RECT 3387.410 2200.225 3387.580 2200.810 ;
        RECT 3386.560 2200.055 3387.580 2200.225 ;
        RECT 3387.410 2199.385 3387.580 2200.055 ;
        RECT 3386.560 2199.215 3387.580 2199.385 ;
        RECT 3387.410 2198.545 3387.580 2199.215 ;
        RECT 3386.560 2198.375 3387.580 2198.545 ;
        RECT 3388.120 2200.225 3388.290 2200.810 ;
        RECT 3388.120 2200.055 3388.770 2200.225 ;
        RECT 3388.120 2199.385 3388.290 2200.055 ;
        RECT 3388.120 2199.215 3388.770 2199.385 ;
        RECT 3388.120 2198.545 3388.290 2199.215 ;
        RECT 3388.120 2198.375 3388.770 2198.545 ;
      LAYER met1 ;
        RECT 3378.120 2201.115 3378.260 2270.275 ;
        RECT 3378.120 2200.795 3378.380 2201.115 ;
        RECT 3387.350 2200.760 3388.320 2201.020 ;
      LAYER via ;
        RECT 3378.120 2200.825 3378.380 2201.085 ;
        RECT 3387.410 2200.760 3388.260 2201.020 ;
      LAYER met2 ;
        RECT 3378.090 2200.965 3378.410 2201.085 ;
        RECT 3387.410 2200.965 3388.260 2201.050 ;
        RECT 3377.950 2200.825 3388.260 2200.965 ;
        RECT 3387.410 2200.730 3388.260 2200.825 ;
    END
  END mgmt_io_out_buf[7]
  PIN mgmt_io_out_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2206.875 3388.770 2207.045 ;
        RECT 3387.410 2206.790 3388.290 2206.875 ;
        RECT 3387.410 2206.205 3387.580 2206.790 ;
        RECT 3386.560 2206.035 3387.580 2206.205 ;
        RECT 3387.410 2205.365 3387.580 2206.035 ;
        RECT 3386.560 2205.195 3387.580 2205.365 ;
        RECT 3387.410 2204.525 3387.580 2205.195 ;
        RECT 3386.560 2204.355 3387.580 2204.525 ;
        RECT 3388.120 2206.205 3388.290 2206.790 ;
        RECT 3388.120 2206.035 3388.770 2206.205 ;
        RECT 3388.120 2205.365 3388.290 2206.035 ;
        RECT 3388.120 2205.195 3388.770 2205.365 ;
        RECT 3388.120 2204.525 3388.290 2205.195 ;
        RECT 3388.120 2204.355 3388.770 2204.525 ;
      LAYER met1 ;
        RECT 3378.680 2207.095 3378.820 2272.275 ;
        RECT 3378.680 2206.775 3378.940 2207.095 ;
        RECT 3387.350 2206.740 3388.320 2207.000 ;
      LAYER via ;
        RECT 3378.680 2206.805 3378.940 2207.065 ;
        RECT 3387.410 2206.740 3388.260 2207.000 ;
      LAYER met2 ;
        RECT 3378.650 2206.945 3378.970 2207.065 ;
        RECT 3387.410 2206.945 3388.260 2207.030 ;
        RECT 3377.950 2206.805 3388.260 2206.945 ;
        RECT 3387.410 2206.710 3388.260 2206.805 ;
    END
  END mgmt_io_out_buf[8]
  PIN mgmt_io_out_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2212.855 3388.770 2213.025 ;
        RECT 3387.410 2212.770 3388.290 2212.855 ;
        RECT 3387.410 2212.185 3387.580 2212.770 ;
        RECT 3386.560 2212.015 3387.580 2212.185 ;
        RECT 3387.410 2211.345 3387.580 2212.015 ;
        RECT 3386.560 2211.175 3387.580 2211.345 ;
        RECT 3387.410 2210.505 3387.580 2211.175 ;
        RECT 3386.560 2210.335 3387.580 2210.505 ;
        RECT 3388.120 2212.185 3388.290 2212.770 ;
        RECT 3388.120 2212.015 3388.770 2212.185 ;
        RECT 3388.120 2211.345 3388.290 2212.015 ;
        RECT 3388.120 2211.175 3388.770 2211.345 ;
        RECT 3388.120 2210.505 3388.290 2211.175 ;
        RECT 3388.120 2210.335 3388.770 2210.505 ;
      LAYER met1 ;
        RECT 3379.240 2213.075 3379.380 2274.275 ;
        RECT 3379.240 2212.755 3379.500 2213.075 ;
        RECT 3387.350 2212.720 3388.320 2212.980 ;
      LAYER via ;
        RECT 3379.240 2212.785 3379.500 2213.045 ;
        RECT 3387.410 2212.720 3388.260 2212.980 ;
      LAYER met2 ;
        RECT 3379.210 2212.925 3379.530 2213.045 ;
        RECT 3387.410 2212.925 3388.260 2213.010 ;
        RECT 3377.950 2212.785 3388.260 2212.925 ;
        RECT 3387.410 2212.690 3388.260 2212.785 ;
    END
  END mgmt_io_out_buf[9]
  PIN mgmt_io_out_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2218.835 3388.770 2219.005 ;
        RECT 3387.410 2218.750 3388.290 2218.835 ;
        RECT 3387.410 2218.165 3387.580 2218.750 ;
        RECT 3386.560 2217.995 3387.580 2218.165 ;
        RECT 3387.410 2217.325 3387.580 2217.995 ;
        RECT 3386.560 2217.155 3387.580 2217.325 ;
        RECT 3387.410 2216.485 3387.580 2217.155 ;
        RECT 3386.560 2216.315 3387.580 2216.485 ;
        RECT 3388.120 2218.165 3388.290 2218.750 ;
        RECT 3388.120 2217.995 3388.770 2218.165 ;
        RECT 3388.120 2217.325 3388.290 2217.995 ;
        RECT 3388.120 2217.155 3388.770 2217.325 ;
        RECT 3388.120 2216.485 3388.290 2217.155 ;
        RECT 3388.120 2216.315 3388.770 2216.485 ;
      LAYER met1 ;
        RECT 3379.800 2219.055 3379.940 2276.275 ;
        RECT 3379.800 2218.735 3380.060 2219.055 ;
        RECT 3387.350 2218.700 3388.320 2218.960 ;
      LAYER via ;
        RECT 3379.800 2218.765 3380.060 2219.025 ;
        RECT 3387.410 2218.700 3388.260 2218.960 ;
      LAYER met2 ;
        RECT 3379.770 2218.905 3380.090 2219.025 ;
        RECT 3387.410 2218.905 3388.260 2218.990 ;
        RECT 3377.950 2218.765 3388.260 2218.905 ;
        RECT 3387.410 2218.670 3388.260 2218.765 ;
    END
  END mgmt_io_out_buf[10]
  PIN mgmt_io_out_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2224.815 3388.770 2224.985 ;
        RECT 3387.410 2224.730 3388.290 2224.815 ;
        RECT 3387.410 2224.145 3387.580 2224.730 ;
        RECT 3386.560 2223.975 3387.580 2224.145 ;
        RECT 3387.410 2223.305 3387.580 2223.975 ;
        RECT 3386.560 2223.135 3387.580 2223.305 ;
        RECT 3387.410 2222.465 3387.580 2223.135 ;
        RECT 3386.560 2222.295 3387.580 2222.465 ;
        RECT 3388.120 2224.145 3388.290 2224.730 ;
        RECT 3388.120 2223.975 3388.770 2224.145 ;
        RECT 3388.120 2223.305 3388.290 2223.975 ;
        RECT 3388.120 2223.135 3388.770 2223.305 ;
        RECT 3388.120 2222.465 3388.290 2223.135 ;
        RECT 3388.120 2222.295 3388.770 2222.465 ;
      LAYER met1 ;
        RECT 3380.360 2225.035 3380.500 2278.275 ;
        RECT 3380.360 2224.715 3380.620 2225.035 ;
        RECT 3387.350 2224.680 3388.320 2224.940 ;
      LAYER via ;
        RECT 3380.360 2224.745 3380.620 2225.005 ;
        RECT 3387.410 2224.680 3388.260 2224.940 ;
      LAYER met2 ;
        RECT 3380.330 2224.885 3380.650 2225.005 ;
        RECT 3387.410 2224.885 3388.260 2224.970 ;
        RECT 3377.950 2224.745 3388.260 2224.885 ;
        RECT 3387.410 2224.650 3388.260 2224.745 ;
    END
  END mgmt_io_out_buf[11]
  PIN mgmt_io_out_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2230.795 3388.770 2230.965 ;
        RECT 3387.410 2230.710 3388.290 2230.795 ;
        RECT 3387.410 2230.125 3387.580 2230.710 ;
        RECT 3386.560 2229.955 3387.580 2230.125 ;
        RECT 3387.410 2229.285 3387.580 2229.955 ;
        RECT 3386.560 2229.115 3387.580 2229.285 ;
        RECT 3387.410 2228.445 3387.580 2229.115 ;
        RECT 3386.560 2228.275 3387.580 2228.445 ;
        RECT 3388.120 2230.125 3388.290 2230.710 ;
        RECT 3388.120 2229.955 3388.770 2230.125 ;
        RECT 3388.120 2229.285 3388.290 2229.955 ;
        RECT 3388.120 2229.115 3388.770 2229.285 ;
        RECT 3388.120 2228.445 3388.290 2229.115 ;
        RECT 3388.120 2228.275 3388.770 2228.445 ;
      LAYER met1 ;
        RECT 3380.920 2231.015 3381.060 2280.275 ;
        RECT 3380.920 2230.695 3381.180 2231.015 ;
        RECT 3387.350 2230.660 3388.320 2230.920 ;
      LAYER via ;
        RECT 3380.920 2230.725 3381.180 2230.985 ;
        RECT 3387.410 2230.660 3388.260 2230.920 ;
      LAYER met2 ;
        RECT 3380.890 2230.865 3381.210 2230.985 ;
        RECT 3387.410 2230.865 3388.260 2230.950 ;
        RECT 3377.950 2230.725 3388.260 2230.865 ;
        RECT 3387.410 2230.630 3388.260 2230.725 ;
    END
  END mgmt_io_out_buf[12]
  PIN mgmt_io_out_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2196.660 3387.950 2197.760 ;
      LAYER mcon ;
        RECT 3387.750 2196.670 3387.920 2197.760 ;
      LAYER met1 ;
        RECT 3378.140 2196.930 3378.400 2197.250 ;
        RECT 3378.260 1075.250 3378.400 2196.930 ;
        RECT 3387.700 2196.610 3387.960 2197.820 ;
      LAYER via ;
        RECT 3378.140 2196.960 3378.400 2197.220 ;
        RECT 3387.700 2196.670 3387.960 2197.760 ;
      LAYER met2 ;
        RECT 3378.110 2197.100 3378.430 2197.220 ;
        RECT 3387.670 2197.100 3387.990 2197.760 ;
        RECT 3377.950 2196.960 3387.990 2197.100 ;
        RECT 3387.670 2196.670 3387.990 2196.960 ;
    END
  END mgmt_io_out_unbuf[7]
  PIN mgmt_io_out_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2202.640 3387.950 2203.740 ;
      LAYER mcon ;
        RECT 3387.750 2202.650 3387.920 2203.740 ;
      LAYER met1 ;
        RECT 3378.700 2202.910 3378.960 2203.230 ;
        RECT 3378.820 1073.250 3378.960 2202.910 ;
        RECT 3387.700 2202.590 3387.960 2203.800 ;
      LAYER via ;
        RECT 3378.700 2202.940 3378.960 2203.200 ;
        RECT 3387.700 2202.650 3387.960 2203.740 ;
      LAYER met2 ;
        RECT 3378.670 2203.080 3378.990 2203.200 ;
        RECT 3387.670 2203.080 3387.990 2203.740 ;
        RECT 3377.950 2202.940 3387.990 2203.080 ;
        RECT 3387.670 2202.650 3387.990 2202.940 ;
    END
  END mgmt_io_out_unbuf[8]
  PIN mgmt_io_out_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2208.620 3387.950 2209.720 ;
      LAYER mcon ;
        RECT 3387.750 2208.630 3387.920 2209.720 ;
      LAYER met1 ;
        RECT 3379.260 2208.890 3379.520 2209.210 ;
        RECT 3379.380 1071.250 3379.520 2208.890 ;
        RECT 3387.700 2208.570 3387.960 2209.780 ;
      LAYER via ;
        RECT 3379.260 2208.920 3379.520 2209.180 ;
        RECT 3387.700 2208.630 3387.960 2209.720 ;
      LAYER met2 ;
        RECT 3379.230 2209.060 3379.550 2209.180 ;
        RECT 3387.670 2209.060 3387.990 2209.720 ;
        RECT 3377.950 2208.920 3387.990 2209.060 ;
        RECT 3387.670 2208.630 3387.990 2208.920 ;
    END
  END mgmt_io_out_unbuf[9]
  PIN mgmt_io_out_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2214.600 3387.950 2215.700 ;
      LAYER mcon ;
        RECT 3387.750 2214.610 3387.920 2215.700 ;
      LAYER met1 ;
        RECT 3379.820 2214.870 3380.080 2215.190 ;
        RECT 3379.940 1069.250 3380.080 2214.870 ;
        RECT 3387.700 2214.550 3387.960 2215.760 ;
      LAYER via ;
        RECT 3379.820 2214.900 3380.080 2215.160 ;
        RECT 3387.700 2214.610 3387.960 2215.700 ;
      LAYER met2 ;
        RECT 3379.790 2215.040 3380.110 2215.160 ;
        RECT 3387.670 2215.040 3387.990 2215.700 ;
        RECT 3377.950 2214.900 3387.990 2215.040 ;
        RECT 3387.670 2214.610 3387.990 2214.900 ;
    END
  END mgmt_io_out_unbuf[10]
  PIN mgmt_io_out_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2220.580 3387.950 2221.680 ;
      LAYER mcon ;
        RECT 3387.750 2220.590 3387.920 2221.680 ;
      LAYER met1 ;
        RECT 3380.380 2220.850 3380.640 2221.170 ;
        RECT 3380.500 1067.250 3380.640 2220.850 ;
        RECT 3387.700 2220.530 3387.960 2221.740 ;
      LAYER via ;
        RECT 3380.380 2220.880 3380.640 2221.140 ;
        RECT 3387.700 2220.590 3387.960 2221.680 ;
      LAYER met2 ;
        RECT 3380.350 2221.020 3380.670 2221.140 ;
        RECT 3387.670 2221.020 3387.990 2221.680 ;
        RECT 3377.950 2220.880 3387.990 2221.020 ;
        RECT 3387.670 2220.590 3387.990 2220.880 ;
    END
  END mgmt_io_out_unbuf[11]
  PIN mgmt_io_out_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2226.560 3387.950 2227.660 ;
      LAYER mcon ;
        RECT 3387.750 2226.570 3387.920 2227.660 ;
      LAYER met1 ;
        RECT 3380.940 2226.830 3381.200 2227.150 ;
        RECT 3381.060 1065.250 3381.200 2226.830 ;
        RECT 3387.700 2226.510 3387.960 2227.720 ;
      LAYER via ;
        RECT 3380.940 2226.860 3381.200 2227.120 ;
        RECT 3387.700 2226.570 3387.960 2227.660 ;
      LAYER met2 ;
        RECT 3380.910 2227.000 3381.230 2227.120 ;
        RECT 3387.670 2227.000 3387.990 2227.660 ;
        RECT 3377.950 2226.860 3387.990 2227.000 ;
        RECT 3387.670 2226.570 3387.990 2226.860 ;
    END
  END mgmt_io_out_unbuf[12]
  PIN mgmt_io_out_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2232.540 3387.950 2233.640 ;
      LAYER mcon ;
        RECT 3387.750 2232.550 3387.920 2233.640 ;
      LAYER met1 ;
        RECT 3381.500 2232.810 3381.760 2233.130 ;
        RECT 3381.620 1063.250 3381.760 2232.810 ;
        RECT 3387.700 2232.490 3387.960 2233.700 ;
      LAYER via ;
        RECT 3381.500 2232.840 3381.760 2233.100 ;
        RECT 3387.700 2232.550 3387.960 2233.640 ;
      LAYER met2 ;
        RECT 3381.470 2232.980 3381.790 2233.100 ;
        RECT 3387.670 2232.980 3387.990 2233.640 ;
        RECT 3377.950 2232.840 3387.990 2232.980 ;
        RECT 3387.670 2232.550 3387.990 2232.840 ;
    END
  END mgmt_io_out_unbuf[13]
  PIN mgmt_io_in_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2235.895 3384.490 2236.065 ;
        RECT 3384.320 2235.225 3384.490 2235.895 ;
        RECT 3383.840 2235.055 3384.490 2235.225 ;
        RECT 3384.320 2234.385 3384.490 2235.055 ;
        RECT 3383.840 2234.215 3384.490 2234.385 ;
        RECT 3384.320 2233.630 3384.490 2234.215 ;
        RECT 3385.030 2235.895 3386.050 2236.065 ;
        RECT 3385.030 2235.225 3385.200 2235.895 ;
        RECT 3385.030 2235.055 3386.050 2235.225 ;
        RECT 3385.030 2234.385 3385.200 2235.055 ;
        RECT 3385.030 2234.215 3386.050 2234.385 ;
        RECT 3385.030 2233.630 3385.200 2234.215 ;
        RECT 3384.320 2233.545 3385.200 2233.630 ;
        RECT 3383.840 2233.375 3386.050 2233.545 ;
      LAYER mcon ;
        RECT 3384.350 2233.460 3385.200 2233.630 ;
      LAYER met1 ;
        RECT 3381.780 2233.430 3382.040 2233.750 ;
        RECT 3381.900 1062.250 3382.040 2233.430 ;
        RECT 3384.290 2233.410 3385.260 2233.670 ;
      LAYER via ;
        RECT 3381.780 2233.460 3382.040 2233.720 ;
        RECT 3384.350 2233.410 3385.200 2233.670 ;
      LAYER met2 ;
        RECT 3381.750 2233.600 3382.070 2233.720 ;
        RECT 3384.350 2233.600 3385.200 2233.700 ;
        RECT 3377.950 2233.460 3385.200 2233.600 ;
        RECT 3384.350 2233.380 3385.200 2233.460 ;
    END
  END mgmt_io_in_buf[13]
  PIN mgmt_io_in_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2229.915 3384.490 2230.085 ;
        RECT 3384.320 2229.245 3384.490 2229.915 ;
        RECT 3383.840 2229.075 3384.490 2229.245 ;
        RECT 3384.320 2228.405 3384.490 2229.075 ;
        RECT 3383.840 2228.235 3384.490 2228.405 ;
        RECT 3384.320 2227.650 3384.490 2228.235 ;
        RECT 3385.030 2229.915 3386.050 2230.085 ;
        RECT 3385.030 2229.245 3385.200 2229.915 ;
        RECT 3385.030 2229.075 3386.050 2229.245 ;
        RECT 3385.030 2228.405 3385.200 2229.075 ;
        RECT 3385.030 2228.235 3386.050 2228.405 ;
        RECT 3385.030 2227.650 3385.200 2228.235 ;
        RECT 3384.320 2227.565 3385.200 2227.650 ;
        RECT 3383.840 2227.395 3386.050 2227.565 ;
      LAYER mcon ;
        RECT 3384.350 2227.480 3385.200 2227.650 ;
      LAYER met1 ;
        RECT 3381.220 2227.450 3381.480 2227.770 ;
        RECT 3381.340 1064.250 3381.480 2227.450 ;
        RECT 3384.290 2227.430 3385.260 2227.690 ;
      LAYER via ;
        RECT 3381.220 2227.480 3381.480 2227.740 ;
        RECT 3384.350 2227.430 3385.200 2227.690 ;
      LAYER met2 ;
        RECT 3381.190 2227.620 3381.510 2227.740 ;
        RECT 3384.350 2227.620 3385.200 2227.720 ;
        RECT 3377.950 2227.480 3385.200 2227.620 ;
        RECT 3384.350 2227.400 3385.200 2227.480 ;
    END
  END mgmt_io_in_buf[12]
  PIN mgmt_io_in_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2223.935 3384.490 2224.105 ;
        RECT 3384.320 2223.265 3384.490 2223.935 ;
        RECT 3383.840 2223.095 3384.490 2223.265 ;
        RECT 3384.320 2222.425 3384.490 2223.095 ;
        RECT 3383.840 2222.255 3384.490 2222.425 ;
        RECT 3384.320 2221.670 3384.490 2222.255 ;
        RECT 3385.030 2223.935 3386.050 2224.105 ;
        RECT 3385.030 2223.265 3385.200 2223.935 ;
        RECT 3385.030 2223.095 3386.050 2223.265 ;
        RECT 3385.030 2222.425 3385.200 2223.095 ;
        RECT 3385.030 2222.255 3386.050 2222.425 ;
        RECT 3385.030 2221.670 3385.200 2222.255 ;
        RECT 3384.320 2221.585 3385.200 2221.670 ;
        RECT 3383.840 2221.415 3386.050 2221.585 ;
      LAYER mcon ;
        RECT 3384.350 2221.500 3385.200 2221.670 ;
      LAYER met1 ;
        RECT 3380.660 2221.470 3380.920 2221.790 ;
        RECT 3380.780 1066.250 3380.920 2221.470 ;
        RECT 3384.290 2221.450 3385.260 2221.710 ;
      LAYER via ;
        RECT 3380.660 2221.500 3380.920 2221.760 ;
        RECT 3384.350 2221.450 3385.200 2221.710 ;
      LAYER met2 ;
        RECT 3380.630 2221.640 3380.950 2221.760 ;
        RECT 3384.350 2221.640 3385.200 2221.740 ;
        RECT 3377.950 2221.500 3385.200 2221.640 ;
        RECT 3384.350 2221.420 3385.200 2221.500 ;
    END
  END mgmt_io_in_buf[11]
  PIN mgmt_io_in_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2217.955 3384.490 2218.125 ;
        RECT 3384.320 2217.285 3384.490 2217.955 ;
        RECT 3383.840 2217.115 3384.490 2217.285 ;
        RECT 3384.320 2216.445 3384.490 2217.115 ;
        RECT 3383.840 2216.275 3384.490 2216.445 ;
        RECT 3384.320 2215.690 3384.490 2216.275 ;
        RECT 3385.030 2217.955 3386.050 2218.125 ;
        RECT 3385.030 2217.285 3385.200 2217.955 ;
        RECT 3385.030 2217.115 3386.050 2217.285 ;
        RECT 3385.030 2216.445 3385.200 2217.115 ;
        RECT 3385.030 2216.275 3386.050 2216.445 ;
        RECT 3385.030 2215.690 3385.200 2216.275 ;
        RECT 3384.320 2215.605 3385.200 2215.690 ;
        RECT 3383.840 2215.435 3386.050 2215.605 ;
      LAYER mcon ;
        RECT 3384.350 2215.520 3385.200 2215.690 ;
      LAYER met1 ;
        RECT 3380.100 2215.490 3380.360 2215.810 ;
        RECT 3380.220 1068.250 3380.360 2215.490 ;
        RECT 3384.290 2215.470 3385.260 2215.730 ;
      LAYER via ;
        RECT 3380.100 2215.520 3380.360 2215.780 ;
        RECT 3384.350 2215.470 3385.200 2215.730 ;
      LAYER met2 ;
        RECT 3380.070 2215.660 3380.390 2215.780 ;
        RECT 3384.350 2215.660 3385.200 2215.760 ;
        RECT 3377.950 2215.520 3385.200 2215.660 ;
        RECT 3384.350 2215.440 3385.200 2215.520 ;
    END
  END mgmt_io_in_buf[10]
  PIN mgmt_io_in_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2211.975 3384.490 2212.145 ;
        RECT 3384.320 2211.305 3384.490 2211.975 ;
        RECT 3383.840 2211.135 3384.490 2211.305 ;
        RECT 3384.320 2210.465 3384.490 2211.135 ;
        RECT 3383.840 2210.295 3384.490 2210.465 ;
        RECT 3384.320 2209.710 3384.490 2210.295 ;
        RECT 3385.030 2211.975 3386.050 2212.145 ;
        RECT 3385.030 2211.305 3385.200 2211.975 ;
        RECT 3385.030 2211.135 3386.050 2211.305 ;
        RECT 3385.030 2210.465 3385.200 2211.135 ;
        RECT 3385.030 2210.295 3386.050 2210.465 ;
        RECT 3385.030 2209.710 3385.200 2210.295 ;
        RECT 3384.320 2209.625 3385.200 2209.710 ;
        RECT 3383.840 2209.455 3386.050 2209.625 ;
      LAYER mcon ;
        RECT 3384.350 2209.540 3385.200 2209.710 ;
      LAYER met1 ;
        RECT 3379.540 2209.510 3379.800 2209.830 ;
        RECT 3379.660 1070.250 3379.800 2209.510 ;
        RECT 3384.290 2209.490 3385.260 2209.750 ;
      LAYER via ;
        RECT 3379.540 2209.540 3379.800 2209.800 ;
        RECT 3384.350 2209.490 3385.200 2209.750 ;
      LAYER met2 ;
        RECT 3379.510 2209.680 3379.830 2209.800 ;
        RECT 3384.350 2209.680 3385.200 2209.780 ;
        RECT 3377.950 2209.540 3385.200 2209.680 ;
        RECT 3384.350 2209.460 3385.200 2209.540 ;
    END
  END mgmt_io_in_buf[9]
  PIN mgmt_io_in_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2205.995 3384.490 2206.165 ;
        RECT 3384.320 2205.325 3384.490 2205.995 ;
        RECT 3383.840 2205.155 3384.490 2205.325 ;
        RECT 3384.320 2204.485 3384.490 2205.155 ;
        RECT 3383.840 2204.315 3384.490 2204.485 ;
        RECT 3384.320 2203.730 3384.490 2204.315 ;
        RECT 3385.030 2205.995 3386.050 2206.165 ;
        RECT 3385.030 2205.325 3385.200 2205.995 ;
        RECT 3385.030 2205.155 3386.050 2205.325 ;
        RECT 3385.030 2204.485 3385.200 2205.155 ;
        RECT 3385.030 2204.315 3386.050 2204.485 ;
        RECT 3385.030 2203.730 3385.200 2204.315 ;
        RECT 3384.320 2203.645 3385.200 2203.730 ;
        RECT 3383.840 2203.475 3386.050 2203.645 ;
      LAYER mcon ;
        RECT 3384.350 2203.560 3385.200 2203.730 ;
      LAYER met1 ;
        RECT 3378.980 2203.530 3379.240 2203.850 ;
        RECT 3379.100 1072.250 3379.240 2203.530 ;
        RECT 3384.290 2203.510 3385.260 2203.770 ;
      LAYER via ;
        RECT 3378.980 2203.560 3379.240 2203.820 ;
        RECT 3384.350 2203.510 3385.200 2203.770 ;
      LAYER met2 ;
        RECT 3378.950 2203.700 3379.270 2203.820 ;
        RECT 3384.350 2203.700 3385.200 2203.800 ;
        RECT 3377.950 2203.560 3385.200 2203.700 ;
        RECT 3384.350 2203.480 3385.200 2203.560 ;
    END
  END mgmt_io_in_buf[8]
  PIN mgmt_io_in_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2200.015 3384.490 2200.185 ;
        RECT 3384.320 2199.345 3384.490 2200.015 ;
        RECT 3383.840 2199.175 3384.490 2199.345 ;
        RECT 3384.320 2198.505 3384.490 2199.175 ;
        RECT 3383.840 2198.335 3384.490 2198.505 ;
        RECT 3384.320 2197.750 3384.490 2198.335 ;
        RECT 3385.030 2200.015 3386.050 2200.185 ;
        RECT 3385.030 2199.345 3385.200 2200.015 ;
        RECT 3385.030 2199.175 3386.050 2199.345 ;
        RECT 3385.030 2198.505 3385.200 2199.175 ;
        RECT 3385.030 2198.335 3386.050 2198.505 ;
        RECT 3385.030 2197.750 3385.200 2198.335 ;
        RECT 3384.320 2197.665 3385.200 2197.750 ;
        RECT 3383.840 2197.495 3386.050 2197.665 ;
      LAYER mcon ;
        RECT 3384.350 2197.580 3385.200 2197.750 ;
      LAYER met1 ;
        RECT 3378.420 2197.550 3378.680 2197.870 ;
        RECT 3378.540 1074.250 3378.680 2197.550 ;
        RECT 3384.290 2197.530 3385.260 2197.790 ;
      LAYER via ;
        RECT 3378.420 2197.580 3378.680 2197.840 ;
        RECT 3384.350 2197.530 3385.200 2197.790 ;
      LAYER met2 ;
        RECT 3378.390 2197.720 3378.710 2197.840 ;
        RECT 3384.350 2197.720 3385.200 2197.820 ;
        RECT 3377.950 2197.580 3385.200 2197.720 ;
        RECT 3384.350 2197.500 3385.200 2197.580 ;
    END
  END mgmt_io_in_buf[7]
  PIN mgmt_io_out_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3022.465 201.235 3022.635 ;
        RECT 199.505 3022.380 200.385 3022.465 ;
        RECT 199.505 3021.795 199.675 3022.380 ;
        RECT 199.025 3021.625 199.675 3021.795 ;
        RECT 199.505 3020.955 199.675 3021.625 ;
        RECT 199.025 3020.785 199.675 3020.955 ;
        RECT 199.505 3020.115 199.675 3020.785 ;
        RECT 199.025 3019.945 199.675 3020.115 ;
        RECT 200.215 3021.795 200.385 3022.380 ;
        RECT 200.215 3021.625 201.235 3021.795 ;
        RECT 200.215 3020.955 200.385 3021.625 ;
        RECT 200.215 3020.785 201.235 3020.955 ;
        RECT 200.215 3020.115 200.385 3020.785 ;
        RECT 200.215 3019.945 201.235 3020.115 ;
      LAYER mcon ;
        RECT 199.535 3022.380 200.385 3022.550 ;
      LAYER met1 ;
        RECT 206.295 3022.685 206.435 3066.780 ;
        RECT 199.475 3022.330 200.445 3022.590 ;
        RECT 206.175 3022.365 206.435 3022.685 ;
      LAYER via ;
        RECT 199.535 3022.330 200.385 3022.590 ;
        RECT 206.175 3022.395 206.435 3022.655 ;
      LAYER met2 ;
        RECT 199.535 3022.535 200.385 3022.620 ;
        RECT 206.145 3022.535 206.465 3022.655 ;
        RECT 199.535 3022.395 209.300 3022.535 ;
        RECT 199.535 3022.300 200.385 3022.395 ;
    END
  END mgmt_io_out_buf[24]
  PIN mgmt_io_out_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3016.485 201.235 3016.655 ;
        RECT 199.505 3016.400 200.385 3016.485 ;
        RECT 199.505 3015.815 199.675 3016.400 ;
        RECT 199.025 3015.645 199.675 3015.815 ;
        RECT 199.505 3014.975 199.675 3015.645 ;
        RECT 199.025 3014.805 199.675 3014.975 ;
        RECT 199.505 3014.135 199.675 3014.805 ;
        RECT 199.025 3013.965 199.675 3014.135 ;
        RECT 200.215 3015.815 200.385 3016.400 ;
        RECT 200.215 3015.645 201.235 3015.815 ;
        RECT 200.215 3014.975 200.385 3015.645 ;
        RECT 200.215 3014.805 201.235 3014.975 ;
        RECT 200.215 3014.135 200.385 3014.805 ;
        RECT 200.215 3013.965 201.235 3014.135 ;
      LAYER mcon ;
        RECT 199.535 3016.400 200.385 3016.570 ;
      LAYER met1 ;
        RECT 206.855 3016.705 206.995 3064.780 ;
        RECT 199.475 3016.350 200.445 3016.610 ;
        RECT 206.735 3016.385 206.995 3016.705 ;
      LAYER via ;
        RECT 199.535 3016.350 200.385 3016.610 ;
        RECT 206.735 3016.415 206.995 3016.675 ;
      LAYER met2 ;
        RECT 199.535 3016.555 200.385 3016.640 ;
        RECT 206.705 3016.555 207.025 3016.675 ;
        RECT 199.535 3016.415 209.300 3016.555 ;
        RECT 199.535 3016.320 200.385 3016.415 ;
    END
  END mgmt_io_out_buf[25]
  PIN mgmt_io_out_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3010.505 201.235 3010.675 ;
        RECT 199.505 3010.420 200.385 3010.505 ;
        RECT 199.505 3009.835 199.675 3010.420 ;
        RECT 199.025 3009.665 199.675 3009.835 ;
        RECT 199.505 3008.995 199.675 3009.665 ;
        RECT 199.025 3008.825 199.675 3008.995 ;
        RECT 199.505 3008.155 199.675 3008.825 ;
        RECT 199.025 3007.985 199.675 3008.155 ;
        RECT 200.215 3009.835 200.385 3010.420 ;
        RECT 200.215 3009.665 201.235 3009.835 ;
        RECT 200.215 3008.995 200.385 3009.665 ;
        RECT 200.215 3008.825 201.235 3008.995 ;
        RECT 200.215 3008.155 200.385 3008.825 ;
        RECT 200.215 3007.985 201.235 3008.155 ;
      LAYER mcon ;
        RECT 199.535 3010.420 200.385 3010.590 ;
      LAYER met1 ;
        RECT 207.415 3010.725 207.555 3062.780 ;
        RECT 199.475 3010.370 200.445 3010.630 ;
        RECT 207.295 3010.405 207.555 3010.725 ;
      LAYER via ;
        RECT 199.535 3010.370 200.385 3010.630 ;
        RECT 207.295 3010.435 207.555 3010.695 ;
      LAYER met2 ;
        RECT 199.535 3010.575 200.385 3010.660 ;
        RECT 207.265 3010.575 207.585 3010.695 ;
        RECT 199.535 3010.435 209.300 3010.575 ;
        RECT 199.535 3010.340 200.385 3010.435 ;
    END
  END mgmt_io_out_buf[26]
  PIN mgmt_io_out_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3004.525 201.235 3004.695 ;
        RECT 199.505 3004.440 200.385 3004.525 ;
        RECT 199.505 3003.855 199.675 3004.440 ;
        RECT 199.025 3003.685 199.675 3003.855 ;
        RECT 199.505 3003.015 199.675 3003.685 ;
        RECT 199.025 3002.845 199.675 3003.015 ;
        RECT 199.505 3002.175 199.675 3002.845 ;
        RECT 199.025 3002.005 199.675 3002.175 ;
        RECT 200.215 3003.855 200.385 3004.440 ;
        RECT 200.215 3003.685 201.235 3003.855 ;
        RECT 200.215 3003.015 200.385 3003.685 ;
        RECT 200.215 3002.845 201.235 3003.015 ;
        RECT 200.215 3002.175 200.385 3002.845 ;
        RECT 200.215 3002.005 201.235 3002.175 ;
      LAYER mcon ;
        RECT 199.535 3004.440 200.385 3004.610 ;
      LAYER met1 ;
        RECT 207.975 3004.745 208.115 3060.780 ;
        RECT 199.475 3004.390 200.445 3004.650 ;
        RECT 207.855 3004.425 208.115 3004.745 ;
      LAYER via ;
        RECT 199.535 3004.390 200.385 3004.650 ;
        RECT 207.855 3004.455 208.115 3004.715 ;
      LAYER met2 ;
        RECT 199.535 3004.595 200.385 3004.680 ;
        RECT 207.825 3004.595 208.145 3004.715 ;
        RECT 199.535 3004.455 209.300 3004.595 ;
        RECT 199.535 3004.360 200.385 3004.455 ;
    END
  END mgmt_io_out_buf[27]
  PIN mgmt_io_out_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 2998.545 201.235 2998.715 ;
        RECT 199.505 2998.460 200.385 2998.545 ;
        RECT 199.505 2997.875 199.675 2998.460 ;
        RECT 199.025 2997.705 199.675 2997.875 ;
        RECT 199.505 2997.035 199.675 2997.705 ;
        RECT 199.025 2996.865 199.675 2997.035 ;
        RECT 199.505 2996.195 199.675 2996.865 ;
        RECT 199.025 2996.025 199.675 2996.195 ;
        RECT 200.215 2997.875 200.385 2998.460 ;
        RECT 200.215 2997.705 201.235 2997.875 ;
        RECT 200.215 2997.035 200.385 2997.705 ;
        RECT 200.215 2996.865 201.235 2997.035 ;
        RECT 200.215 2996.195 200.385 2996.865 ;
        RECT 200.215 2996.025 201.235 2996.195 ;
      LAYER mcon ;
        RECT 199.535 2998.460 200.385 2998.630 ;
      LAYER met1 ;
        RECT 208.535 2998.765 208.675 3058.780 ;
        RECT 199.475 2998.410 200.445 2998.670 ;
        RECT 208.415 2998.445 208.675 2998.765 ;
      LAYER via ;
        RECT 199.535 2998.410 200.385 2998.670 ;
        RECT 208.415 2998.475 208.675 2998.735 ;
      LAYER met2 ;
        RECT 199.535 2998.615 200.385 2998.700 ;
        RECT 208.385 2998.615 208.705 2998.735 ;
        RECT 199.535 2998.475 209.300 2998.615 ;
        RECT 199.535 2998.380 200.385 2998.475 ;
    END
  END mgmt_io_out_buf[28]
  PIN mgmt_io_out_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 2992.565 201.235 2992.735 ;
        RECT 199.505 2992.480 200.385 2992.565 ;
        RECT 199.505 2991.895 199.675 2992.480 ;
        RECT 199.025 2991.725 199.675 2991.895 ;
        RECT 199.505 2991.055 199.675 2991.725 ;
        RECT 199.025 2990.885 199.675 2991.055 ;
        RECT 199.505 2990.215 199.675 2990.885 ;
        RECT 199.025 2990.045 199.675 2990.215 ;
        RECT 200.215 2991.895 200.385 2992.480 ;
        RECT 200.215 2991.725 201.235 2991.895 ;
        RECT 200.215 2991.055 200.385 2991.725 ;
        RECT 200.215 2990.885 201.235 2991.055 ;
        RECT 200.215 2990.215 200.385 2990.885 ;
        RECT 200.215 2990.045 201.235 2990.215 ;
      LAYER mcon ;
        RECT 199.535 2992.480 200.385 2992.650 ;
      LAYER met1 ;
        RECT 209.095 2992.785 209.235 3056.780 ;
        RECT 199.475 2992.430 200.445 2992.690 ;
        RECT 208.975 2992.465 209.235 2992.785 ;
      LAYER via ;
        RECT 199.535 2992.430 200.385 2992.690 ;
        RECT 208.975 2992.495 209.235 2992.755 ;
      LAYER met2 ;
        RECT 199.535 2992.635 200.385 2992.720 ;
        RECT 208.945 2992.635 209.265 2992.755 ;
        RECT 199.535 2992.495 209.300 2992.635 ;
        RECT 199.535 2992.400 200.385 2992.495 ;
    END
  END mgmt_io_out_buf[29]
  PIN mgmt_io_in_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 2992.470 203.135 2994.060 ;
      LAYER mcon ;
        RECT 202.935 2992.970 203.105 2994.060 ;
      LAYER met1 ;
        RECT 202.895 2992.910 203.155 2994.120 ;
        RECT 208.815 2993.755 208.955 3057.780 ;
        RECT 208.695 2993.435 208.955 2993.755 ;
      LAYER via ;
        RECT 202.895 2992.970 203.155 2994.060 ;
        RECT 208.695 2993.465 208.955 2993.725 ;
      LAYER met2 ;
        RECT 202.865 2993.605 203.185 2994.060 ;
        RECT 208.665 2993.605 208.985 2993.725 ;
        RECT 202.865 2993.465 209.300 2993.605 ;
        RECT 202.865 2992.970 203.185 2993.465 ;
    END
  END mgmt_io_in_unbuf[29]
  PIN mgmt_io_in_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 2998.450 203.135 3000.040 ;
      LAYER mcon ;
        RECT 202.935 2998.950 203.105 3000.040 ;
      LAYER met1 ;
        RECT 202.895 2998.890 203.155 3000.100 ;
        RECT 208.255 2999.735 208.395 3059.780 ;
        RECT 208.135 2999.415 208.395 2999.735 ;
      LAYER via ;
        RECT 202.895 2998.950 203.155 3000.040 ;
        RECT 208.135 2999.445 208.395 2999.705 ;
      LAYER met2 ;
        RECT 202.865 2999.585 203.185 3000.040 ;
        RECT 208.105 2999.585 208.425 2999.705 ;
        RECT 202.865 2999.445 209.300 2999.585 ;
        RECT 202.865 2998.950 203.185 2999.445 ;
    END
  END mgmt_io_in_unbuf[28]
  PIN mgmt_io_in_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3004.430 203.135 3006.020 ;
      LAYER mcon ;
        RECT 202.935 3004.930 203.105 3006.020 ;
      LAYER met1 ;
        RECT 202.895 3004.870 203.155 3006.080 ;
        RECT 207.695 3005.715 207.835 3061.780 ;
        RECT 207.575 3005.395 207.835 3005.715 ;
      LAYER via ;
        RECT 202.895 3004.930 203.155 3006.020 ;
        RECT 207.575 3005.425 207.835 3005.685 ;
      LAYER met2 ;
        RECT 202.865 3005.565 203.185 3006.020 ;
        RECT 207.545 3005.565 207.865 3005.685 ;
        RECT 202.865 3005.425 209.300 3005.565 ;
        RECT 202.865 3004.930 203.185 3005.425 ;
    END
  END mgmt_io_in_unbuf[27]
  PIN mgmt_io_in_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3010.410 203.135 3012.000 ;
      LAYER mcon ;
        RECT 202.935 3010.910 203.105 3012.000 ;
      LAYER met1 ;
        RECT 202.895 3010.850 203.155 3012.060 ;
        RECT 207.135 3011.695 207.275 3063.780 ;
        RECT 207.015 3011.375 207.275 3011.695 ;
      LAYER via ;
        RECT 202.895 3010.910 203.155 3012.000 ;
        RECT 207.015 3011.405 207.275 3011.665 ;
      LAYER met2 ;
        RECT 202.865 3011.545 203.185 3012.000 ;
        RECT 206.985 3011.545 207.305 3011.665 ;
        RECT 202.865 3011.405 209.300 3011.545 ;
        RECT 202.865 3010.910 203.185 3011.405 ;
    END
  END mgmt_io_in_unbuf[26]
  PIN mgmt_io_in_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3016.390 203.135 3017.980 ;
      LAYER mcon ;
        RECT 202.935 3016.890 203.105 3017.980 ;
      LAYER met1 ;
        RECT 202.895 3016.830 203.155 3018.040 ;
        RECT 206.575 3017.675 206.715 3065.780 ;
        RECT 206.455 3017.355 206.715 3017.675 ;
      LAYER via ;
        RECT 202.895 3016.890 203.155 3017.980 ;
        RECT 206.455 3017.385 206.715 3017.645 ;
      LAYER met2 ;
        RECT 202.865 3017.525 203.185 3017.980 ;
        RECT 206.425 3017.525 206.745 3017.645 ;
        RECT 202.865 3017.385 209.300 3017.525 ;
        RECT 202.865 3016.890 203.185 3017.385 ;
    END
  END mgmt_io_in_unbuf[25]
  PIN mgmt_io_in_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3022.370 203.135 3023.960 ;
      LAYER mcon ;
        RECT 202.935 3022.870 203.105 3023.960 ;
      LAYER met1 ;
        RECT 202.895 3022.810 203.155 3024.020 ;
        RECT 206.015 3023.655 206.155 3067.780 ;
        RECT 205.895 3023.335 206.155 3023.655 ;
      LAYER via ;
        RECT 202.895 3022.870 203.155 3023.960 ;
        RECT 205.895 3023.365 206.155 3023.625 ;
      LAYER met2 ;
        RECT 202.865 3023.505 203.185 3023.960 ;
        RECT 205.865 3023.505 206.185 3023.625 ;
        RECT 202.865 3023.365 209.300 3023.505 ;
        RECT 202.865 3022.870 203.185 3023.365 ;
    END
  END mgmt_io_in_unbuf[24]
  PIN mgmt_io_out_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1695.680 201.345 1695.850 ;
        RECT 199.615 1695.595 200.495 1695.680 ;
        RECT 199.615 1695.010 199.785 1695.595 ;
        RECT 199.135 1694.840 199.785 1695.010 ;
        RECT 199.615 1694.170 199.785 1694.840 ;
        RECT 199.135 1694.000 199.785 1694.170 ;
        RECT 199.615 1693.330 199.785 1694.000 ;
        RECT 199.135 1693.160 199.785 1693.330 ;
        RECT 200.325 1695.010 200.495 1695.595 ;
        RECT 200.325 1694.840 201.345 1695.010 ;
        RECT 200.325 1694.170 200.495 1694.840 ;
        RECT 200.325 1694.000 201.345 1694.170 ;
        RECT 200.325 1693.330 200.495 1694.000 ;
        RECT 200.325 1693.160 201.345 1693.330 ;
      LAYER mcon ;
        RECT 199.645 1695.595 200.495 1695.765 ;
      LAYER met1 ;
        RECT 209.515 1695.900 209.655 1772.650 ;
        RECT 199.585 1695.545 200.555 1695.805 ;
        RECT 209.395 1695.580 209.655 1695.900 ;
      LAYER via ;
        RECT 199.645 1695.545 200.495 1695.805 ;
        RECT 209.395 1695.610 209.655 1695.870 ;
      LAYER met2 ;
        RECT 199.645 1695.750 200.495 1695.835 ;
        RECT 209.365 1695.750 209.685 1695.870 ;
        RECT 199.645 1695.610 211.440 1695.750 ;
        RECT 199.645 1695.515 200.495 1695.610 ;
    END
  END mgmt_io_out_buf[30]
  PIN mgmt_io_out_buf[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1689.700 201.345 1689.870 ;
        RECT 199.615 1689.615 200.495 1689.700 ;
        RECT 199.615 1689.030 199.785 1689.615 ;
        RECT 199.135 1688.860 199.785 1689.030 ;
        RECT 199.615 1688.190 199.785 1688.860 ;
        RECT 199.135 1688.020 199.785 1688.190 ;
        RECT 199.615 1687.350 199.785 1688.020 ;
        RECT 199.135 1687.180 199.785 1687.350 ;
        RECT 200.325 1689.030 200.495 1689.615 ;
        RECT 200.325 1688.860 201.345 1689.030 ;
        RECT 200.325 1688.190 200.495 1688.860 ;
        RECT 200.325 1688.020 201.345 1688.190 ;
        RECT 200.325 1687.350 200.495 1688.020 ;
        RECT 200.325 1687.180 201.345 1687.350 ;
      LAYER mcon ;
        RECT 199.645 1689.615 200.495 1689.785 ;
      LAYER met1 ;
        RECT 210.075 1689.920 210.215 1770.650 ;
        RECT 199.585 1689.565 200.555 1689.825 ;
        RECT 209.955 1689.600 210.215 1689.920 ;
      LAYER via ;
        RECT 199.645 1689.565 200.495 1689.825 ;
        RECT 209.955 1689.630 210.215 1689.890 ;
      LAYER met2 ;
        RECT 199.645 1689.770 200.495 1689.855 ;
        RECT 209.925 1689.770 210.245 1689.890 ;
        RECT 199.645 1689.630 211.440 1689.770 ;
        RECT 199.645 1689.535 200.495 1689.630 ;
    END
  END mgmt_io_out_buf[31]
  PIN mgmt_io_out_buf[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1683.720 201.345 1683.890 ;
        RECT 199.615 1683.635 200.495 1683.720 ;
        RECT 199.615 1683.050 199.785 1683.635 ;
        RECT 199.135 1682.880 199.785 1683.050 ;
        RECT 199.615 1682.210 199.785 1682.880 ;
        RECT 199.135 1682.040 199.785 1682.210 ;
        RECT 199.615 1681.370 199.785 1682.040 ;
        RECT 199.135 1681.200 199.785 1681.370 ;
        RECT 200.325 1683.050 200.495 1683.635 ;
        RECT 200.325 1682.880 201.345 1683.050 ;
        RECT 200.325 1682.210 200.495 1682.880 ;
        RECT 200.325 1682.040 201.345 1682.210 ;
        RECT 200.325 1681.370 200.495 1682.040 ;
        RECT 200.325 1681.200 201.345 1681.370 ;
      LAYER mcon ;
        RECT 199.645 1683.635 200.495 1683.805 ;
      LAYER met1 ;
        RECT 210.635 1683.940 210.775 1768.650 ;
        RECT 199.585 1683.585 200.555 1683.845 ;
        RECT 210.515 1683.620 210.775 1683.940 ;
      LAYER via ;
        RECT 199.645 1683.585 200.495 1683.845 ;
        RECT 210.515 1683.650 210.775 1683.910 ;
      LAYER met2 ;
        RECT 199.645 1683.790 200.495 1683.875 ;
        RECT 210.485 1683.790 210.805 1683.910 ;
        RECT 199.645 1683.650 211.440 1683.790 ;
        RECT 199.645 1683.555 200.495 1683.650 ;
    END
  END mgmt_io_out_buf[32]
  PIN mgmt_io_out_buf[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1677.740 201.345 1677.910 ;
        RECT 199.615 1677.655 200.495 1677.740 ;
        RECT 199.615 1677.070 199.785 1677.655 ;
        RECT 199.135 1676.900 199.785 1677.070 ;
        RECT 199.615 1676.230 199.785 1676.900 ;
        RECT 199.135 1676.060 199.785 1676.230 ;
        RECT 199.615 1675.390 199.785 1676.060 ;
        RECT 199.135 1675.220 199.785 1675.390 ;
        RECT 200.325 1677.070 200.495 1677.655 ;
        RECT 200.325 1676.900 201.345 1677.070 ;
        RECT 200.325 1676.230 200.495 1676.900 ;
        RECT 200.325 1676.060 201.345 1676.230 ;
        RECT 200.325 1675.390 200.495 1676.060 ;
        RECT 200.325 1675.220 201.345 1675.390 ;
      LAYER mcon ;
        RECT 199.645 1677.655 200.495 1677.825 ;
      LAYER met1 ;
        RECT 211.195 1677.960 211.335 1766.650 ;
        RECT 199.585 1677.605 200.555 1677.865 ;
        RECT 211.075 1677.640 211.335 1677.960 ;
      LAYER via ;
        RECT 199.645 1677.605 200.495 1677.865 ;
        RECT 211.075 1677.670 211.335 1677.930 ;
      LAYER met2 ;
        RECT 199.645 1677.810 200.495 1677.895 ;
        RECT 211.045 1677.810 211.365 1677.930 ;
        RECT 199.645 1677.670 211.440 1677.810 ;
        RECT 199.645 1677.575 200.495 1677.670 ;
    END
  END mgmt_io_out_buf[33]
  PIN mgmt_io_in_unbuf[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1677.645 203.245 1679.235 ;
      LAYER mcon ;
        RECT 203.045 1678.145 203.215 1679.235 ;
      LAYER met1 ;
        RECT 203.005 1678.085 203.265 1679.295 ;
        RECT 210.915 1678.930 211.055 1767.650 ;
        RECT 210.795 1678.610 211.055 1678.930 ;
      LAYER via ;
        RECT 203.005 1678.145 203.265 1679.235 ;
        RECT 210.795 1678.640 211.055 1678.900 ;
      LAYER met2 ;
        RECT 202.975 1678.780 203.295 1679.235 ;
        RECT 210.765 1678.780 211.085 1678.900 ;
        RECT 202.975 1678.640 211.440 1678.780 ;
        RECT 202.975 1678.145 203.295 1678.640 ;
    END
  END mgmt_io_in_unbuf[33]
  PIN mgmt_io_in_unbuf[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1683.625 203.245 1685.215 ;
      LAYER mcon ;
        RECT 203.045 1684.125 203.215 1685.215 ;
      LAYER met1 ;
        RECT 203.005 1684.065 203.265 1685.275 ;
        RECT 210.355 1684.790 210.495 1769.650 ;
        RECT 210.235 1684.470 210.495 1684.790 ;
      LAYER via ;
        RECT 203.005 1684.125 203.265 1685.215 ;
        RECT 210.235 1684.500 210.495 1684.760 ;
      LAYER met2 ;
        RECT 202.975 1684.760 203.295 1685.215 ;
        RECT 202.975 1684.620 211.440 1684.760 ;
        RECT 202.975 1684.125 203.295 1684.620 ;
        RECT 210.205 1684.500 210.525 1684.620 ;
    END
  END mgmt_io_in_unbuf[32]
  PIN mgmt_io_in_unbuf[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1689.605 203.245 1691.195 ;
      LAYER mcon ;
        RECT 203.045 1690.105 203.215 1691.195 ;
      LAYER met1 ;
        RECT 203.005 1690.045 203.265 1691.255 ;
        RECT 209.795 1690.890 209.935 1771.650 ;
        RECT 209.675 1690.570 209.935 1690.890 ;
      LAYER via ;
        RECT 203.005 1690.105 203.265 1691.195 ;
        RECT 209.675 1690.600 209.935 1690.860 ;
      LAYER met2 ;
        RECT 202.975 1690.740 203.295 1691.195 ;
        RECT 209.645 1690.740 209.965 1690.860 ;
        RECT 202.975 1690.600 211.440 1690.740 ;
        RECT 202.975 1690.105 203.295 1690.600 ;
    END
  END mgmt_io_in_unbuf[31]
  PIN mgmt_io_in_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1695.585 203.245 1697.175 ;
      LAYER mcon ;
        RECT 203.045 1696.085 203.215 1697.175 ;
      LAYER met1 ;
        RECT 203.005 1696.025 203.265 1697.235 ;
        RECT 209.235 1696.870 209.375 1773.650 ;
        RECT 209.115 1696.550 209.375 1696.870 ;
      LAYER via ;
        RECT 203.005 1696.085 203.265 1697.175 ;
        RECT 209.115 1696.580 209.375 1696.840 ;
      LAYER met2 ;
        RECT 202.975 1696.720 203.295 1697.175 ;
        RECT 209.085 1696.720 209.405 1696.840 ;
        RECT 202.975 1696.580 211.440 1696.720 ;
        RECT 202.975 1696.085 203.295 1696.580 ;
    END
  END mgmt_io_in_unbuf[30]
  PIN mgmt_io_out_buf[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 736.215 1116.390 736.385 1116.870 ;
        RECT 737.055 1116.390 737.225 1116.870 ;
        RECT 737.895 1116.390 738.065 1116.870 ;
        RECT 738.735 1116.390 738.905 1116.870 ;
        RECT 736.215 1116.220 738.905 1116.390 ;
        RECT 736.215 1115.680 736.470 1116.220 ;
        RECT 736.215 1115.510 738.905 1115.680 ;
        RECT 736.215 1114.660 736.385 1115.510 ;
        RECT 737.055 1114.660 737.225 1115.510 ;
        RECT 737.895 1114.660 738.065 1115.510 ;
        RECT 738.735 1114.660 738.905 1115.510 ;
      LAYER mcon ;
        RECT 736.300 1115.510 736.470 1116.360 ;
      LAYER met1 ;
        RECT 736.270 1120.980 736.590 1121.100 ;
        RECT 655.615 1120.840 736.590 1120.980 ;
        RECT 736.250 1115.450 736.510 1116.420 ;
      LAYER via ;
        RECT 736.300 1120.840 736.560 1121.100 ;
        RECT 736.250 1115.510 736.510 1116.360 ;
      LAYER met2 ;
        RECT 736.300 1121.130 736.440 1126.825 ;
        RECT 736.300 1120.810 736.560 1121.130 ;
        RECT 736.300 1116.360 736.440 1120.810 ;
        RECT 736.220 1115.510 736.540 1116.360 ;
    END
  END mgmt_io_out_buf[34]
  PIN mgmt_io_out_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 742.195 1116.390 742.365 1116.870 ;
        RECT 743.035 1116.390 743.205 1116.870 ;
        RECT 743.875 1116.390 744.045 1116.870 ;
        RECT 744.715 1116.390 744.885 1116.870 ;
        RECT 742.195 1116.220 744.885 1116.390 ;
        RECT 742.195 1115.680 742.450 1116.220 ;
        RECT 742.195 1115.510 744.885 1115.680 ;
        RECT 742.195 1114.660 742.365 1115.510 ;
        RECT 743.035 1114.660 743.205 1115.510 ;
        RECT 743.875 1114.660 744.045 1115.510 ;
        RECT 744.715 1114.660 744.885 1115.510 ;
      LAYER mcon ;
        RECT 742.280 1115.510 742.450 1116.360 ;
      LAYER met1 ;
        RECT 742.250 1120.420 742.570 1120.540 ;
        RECT 657.615 1120.280 742.570 1120.420 ;
        RECT 742.230 1115.450 742.490 1116.420 ;
      LAYER via ;
        RECT 742.280 1120.280 742.540 1120.540 ;
        RECT 742.230 1115.510 742.490 1116.360 ;
      LAYER met2 ;
        RECT 742.280 1120.570 742.420 1126.825 ;
        RECT 742.280 1120.250 742.540 1120.570 ;
        RECT 742.280 1116.360 742.420 1120.250 ;
        RECT 742.200 1115.510 742.520 1116.360 ;
    END
  END mgmt_io_out_buf[35]
  PIN mgmt_io_out_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 748.175 1116.390 748.345 1116.870 ;
        RECT 749.015 1116.390 749.185 1116.870 ;
        RECT 749.855 1116.390 750.025 1116.870 ;
        RECT 750.695 1116.390 750.865 1116.870 ;
        RECT 748.175 1116.220 750.865 1116.390 ;
        RECT 748.175 1115.680 748.430 1116.220 ;
        RECT 748.175 1115.510 750.865 1115.680 ;
        RECT 748.175 1114.660 748.345 1115.510 ;
        RECT 749.015 1114.660 749.185 1115.510 ;
        RECT 749.855 1114.660 750.025 1115.510 ;
        RECT 750.695 1114.660 750.865 1115.510 ;
      LAYER mcon ;
        RECT 748.260 1115.510 748.430 1116.360 ;
      LAYER met1 ;
        RECT 748.230 1119.860 748.550 1119.980 ;
        RECT 659.615 1119.720 748.550 1119.860 ;
        RECT 748.210 1115.450 748.470 1116.420 ;
      LAYER via ;
        RECT 748.260 1119.720 748.520 1119.980 ;
        RECT 748.210 1115.510 748.470 1116.360 ;
      LAYER met2 ;
        RECT 748.260 1120.010 748.400 1126.825 ;
        RECT 748.260 1119.690 748.520 1120.010 ;
        RECT 748.260 1116.360 748.400 1119.690 ;
        RECT 748.180 1115.510 748.500 1116.360 ;
    END
  END mgmt_io_out_buf[36]
  PIN mgmt_io_out_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 754.155 1116.390 754.325 1116.870 ;
        RECT 754.995 1116.390 755.165 1116.870 ;
        RECT 755.835 1116.390 756.005 1116.870 ;
        RECT 756.675 1116.390 756.845 1116.870 ;
        RECT 754.155 1116.220 756.845 1116.390 ;
        RECT 754.155 1115.680 754.410 1116.220 ;
        RECT 754.155 1115.510 756.845 1115.680 ;
        RECT 754.155 1114.660 754.325 1115.510 ;
        RECT 754.995 1114.660 755.165 1115.510 ;
        RECT 755.835 1114.660 756.005 1115.510 ;
        RECT 756.675 1114.660 756.845 1115.510 ;
      LAYER mcon ;
        RECT 754.240 1115.510 754.410 1116.360 ;
      LAYER met1 ;
        RECT 754.210 1119.300 754.530 1119.420 ;
        RECT 661.615 1119.160 754.530 1119.300 ;
        RECT 754.190 1115.450 754.450 1116.420 ;
      LAYER via ;
        RECT 754.240 1119.160 754.500 1119.420 ;
        RECT 754.190 1115.510 754.450 1116.360 ;
      LAYER met2 ;
        RECT 754.240 1119.450 754.380 1126.825 ;
        RECT 754.240 1119.130 754.500 1119.450 ;
        RECT 754.240 1116.360 754.380 1119.130 ;
        RECT 754.160 1115.510 754.480 1116.360 ;
    END
  END mgmt_io_out_buf[37]
  PIN mgmt_io_in_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 759.300 1112.760 760.400 1112.960 ;
      LAYER mcon ;
        RECT 759.310 1112.790 760.400 1112.960 ;
      LAYER met1 ;
        RECT 759.570 1119.020 759.890 1119.140 ;
        RECT 662.615 1118.880 759.890 1119.020 ;
        RECT 759.250 1112.750 760.460 1113.010 ;
      LAYER via ;
        RECT 759.600 1118.880 759.860 1119.140 ;
        RECT 759.310 1112.750 760.400 1113.010 ;
      LAYER met2 ;
        RECT 759.600 1119.170 759.740 1126.825 ;
        RECT 759.600 1118.850 759.860 1119.170 ;
        RECT 759.600 1113.040 759.740 1118.850 ;
        RECT 759.310 1112.720 760.400 1113.040 ;
    END
  END mgmt_io_in_unbuf[37]
  PIN mgmt_io_in_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 753.320 1112.760 754.420 1112.960 ;
      LAYER mcon ;
        RECT 753.330 1112.790 754.420 1112.960 ;
      LAYER met1 ;
        RECT 753.590 1119.580 753.910 1119.700 ;
        RECT 660.615 1119.440 753.910 1119.580 ;
        RECT 753.270 1112.750 754.480 1113.010 ;
      LAYER via ;
        RECT 753.620 1119.440 753.880 1119.700 ;
        RECT 753.330 1112.750 754.420 1113.010 ;
      LAYER met2 ;
        RECT 753.620 1119.730 753.760 1126.825 ;
        RECT 753.620 1119.410 753.880 1119.730 ;
        RECT 753.620 1113.040 753.760 1119.410 ;
        RECT 753.330 1112.720 754.420 1113.040 ;
    END
  END mgmt_io_in_unbuf[36]
  PIN mgmt_io_in_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 747.340 1112.760 748.440 1112.960 ;
      LAYER mcon ;
        RECT 747.350 1112.790 748.440 1112.960 ;
      LAYER met1 ;
        RECT 747.610 1120.140 747.930 1120.260 ;
        RECT 658.615 1120.000 747.930 1120.140 ;
        RECT 747.290 1112.750 748.500 1113.010 ;
      LAYER via ;
        RECT 747.640 1120.000 747.900 1120.260 ;
        RECT 747.350 1112.750 748.440 1113.010 ;
      LAYER met2 ;
        RECT 747.640 1120.290 747.780 1126.825 ;
        RECT 747.640 1119.970 747.900 1120.290 ;
        RECT 747.640 1113.040 747.780 1119.970 ;
        RECT 747.350 1112.720 748.440 1113.040 ;
    END
  END mgmt_io_in_unbuf[35]
  PIN mgmt_io_in_unbuf[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 741.360 1112.760 742.460 1112.960 ;
      LAYER mcon ;
        RECT 741.370 1112.790 742.460 1112.960 ;
      LAYER met1 ;
        RECT 741.630 1120.700 741.950 1120.820 ;
        RECT 656.615 1120.560 741.950 1120.700 ;
        RECT 741.310 1112.750 742.520 1113.010 ;
      LAYER via ;
        RECT 741.660 1120.560 741.920 1120.820 ;
        RECT 741.370 1112.750 742.460 1113.010 ;
      LAYER met2 ;
        RECT 741.660 1120.850 741.800 1126.825 ;
        RECT 741.660 1120.530 741.920 1120.850 ;
        RECT 741.660 1113.040 741.800 1120.530 ;
        RECT 741.370 1112.720 742.460 1113.040 ;
    END
  END mgmt_io_in_unbuf[34]
  PIN mgmt_io_oeb_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 760.135 1116.390 760.305 1116.870 ;
        RECT 760.975 1116.390 761.145 1116.870 ;
        RECT 761.815 1116.390 761.985 1116.870 ;
        RECT 762.655 1116.390 762.825 1116.870 ;
        RECT 760.135 1116.220 762.825 1116.390 ;
        RECT 760.135 1115.680 760.390 1116.220 ;
        RECT 760.135 1115.510 762.825 1115.680 ;
        RECT 760.135 1114.660 760.305 1115.510 ;
        RECT 760.975 1114.660 761.145 1115.510 ;
        RECT 761.815 1114.660 761.985 1115.510 ;
        RECT 762.655 1114.660 762.825 1115.510 ;
      LAYER mcon ;
        RECT 760.220 1115.510 760.390 1116.360 ;
      LAYER met1 ;
        RECT 760.190 1118.740 760.510 1118.860 ;
        RECT 663.615 1118.600 760.510 1118.740 ;
        RECT 760.170 1115.450 760.430 1116.420 ;
      LAYER via ;
        RECT 760.220 1118.600 760.480 1118.860 ;
        RECT 760.170 1115.510 760.430 1116.360 ;
      LAYER met2 ;
        RECT 760.220 1118.890 760.360 1126.825 ;
        RECT 760.220 1118.570 760.480 1118.890 ;
        RECT 760.220 1116.360 760.360 1118.570 ;
        RECT 760.140 1115.510 760.460 1116.360 ;
    END
  END mgmt_io_oeb_buf[35]
  PIN mgmt_io_oeb_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 766.115 1113.300 766.285 1114.150 ;
        RECT 766.955 1113.300 767.125 1114.150 ;
        RECT 767.795 1113.300 767.965 1114.150 ;
        RECT 768.635 1113.300 768.805 1114.150 ;
        RECT 766.115 1113.130 768.805 1113.300 ;
        RECT 766.115 1112.590 766.370 1113.130 ;
        RECT 766.115 1112.420 768.805 1112.590 ;
        RECT 766.115 1111.940 766.285 1112.420 ;
        RECT 766.955 1111.940 767.125 1112.420 ;
        RECT 767.795 1111.940 767.965 1112.420 ;
        RECT 768.635 1111.940 768.805 1112.420 ;
      LAYER mcon ;
        RECT 766.200 1112.450 766.370 1113.300 ;
      LAYER met1 ;
        RECT 765.550 1118.460 765.870 1118.580 ;
        RECT 664.615 1118.320 765.870 1118.460 ;
        RECT 766.160 1112.390 766.420 1113.360 ;
      LAYER via ;
        RECT 765.580 1118.320 765.840 1118.580 ;
        RECT 766.160 1112.450 766.420 1113.300 ;
      LAYER met2 ;
        RECT 765.580 1118.610 765.720 1126.825 ;
        RECT 765.580 1118.290 765.840 1118.610 ;
        RECT 765.580 1114.240 765.720 1118.290 ;
        RECT 765.580 1114.100 766.355 1114.240 ;
        RECT 766.215 1113.300 766.355 1114.100 ;
        RECT 766.130 1112.450 766.450 1113.300 ;
    END
  END mgmt_io_oeb_buf[36]
  PIN mgmt_io_oeb_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 766.115 1116.390 766.285 1116.870 ;
        RECT 766.955 1116.390 767.125 1116.870 ;
        RECT 767.795 1116.390 767.965 1116.870 ;
        RECT 768.635 1116.390 768.805 1116.870 ;
        RECT 766.115 1116.220 768.805 1116.390 ;
        RECT 766.115 1115.680 766.370 1116.220 ;
        RECT 766.115 1115.510 768.805 1115.680 ;
        RECT 766.115 1114.660 766.285 1115.510 ;
        RECT 766.955 1114.660 767.125 1115.510 ;
        RECT 767.795 1114.660 767.965 1115.510 ;
        RECT 768.635 1114.660 768.805 1115.510 ;
      LAYER mcon ;
        RECT 766.200 1115.510 766.370 1116.360 ;
      LAYER met1 ;
        RECT 766.170 1118.180 766.490 1118.300 ;
        RECT 665.615 1118.040 766.490 1118.180 ;
        RECT 766.150 1115.450 766.410 1116.420 ;
      LAYER via ;
        RECT 766.200 1118.040 766.460 1118.300 ;
        RECT 766.150 1115.510 766.410 1116.360 ;
      LAYER met2 ;
        RECT 766.200 1118.330 766.340 1126.825 ;
        RECT 766.200 1118.010 766.460 1118.330 ;
        RECT 766.200 1116.360 766.340 1118.010 ;
        RECT 766.120 1115.510 766.440 1116.360 ;
    END
  END mgmt_io_oeb_buf[37]
  PIN mgmt_io_oeb_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2069.420 1115.850 2071.010 1116.050 ;
      LAYER mcon ;
        RECT 2069.920 1115.850 2071.010 1116.020 ;
      LAYER met1 ;
        RECT 2070.385 1118.320 3369.440 1118.460 ;
        RECT 2070.385 1118.200 2070.705 1118.320 ;
        RECT 2069.860 1115.810 2071.070 1116.070 ;
        RECT 3369.300 1105.250 3369.440 1118.320 ;
      LAYER via ;
        RECT 2070.415 1118.200 2070.675 1118.460 ;
        RECT 2069.920 1115.810 2071.010 1116.070 ;
      LAYER met2 ;
        RECT 2070.415 1118.490 2070.555 1126.965 ;
        RECT 2070.415 1118.170 2070.675 1118.490 ;
        RECT 2070.415 1116.100 2070.555 1118.170 ;
        RECT 2069.920 1115.780 2071.010 1116.100 ;
    END
  END mgmt_io_oeb_unbuf[37]
  PIN mgmt_io_oeb_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2069.420 1112.760 2070.520 1112.960 ;
      LAYER mcon ;
        RECT 2069.420 1112.790 2070.510 1112.960 ;
      LAYER met1 ;
        RECT 2069.415 1118.600 3369.720 1118.740 ;
        RECT 2069.415 1118.480 2069.735 1118.600 ;
        RECT 2069.360 1112.750 2070.570 1113.010 ;
        RECT 3369.580 1104.250 3369.720 1118.600 ;
      LAYER via ;
        RECT 2069.445 1118.480 2069.705 1118.740 ;
        RECT 2069.420 1112.750 2070.510 1113.010 ;
      LAYER met2 ;
        RECT 2069.445 1118.770 2069.585 1126.965 ;
        RECT 2069.445 1118.450 2069.705 1118.770 ;
        RECT 2069.445 1114.170 2069.585 1118.450 ;
        RECT 2069.445 1114.030 2070.220 1114.170 ;
        RECT 2070.080 1113.040 2070.220 1114.030 ;
        RECT 2069.420 1112.720 2070.510 1113.040 ;
    END
  END mgmt_io_oeb_unbuf[36]
  PIN mgmt_io_oeb_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2063.440 1115.850 2065.030 1116.050 ;
      LAYER mcon ;
        RECT 2063.940 1115.850 2065.030 1116.020 ;
      LAYER met1 ;
        RECT 2064.285 1118.880 3370.000 1119.020 ;
        RECT 2064.285 1118.760 2064.605 1118.880 ;
        RECT 2063.880 1115.810 2065.090 1116.070 ;
        RECT 3369.860 1103.250 3370.000 1118.880 ;
      LAYER via ;
        RECT 2064.315 1118.760 2064.575 1119.020 ;
        RECT 2063.940 1115.810 2065.030 1116.070 ;
      LAYER met2 ;
        RECT 2064.435 1119.050 2064.575 1126.965 ;
        RECT 2064.315 1118.730 2064.575 1119.050 ;
        RECT 2064.435 1116.100 2064.575 1118.730 ;
        RECT 2063.940 1115.780 2065.030 1116.100 ;
    END
  END mgmt_io_oeb_unbuf[35]
  PIN mgmt_io_in_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2061.015 1113.300 2061.185 1114.150 ;
        RECT 2061.855 1113.300 2062.025 1114.150 ;
        RECT 2062.695 1113.300 2062.865 1114.150 ;
        RECT 2063.535 1113.300 2063.705 1114.150 ;
        RECT 2061.015 1113.130 2063.705 1113.300 ;
        RECT 2063.450 1112.590 2063.705 1113.130 ;
        RECT 2061.015 1112.420 2063.705 1112.590 ;
        RECT 2061.015 1111.940 2061.185 1112.420 ;
        RECT 2061.855 1111.940 2062.025 1112.420 ;
        RECT 2062.695 1111.940 2062.865 1112.420 ;
        RECT 2063.535 1111.940 2063.705 1112.420 ;
      LAYER mcon ;
        RECT 2063.450 1112.450 2063.620 1113.300 ;
      LAYER met1 ;
        RECT 2063.435 1119.160 3370.280 1119.300 ;
        RECT 2063.435 1119.040 2063.755 1119.160 ;
        RECT 2063.400 1112.390 2063.660 1113.360 ;
        RECT 3370.140 1102.250 3370.280 1119.160 ;
      LAYER via ;
        RECT 2063.465 1119.040 2063.725 1119.300 ;
        RECT 2063.400 1112.450 2063.660 1113.300 ;
      LAYER met2 ;
        RECT 2063.465 1119.330 2063.605 1126.965 ;
        RECT 2063.465 1119.010 2063.725 1119.330 ;
        RECT 2063.465 1113.300 2063.605 1119.010 ;
        RECT 2063.370 1112.450 2063.690 1113.300 ;
    END
  END mgmt_io_in_buf[37]
  PIN mgmt_io_in_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2055.035 1113.300 2055.205 1114.150 ;
        RECT 2055.875 1113.300 2056.045 1114.150 ;
        RECT 2056.715 1113.300 2056.885 1114.150 ;
        RECT 2057.555 1113.300 2057.725 1114.150 ;
        RECT 2055.035 1113.130 2057.725 1113.300 ;
        RECT 2057.470 1112.590 2057.725 1113.130 ;
        RECT 2055.035 1112.420 2057.725 1112.590 ;
        RECT 2055.035 1111.940 2055.205 1112.420 ;
        RECT 2055.875 1111.940 2056.045 1112.420 ;
        RECT 2056.715 1111.940 2056.885 1112.420 ;
        RECT 2057.555 1111.940 2057.725 1112.420 ;
      LAYER mcon ;
        RECT 2057.470 1112.450 2057.640 1113.300 ;
      LAYER met1 ;
        RECT 2057.455 1119.720 3370.840 1119.860 ;
        RECT 2057.455 1119.600 2057.775 1119.720 ;
        RECT 2057.420 1112.390 2057.680 1113.360 ;
        RECT 3370.700 1100.250 3370.840 1119.720 ;
      LAYER via ;
        RECT 2057.485 1119.600 2057.745 1119.860 ;
        RECT 2057.420 1112.450 2057.680 1113.300 ;
      LAYER met2 ;
        RECT 2057.485 1119.890 2057.625 1126.965 ;
        RECT 2057.485 1119.570 2057.745 1119.890 ;
        RECT 2057.485 1113.300 2057.625 1119.570 ;
        RECT 2057.390 1112.450 2057.710 1113.300 ;
    END
  END mgmt_io_in_buf[36]
  PIN mgmt_io_in_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2049.055 1113.300 2049.225 1114.150 ;
        RECT 2049.895 1113.300 2050.065 1114.150 ;
        RECT 2050.735 1113.300 2050.905 1114.150 ;
        RECT 2051.575 1113.300 2051.745 1114.150 ;
        RECT 2049.055 1113.130 2051.745 1113.300 ;
        RECT 2051.490 1112.590 2051.745 1113.130 ;
        RECT 2049.055 1112.420 2051.745 1112.590 ;
        RECT 2049.055 1111.940 2049.225 1112.420 ;
        RECT 2049.895 1111.940 2050.065 1112.420 ;
        RECT 2050.735 1111.940 2050.905 1112.420 ;
        RECT 2051.575 1111.940 2051.745 1112.420 ;
      LAYER mcon ;
        RECT 2051.490 1112.450 2051.660 1113.300 ;
      LAYER met1 ;
        RECT 2051.475 1120.280 3371.400 1120.420 ;
        RECT 2051.475 1120.160 2051.795 1120.280 ;
        RECT 2051.440 1112.390 2051.700 1113.360 ;
        RECT 3371.260 1098.250 3371.400 1120.280 ;
      LAYER via ;
        RECT 2051.505 1120.160 2051.765 1120.420 ;
        RECT 2051.440 1112.450 2051.700 1113.300 ;
      LAYER met2 ;
        RECT 2051.505 1120.450 2051.645 1126.965 ;
        RECT 2051.505 1120.130 2051.765 1120.450 ;
        RECT 2051.505 1113.300 2051.645 1120.130 ;
        RECT 2051.410 1112.450 2051.730 1113.300 ;
    END
  END mgmt_io_in_buf[35]
  PIN mgmt_io_in_buf[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2043.075 1113.300 2043.245 1114.150 ;
        RECT 2043.915 1113.300 2044.085 1114.150 ;
        RECT 2044.755 1113.300 2044.925 1114.150 ;
        RECT 2045.595 1113.300 2045.765 1114.150 ;
        RECT 2043.075 1113.130 2045.765 1113.300 ;
        RECT 2045.510 1112.590 2045.765 1113.130 ;
        RECT 2043.075 1112.420 2045.765 1112.590 ;
        RECT 2043.075 1111.940 2043.245 1112.420 ;
        RECT 2043.915 1111.940 2044.085 1112.420 ;
        RECT 2044.755 1111.940 2044.925 1112.420 ;
        RECT 2045.595 1111.940 2045.765 1112.420 ;
      LAYER mcon ;
        RECT 2045.510 1112.450 2045.680 1113.300 ;
      LAYER met1 ;
        RECT 2045.495 1120.840 3371.960 1120.980 ;
        RECT 2045.495 1120.720 2045.815 1120.840 ;
        RECT 2045.460 1112.390 2045.720 1113.360 ;
        RECT 3371.820 1096.250 3371.960 1120.840 ;
      LAYER via ;
        RECT 2045.525 1120.720 2045.785 1120.980 ;
        RECT 2045.460 1112.450 2045.720 1113.300 ;
      LAYER met2 ;
        RECT 2045.525 1121.010 2045.665 1126.965 ;
        RECT 2045.525 1120.690 2045.785 1121.010 ;
        RECT 2045.525 1113.300 2045.665 1120.690 ;
        RECT 2045.430 1112.450 2045.750 1113.300 ;
    END
  END mgmt_io_in_buf[34]
  PIN mgmt_io_out_unbuf[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2039.520 1115.850 2041.110 1116.050 ;
      LAYER mcon ;
        RECT 2040.020 1115.850 2041.110 1116.020 ;
      LAYER met1 ;
        RECT 2040.485 1121.120 3372.240 1121.260 ;
        RECT 2040.485 1121.000 2040.805 1121.120 ;
        RECT 2039.960 1115.810 2041.170 1116.070 ;
        RECT 3372.100 1095.250 3372.240 1121.120 ;
      LAYER via ;
        RECT 2040.515 1121.000 2040.775 1121.260 ;
        RECT 2040.020 1115.810 2041.110 1116.070 ;
      LAYER met2 ;
        RECT 2040.515 1121.290 2040.655 1126.965 ;
        RECT 2040.515 1120.970 2040.775 1121.290 ;
        RECT 2040.515 1116.100 2040.655 1120.970 ;
        RECT 2040.020 1115.780 2041.110 1116.100 ;
    END
  END mgmt_io_out_unbuf[34]
  PIN mgmt_io_out_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2045.500 1115.850 2047.090 1116.050 ;
      LAYER mcon ;
        RECT 2046.000 1115.850 2047.090 1116.020 ;
      LAYER met1 ;
        RECT 2046.465 1120.560 3371.680 1120.700 ;
        RECT 2046.465 1120.440 2046.785 1120.560 ;
        RECT 2045.940 1115.810 2047.150 1116.070 ;
        RECT 3371.540 1097.250 3371.680 1120.560 ;
      LAYER via ;
        RECT 2046.495 1120.440 2046.755 1120.700 ;
        RECT 2046.000 1115.810 2047.090 1116.070 ;
      LAYER met2 ;
        RECT 2046.495 1120.730 2046.635 1126.965 ;
        RECT 2046.495 1120.410 2046.755 1120.730 ;
        RECT 2046.495 1116.100 2046.635 1120.410 ;
        RECT 2046.000 1115.780 2047.090 1116.100 ;
    END
  END mgmt_io_out_unbuf[35]
  PIN mgmt_io_out_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2051.480 1115.850 2053.070 1116.050 ;
      LAYER mcon ;
        RECT 2051.980 1115.850 2053.070 1116.020 ;
      LAYER met1 ;
        RECT 2052.325 1120.000 3371.120 1120.140 ;
        RECT 2052.325 1119.880 2052.645 1120.000 ;
        RECT 2051.920 1115.810 2053.130 1116.070 ;
        RECT 3370.980 1099.250 3371.120 1120.000 ;
      LAYER via ;
        RECT 2052.355 1119.880 2052.615 1120.140 ;
        RECT 2051.980 1115.810 2053.070 1116.070 ;
      LAYER met2 ;
        RECT 2052.475 1120.170 2052.615 1126.965 ;
        RECT 2052.355 1119.850 2052.615 1120.170 ;
        RECT 2052.475 1116.100 2052.615 1119.850 ;
        RECT 2051.980 1115.780 2053.070 1116.100 ;
    END
  END mgmt_io_out_unbuf[36]
  PIN mgmt_io_out_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2057.460 1115.850 2059.050 1116.050 ;
      LAYER mcon ;
        RECT 2057.960 1115.850 2059.050 1116.020 ;
      LAYER met1 ;
        RECT 2058.425 1119.440 3370.560 1119.580 ;
        RECT 2058.425 1119.320 2058.745 1119.440 ;
        RECT 2057.900 1115.810 2059.110 1116.070 ;
        RECT 3370.420 1101.250 3370.560 1119.440 ;
      LAYER via ;
        RECT 2058.455 1119.320 2058.715 1119.580 ;
        RECT 2057.960 1115.810 2059.050 1116.070 ;
      LAYER met2 ;
        RECT 2058.455 1119.610 2058.595 1126.965 ;
        RECT 2058.455 1119.290 2058.715 1119.610 ;
        RECT 2058.455 1116.100 2058.595 1119.290 ;
        RECT 2057.960 1115.780 2059.050 1116.100 ;
    END
  END mgmt_io_out_unbuf[37]
  PIN mgmt_io_out_unbuf[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1973.740 1115.850 1975.330 1116.050 ;
      LAYER mcon ;
        RECT 1974.240 1115.850 1975.330 1116.020 ;
      LAYER met1 ;
        RECT 1974.705 1126.720 3377.840 1126.860 ;
        RECT 1974.705 1126.600 1975.025 1126.720 ;
        RECT 1974.180 1115.810 1975.390 1116.070 ;
        RECT 3377.700 1075.250 3377.840 1126.720 ;
      LAYER via ;
        RECT 1974.735 1126.600 1974.995 1126.860 ;
        RECT 1974.240 1115.810 1975.330 1116.070 ;
      LAYER met2 ;
        RECT 1974.735 1126.890 1974.875 1126.965 ;
        RECT 1974.735 1126.570 1974.995 1126.890 ;
        RECT 1974.735 1116.100 1974.875 1126.570 ;
        RECT 1974.240 1115.780 1975.330 1116.100 ;
    END
  END mgmt_io_out_unbuf[33]
  PIN mgmt_io_out_unbuf[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1979.720 1115.850 1981.310 1116.050 ;
      LAYER mcon ;
        RECT 1980.220 1115.850 1981.310 1116.020 ;
      LAYER met1 ;
        RECT 1980.685 1126.160 3377.280 1126.300 ;
        RECT 1980.685 1126.040 1981.005 1126.160 ;
        RECT 1980.160 1115.810 1981.370 1116.070 ;
        RECT 3377.140 1077.250 3377.280 1126.160 ;
      LAYER via ;
        RECT 1980.715 1126.040 1980.975 1126.300 ;
        RECT 1980.220 1115.810 1981.310 1116.070 ;
      LAYER met2 ;
        RECT 1980.715 1126.330 1980.855 1126.965 ;
        RECT 1980.715 1126.010 1980.975 1126.330 ;
        RECT 1980.715 1116.100 1980.855 1126.010 ;
        RECT 1980.220 1115.780 1981.310 1116.100 ;
    END
  END mgmt_io_out_unbuf[32]
  PIN mgmt_io_out_unbuf[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1985.700 1115.850 1987.290 1116.050 ;
      LAYER mcon ;
        RECT 1986.200 1115.850 1987.290 1116.020 ;
      LAYER met1 ;
        RECT 1986.665 1125.600 3376.720 1125.740 ;
        RECT 1986.665 1125.480 1986.985 1125.600 ;
        RECT 1986.140 1115.810 1987.350 1116.070 ;
        RECT 3376.580 1079.250 3376.720 1125.600 ;
      LAYER via ;
        RECT 1986.695 1125.480 1986.955 1125.740 ;
        RECT 1986.200 1115.810 1987.290 1116.070 ;
      LAYER met2 ;
        RECT 1986.695 1125.770 1986.835 1126.965 ;
        RECT 1986.695 1125.450 1986.955 1125.770 ;
        RECT 1986.695 1116.100 1986.835 1125.450 ;
        RECT 1986.200 1115.780 1987.290 1116.100 ;
    END
  END mgmt_io_out_unbuf[31]
  PIN mgmt_io_out_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1991.680 1115.850 1993.270 1116.050 ;
      LAYER mcon ;
        RECT 1992.180 1115.850 1993.270 1116.020 ;
      LAYER met1 ;
        RECT 1992.645 1125.040 3376.160 1125.180 ;
        RECT 1992.645 1124.920 1992.965 1125.040 ;
        RECT 1992.120 1115.810 1993.330 1116.070 ;
        RECT 3376.020 1081.250 3376.160 1125.040 ;
      LAYER via ;
        RECT 1992.675 1124.920 1992.935 1125.180 ;
        RECT 1992.180 1115.810 1993.270 1116.070 ;
      LAYER met2 ;
        RECT 1992.675 1125.210 1992.815 1126.965 ;
        RECT 1992.675 1124.890 1992.935 1125.210 ;
        RECT 1992.675 1116.100 1992.815 1124.890 ;
        RECT 1992.180 1115.780 1993.270 1116.100 ;
    END
  END mgmt_io_out_unbuf[30]
  PIN mgmt_io_out_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1997.660 1115.850 1999.250 1116.050 ;
      LAYER mcon ;
        RECT 1998.160 1115.850 1999.250 1116.020 ;
      LAYER met1 ;
        RECT 1998.625 1124.480 3375.600 1124.620 ;
        RECT 1998.625 1124.360 1998.945 1124.480 ;
        RECT 1998.100 1115.810 1999.310 1116.070 ;
        RECT 3375.460 1083.250 3375.600 1124.480 ;
      LAYER via ;
        RECT 1998.655 1124.360 1998.915 1124.620 ;
        RECT 1998.160 1115.810 1999.250 1116.070 ;
      LAYER met2 ;
        RECT 1998.655 1124.650 1998.795 1126.965 ;
        RECT 1998.655 1124.330 1998.915 1124.650 ;
        RECT 1998.655 1116.100 1998.795 1124.330 ;
        RECT 1998.160 1115.780 1999.250 1116.100 ;
    END
  END mgmt_io_out_unbuf[29]
  PIN mgmt_io_out_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2003.640 1115.850 2005.230 1116.050 ;
      LAYER mcon ;
        RECT 2004.140 1115.850 2005.230 1116.020 ;
      LAYER met1 ;
        RECT 2004.485 1123.920 3375.040 1124.060 ;
        RECT 2004.485 1123.800 2004.805 1123.920 ;
        RECT 2004.080 1115.810 2005.290 1116.070 ;
        RECT 3374.900 1085.250 3375.040 1123.920 ;
      LAYER via ;
        RECT 2004.515 1123.800 2004.775 1124.060 ;
        RECT 2004.140 1115.810 2005.230 1116.070 ;
      LAYER met2 ;
        RECT 2004.635 1124.090 2004.775 1126.965 ;
        RECT 2004.515 1123.770 2004.775 1124.090 ;
        RECT 2004.635 1116.100 2004.775 1123.770 ;
        RECT 2004.140 1115.780 2005.230 1116.100 ;
    END
  END mgmt_io_out_unbuf[28]
  PIN mgmt_io_out_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2009.620 1115.850 2011.210 1116.050 ;
      LAYER mcon ;
        RECT 2010.120 1115.850 2011.210 1116.020 ;
      LAYER met1 ;
        RECT 2010.585 1123.360 3374.480 1123.500 ;
        RECT 2010.585 1123.240 2010.905 1123.360 ;
        RECT 2010.060 1115.810 2011.270 1116.070 ;
        RECT 3374.340 1087.250 3374.480 1123.360 ;
      LAYER via ;
        RECT 2010.615 1123.240 2010.875 1123.500 ;
        RECT 2010.120 1115.810 2011.210 1116.070 ;
      LAYER met2 ;
        RECT 2010.615 1123.530 2010.755 1126.965 ;
        RECT 2010.615 1123.210 2010.875 1123.530 ;
        RECT 2010.615 1116.100 2010.755 1123.210 ;
        RECT 2010.120 1115.780 2011.210 1116.100 ;
    END
  END mgmt_io_out_unbuf[27]
  PIN mgmt_io_out_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2015.600 1115.850 2017.190 1116.050 ;
      LAYER mcon ;
        RECT 2016.100 1115.850 2017.190 1116.020 ;
      LAYER met1 ;
        RECT 2016.445 1122.800 3373.920 1122.940 ;
        RECT 2016.445 1122.680 2016.765 1122.800 ;
        RECT 2016.040 1115.810 2017.250 1116.070 ;
        RECT 3373.780 1089.250 3373.920 1122.800 ;
      LAYER via ;
        RECT 2016.475 1122.680 2016.735 1122.940 ;
        RECT 2016.100 1115.810 2017.190 1116.070 ;
      LAYER met2 ;
        RECT 2016.595 1122.970 2016.735 1126.965 ;
        RECT 2016.475 1122.650 2016.735 1122.970 ;
        RECT 2016.595 1116.100 2016.735 1122.650 ;
        RECT 2016.100 1115.780 2017.190 1116.100 ;
    END
  END mgmt_io_out_unbuf[26]
  PIN mgmt_io_out_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2021.580 1115.850 2023.170 1116.050 ;
      LAYER mcon ;
        RECT 2022.080 1115.850 2023.170 1116.020 ;
      LAYER met1 ;
        RECT 2022.545 1122.240 3373.360 1122.380 ;
        RECT 2022.545 1122.120 2022.865 1122.240 ;
        RECT 2022.020 1115.810 2023.230 1116.070 ;
        RECT 3373.220 1091.250 3373.360 1122.240 ;
      LAYER via ;
        RECT 2022.575 1122.120 2022.835 1122.380 ;
        RECT 2022.080 1115.810 2023.170 1116.070 ;
      LAYER met2 ;
        RECT 2022.575 1122.410 2022.715 1126.965 ;
        RECT 2022.575 1122.090 2022.835 1122.410 ;
        RECT 2022.575 1116.100 2022.715 1122.090 ;
        RECT 2022.080 1115.780 2023.170 1116.100 ;
    END
  END mgmt_io_out_unbuf[25]
  PIN mgmt_io_out_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2027.560 1115.850 2029.150 1116.050 ;
      LAYER mcon ;
        RECT 2028.060 1115.850 2029.150 1116.020 ;
      LAYER met1 ;
        RECT 2028.525 1121.680 3372.800 1121.820 ;
        RECT 2028.525 1121.560 2028.845 1121.680 ;
        RECT 2028.000 1115.810 2029.210 1116.070 ;
        RECT 3372.660 1093.250 3372.800 1121.680 ;
      LAYER via ;
        RECT 2028.555 1121.560 2028.815 1121.820 ;
        RECT 2028.060 1115.810 2029.150 1116.070 ;
      LAYER met2 ;
        RECT 2028.555 1121.850 2028.695 1126.965 ;
        RECT 2028.555 1121.530 2028.815 1121.850 ;
        RECT 2028.555 1116.100 2028.695 1121.530 ;
        RECT 2028.060 1115.780 2029.150 1116.100 ;
    END
  END mgmt_io_out_unbuf[24]
  PIN mgmt_io_in_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2031.115 1113.300 2031.285 1114.150 ;
        RECT 2031.955 1113.300 2032.125 1114.150 ;
        RECT 2032.795 1113.300 2032.965 1114.150 ;
        RECT 2033.635 1113.300 2033.805 1114.150 ;
        RECT 2031.115 1113.130 2033.805 1113.300 ;
        RECT 2033.550 1112.590 2033.805 1113.130 ;
        RECT 2031.115 1112.420 2033.805 1112.590 ;
        RECT 2031.115 1111.940 2031.285 1112.420 ;
        RECT 2031.955 1111.940 2032.125 1112.420 ;
        RECT 2032.795 1111.940 2032.965 1112.420 ;
        RECT 2033.635 1111.940 2033.805 1112.420 ;
      LAYER mcon ;
        RECT 2033.550 1112.450 2033.720 1113.300 ;
      LAYER met1 ;
        RECT 2033.535 1121.400 3372.520 1121.540 ;
        RECT 2033.535 1121.280 2033.855 1121.400 ;
        RECT 2033.500 1112.390 2033.760 1113.360 ;
        RECT 3372.380 1094.250 3372.520 1121.400 ;
      LAYER via ;
        RECT 2033.565 1121.280 2033.825 1121.540 ;
        RECT 2033.500 1112.450 2033.760 1113.300 ;
      LAYER met2 ;
        RECT 2033.565 1121.570 2033.705 1126.965 ;
        RECT 2033.565 1121.250 2033.825 1121.570 ;
        RECT 2033.565 1113.300 2033.705 1121.250 ;
        RECT 2033.470 1112.450 2033.790 1113.300 ;
    END
  END mgmt_io_in_buf[24]
  PIN mgmt_io_in_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2025.135 1113.300 2025.305 1114.150 ;
        RECT 2025.975 1113.300 2026.145 1114.150 ;
        RECT 2026.815 1113.300 2026.985 1114.150 ;
        RECT 2027.655 1113.300 2027.825 1114.150 ;
        RECT 2025.135 1113.130 2027.825 1113.300 ;
        RECT 2027.570 1112.590 2027.825 1113.130 ;
        RECT 2025.135 1112.420 2027.825 1112.590 ;
        RECT 2025.135 1111.940 2025.305 1112.420 ;
        RECT 2025.975 1111.940 2026.145 1112.420 ;
        RECT 2026.815 1111.940 2026.985 1112.420 ;
        RECT 2027.655 1111.940 2027.825 1112.420 ;
      LAYER mcon ;
        RECT 2027.570 1112.450 2027.740 1113.300 ;
      LAYER met1 ;
        RECT 2027.555 1121.960 3373.080 1122.100 ;
        RECT 2027.555 1121.840 2027.875 1121.960 ;
        RECT 2027.520 1112.390 2027.780 1113.360 ;
        RECT 3372.940 1092.250 3373.080 1121.960 ;
      LAYER via ;
        RECT 2027.585 1121.840 2027.845 1122.100 ;
        RECT 2027.520 1112.450 2027.780 1113.300 ;
      LAYER met2 ;
        RECT 2027.585 1122.130 2027.725 1126.965 ;
        RECT 2027.585 1121.810 2027.845 1122.130 ;
        RECT 2027.585 1113.300 2027.725 1121.810 ;
        RECT 2027.490 1112.450 2027.810 1113.300 ;
    END
  END mgmt_io_in_buf[25]
  PIN mgmt_io_in_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2019.155 1113.300 2019.325 1114.150 ;
        RECT 2019.995 1113.300 2020.165 1114.150 ;
        RECT 2020.835 1113.300 2021.005 1114.150 ;
        RECT 2021.675 1113.300 2021.845 1114.150 ;
        RECT 2019.155 1113.130 2021.845 1113.300 ;
        RECT 2021.590 1112.590 2021.845 1113.130 ;
        RECT 2019.155 1112.420 2021.845 1112.590 ;
        RECT 2019.155 1111.940 2019.325 1112.420 ;
        RECT 2019.995 1111.940 2020.165 1112.420 ;
        RECT 2020.835 1111.940 2021.005 1112.420 ;
        RECT 2021.675 1111.940 2021.845 1112.420 ;
      LAYER mcon ;
        RECT 2021.590 1112.450 2021.760 1113.300 ;
      LAYER met1 ;
        RECT 2021.575 1122.520 3373.640 1122.660 ;
        RECT 2021.575 1122.400 2021.895 1122.520 ;
        RECT 2021.540 1112.390 2021.800 1113.360 ;
        RECT 3373.500 1090.250 3373.640 1122.520 ;
      LAYER via ;
        RECT 2021.605 1122.400 2021.865 1122.660 ;
        RECT 2021.540 1112.450 2021.800 1113.300 ;
      LAYER met2 ;
        RECT 2021.605 1122.690 2021.745 1126.965 ;
        RECT 2021.605 1122.370 2021.865 1122.690 ;
        RECT 2021.605 1113.300 2021.745 1122.370 ;
        RECT 2021.510 1112.450 2021.830 1113.300 ;
    END
  END mgmt_io_in_buf[26]
  PIN mgmt_io_in_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2013.175 1113.300 2013.345 1114.150 ;
        RECT 2014.015 1113.300 2014.185 1114.150 ;
        RECT 2014.855 1113.300 2015.025 1114.150 ;
        RECT 2015.695 1113.300 2015.865 1114.150 ;
        RECT 2013.175 1113.130 2015.865 1113.300 ;
        RECT 2015.610 1112.590 2015.865 1113.130 ;
        RECT 2013.175 1112.420 2015.865 1112.590 ;
        RECT 2013.175 1111.940 2013.345 1112.420 ;
        RECT 2014.015 1111.940 2014.185 1112.420 ;
        RECT 2014.855 1111.940 2015.025 1112.420 ;
        RECT 2015.695 1111.940 2015.865 1112.420 ;
      LAYER mcon ;
        RECT 2015.610 1112.450 2015.780 1113.300 ;
      LAYER met1 ;
        RECT 2015.595 1123.080 3374.200 1123.220 ;
        RECT 2015.595 1122.960 2015.915 1123.080 ;
        RECT 2015.560 1112.390 2015.820 1113.360 ;
        RECT 3374.060 1088.250 3374.200 1123.080 ;
      LAYER via ;
        RECT 2015.625 1122.960 2015.885 1123.220 ;
        RECT 2015.560 1112.450 2015.820 1113.300 ;
      LAYER met2 ;
        RECT 2015.625 1123.250 2015.765 1126.965 ;
        RECT 2015.625 1122.930 2015.885 1123.250 ;
        RECT 2015.625 1113.300 2015.765 1122.930 ;
        RECT 2015.530 1112.450 2015.850 1113.300 ;
    END
  END mgmt_io_in_buf[27]
  PIN mgmt_io_in_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2007.195 1113.300 2007.365 1114.150 ;
        RECT 2008.035 1113.300 2008.205 1114.150 ;
        RECT 2008.875 1113.300 2009.045 1114.150 ;
        RECT 2009.715 1113.300 2009.885 1114.150 ;
        RECT 2007.195 1113.130 2009.885 1113.300 ;
        RECT 2009.630 1112.590 2009.885 1113.130 ;
        RECT 2007.195 1112.420 2009.885 1112.590 ;
        RECT 2007.195 1111.940 2007.365 1112.420 ;
        RECT 2008.035 1111.940 2008.205 1112.420 ;
        RECT 2008.875 1111.940 2009.045 1112.420 ;
        RECT 2009.715 1111.940 2009.885 1112.420 ;
      LAYER mcon ;
        RECT 2009.630 1112.450 2009.800 1113.300 ;
      LAYER met1 ;
        RECT 2009.615 1123.640 3374.760 1123.780 ;
        RECT 2009.615 1123.520 2009.935 1123.640 ;
        RECT 2009.580 1112.390 2009.840 1113.360 ;
        RECT 3374.620 1086.250 3374.760 1123.640 ;
      LAYER via ;
        RECT 2009.645 1123.520 2009.905 1123.780 ;
        RECT 2009.580 1112.450 2009.840 1113.300 ;
      LAYER met2 ;
        RECT 2009.645 1123.810 2009.785 1126.965 ;
        RECT 2009.645 1123.490 2009.905 1123.810 ;
        RECT 2009.645 1113.300 2009.785 1123.490 ;
        RECT 2009.550 1112.450 2009.870 1113.300 ;
    END
  END mgmt_io_in_buf[28]
  PIN mgmt_io_in_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2001.215 1113.300 2001.385 1114.150 ;
        RECT 2002.055 1113.300 2002.225 1114.150 ;
        RECT 2002.895 1113.300 2003.065 1114.150 ;
        RECT 2003.735 1113.300 2003.905 1114.150 ;
        RECT 2001.215 1113.130 2003.905 1113.300 ;
        RECT 2003.650 1112.590 2003.905 1113.130 ;
        RECT 2001.215 1112.420 2003.905 1112.590 ;
        RECT 2001.215 1111.940 2001.385 1112.420 ;
        RECT 2002.055 1111.940 2002.225 1112.420 ;
        RECT 2002.895 1111.940 2003.065 1112.420 ;
        RECT 2003.735 1111.940 2003.905 1112.420 ;
      LAYER mcon ;
        RECT 2003.650 1112.450 2003.820 1113.300 ;
      LAYER met1 ;
        RECT 2003.635 1124.200 3375.320 1124.340 ;
        RECT 2003.635 1124.080 2003.955 1124.200 ;
        RECT 2003.600 1112.390 2003.860 1113.360 ;
        RECT 3375.180 1084.250 3375.320 1124.200 ;
      LAYER via ;
        RECT 2003.665 1124.080 2003.925 1124.340 ;
        RECT 2003.600 1112.450 2003.860 1113.300 ;
      LAYER met2 ;
        RECT 2003.665 1124.370 2003.805 1126.965 ;
        RECT 2003.665 1124.050 2003.925 1124.370 ;
        RECT 2003.665 1113.300 2003.805 1124.050 ;
        RECT 2003.570 1112.450 2003.890 1113.300 ;
    END
  END mgmt_io_in_buf[29]
  PIN mgmt_io_in_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1995.235 1113.300 1995.405 1114.150 ;
        RECT 1996.075 1113.300 1996.245 1114.150 ;
        RECT 1996.915 1113.300 1997.085 1114.150 ;
        RECT 1997.755 1113.300 1997.925 1114.150 ;
        RECT 1995.235 1113.130 1997.925 1113.300 ;
        RECT 1997.670 1112.590 1997.925 1113.130 ;
        RECT 1995.235 1112.420 1997.925 1112.590 ;
        RECT 1995.235 1111.940 1995.405 1112.420 ;
        RECT 1996.075 1111.940 1996.245 1112.420 ;
        RECT 1996.915 1111.940 1997.085 1112.420 ;
        RECT 1997.755 1111.940 1997.925 1112.420 ;
      LAYER mcon ;
        RECT 1997.670 1112.450 1997.840 1113.300 ;
      LAYER met1 ;
        RECT 1997.655 1124.760 3375.880 1124.900 ;
        RECT 1997.655 1124.640 1997.975 1124.760 ;
        RECT 1997.620 1112.390 1997.880 1113.360 ;
        RECT 3375.740 1082.250 3375.880 1124.760 ;
      LAYER via ;
        RECT 1997.685 1124.640 1997.945 1124.900 ;
        RECT 1997.620 1112.450 1997.880 1113.300 ;
      LAYER met2 ;
        RECT 1997.685 1124.930 1997.825 1126.965 ;
        RECT 1997.685 1124.610 1997.945 1124.930 ;
        RECT 1997.685 1113.300 1997.825 1124.610 ;
        RECT 1997.590 1112.450 1997.910 1113.300 ;
    END
  END mgmt_io_in_buf[30]
  PIN mgmt_io_in_buf[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1989.255 1113.300 1989.425 1114.150 ;
        RECT 1990.095 1113.300 1990.265 1114.150 ;
        RECT 1990.935 1113.300 1991.105 1114.150 ;
        RECT 1991.775 1113.300 1991.945 1114.150 ;
        RECT 1989.255 1113.130 1991.945 1113.300 ;
        RECT 1991.690 1112.590 1991.945 1113.130 ;
        RECT 1989.255 1112.420 1991.945 1112.590 ;
        RECT 1989.255 1111.940 1989.425 1112.420 ;
        RECT 1990.095 1111.940 1990.265 1112.420 ;
        RECT 1990.935 1111.940 1991.105 1112.420 ;
        RECT 1991.775 1111.940 1991.945 1112.420 ;
      LAYER mcon ;
        RECT 1991.690 1112.450 1991.860 1113.300 ;
      LAYER met1 ;
        RECT 1991.675 1125.320 3376.440 1125.460 ;
        RECT 1991.675 1125.200 1991.995 1125.320 ;
        RECT 1991.640 1112.390 1991.900 1113.360 ;
        RECT 3376.300 1080.250 3376.440 1125.320 ;
      LAYER via ;
        RECT 1991.705 1125.200 1991.965 1125.460 ;
        RECT 1991.640 1112.450 1991.900 1113.300 ;
      LAYER met2 ;
        RECT 1991.705 1125.490 1991.845 1126.965 ;
        RECT 1991.705 1125.170 1991.965 1125.490 ;
        RECT 1991.705 1113.300 1991.845 1125.170 ;
        RECT 1991.610 1112.450 1991.930 1113.300 ;
    END
  END mgmt_io_in_buf[31]
  PIN mgmt_io_in_buf[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1983.275 1113.300 1983.445 1114.150 ;
        RECT 1984.115 1113.300 1984.285 1114.150 ;
        RECT 1984.955 1113.300 1985.125 1114.150 ;
        RECT 1985.795 1113.300 1985.965 1114.150 ;
        RECT 1983.275 1113.130 1985.965 1113.300 ;
        RECT 1985.710 1112.590 1985.965 1113.130 ;
        RECT 1983.275 1112.420 1985.965 1112.590 ;
        RECT 1983.275 1111.940 1983.445 1112.420 ;
        RECT 1984.115 1111.940 1984.285 1112.420 ;
        RECT 1984.955 1111.940 1985.125 1112.420 ;
        RECT 1985.795 1111.940 1985.965 1112.420 ;
      LAYER mcon ;
        RECT 1985.710 1112.450 1985.880 1113.300 ;
      LAYER met1 ;
        RECT 1985.695 1125.880 3377.000 1126.020 ;
        RECT 1985.695 1125.760 1986.015 1125.880 ;
        RECT 1985.660 1112.390 1985.920 1113.360 ;
        RECT 3376.860 1078.250 3377.000 1125.880 ;
      LAYER via ;
        RECT 1985.725 1125.760 1985.985 1126.020 ;
        RECT 1985.660 1112.450 1985.920 1113.300 ;
      LAYER met2 ;
        RECT 1985.725 1126.050 1985.865 1126.965 ;
        RECT 1985.725 1125.730 1985.985 1126.050 ;
        RECT 1985.725 1113.300 1985.865 1125.730 ;
        RECT 1985.630 1112.450 1985.950 1113.300 ;
    END
  END mgmt_io_in_buf[32]
  PIN mgmt_io_in_buf[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1977.295 1113.300 1977.465 1114.150 ;
        RECT 1978.135 1113.300 1978.305 1114.150 ;
        RECT 1978.975 1113.300 1979.145 1114.150 ;
        RECT 1979.815 1113.300 1979.985 1114.150 ;
        RECT 1977.295 1113.130 1979.985 1113.300 ;
        RECT 1979.730 1112.590 1979.985 1113.130 ;
        RECT 1977.295 1112.420 1979.985 1112.590 ;
        RECT 1977.295 1111.940 1977.465 1112.420 ;
        RECT 1978.135 1111.940 1978.305 1112.420 ;
        RECT 1978.975 1111.940 1979.145 1112.420 ;
        RECT 1979.815 1111.940 1979.985 1112.420 ;
      LAYER mcon ;
        RECT 1979.730 1112.450 1979.900 1113.300 ;
      LAYER met1 ;
        RECT 1979.715 1126.440 3377.560 1126.580 ;
        RECT 1979.715 1126.320 1980.035 1126.440 ;
        RECT 1979.680 1112.390 1979.940 1113.360 ;
        RECT 3377.420 1076.250 3377.560 1126.440 ;
      LAYER via ;
        RECT 1979.745 1126.320 1980.005 1126.580 ;
        RECT 1979.680 1112.450 1979.940 1113.300 ;
      LAYER met2 ;
        RECT 1979.745 1126.610 1979.885 1126.965 ;
        RECT 1979.745 1126.290 1980.005 1126.610 ;
        RECT 1979.745 1113.300 1979.885 1126.290 ;
        RECT 1979.650 1112.450 1979.970 1113.300 ;
    END
  END mgmt_io_in_buf[33]
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 669.145 1117.040 669.315 1117.210 ;
        RECT 669.605 1117.040 669.775 1117.210 ;
        RECT 670.065 1117.040 670.235 1117.210 ;
        RECT 670.525 1117.040 670.695 1117.210 ;
        RECT 670.985 1117.040 671.155 1117.210 ;
        RECT 671.445 1117.040 671.615 1117.210 ;
        RECT 671.905 1117.040 672.075 1117.210 ;
        RECT 672.365 1117.040 672.535 1117.210 ;
        RECT 672.825 1117.040 672.995 1117.210 ;
        RECT 673.285 1117.040 673.455 1117.210 ;
        RECT 673.745 1117.040 673.915 1117.210 ;
        RECT 674.205 1117.040 674.375 1117.210 ;
        RECT 674.665 1117.040 674.835 1117.210 ;
        RECT 675.125 1117.040 675.295 1117.210 ;
        RECT 675.585 1117.040 675.755 1117.210 ;
        RECT 676.045 1117.040 676.215 1117.210 ;
        RECT 676.505 1117.040 676.675 1117.210 ;
        RECT 676.965 1117.040 677.135 1117.210 ;
        RECT 677.425 1117.040 677.595 1117.210 ;
        RECT 677.885 1117.040 678.055 1117.210 ;
        RECT 678.345 1117.040 678.515 1117.210 ;
        RECT 678.805 1117.040 678.975 1117.210 ;
        RECT 679.265 1117.040 679.435 1117.210 ;
        RECT 679.725 1117.040 679.895 1117.210 ;
        RECT 680.185 1117.040 680.355 1117.210 ;
        RECT 680.645 1117.040 680.815 1117.210 ;
        RECT 681.105 1117.040 681.275 1117.210 ;
        RECT 681.565 1117.040 681.735 1117.210 ;
        RECT 682.025 1117.040 682.195 1117.210 ;
        RECT 682.485 1117.040 682.655 1117.210 ;
        RECT 682.945 1117.040 683.115 1117.210 ;
        RECT 683.405 1117.040 683.575 1117.210 ;
        RECT 683.865 1117.040 684.035 1117.210 ;
        RECT 684.325 1117.040 684.495 1117.210 ;
        RECT 684.785 1117.040 684.955 1117.210 ;
        RECT 685.245 1117.040 685.415 1117.210 ;
        RECT 685.705 1117.040 685.875 1117.210 ;
        RECT 686.165 1117.040 686.335 1117.210 ;
        RECT 686.625 1117.040 686.795 1117.210 ;
        RECT 687.085 1117.040 687.255 1117.210 ;
        RECT 687.545 1117.040 687.715 1117.210 ;
        RECT 688.005 1117.040 688.175 1117.210 ;
        RECT 688.465 1117.040 688.635 1117.210 ;
        RECT 688.925 1117.040 689.095 1117.210 ;
        RECT 689.385 1117.040 689.555 1117.210 ;
        RECT 689.845 1117.040 690.015 1117.210 ;
        RECT 690.305 1117.040 690.475 1117.210 ;
        RECT 690.765 1117.040 690.935 1117.210 ;
        RECT 691.225 1117.040 691.395 1117.210 ;
        RECT 691.685 1117.040 691.855 1117.210 ;
        RECT 692.145 1117.040 692.315 1117.210 ;
        RECT 692.605 1117.040 692.775 1117.210 ;
        RECT 693.065 1117.040 693.235 1117.210 ;
        RECT 693.525 1117.040 693.695 1117.210 ;
        RECT 693.985 1117.040 694.155 1117.210 ;
        RECT 694.445 1117.040 694.615 1117.210 ;
        RECT 694.905 1117.040 695.075 1117.210 ;
        RECT 695.365 1117.040 695.535 1117.210 ;
        RECT 695.825 1117.040 695.995 1117.210 ;
        RECT 696.285 1117.040 696.455 1117.210 ;
        RECT 696.745 1117.040 696.915 1117.210 ;
        RECT 697.205 1117.040 697.375 1117.210 ;
        RECT 697.665 1117.040 697.835 1117.210 ;
        RECT 698.125 1117.040 698.295 1117.210 ;
        RECT 698.585 1117.040 698.755 1117.210 ;
        RECT 699.045 1117.040 699.215 1117.210 ;
        RECT 699.505 1117.040 699.675 1117.210 ;
        RECT 699.965 1117.040 700.135 1117.210 ;
        RECT 700.425 1117.040 700.595 1117.210 ;
        RECT 700.885 1117.040 701.055 1117.210 ;
        RECT 701.345 1117.040 701.515 1117.210 ;
        RECT 701.805 1117.040 701.975 1117.210 ;
        RECT 702.265 1117.040 702.435 1117.210 ;
        RECT 702.725 1117.040 702.895 1117.210 ;
        RECT 703.185 1117.040 703.355 1117.210 ;
        RECT 703.645 1117.040 703.815 1117.210 ;
        RECT 704.105 1117.040 704.275 1117.210 ;
        RECT 704.565 1117.040 704.735 1117.210 ;
        RECT 705.025 1117.040 705.195 1117.210 ;
        RECT 705.485 1117.040 705.655 1117.210 ;
        RECT 705.945 1117.040 706.115 1117.210 ;
        RECT 706.405 1117.040 706.575 1117.210 ;
        RECT 706.865 1117.040 707.035 1117.210 ;
        RECT 707.325 1117.040 707.495 1117.210 ;
        RECT 707.785 1117.040 707.955 1117.210 ;
        RECT 708.245 1117.040 708.415 1117.210 ;
        RECT 708.705 1117.040 708.875 1117.210 ;
        RECT 709.165 1117.040 709.335 1117.210 ;
        RECT 709.625 1117.040 709.795 1117.210 ;
        RECT 710.085 1117.040 710.255 1117.210 ;
        RECT 710.545 1117.040 710.715 1117.210 ;
        RECT 711.005 1117.040 711.175 1117.210 ;
        RECT 711.465 1117.040 711.635 1117.210 ;
        RECT 711.925 1117.040 712.095 1117.210 ;
        RECT 712.385 1117.040 712.555 1117.210 ;
        RECT 712.845 1117.040 713.015 1117.210 ;
        RECT 713.305 1117.040 713.475 1117.210 ;
        RECT 713.765 1117.040 713.935 1117.210 ;
        RECT 714.225 1117.040 714.395 1117.210 ;
        RECT 714.685 1117.040 714.855 1117.210 ;
        RECT 715.145 1117.040 715.315 1117.210 ;
        RECT 715.605 1117.040 715.775 1117.210 ;
        RECT 716.065 1117.040 716.235 1117.210 ;
        RECT 716.525 1117.040 716.695 1117.210 ;
        RECT 716.985 1117.040 717.155 1117.210 ;
        RECT 717.445 1117.040 717.615 1117.210 ;
        RECT 717.905 1117.040 718.075 1117.210 ;
        RECT 718.365 1117.040 718.535 1117.210 ;
        RECT 718.825 1117.040 718.995 1117.210 ;
        RECT 719.285 1117.040 719.455 1117.210 ;
        RECT 719.745 1117.040 719.915 1117.210 ;
        RECT 720.205 1117.040 720.375 1117.210 ;
        RECT 720.665 1117.040 720.835 1117.210 ;
        RECT 721.125 1117.040 721.295 1117.210 ;
        RECT 721.585 1117.040 721.755 1117.210 ;
        RECT 722.045 1117.040 722.215 1117.210 ;
        RECT 722.505 1117.040 722.675 1117.210 ;
        RECT 722.965 1117.040 723.135 1117.210 ;
        RECT 723.425 1117.040 723.595 1117.210 ;
        RECT 723.885 1117.040 724.055 1117.210 ;
        RECT 724.345 1117.040 724.515 1117.210 ;
        RECT 724.805 1117.040 724.975 1117.210 ;
        RECT 725.265 1117.040 725.435 1117.210 ;
        RECT 725.725 1117.040 725.895 1117.210 ;
        RECT 726.185 1117.040 726.355 1117.210 ;
        RECT 726.645 1117.040 726.815 1117.210 ;
        RECT 727.105 1117.040 727.275 1117.210 ;
        RECT 727.565 1117.040 727.735 1117.210 ;
        RECT 728.025 1117.040 728.195 1117.210 ;
        RECT 728.485 1117.040 728.655 1117.210 ;
        RECT 728.945 1117.040 729.115 1117.210 ;
        RECT 729.405 1117.040 729.575 1117.210 ;
        RECT 729.865 1117.040 730.035 1117.210 ;
        RECT 730.325 1117.040 730.495 1117.210 ;
        RECT 730.785 1117.040 730.955 1117.210 ;
        RECT 731.245 1117.040 731.415 1117.210 ;
        RECT 731.705 1117.040 731.875 1117.210 ;
        RECT 732.165 1117.040 732.335 1117.210 ;
        RECT 732.625 1117.040 732.795 1117.210 ;
        RECT 733.085 1117.040 733.255 1117.210 ;
        RECT 733.545 1117.040 733.715 1117.210 ;
        RECT 734.005 1117.040 734.175 1117.210 ;
        RECT 734.465 1117.040 734.635 1117.210 ;
        RECT 734.925 1117.040 735.095 1117.210 ;
        RECT 735.385 1117.040 735.555 1117.210 ;
        RECT 735.845 1117.040 736.015 1117.210 ;
        RECT 736.305 1117.040 736.475 1117.210 ;
        RECT 736.765 1117.040 736.935 1117.210 ;
        RECT 737.225 1117.040 737.395 1117.210 ;
        RECT 737.685 1117.040 737.855 1117.210 ;
        RECT 738.145 1117.040 738.315 1117.210 ;
        RECT 738.605 1117.040 738.775 1117.210 ;
        RECT 739.065 1117.040 739.235 1117.210 ;
        RECT 739.525 1117.040 739.695 1117.210 ;
        RECT 739.985 1117.040 740.155 1117.210 ;
        RECT 740.445 1117.040 740.615 1117.210 ;
        RECT 740.905 1117.040 741.075 1117.210 ;
        RECT 741.365 1117.040 741.535 1117.210 ;
        RECT 741.825 1117.040 741.995 1117.210 ;
        RECT 742.285 1117.040 742.455 1117.210 ;
        RECT 742.745 1117.040 742.915 1117.210 ;
        RECT 743.205 1117.040 743.375 1117.210 ;
        RECT 743.665 1117.040 743.835 1117.210 ;
        RECT 744.125 1117.040 744.295 1117.210 ;
        RECT 744.585 1117.040 744.755 1117.210 ;
        RECT 745.045 1117.040 745.215 1117.210 ;
        RECT 745.505 1117.040 745.675 1117.210 ;
        RECT 745.965 1117.040 746.135 1117.210 ;
        RECT 746.425 1117.040 746.595 1117.210 ;
        RECT 746.885 1117.040 747.055 1117.210 ;
        RECT 747.345 1117.040 747.515 1117.210 ;
        RECT 747.805 1117.040 747.975 1117.210 ;
        RECT 748.265 1117.040 748.435 1117.210 ;
        RECT 748.725 1117.040 748.895 1117.210 ;
        RECT 749.185 1117.040 749.355 1117.210 ;
        RECT 749.645 1117.040 749.815 1117.210 ;
        RECT 750.105 1117.040 750.275 1117.210 ;
        RECT 750.565 1117.040 750.735 1117.210 ;
        RECT 751.025 1117.040 751.195 1117.210 ;
        RECT 751.485 1117.040 751.655 1117.210 ;
        RECT 751.945 1117.040 752.115 1117.210 ;
        RECT 752.405 1117.040 752.575 1117.210 ;
        RECT 752.865 1117.040 753.035 1117.210 ;
        RECT 753.325 1117.040 753.495 1117.210 ;
        RECT 753.785 1117.040 753.955 1117.210 ;
        RECT 754.245 1117.040 754.415 1117.210 ;
        RECT 754.705 1117.040 754.875 1117.210 ;
        RECT 755.165 1117.040 755.335 1117.210 ;
        RECT 755.625 1117.040 755.795 1117.210 ;
        RECT 756.085 1117.040 756.255 1117.210 ;
        RECT 756.545 1117.040 756.715 1117.210 ;
        RECT 757.005 1117.040 757.175 1117.210 ;
        RECT 757.465 1117.040 757.635 1117.210 ;
        RECT 757.925 1117.040 758.095 1117.210 ;
        RECT 758.385 1117.040 758.555 1117.210 ;
        RECT 758.845 1117.040 759.015 1117.210 ;
        RECT 759.305 1117.040 759.475 1117.210 ;
        RECT 759.765 1117.040 759.935 1117.210 ;
        RECT 760.225 1117.040 760.395 1117.210 ;
        RECT 760.685 1117.040 760.855 1117.210 ;
        RECT 761.145 1117.040 761.315 1117.210 ;
        RECT 761.605 1117.040 761.775 1117.210 ;
        RECT 762.065 1117.040 762.235 1117.210 ;
        RECT 762.525 1117.040 762.695 1117.210 ;
        RECT 762.985 1117.040 763.155 1117.210 ;
        RECT 763.445 1117.040 763.615 1117.210 ;
        RECT 763.905 1117.040 764.075 1117.210 ;
        RECT 764.365 1117.040 764.535 1117.210 ;
        RECT 764.825 1117.040 764.995 1117.210 ;
        RECT 765.285 1117.040 765.455 1117.210 ;
        RECT 765.745 1117.040 765.915 1117.210 ;
        RECT 766.205 1117.040 766.375 1117.210 ;
        RECT 766.665 1117.040 766.835 1117.210 ;
        RECT 767.125 1117.040 767.295 1117.210 ;
        RECT 767.585 1117.040 767.755 1117.210 ;
        RECT 768.045 1117.040 768.215 1117.210 ;
        RECT 768.505 1117.040 768.675 1117.210 ;
        RECT 768.965 1117.040 769.135 1117.210 ;
        RECT 769.425 1117.040 769.595 1117.210 ;
        RECT 769.885 1117.040 770.055 1117.210 ;
        RECT 770.345 1117.040 770.515 1117.210 ;
        RECT 770.805 1117.040 770.975 1117.210 ;
        RECT 675.125 1111.600 675.295 1111.770 ;
        RECT 675.585 1111.600 675.755 1111.770 ;
        RECT 676.045 1111.600 676.215 1111.770 ;
        RECT 676.505 1111.600 676.675 1111.770 ;
        RECT 676.965 1111.600 677.135 1111.770 ;
        RECT 677.425 1111.600 677.595 1111.770 ;
        RECT 677.885 1111.600 678.055 1111.770 ;
        RECT 678.345 1111.600 678.515 1111.770 ;
        RECT 678.805 1111.600 678.975 1111.770 ;
        RECT 679.265 1111.600 679.435 1111.770 ;
        RECT 679.725 1111.600 679.895 1111.770 ;
        RECT 680.185 1111.600 680.355 1111.770 ;
        RECT 680.645 1111.600 680.815 1111.770 ;
        RECT 681.105 1111.600 681.275 1111.770 ;
        RECT 681.565 1111.600 681.735 1111.770 ;
        RECT 682.025 1111.600 682.195 1111.770 ;
        RECT 682.485 1111.600 682.655 1111.770 ;
        RECT 682.945 1111.600 683.115 1111.770 ;
        RECT 683.405 1111.600 683.575 1111.770 ;
        RECT 683.865 1111.600 684.035 1111.770 ;
        RECT 684.325 1111.600 684.495 1111.770 ;
        RECT 684.785 1111.600 684.955 1111.770 ;
        RECT 685.245 1111.600 685.415 1111.770 ;
        RECT 685.705 1111.600 685.875 1111.770 ;
        RECT 686.165 1111.600 686.335 1111.770 ;
        RECT 686.625 1111.600 686.795 1111.770 ;
        RECT 687.085 1111.600 687.255 1111.770 ;
        RECT 687.545 1111.600 687.715 1111.770 ;
        RECT 688.005 1111.600 688.175 1111.770 ;
        RECT 688.465 1111.600 688.635 1111.770 ;
        RECT 688.925 1111.600 689.095 1111.770 ;
        RECT 689.385 1111.600 689.555 1111.770 ;
        RECT 689.845 1111.600 690.015 1111.770 ;
        RECT 690.305 1111.600 690.475 1111.770 ;
        RECT 690.765 1111.600 690.935 1111.770 ;
        RECT 691.225 1111.600 691.395 1111.770 ;
        RECT 691.685 1111.600 691.855 1111.770 ;
        RECT 692.145 1111.600 692.315 1111.770 ;
        RECT 692.605 1111.600 692.775 1111.770 ;
        RECT 693.065 1111.600 693.235 1111.770 ;
        RECT 693.525 1111.600 693.695 1111.770 ;
        RECT 693.985 1111.600 694.155 1111.770 ;
        RECT 694.445 1111.600 694.615 1111.770 ;
        RECT 694.905 1111.600 695.075 1111.770 ;
        RECT 695.365 1111.600 695.535 1111.770 ;
        RECT 695.825 1111.600 695.995 1111.770 ;
        RECT 696.285 1111.600 696.455 1111.770 ;
        RECT 696.745 1111.600 696.915 1111.770 ;
        RECT 697.205 1111.600 697.375 1111.770 ;
        RECT 697.665 1111.600 697.835 1111.770 ;
        RECT 698.125 1111.600 698.295 1111.770 ;
        RECT 698.585 1111.600 698.755 1111.770 ;
        RECT 699.045 1111.600 699.215 1111.770 ;
        RECT 699.505 1111.600 699.675 1111.770 ;
        RECT 699.965 1111.600 700.135 1111.770 ;
        RECT 700.425 1111.600 700.595 1111.770 ;
        RECT 700.885 1111.600 701.055 1111.770 ;
        RECT 701.345 1111.600 701.515 1111.770 ;
        RECT 701.805 1111.600 701.975 1111.770 ;
        RECT 702.265 1111.600 702.435 1111.770 ;
        RECT 702.725 1111.600 702.895 1111.770 ;
        RECT 703.185 1111.600 703.355 1111.770 ;
        RECT 703.645 1111.600 703.815 1111.770 ;
        RECT 704.105 1111.600 704.275 1111.770 ;
        RECT 704.565 1111.600 704.735 1111.770 ;
        RECT 705.025 1111.600 705.195 1111.770 ;
        RECT 705.485 1111.600 705.655 1111.770 ;
        RECT 705.945 1111.600 706.115 1111.770 ;
        RECT 706.405 1111.600 706.575 1111.770 ;
        RECT 706.865 1111.600 707.035 1111.770 ;
        RECT 707.325 1111.600 707.495 1111.770 ;
        RECT 707.785 1111.600 707.955 1111.770 ;
        RECT 708.245 1111.600 708.415 1111.770 ;
        RECT 708.705 1111.600 708.875 1111.770 ;
        RECT 709.165 1111.600 709.335 1111.770 ;
        RECT 709.625 1111.600 709.795 1111.770 ;
        RECT 710.085 1111.600 710.255 1111.770 ;
        RECT 710.545 1111.600 710.715 1111.770 ;
        RECT 711.005 1111.600 711.175 1111.770 ;
        RECT 711.465 1111.600 711.635 1111.770 ;
        RECT 711.925 1111.600 712.095 1111.770 ;
        RECT 712.385 1111.600 712.555 1111.770 ;
        RECT 712.845 1111.600 713.015 1111.770 ;
        RECT 713.305 1111.600 713.475 1111.770 ;
        RECT 713.765 1111.600 713.935 1111.770 ;
        RECT 714.225 1111.600 714.395 1111.770 ;
        RECT 714.685 1111.600 714.855 1111.770 ;
        RECT 715.145 1111.600 715.315 1111.770 ;
        RECT 715.605 1111.600 715.775 1111.770 ;
        RECT 716.065 1111.600 716.235 1111.770 ;
        RECT 716.525 1111.600 716.695 1111.770 ;
        RECT 716.985 1111.600 717.155 1111.770 ;
        RECT 717.445 1111.600 717.615 1111.770 ;
        RECT 717.905 1111.600 718.075 1111.770 ;
        RECT 718.365 1111.600 718.535 1111.770 ;
        RECT 718.825 1111.600 718.995 1111.770 ;
        RECT 719.285 1111.600 719.455 1111.770 ;
        RECT 719.745 1111.600 719.915 1111.770 ;
        RECT 720.205 1111.600 720.375 1111.770 ;
        RECT 720.665 1111.600 720.835 1111.770 ;
        RECT 721.125 1111.600 721.295 1111.770 ;
        RECT 721.585 1111.600 721.755 1111.770 ;
        RECT 722.045 1111.600 722.215 1111.770 ;
        RECT 722.505 1111.600 722.675 1111.770 ;
        RECT 722.965 1111.600 723.135 1111.770 ;
        RECT 723.425 1111.600 723.595 1111.770 ;
        RECT 723.885 1111.600 724.055 1111.770 ;
        RECT 724.345 1111.600 724.515 1111.770 ;
        RECT 724.805 1111.600 724.975 1111.770 ;
        RECT 725.265 1111.600 725.435 1111.770 ;
        RECT 725.725 1111.600 725.895 1111.770 ;
        RECT 726.185 1111.600 726.355 1111.770 ;
        RECT 726.645 1111.600 726.815 1111.770 ;
        RECT 727.105 1111.600 727.275 1111.770 ;
        RECT 727.565 1111.600 727.735 1111.770 ;
        RECT 728.025 1111.600 728.195 1111.770 ;
        RECT 728.485 1111.600 728.655 1111.770 ;
        RECT 728.945 1111.600 729.115 1111.770 ;
        RECT 729.405 1111.600 729.575 1111.770 ;
        RECT 729.865 1111.600 730.035 1111.770 ;
        RECT 730.325 1111.600 730.495 1111.770 ;
        RECT 730.785 1111.600 730.955 1111.770 ;
        RECT 731.245 1111.600 731.415 1111.770 ;
        RECT 731.705 1111.600 731.875 1111.770 ;
        RECT 732.165 1111.600 732.335 1111.770 ;
        RECT 732.625 1111.600 732.795 1111.770 ;
        RECT 733.085 1111.600 733.255 1111.770 ;
        RECT 733.545 1111.600 733.715 1111.770 ;
        RECT 734.005 1111.600 734.175 1111.770 ;
        RECT 734.465 1111.600 734.635 1111.770 ;
        RECT 734.925 1111.600 735.095 1111.770 ;
        RECT 735.385 1111.600 735.555 1111.770 ;
        RECT 735.845 1111.600 736.015 1111.770 ;
        RECT 736.305 1111.600 736.475 1111.770 ;
        RECT 736.765 1111.600 736.935 1111.770 ;
        RECT 737.225 1111.600 737.395 1111.770 ;
        RECT 737.685 1111.600 737.855 1111.770 ;
        RECT 738.145 1111.600 738.315 1111.770 ;
        RECT 738.605 1111.600 738.775 1111.770 ;
        RECT 739.065 1111.600 739.235 1111.770 ;
        RECT 739.525 1111.600 739.695 1111.770 ;
        RECT 739.985 1111.600 740.155 1111.770 ;
        RECT 740.445 1111.600 740.615 1111.770 ;
        RECT 740.905 1111.600 741.075 1111.770 ;
        RECT 741.365 1111.600 741.535 1111.770 ;
        RECT 741.825 1111.600 741.995 1111.770 ;
        RECT 742.285 1111.600 742.455 1111.770 ;
        RECT 742.745 1111.600 742.915 1111.770 ;
        RECT 743.205 1111.600 743.375 1111.770 ;
        RECT 743.665 1111.600 743.835 1111.770 ;
        RECT 744.125 1111.600 744.295 1111.770 ;
        RECT 744.585 1111.600 744.755 1111.770 ;
        RECT 745.045 1111.600 745.215 1111.770 ;
        RECT 745.505 1111.600 745.675 1111.770 ;
        RECT 745.965 1111.600 746.135 1111.770 ;
        RECT 746.425 1111.600 746.595 1111.770 ;
        RECT 746.885 1111.600 747.055 1111.770 ;
        RECT 747.345 1111.600 747.515 1111.770 ;
        RECT 747.805 1111.600 747.975 1111.770 ;
        RECT 748.265 1111.600 748.435 1111.770 ;
        RECT 748.725 1111.600 748.895 1111.770 ;
        RECT 749.185 1111.600 749.355 1111.770 ;
        RECT 749.645 1111.600 749.815 1111.770 ;
        RECT 750.105 1111.600 750.275 1111.770 ;
        RECT 750.565 1111.600 750.735 1111.770 ;
        RECT 751.025 1111.600 751.195 1111.770 ;
        RECT 751.485 1111.600 751.655 1111.770 ;
        RECT 751.945 1111.600 752.115 1111.770 ;
        RECT 752.405 1111.600 752.575 1111.770 ;
        RECT 752.865 1111.600 753.035 1111.770 ;
        RECT 753.325 1111.600 753.495 1111.770 ;
        RECT 753.785 1111.600 753.955 1111.770 ;
        RECT 754.245 1111.600 754.415 1111.770 ;
        RECT 754.705 1111.600 754.875 1111.770 ;
        RECT 755.165 1111.600 755.335 1111.770 ;
        RECT 755.625 1111.600 755.795 1111.770 ;
        RECT 756.085 1111.600 756.255 1111.770 ;
        RECT 756.545 1111.600 756.715 1111.770 ;
        RECT 757.005 1111.600 757.175 1111.770 ;
        RECT 757.465 1111.600 757.635 1111.770 ;
        RECT 757.925 1111.600 758.095 1111.770 ;
        RECT 758.385 1111.600 758.555 1111.770 ;
        RECT 758.845 1111.600 759.015 1111.770 ;
        RECT 759.305 1111.600 759.475 1111.770 ;
        RECT 759.765 1111.600 759.935 1111.770 ;
        RECT 760.225 1111.600 760.395 1111.770 ;
        RECT 760.685 1111.600 760.855 1111.770 ;
        RECT 761.145 1111.600 761.315 1111.770 ;
        RECT 761.605 1111.600 761.775 1111.770 ;
        RECT 762.065 1111.600 762.235 1111.770 ;
        RECT 762.525 1111.600 762.695 1111.770 ;
        RECT 762.985 1111.600 763.155 1111.770 ;
        RECT 763.445 1111.600 763.615 1111.770 ;
        RECT 763.905 1111.600 764.075 1111.770 ;
        RECT 764.365 1111.600 764.535 1111.770 ;
        RECT 764.825 1111.600 764.995 1111.770 ;
        RECT 765.285 1111.600 765.455 1111.770 ;
        RECT 765.745 1111.600 765.915 1111.770 ;
        RECT 766.205 1111.600 766.375 1111.770 ;
        RECT 766.665 1111.600 766.835 1111.770 ;
        RECT 767.125 1111.600 767.295 1111.770 ;
        RECT 767.585 1111.600 767.755 1111.770 ;
        RECT 768.045 1111.600 768.215 1111.770 ;
        RECT 768.505 1111.600 768.675 1111.770 ;
        RECT 768.965 1111.600 769.135 1111.770 ;
        RECT 769.425 1111.600 769.595 1111.770 ;
        RECT 769.885 1111.600 770.055 1111.770 ;
        RECT 770.345 1111.600 770.515 1111.770 ;
        RECT 770.805 1111.600 770.975 1111.770 ;
      LAYER met1 ;
        RECT 669.000 1116.885 771.120 1117.365 ;
        RECT 674.980 1111.445 771.120 1111.925 ;
      LAYER via ;
        RECT 736.975 1116.985 738.760 1117.285 ;
        RECT 736.975 1111.575 738.760 1111.875 ;
      LAYER met2 ;
        RECT 736.975 1116.985 738.760 1117.285 ;
        RECT 736.935 1111.490 738.800 1111.920 ;
      LAYER via2 ;
        RECT 736.975 1111.575 738.760 1111.875 ;
      LAYER met3 ;
        RECT 736.940 1109.835 738.805 1117.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 1969.145 1117.040 1969.315 1117.210 ;
        RECT 1969.605 1117.040 1969.775 1117.210 ;
        RECT 1970.065 1117.040 1970.235 1117.210 ;
        RECT 1970.525 1117.040 1970.695 1117.210 ;
        RECT 1970.985 1117.040 1971.155 1117.210 ;
        RECT 1971.445 1117.040 1971.615 1117.210 ;
        RECT 1971.905 1117.040 1972.075 1117.210 ;
        RECT 1972.365 1117.040 1972.535 1117.210 ;
        RECT 1972.825 1117.040 1972.995 1117.210 ;
        RECT 1973.285 1117.040 1973.455 1117.210 ;
        RECT 1973.745 1117.040 1973.915 1117.210 ;
        RECT 1974.205 1117.040 1974.375 1117.210 ;
        RECT 1974.665 1117.040 1974.835 1117.210 ;
        RECT 1975.125 1117.040 1975.295 1117.210 ;
        RECT 1975.585 1117.040 1975.755 1117.210 ;
        RECT 1976.045 1117.040 1976.215 1117.210 ;
        RECT 1976.505 1117.040 1976.675 1117.210 ;
        RECT 1976.965 1117.040 1977.135 1117.210 ;
        RECT 1977.425 1117.040 1977.595 1117.210 ;
        RECT 1977.885 1117.040 1978.055 1117.210 ;
        RECT 1978.345 1117.040 1978.515 1117.210 ;
        RECT 1978.805 1117.040 1978.975 1117.210 ;
        RECT 1979.265 1117.040 1979.435 1117.210 ;
        RECT 1979.725 1117.040 1979.895 1117.210 ;
        RECT 1980.185 1117.040 1980.355 1117.210 ;
        RECT 1980.645 1117.040 1980.815 1117.210 ;
        RECT 1981.105 1117.040 1981.275 1117.210 ;
        RECT 1981.565 1117.040 1981.735 1117.210 ;
        RECT 1982.025 1117.040 1982.195 1117.210 ;
        RECT 1982.485 1117.040 1982.655 1117.210 ;
        RECT 1982.945 1117.040 1983.115 1117.210 ;
        RECT 1983.405 1117.040 1983.575 1117.210 ;
        RECT 1983.865 1117.040 1984.035 1117.210 ;
        RECT 1984.325 1117.040 1984.495 1117.210 ;
        RECT 1984.785 1117.040 1984.955 1117.210 ;
        RECT 1985.245 1117.040 1985.415 1117.210 ;
        RECT 1985.705 1117.040 1985.875 1117.210 ;
        RECT 1986.165 1117.040 1986.335 1117.210 ;
        RECT 1986.625 1117.040 1986.795 1117.210 ;
        RECT 1987.085 1117.040 1987.255 1117.210 ;
        RECT 1987.545 1117.040 1987.715 1117.210 ;
        RECT 1988.005 1117.040 1988.175 1117.210 ;
        RECT 1988.465 1117.040 1988.635 1117.210 ;
        RECT 1988.925 1117.040 1989.095 1117.210 ;
        RECT 1989.385 1117.040 1989.555 1117.210 ;
        RECT 1989.845 1117.040 1990.015 1117.210 ;
        RECT 1990.305 1117.040 1990.475 1117.210 ;
        RECT 1990.765 1117.040 1990.935 1117.210 ;
        RECT 1991.225 1117.040 1991.395 1117.210 ;
        RECT 1991.685 1117.040 1991.855 1117.210 ;
        RECT 1992.145 1117.040 1992.315 1117.210 ;
        RECT 1992.605 1117.040 1992.775 1117.210 ;
        RECT 1993.065 1117.040 1993.235 1117.210 ;
        RECT 1993.525 1117.040 1993.695 1117.210 ;
        RECT 1993.985 1117.040 1994.155 1117.210 ;
        RECT 1994.445 1117.040 1994.615 1117.210 ;
        RECT 1994.905 1117.040 1995.075 1117.210 ;
        RECT 1995.365 1117.040 1995.535 1117.210 ;
        RECT 1995.825 1117.040 1995.995 1117.210 ;
        RECT 1996.285 1117.040 1996.455 1117.210 ;
        RECT 1996.745 1117.040 1996.915 1117.210 ;
        RECT 1997.205 1117.040 1997.375 1117.210 ;
        RECT 1997.665 1117.040 1997.835 1117.210 ;
        RECT 1998.125 1117.040 1998.295 1117.210 ;
        RECT 1998.585 1117.040 1998.755 1117.210 ;
        RECT 1999.045 1117.040 1999.215 1117.210 ;
        RECT 1999.505 1117.040 1999.675 1117.210 ;
        RECT 1999.965 1117.040 2000.135 1117.210 ;
        RECT 2000.425 1117.040 2000.595 1117.210 ;
        RECT 2000.885 1117.040 2001.055 1117.210 ;
        RECT 2001.345 1117.040 2001.515 1117.210 ;
        RECT 2001.805 1117.040 2001.975 1117.210 ;
        RECT 2002.265 1117.040 2002.435 1117.210 ;
        RECT 2002.725 1117.040 2002.895 1117.210 ;
        RECT 2003.185 1117.040 2003.355 1117.210 ;
        RECT 2003.645 1117.040 2003.815 1117.210 ;
        RECT 2004.105 1117.040 2004.275 1117.210 ;
        RECT 2004.565 1117.040 2004.735 1117.210 ;
        RECT 2005.025 1117.040 2005.195 1117.210 ;
        RECT 2005.485 1117.040 2005.655 1117.210 ;
        RECT 2005.945 1117.040 2006.115 1117.210 ;
        RECT 2006.405 1117.040 2006.575 1117.210 ;
        RECT 2006.865 1117.040 2007.035 1117.210 ;
        RECT 2007.325 1117.040 2007.495 1117.210 ;
        RECT 2007.785 1117.040 2007.955 1117.210 ;
        RECT 2008.245 1117.040 2008.415 1117.210 ;
        RECT 2008.705 1117.040 2008.875 1117.210 ;
        RECT 2009.165 1117.040 2009.335 1117.210 ;
        RECT 2009.625 1117.040 2009.795 1117.210 ;
        RECT 2010.085 1117.040 2010.255 1117.210 ;
        RECT 2010.545 1117.040 2010.715 1117.210 ;
        RECT 2011.005 1117.040 2011.175 1117.210 ;
        RECT 2011.465 1117.040 2011.635 1117.210 ;
        RECT 2011.925 1117.040 2012.095 1117.210 ;
        RECT 2012.385 1117.040 2012.555 1117.210 ;
        RECT 2012.845 1117.040 2013.015 1117.210 ;
        RECT 2013.305 1117.040 2013.475 1117.210 ;
        RECT 2013.765 1117.040 2013.935 1117.210 ;
        RECT 2014.225 1117.040 2014.395 1117.210 ;
        RECT 2014.685 1117.040 2014.855 1117.210 ;
        RECT 2015.145 1117.040 2015.315 1117.210 ;
        RECT 2015.605 1117.040 2015.775 1117.210 ;
        RECT 2016.065 1117.040 2016.235 1117.210 ;
        RECT 2016.525 1117.040 2016.695 1117.210 ;
        RECT 2016.985 1117.040 2017.155 1117.210 ;
        RECT 2017.445 1117.040 2017.615 1117.210 ;
        RECT 2017.905 1117.040 2018.075 1117.210 ;
        RECT 2018.365 1117.040 2018.535 1117.210 ;
        RECT 2018.825 1117.040 2018.995 1117.210 ;
        RECT 2019.285 1117.040 2019.455 1117.210 ;
        RECT 2019.745 1117.040 2019.915 1117.210 ;
        RECT 2020.205 1117.040 2020.375 1117.210 ;
        RECT 2020.665 1117.040 2020.835 1117.210 ;
        RECT 2021.125 1117.040 2021.295 1117.210 ;
        RECT 2021.585 1117.040 2021.755 1117.210 ;
        RECT 2022.045 1117.040 2022.215 1117.210 ;
        RECT 2022.505 1117.040 2022.675 1117.210 ;
        RECT 2022.965 1117.040 2023.135 1117.210 ;
        RECT 2023.425 1117.040 2023.595 1117.210 ;
        RECT 2023.885 1117.040 2024.055 1117.210 ;
        RECT 2024.345 1117.040 2024.515 1117.210 ;
        RECT 2024.805 1117.040 2024.975 1117.210 ;
        RECT 2025.265 1117.040 2025.435 1117.210 ;
        RECT 2025.725 1117.040 2025.895 1117.210 ;
        RECT 2026.185 1117.040 2026.355 1117.210 ;
        RECT 2026.645 1117.040 2026.815 1117.210 ;
        RECT 2027.105 1117.040 2027.275 1117.210 ;
        RECT 2027.565 1117.040 2027.735 1117.210 ;
        RECT 2028.025 1117.040 2028.195 1117.210 ;
        RECT 2028.485 1117.040 2028.655 1117.210 ;
        RECT 2028.945 1117.040 2029.115 1117.210 ;
        RECT 2029.405 1117.040 2029.575 1117.210 ;
        RECT 2029.865 1117.040 2030.035 1117.210 ;
        RECT 2030.325 1117.040 2030.495 1117.210 ;
        RECT 2030.785 1117.040 2030.955 1117.210 ;
        RECT 2031.245 1117.040 2031.415 1117.210 ;
        RECT 2031.705 1117.040 2031.875 1117.210 ;
        RECT 2032.165 1117.040 2032.335 1117.210 ;
        RECT 2032.625 1117.040 2032.795 1117.210 ;
        RECT 2033.085 1117.040 2033.255 1117.210 ;
        RECT 2033.545 1117.040 2033.715 1117.210 ;
        RECT 2034.005 1117.040 2034.175 1117.210 ;
        RECT 2034.465 1117.040 2034.635 1117.210 ;
        RECT 2034.925 1117.040 2035.095 1117.210 ;
        RECT 2035.385 1117.040 2035.555 1117.210 ;
        RECT 2035.845 1117.040 2036.015 1117.210 ;
        RECT 2036.305 1117.040 2036.475 1117.210 ;
        RECT 2036.765 1117.040 2036.935 1117.210 ;
        RECT 2037.225 1117.040 2037.395 1117.210 ;
        RECT 2037.685 1117.040 2037.855 1117.210 ;
        RECT 2038.145 1117.040 2038.315 1117.210 ;
        RECT 2038.605 1117.040 2038.775 1117.210 ;
        RECT 2039.065 1117.040 2039.235 1117.210 ;
        RECT 2039.525 1117.040 2039.695 1117.210 ;
        RECT 2039.985 1117.040 2040.155 1117.210 ;
        RECT 2040.445 1117.040 2040.615 1117.210 ;
        RECT 2040.905 1117.040 2041.075 1117.210 ;
        RECT 2041.365 1117.040 2041.535 1117.210 ;
        RECT 2041.825 1117.040 2041.995 1117.210 ;
        RECT 2042.285 1117.040 2042.455 1117.210 ;
        RECT 2042.745 1117.040 2042.915 1117.210 ;
        RECT 2043.205 1117.040 2043.375 1117.210 ;
        RECT 2043.665 1117.040 2043.835 1117.210 ;
        RECT 2044.125 1117.040 2044.295 1117.210 ;
        RECT 2044.585 1117.040 2044.755 1117.210 ;
        RECT 2045.045 1117.040 2045.215 1117.210 ;
        RECT 2045.505 1117.040 2045.675 1117.210 ;
        RECT 2045.965 1117.040 2046.135 1117.210 ;
        RECT 2046.425 1117.040 2046.595 1117.210 ;
        RECT 2046.885 1117.040 2047.055 1117.210 ;
        RECT 2047.345 1117.040 2047.515 1117.210 ;
        RECT 2047.805 1117.040 2047.975 1117.210 ;
        RECT 2048.265 1117.040 2048.435 1117.210 ;
        RECT 2048.725 1117.040 2048.895 1117.210 ;
        RECT 2049.185 1117.040 2049.355 1117.210 ;
        RECT 2049.645 1117.040 2049.815 1117.210 ;
        RECT 2050.105 1117.040 2050.275 1117.210 ;
        RECT 2050.565 1117.040 2050.735 1117.210 ;
        RECT 2051.025 1117.040 2051.195 1117.210 ;
        RECT 2051.485 1117.040 2051.655 1117.210 ;
        RECT 2051.945 1117.040 2052.115 1117.210 ;
        RECT 2052.405 1117.040 2052.575 1117.210 ;
        RECT 2052.865 1117.040 2053.035 1117.210 ;
        RECT 2053.325 1117.040 2053.495 1117.210 ;
        RECT 2053.785 1117.040 2053.955 1117.210 ;
        RECT 2054.245 1117.040 2054.415 1117.210 ;
        RECT 2054.705 1117.040 2054.875 1117.210 ;
        RECT 2055.165 1117.040 2055.335 1117.210 ;
        RECT 2055.625 1117.040 2055.795 1117.210 ;
        RECT 2056.085 1117.040 2056.255 1117.210 ;
        RECT 2056.545 1117.040 2056.715 1117.210 ;
        RECT 2057.005 1117.040 2057.175 1117.210 ;
        RECT 2057.465 1117.040 2057.635 1117.210 ;
        RECT 2057.925 1117.040 2058.095 1117.210 ;
        RECT 2058.385 1117.040 2058.555 1117.210 ;
        RECT 2058.845 1117.040 2059.015 1117.210 ;
        RECT 2059.305 1117.040 2059.475 1117.210 ;
        RECT 2059.765 1117.040 2059.935 1117.210 ;
        RECT 2060.225 1117.040 2060.395 1117.210 ;
        RECT 2060.685 1117.040 2060.855 1117.210 ;
        RECT 2061.145 1117.040 2061.315 1117.210 ;
        RECT 2061.605 1117.040 2061.775 1117.210 ;
        RECT 2062.065 1117.040 2062.235 1117.210 ;
        RECT 2062.525 1117.040 2062.695 1117.210 ;
        RECT 2062.985 1117.040 2063.155 1117.210 ;
        RECT 2063.445 1117.040 2063.615 1117.210 ;
        RECT 2063.905 1117.040 2064.075 1117.210 ;
        RECT 2064.365 1117.040 2064.535 1117.210 ;
        RECT 2064.825 1117.040 2064.995 1117.210 ;
        RECT 2065.285 1117.040 2065.455 1117.210 ;
        RECT 2065.745 1117.040 2065.915 1117.210 ;
        RECT 2066.205 1117.040 2066.375 1117.210 ;
        RECT 2066.665 1117.040 2066.835 1117.210 ;
        RECT 2067.125 1117.040 2067.295 1117.210 ;
        RECT 2067.585 1117.040 2067.755 1117.210 ;
        RECT 2068.045 1117.040 2068.215 1117.210 ;
        RECT 2068.505 1117.040 2068.675 1117.210 ;
        RECT 2068.965 1117.040 2069.135 1117.210 ;
        RECT 2069.425 1117.040 2069.595 1117.210 ;
        RECT 2069.885 1117.040 2070.055 1117.210 ;
        RECT 2070.345 1117.040 2070.515 1117.210 ;
        RECT 2070.805 1117.040 2070.975 1117.210 ;
        RECT 1975.125 1111.600 1975.295 1111.770 ;
        RECT 1975.585 1111.600 1975.755 1111.770 ;
        RECT 1976.045 1111.600 1976.215 1111.770 ;
        RECT 1976.505 1111.600 1976.675 1111.770 ;
        RECT 1976.965 1111.600 1977.135 1111.770 ;
        RECT 1977.425 1111.600 1977.595 1111.770 ;
        RECT 1977.885 1111.600 1978.055 1111.770 ;
        RECT 1978.345 1111.600 1978.515 1111.770 ;
        RECT 1978.805 1111.600 1978.975 1111.770 ;
        RECT 1979.265 1111.600 1979.435 1111.770 ;
        RECT 1979.725 1111.600 1979.895 1111.770 ;
        RECT 1980.185 1111.600 1980.355 1111.770 ;
        RECT 1980.645 1111.600 1980.815 1111.770 ;
        RECT 1981.105 1111.600 1981.275 1111.770 ;
        RECT 1981.565 1111.600 1981.735 1111.770 ;
        RECT 1982.025 1111.600 1982.195 1111.770 ;
        RECT 1982.485 1111.600 1982.655 1111.770 ;
        RECT 1982.945 1111.600 1983.115 1111.770 ;
        RECT 1983.405 1111.600 1983.575 1111.770 ;
        RECT 1983.865 1111.600 1984.035 1111.770 ;
        RECT 1984.325 1111.600 1984.495 1111.770 ;
        RECT 1984.785 1111.600 1984.955 1111.770 ;
        RECT 1985.245 1111.600 1985.415 1111.770 ;
        RECT 1985.705 1111.600 1985.875 1111.770 ;
        RECT 1986.165 1111.600 1986.335 1111.770 ;
        RECT 1986.625 1111.600 1986.795 1111.770 ;
        RECT 1987.085 1111.600 1987.255 1111.770 ;
        RECT 1987.545 1111.600 1987.715 1111.770 ;
        RECT 1988.005 1111.600 1988.175 1111.770 ;
        RECT 1988.465 1111.600 1988.635 1111.770 ;
        RECT 1988.925 1111.600 1989.095 1111.770 ;
        RECT 1989.385 1111.600 1989.555 1111.770 ;
        RECT 1989.845 1111.600 1990.015 1111.770 ;
        RECT 1990.305 1111.600 1990.475 1111.770 ;
        RECT 1990.765 1111.600 1990.935 1111.770 ;
        RECT 1991.225 1111.600 1991.395 1111.770 ;
        RECT 1991.685 1111.600 1991.855 1111.770 ;
        RECT 1992.145 1111.600 1992.315 1111.770 ;
        RECT 1992.605 1111.600 1992.775 1111.770 ;
        RECT 1993.065 1111.600 1993.235 1111.770 ;
        RECT 1993.525 1111.600 1993.695 1111.770 ;
        RECT 1993.985 1111.600 1994.155 1111.770 ;
        RECT 1994.445 1111.600 1994.615 1111.770 ;
        RECT 1994.905 1111.600 1995.075 1111.770 ;
        RECT 1995.365 1111.600 1995.535 1111.770 ;
        RECT 1995.825 1111.600 1995.995 1111.770 ;
        RECT 1996.285 1111.600 1996.455 1111.770 ;
        RECT 1996.745 1111.600 1996.915 1111.770 ;
        RECT 1997.205 1111.600 1997.375 1111.770 ;
        RECT 1997.665 1111.600 1997.835 1111.770 ;
        RECT 1998.125 1111.600 1998.295 1111.770 ;
        RECT 1998.585 1111.600 1998.755 1111.770 ;
        RECT 1999.045 1111.600 1999.215 1111.770 ;
        RECT 1999.505 1111.600 1999.675 1111.770 ;
        RECT 1999.965 1111.600 2000.135 1111.770 ;
        RECT 2000.425 1111.600 2000.595 1111.770 ;
        RECT 2000.885 1111.600 2001.055 1111.770 ;
        RECT 2001.345 1111.600 2001.515 1111.770 ;
        RECT 2001.805 1111.600 2001.975 1111.770 ;
        RECT 2002.265 1111.600 2002.435 1111.770 ;
        RECT 2002.725 1111.600 2002.895 1111.770 ;
        RECT 2003.185 1111.600 2003.355 1111.770 ;
        RECT 2003.645 1111.600 2003.815 1111.770 ;
        RECT 2004.105 1111.600 2004.275 1111.770 ;
        RECT 2004.565 1111.600 2004.735 1111.770 ;
        RECT 2005.025 1111.600 2005.195 1111.770 ;
        RECT 2005.485 1111.600 2005.655 1111.770 ;
        RECT 2005.945 1111.600 2006.115 1111.770 ;
        RECT 2006.405 1111.600 2006.575 1111.770 ;
        RECT 2006.865 1111.600 2007.035 1111.770 ;
        RECT 2007.325 1111.600 2007.495 1111.770 ;
        RECT 2007.785 1111.600 2007.955 1111.770 ;
        RECT 2008.245 1111.600 2008.415 1111.770 ;
        RECT 2008.705 1111.600 2008.875 1111.770 ;
        RECT 2009.165 1111.600 2009.335 1111.770 ;
        RECT 2009.625 1111.600 2009.795 1111.770 ;
        RECT 2010.085 1111.600 2010.255 1111.770 ;
        RECT 2010.545 1111.600 2010.715 1111.770 ;
        RECT 2011.005 1111.600 2011.175 1111.770 ;
        RECT 2011.465 1111.600 2011.635 1111.770 ;
        RECT 2011.925 1111.600 2012.095 1111.770 ;
        RECT 2012.385 1111.600 2012.555 1111.770 ;
        RECT 2012.845 1111.600 2013.015 1111.770 ;
        RECT 2013.305 1111.600 2013.475 1111.770 ;
        RECT 2013.765 1111.600 2013.935 1111.770 ;
        RECT 2014.225 1111.600 2014.395 1111.770 ;
        RECT 2014.685 1111.600 2014.855 1111.770 ;
        RECT 2015.145 1111.600 2015.315 1111.770 ;
        RECT 2015.605 1111.600 2015.775 1111.770 ;
        RECT 2016.065 1111.600 2016.235 1111.770 ;
        RECT 2016.525 1111.600 2016.695 1111.770 ;
        RECT 2016.985 1111.600 2017.155 1111.770 ;
        RECT 2017.445 1111.600 2017.615 1111.770 ;
        RECT 2017.905 1111.600 2018.075 1111.770 ;
        RECT 2018.365 1111.600 2018.535 1111.770 ;
        RECT 2018.825 1111.600 2018.995 1111.770 ;
        RECT 2019.285 1111.600 2019.455 1111.770 ;
        RECT 2019.745 1111.600 2019.915 1111.770 ;
        RECT 2020.205 1111.600 2020.375 1111.770 ;
        RECT 2020.665 1111.600 2020.835 1111.770 ;
        RECT 2021.125 1111.600 2021.295 1111.770 ;
        RECT 2021.585 1111.600 2021.755 1111.770 ;
        RECT 2022.045 1111.600 2022.215 1111.770 ;
        RECT 2022.505 1111.600 2022.675 1111.770 ;
        RECT 2022.965 1111.600 2023.135 1111.770 ;
        RECT 2023.425 1111.600 2023.595 1111.770 ;
        RECT 2023.885 1111.600 2024.055 1111.770 ;
        RECT 2024.345 1111.600 2024.515 1111.770 ;
        RECT 2024.805 1111.600 2024.975 1111.770 ;
        RECT 2025.265 1111.600 2025.435 1111.770 ;
        RECT 2025.725 1111.600 2025.895 1111.770 ;
        RECT 2026.185 1111.600 2026.355 1111.770 ;
        RECT 2026.645 1111.600 2026.815 1111.770 ;
        RECT 2027.105 1111.600 2027.275 1111.770 ;
        RECT 2027.565 1111.600 2027.735 1111.770 ;
        RECT 2028.025 1111.600 2028.195 1111.770 ;
        RECT 2028.485 1111.600 2028.655 1111.770 ;
        RECT 2028.945 1111.600 2029.115 1111.770 ;
        RECT 2029.405 1111.600 2029.575 1111.770 ;
        RECT 2029.865 1111.600 2030.035 1111.770 ;
        RECT 2030.325 1111.600 2030.495 1111.770 ;
        RECT 2030.785 1111.600 2030.955 1111.770 ;
        RECT 2031.245 1111.600 2031.415 1111.770 ;
        RECT 2031.705 1111.600 2031.875 1111.770 ;
        RECT 2032.165 1111.600 2032.335 1111.770 ;
        RECT 2032.625 1111.600 2032.795 1111.770 ;
        RECT 2033.085 1111.600 2033.255 1111.770 ;
        RECT 2033.545 1111.600 2033.715 1111.770 ;
        RECT 2034.005 1111.600 2034.175 1111.770 ;
        RECT 2034.465 1111.600 2034.635 1111.770 ;
        RECT 2034.925 1111.600 2035.095 1111.770 ;
        RECT 2035.385 1111.600 2035.555 1111.770 ;
        RECT 2035.845 1111.600 2036.015 1111.770 ;
        RECT 2036.305 1111.600 2036.475 1111.770 ;
        RECT 2036.765 1111.600 2036.935 1111.770 ;
        RECT 2037.225 1111.600 2037.395 1111.770 ;
        RECT 2037.685 1111.600 2037.855 1111.770 ;
        RECT 2038.145 1111.600 2038.315 1111.770 ;
        RECT 2038.605 1111.600 2038.775 1111.770 ;
        RECT 2039.065 1111.600 2039.235 1111.770 ;
        RECT 2039.525 1111.600 2039.695 1111.770 ;
        RECT 2039.985 1111.600 2040.155 1111.770 ;
        RECT 2040.445 1111.600 2040.615 1111.770 ;
        RECT 2040.905 1111.600 2041.075 1111.770 ;
        RECT 2041.365 1111.600 2041.535 1111.770 ;
        RECT 2041.825 1111.600 2041.995 1111.770 ;
        RECT 2042.285 1111.600 2042.455 1111.770 ;
        RECT 2042.745 1111.600 2042.915 1111.770 ;
        RECT 2043.205 1111.600 2043.375 1111.770 ;
        RECT 2043.665 1111.600 2043.835 1111.770 ;
        RECT 2044.125 1111.600 2044.295 1111.770 ;
        RECT 2044.585 1111.600 2044.755 1111.770 ;
        RECT 2045.045 1111.600 2045.215 1111.770 ;
        RECT 2045.505 1111.600 2045.675 1111.770 ;
        RECT 2045.965 1111.600 2046.135 1111.770 ;
        RECT 2046.425 1111.600 2046.595 1111.770 ;
        RECT 2046.885 1111.600 2047.055 1111.770 ;
        RECT 2047.345 1111.600 2047.515 1111.770 ;
        RECT 2047.805 1111.600 2047.975 1111.770 ;
        RECT 2048.265 1111.600 2048.435 1111.770 ;
        RECT 2048.725 1111.600 2048.895 1111.770 ;
        RECT 2049.185 1111.600 2049.355 1111.770 ;
        RECT 2049.645 1111.600 2049.815 1111.770 ;
        RECT 2050.105 1111.600 2050.275 1111.770 ;
        RECT 2050.565 1111.600 2050.735 1111.770 ;
        RECT 2051.025 1111.600 2051.195 1111.770 ;
        RECT 2051.485 1111.600 2051.655 1111.770 ;
        RECT 2051.945 1111.600 2052.115 1111.770 ;
        RECT 2052.405 1111.600 2052.575 1111.770 ;
        RECT 2052.865 1111.600 2053.035 1111.770 ;
        RECT 2053.325 1111.600 2053.495 1111.770 ;
        RECT 2053.785 1111.600 2053.955 1111.770 ;
        RECT 2054.245 1111.600 2054.415 1111.770 ;
        RECT 2054.705 1111.600 2054.875 1111.770 ;
        RECT 2055.165 1111.600 2055.335 1111.770 ;
        RECT 2055.625 1111.600 2055.795 1111.770 ;
        RECT 2056.085 1111.600 2056.255 1111.770 ;
        RECT 2056.545 1111.600 2056.715 1111.770 ;
        RECT 2057.005 1111.600 2057.175 1111.770 ;
        RECT 2057.465 1111.600 2057.635 1111.770 ;
        RECT 2057.925 1111.600 2058.095 1111.770 ;
        RECT 2058.385 1111.600 2058.555 1111.770 ;
        RECT 2058.845 1111.600 2059.015 1111.770 ;
        RECT 2059.305 1111.600 2059.475 1111.770 ;
        RECT 2059.765 1111.600 2059.935 1111.770 ;
        RECT 2060.225 1111.600 2060.395 1111.770 ;
        RECT 2060.685 1111.600 2060.855 1111.770 ;
        RECT 2061.145 1111.600 2061.315 1111.770 ;
        RECT 2061.605 1111.600 2061.775 1111.770 ;
        RECT 2062.065 1111.600 2062.235 1111.770 ;
        RECT 2062.525 1111.600 2062.695 1111.770 ;
        RECT 2062.985 1111.600 2063.155 1111.770 ;
        RECT 2063.445 1111.600 2063.615 1111.770 ;
        RECT 2063.905 1111.600 2064.075 1111.770 ;
        RECT 2064.365 1111.600 2064.535 1111.770 ;
        RECT 2064.825 1111.600 2064.995 1111.770 ;
        RECT 2065.285 1111.600 2065.455 1111.770 ;
        RECT 2065.745 1111.600 2065.915 1111.770 ;
        RECT 2066.205 1111.600 2066.375 1111.770 ;
        RECT 2066.665 1111.600 2066.835 1111.770 ;
        RECT 2067.125 1111.600 2067.295 1111.770 ;
        RECT 2067.585 1111.600 2067.755 1111.770 ;
        RECT 2068.045 1111.600 2068.215 1111.770 ;
        RECT 2068.505 1111.600 2068.675 1111.770 ;
        RECT 2068.965 1111.600 2069.135 1111.770 ;
        RECT 2069.425 1111.600 2069.595 1111.770 ;
        RECT 2069.885 1111.600 2070.055 1111.770 ;
        RECT 2070.345 1111.600 2070.515 1111.770 ;
        RECT 2070.805 1111.600 2070.975 1111.770 ;
      LAYER met1 ;
        RECT 1969.000 1116.885 2071.120 1117.365 ;
        RECT 1974.980 1111.445 2071.120 1111.925 ;
      LAYER via ;
        RECT 2031.130 1116.950 2032.915 1117.250 ;
        RECT 2031.130 1111.540 2032.915 1111.840 ;
      LAYER met2 ;
        RECT 2031.090 1116.880 2032.955 1117.310 ;
        RECT 2031.090 1111.455 2032.955 1111.885 ;
      LAYER via2 ;
        RECT 2031.130 1116.950 2032.915 1117.250 ;
        RECT 2031.130 1111.540 2032.915 1111.840 ;
      LAYER met3 ;
        RECT 2031.095 1109.800 2032.960 1117.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 198.795 1732.850 198.965 1733.020 ;
        RECT 204.235 1732.850 204.405 1733.020 ;
        RECT 198.795 1732.390 198.965 1732.560 ;
        RECT 204.235 1732.390 204.405 1732.560 ;
        RECT 198.795 1731.930 198.965 1732.100 ;
        RECT 204.235 1731.930 204.405 1732.100 ;
        RECT 198.795 1731.470 198.965 1731.640 ;
        RECT 204.235 1731.470 204.405 1731.640 ;
        RECT 198.795 1731.010 198.965 1731.180 ;
        RECT 204.235 1731.010 204.405 1731.180 ;
        RECT 198.795 1730.550 198.965 1730.720 ;
        RECT 204.235 1730.550 204.405 1730.720 ;
        RECT 198.795 1730.090 198.965 1730.260 ;
        RECT 204.235 1730.090 204.405 1730.260 ;
        RECT 198.795 1729.630 198.965 1729.800 ;
        RECT 204.235 1729.630 204.405 1729.800 ;
        RECT 198.795 1729.170 198.965 1729.340 ;
        RECT 204.235 1729.170 204.405 1729.340 ;
        RECT 198.795 1728.710 198.965 1728.880 ;
        RECT 204.235 1728.710 204.405 1728.880 ;
        RECT 198.795 1728.250 198.965 1728.420 ;
        RECT 204.235 1728.250 204.405 1728.420 ;
        RECT 198.795 1727.790 198.965 1727.960 ;
        RECT 204.235 1727.790 204.405 1727.960 ;
        RECT 198.795 1727.330 198.965 1727.500 ;
        RECT 204.235 1727.330 204.405 1727.500 ;
        RECT 198.795 1726.870 198.965 1727.040 ;
        RECT 204.235 1726.870 204.405 1727.040 ;
        RECT 198.795 1726.410 198.965 1726.580 ;
        RECT 204.235 1726.410 204.405 1726.580 ;
        RECT 198.795 1725.950 198.965 1726.120 ;
        RECT 204.235 1725.950 204.405 1726.120 ;
        RECT 198.795 1725.490 198.965 1725.660 ;
        RECT 204.235 1725.490 204.405 1725.660 ;
        RECT 198.795 1725.030 198.965 1725.200 ;
        RECT 204.235 1725.030 204.405 1725.200 ;
        RECT 198.795 1724.570 198.965 1724.740 ;
        RECT 204.235 1724.570 204.405 1724.740 ;
        RECT 198.795 1724.110 198.965 1724.280 ;
        RECT 204.235 1724.110 204.405 1724.280 ;
        RECT 198.795 1723.650 198.965 1723.820 ;
        RECT 204.235 1723.650 204.405 1723.820 ;
        RECT 198.795 1723.190 198.965 1723.360 ;
        RECT 204.235 1723.190 204.405 1723.360 ;
        RECT 198.795 1722.730 198.965 1722.900 ;
        RECT 204.235 1722.730 204.405 1722.900 ;
        RECT 198.795 1722.270 198.965 1722.440 ;
        RECT 204.235 1722.270 204.405 1722.440 ;
        RECT 198.795 1721.810 198.965 1721.980 ;
        RECT 204.235 1721.810 204.405 1721.980 ;
        RECT 198.795 1721.350 198.965 1721.520 ;
        RECT 204.235 1721.350 204.405 1721.520 ;
        RECT 198.795 1720.890 198.965 1721.060 ;
        RECT 204.235 1720.890 204.405 1721.060 ;
        RECT 198.795 1720.430 198.965 1720.600 ;
        RECT 204.235 1720.430 204.405 1720.600 ;
        RECT 198.795 1719.970 198.965 1720.140 ;
        RECT 204.235 1719.970 204.405 1720.140 ;
        RECT 198.795 1719.510 198.965 1719.680 ;
        RECT 204.235 1719.510 204.405 1719.680 ;
        RECT 198.795 1719.050 198.965 1719.220 ;
        RECT 204.235 1719.050 204.405 1719.220 ;
        RECT 198.795 1718.590 198.965 1718.760 ;
        RECT 204.235 1718.590 204.405 1718.760 ;
        RECT 198.795 1718.130 198.965 1718.300 ;
        RECT 204.235 1718.130 204.405 1718.300 ;
        RECT 198.795 1717.670 198.965 1717.840 ;
        RECT 204.235 1717.670 204.405 1717.840 ;
        RECT 198.795 1717.210 198.965 1717.380 ;
        RECT 204.235 1717.210 204.405 1717.380 ;
        RECT 198.795 1716.750 198.965 1716.920 ;
        RECT 204.235 1716.750 204.405 1716.920 ;
        RECT 198.795 1716.290 198.965 1716.460 ;
        RECT 204.235 1716.290 204.405 1716.460 ;
        RECT 198.795 1715.830 198.965 1716.000 ;
        RECT 204.235 1715.830 204.405 1716.000 ;
        RECT 198.795 1715.370 198.965 1715.540 ;
        RECT 204.235 1715.370 204.405 1715.540 ;
        RECT 198.795 1714.910 198.965 1715.080 ;
        RECT 204.235 1714.910 204.405 1715.080 ;
        RECT 198.795 1714.450 198.965 1714.620 ;
        RECT 204.235 1714.450 204.405 1714.620 ;
        RECT 198.795 1713.990 198.965 1714.160 ;
        RECT 204.235 1713.990 204.405 1714.160 ;
        RECT 198.795 1713.530 198.965 1713.700 ;
        RECT 204.235 1713.530 204.405 1713.700 ;
        RECT 198.795 1713.070 198.965 1713.240 ;
        RECT 204.235 1713.070 204.405 1713.240 ;
        RECT 198.795 1712.610 198.965 1712.780 ;
        RECT 204.235 1712.610 204.405 1712.780 ;
        RECT 198.795 1712.150 198.965 1712.320 ;
        RECT 204.235 1712.150 204.405 1712.320 ;
        RECT 198.795 1711.690 198.965 1711.860 ;
        RECT 204.235 1711.690 204.405 1711.860 ;
        RECT 198.795 1711.230 198.965 1711.400 ;
        RECT 204.235 1711.230 204.405 1711.400 ;
        RECT 198.795 1710.770 198.965 1710.940 ;
        RECT 204.235 1710.770 204.405 1710.940 ;
        RECT 198.795 1710.310 198.965 1710.480 ;
        RECT 204.235 1710.310 204.405 1710.480 ;
        RECT 198.795 1709.850 198.965 1710.020 ;
        RECT 204.235 1709.850 204.405 1710.020 ;
        RECT 198.795 1709.390 198.965 1709.560 ;
        RECT 204.235 1709.390 204.405 1709.560 ;
        RECT 198.795 1708.930 198.965 1709.100 ;
        RECT 204.235 1708.930 204.405 1709.100 ;
        RECT 198.795 1708.470 198.965 1708.640 ;
        RECT 204.235 1708.470 204.405 1708.640 ;
        RECT 198.795 1708.010 198.965 1708.180 ;
        RECT 204.235 1708.010 204.405 1708.180 ;
        RECT 198.795 1707.550 198.965 1707.720 ;
        RECT 204.235 1707.550 204.405 1707.720 ;
        RECT 198.795 1707.090 198.965 1707.260 ;
        RECT 204.235 1707.090 204.405 1707.260 ;
        RECT 198.795 1706.630 198.965 1706.800 ;
        RECT 204.235 1706.630 204.405 1706.800 ;
        RECT 198.795 1706.170 198.965 1706.340 ;
        RECT 204.235 1706.170 204.405 1706.340 ;
        RECT 198.795 1705.710 198.965 1705.880 ;
        RECT 204.235 1705.710 204.405 1705.880 ;
        RECT 198.795 1705.250 198.965 1705.420 ;
        RECT 204.235 1705.250 204.405 1705.420 ;
        RECT 198.795 1704.790 198.965 1704.960 ;
        RECT 204.235 1704.790 204.405 1704.960 ;
        RECT 198.795 1704.330 198.965 1704.500 ;
        RECT 204.235 1704.330 204.405 1704.500 ;
        RECT 198.795 1703.870 198.965 1704.040 ;
        RECT 204.235 1703.870 204.405 1704.040 ;
        RECT 198.795 1703.410 198.965 1703.580 ;
        RECT 204.235 1703.410 204.405 1703.580 ;
        RECT 198.795 1702.950 198.965 1703.120 ;
        RECT 204.235 1702.950 204.405 1703.120 ;
        RECT 198.795 1702.490 198.965 1702.660 ;
        RECT 204.235 1702.490 204.405 1702.660 ;
        RECT 198.795 1702.030 198.965 1702.200 ;
        RECT 204.235 1702.030 204.405 1702.200 ;
        RECT 198.795 1701.570 198.965 1701.740 ;
        RECT 204.235 1701.570 204.405 1701.740 ;
        RECT 198.795 1701.110 198.965 1701.280 ;
        RECT 204.235 1701.110 204.405 1701.280 ;
        RECT 198.795 1700.650 198.965 1700.820 ;
        RECT 204.235 1700.650 204.405 1700.820 ;
        RECT 198.795 1700.190 198.965 1700.360 ;
        RECT 204.235 1700.190 204.405 1700.360 ;
        RECT 198.795 1699.730 198.965 1699.900 ;
        RECT 204.235 1699.730 204.405 1699.900 ;
        RECT 198.795 1699.270 198.965 1699.440 ;
        RECT 204.235 1699.270 204.405 1699.440 ;
        RECT 198.795 1698.810 198.965 1698.980 ;
        RECT 204.235 1698.810 204.405 1698.980 ;
        RECT 198.795 1698.350 198.965 1698.520 ;
        RECT 204.235 1698.350 204.405 1698.520 ;
        RECT 198.795 1697.890 198.965 1698.060 ;
        RECT 204.235 1697.890 204.405 1698.060 ;
        RECT 198.795 1697.430 198.965 1697.600 ;
        RECT 204.235 1697.430 204.405 1697.600 ;
        RECT 198.795 1696.970 198.965 1697.140 ;
        RECT 204.235 1696.970 204.405 1697.140 ;
        RECT 198.795 1696.510 198.965 1696.680 ;
        RECT 204.235 1696.510 204.405 1696.680 ;
        RECT 198.795 1696.050 198.965 1696.220 ;
        RECT 204.235 1696.050 204.405 1696.220 ;
        RECT 198.795 1695.590 198.965 1695.760 ;
        RECT 204.235 1695.590 204.405 1695.760 ;
        RECT 198.795 1695.130 198.965 1695.300 ;
        RECT 204.235 1695.130 204.405 1695.300 ;
        RECT 198.795 1694.670 198.965 1694.840 ;
        RECT 204.235 1694.670 204.405 1694.840 ;
        RECT 198.795 1694.210 198.965 1694.380 ;
        RECT 204.235 1694.210 204.405 1694.380 ;
        RECT 198.795 1693.750 198.965 1693.920 ;
        RECT 204.235 1693.750 204.405 1693.920 ;
        RECT 198.795 1693.290 198.965 1693.460 ;
        RECT 204.235 1693.290 204.405 1693.460 ;
        RECT 198.795 1692.830 198.965 1693.000 ;
        RECT 204.235 1692.830 204.405 1693.000 ;
        RECT 198.795 1692.370 198.965 1692.540 ;
        RECT 204.235 1692.370 204.405 1692.540 ;
        RECT 198.795 1691.910 198.965 1692.080 ;
        RECT 204.235 1691.910 204.405 1692.080 ;
        RECT 198.795 1691.450 198.965 1691.620 ;
        RECT 204.235 1691.450 204.405 1691.620 ;
        RECT 198.795 1690.990 198.965 1691.160 ;
        RECT 204.235 1690.990 204.405 1691.160 ;
        RECT 198.795 1690.530 198.965 1690.700 ;
        RECT 204.235 1690.530 204.405 1690.700 ;
        RECT 198.795 1690.070 198.965 1690.240 ;
        RECT 204.235 1690.070 204.405 1690.240 ;
        RECT 198.795 1689.610 198.965 1689.780 ;
        RECT 204.235 1689.610 204.405 1689.780 ;
        RECT 198.795 1689.150 198.965 1689.320 ;
        RECT 204.235 1689.150 204.405 1689.320 ;
        RECT 198.795 1688.690 198.965 1688.860 ;
        RECT 204.235 1688.690 204.405 1688.860 ;
        RECT 198.795 1688.230 198.965 1688.400 ;
        RECT 204.235 1688.230 204.405 1688.400 ;
        RECT 198.795 1687.770 198.965 1687.940 ;
        RECT 204.235 1687.770 204.405 1687.940 ;
        RECT 198.795 1687.310 198.965 1687.480 ;
        RECT 204.235 1687.310 204.405 1687.480 ;
        RECT 198.795 1686.850 198.965 1687.020 ;
        RECT 204.235 1686.850 204.405 1687.020 ;
        RECT 198.795 1686.390 198.965 1686.560 ;
        RECT 204.235 1686.390 204.405 1686.560 ;
        RECT 198.795 1685.930 198.965 1686.100 ;
        RECT 204.235 1685.930 204.405 1686.100 ;
        RECT 198.795 1685.470 198.965 1685.640 ;
        RECT 204.235 1685.470 204.405 1685.640 ;
        RECT 198.795 1685.010 198.965 1685.180 ;
        RECT 204.235 1685.010 204.405 1685.180 ;
        RECT 198.795 1684.550 198.965 1684.720 ;
        RECT 204.235 1684.550 204.405 1684.720 ;
        RECT 198.795 1684.090 198.965 1684.260 ;
        RECT 204.235 1684.090 204.405 1684.260 ;
        RECT 198.795 1683.630 198.965 1683.800 ;
        RECT 204.235 1683.630 204.405 1683.800 ;
        RECT 198.795 1683.170 198.965 1683.340 ;
        RECT 204.235 1683.170 204.405 1683.340 ;
        RECT 198.795 1682.710 198.965 1682.880 ;
        RECT 204.235 1682.710 204.405 1682.880 ;
        RECT 198.795 1682.250 198.965 1682.420 ;
        RECT 204.235 1682.250 204.405 1682.420 ;
        RECT 198.795 1681.790 198.965 1681.960 ;
        RECT 204.235 1681.790 204.405 1681.960 ;
        RECT 198.795 1681.330 198.965 1681.500 ;
        RECT 204.235 1681.330 204.405 1681.500 ;
        RECT 198.795 1680.870 198.965 1681.040 ;
        RECT 204.235 1680.870 204.405 1681.040 ;
        RECT 198.795 1680.410 198.965 1680.580 ;
        RECT 204.235 1680.410 204.405 1680.580 ;
        RECT 198.795 1679.950 198.965 1680.120 ;
        RECT 204.235 1679.950 204.405 1680.120 ;
        RECT 198.795 1679.490 198.965 1679.660 ;
        RECT 204.235 1679.490 204.405 1679.660 ;
        RECT 198.795 1679.030 198.965 1679.200 ;
        RECT 204.235 1679.030 204.405 1679.200 ;
        RECT 198.795 1678.570 198.965 1678.740 ;
        RECT 204.235 1678.570 204.405 1678.740 ;
        RECT 198.795 1678.110 198.965 1678.280 ;
        RECT 204.235 1678.110 204.405 1678.280 ;
        RECT 198.795 1677.650 198.965 1677.820 ;
        RECT 204.235 1677.650 204.405 1677.820 ;
        RECT 198.795 1677.190 198.965 1677.360 ;
        RECT 204.235 1677.190 204.405 1677.360 ;
        RECT 198.795 1676.730 198.965 1676.900 ;
        RECT 204.235 1676.730 204.405 1676.900 ;
        RECT 198.795 1676.270 198.965 1676.440 ;
        RECT 204.235 1676.270 204.405 1676.440 ;
        RECT 198.795 1675.810 198.965 1675.980 ;
        RECT 204.235 1675.810 204.405 1675.980 ;
        RECT 198.795 1675.350 198.965 1675.520 ;
        RECT 204.235 1675.350 204.405 1675.520 ;
        RECT 198.795 1674.890 198.965 1675.060 ;
        RECT 204.235 1674.890 204.405 1675.060 ;
        RECT 198.795 1674.430 198.965 1674.600 ;
        RECT 204.235 1674.430 204.405 1674.600 ;
        RECT 198.795 1673.970 198.965 1674.140 ;
        RECT 204.235 1673.970 204.405 1674.140 ;
        RECT 198.795 1673.510 198.965 1673.680 ;
        RECT 204.235 1673.510 204.405 1673.680 ;
        RECT 198.795 1673.050 198.965 1673.220 ;
        RECT 204.235 1673.050 204.405 1673.220 ;
      LAYER met1 ;
        RECT 198.640 1672.905 199.120 1733.165 ;
        RECT 204.080 1672.905 204.560 1733.165 ;
      LAYER via ;
        RECT 198.750 1710.875 199.050 1712.660 ;
        RECT 204.160 1710.875 204.460 1712.660 ;
      LAYER met2 ;
        RECT 198.665 1710.835 199.095 1712.700 ;
        RECT 204.090 1710.835 204.520 1712.700 ;
      LAYER via2 ;
        RECT 198.750 1710.875 199.050 1712.660 ;
        RECT 204.160 1710.875 204.460 1712.660 ;
      LAYER met3 ;
        RECT 197.010 1710.830 204.535 1712.695 ;
    END
    PORT
      LAYER li1 ;
        RECT 198.685 3023.755 198.855 3023.925 ;
        RECT 204.125 3023.755 204.295 3023.925 ;
        RECT 198.685 3023.295 198.855 3023.465 ;
        RECT 204.125 3023.295 204.295 3023.465 ;
        RECT 198.685 3022.835 198.855 3023.005 ;
        RECT 204.125 3022.835 204.295 3023.005 ;
        RECT 198.685 3022.375 198.855 3022.545 ;
        RECT 204.125 3022.375 204.295 3022.545 ;
        RECT 198.685 3021.915 198.855 3022.085 ;
        RECT 204.125 3021.915 204.295 3022.085 ;
        RECT 198.685 3021.455 198.855 3021.625 ;
        RECT 204.125 3021.455 204.295 3021.625 ;
        RECT 198.685 3020.995 198.855 3021.165 ;
        RECT 204.125 3020.995 204.295 3021.165 ;
        RECT 198.685 3020.535 198.855 3020.705 ;
        RECT 204.125 3020.535 204.295 3020.705 ;
        RECT 198.685 3020.075 198.855 3020.245 ;
        RECT 204.125 3020.075 204.295 3020.245 ;
        RECT 198.685 3019.615 198.855 3019.785 ;
        RECT 204.125 3019.615 204.295 3019.785 ;
        RECT 198.685 3019.155 198.855 3019.325 ;
        RECT 204.125 3019.155 204.295 3019.325 ;
        RECT 198.685 3018.695 198.855 3018.865 ;
        RECT 204.125 3018.695 204.295 3018.865 ;
        RECT 198.685 3018.235 198.855 3018.405 ;
        RECT 204.125 3018.235 204.295 3018.405 ;
        RECT 198.685 3017.775 198.855 3017.945 ;
        RECT 204.125 3017.775 204.295 3017.945 ;
        RECT 198.685 3017.315 198.855 3017.485 ;
        RECT 204.125 3017.315 204.295 3017.485 ;
        RECT 198.685 3016.855 198.855 3017.025 ;
        RECT 204.125 3016.855 204.295 3017.025 ;
        RECT 198.685 3016.395 198.855 3016.565 ;
        RECT 204.125 3016.395 204.295 3016.565 ;
        RECT 198.685 3015.935 198.855 3016.105 ;
        RECT 204.125 3015.935 204.295 3016.105 ;
        RECT 198.685 3015.475 198.855 3015.645 ;
        RECT 204.125 3015.475 204.295 3015.645 ;
        RECT 198.685 3015.015 198.855 3015.185 ;
        RECT 204.125 3015.015 204.295 3015.185 ;
        RECT 198.685 3014.555 198.855 3014.725 ;
        RECT 204.125 3014.555 204.295 3014.725 ;
        RECT 198.685 3014.095 198.855 3014.265 ;
        RECT 204.125 3014.095 204.295 3014.265 ;
        RECT 198.685 3013.635 198.855 3013.805 ;
        RECT 204.125 3013.635 204.295 3013.805 ;
        RECT 198.685 3013.175 198.855 3013.345 ;
        RECT 204.125 3013.175 204.295 3013.345 ;
        RECT 198.685 3012.715 198.855 3012.885 ;
        RECT 204.125 3012.715 204.295 3012.885 ;
        RECT 198.685 3012.255 198.855 3012.425 ;
        RECT 204.125 3012.255 204.295 3012.425 ;
        RECT 198.685 3011.795 198.855 3011.965 ;
        RECT 204.125 3011.795 204.295 3011.965 ;
        RECT 198.685 3011.335 198.855 3011.505 ;
        RECT 204.125 3011.335 204.295 3011.505 ;
        RECT 198.685 3010.875 198.855 3011.045 ;
        RECT 204.125 3010.875 204.295 3011.045 ;
        RECT 198.685 3010.415 198.855 3010.585 ;
        RECT 204.125 3010.415 204.295 3010.585 ;
        RECT 198.685 3009.955 198.855 3010.125 ;
        RECT 204.125 3009.955 204.295 3010.125 ;
        RECT 198.685 3009.495 198.855 3009.665 ;
        RECT 204.125 3009.495 204.295 3009.665 ;
        RECT 198.685 3009.035 198.855 3009.205 ;
        RECT 204.125 3009.035 204.295 3009.205 ;
        RECT 198.685 3008.575 198.855 3008.745 ;
        RECT 204.125 3008.575 204.295 3008.745 ;
        RECT 198.685 3008.115 198.855 3008.285 ;
        RECT 204.125 3008.115 204.295 3008.285 ;
        RECT 198.685 3007.655 198.855 3007.825 ;
        RECT 204.125 3007.655 204.295 3007.825 ;
        RECT 198.685 3007.195 198.855 3007.365 ;
        RECT 204.125 3007.195 204.295 3007.365 ;
        RECT 198.685 3006.735 198.855 3006.905 ;
        RECT 204.125 3006.735 204.295 3006.905 ;
        RECT 198.685 3006.275 198.855 3006.445 ;
        RECT 204.125 3006.275 204.295 3006.445 ;
        RECT 198.685 3005.815 198.855 3005.985 ;
        RECT 204.125 3005.815 204.295 3005.985 ;
        RECT 198.685 3005.355 198.855 3005.525 ;
        RECT 204.125 3005.355 204.295 3005.525 ;
        RECT 198.685 3004.895 198.855 3005.065 ;
        RECT 204.125 3004.895 204.295 3005.065 ;
        RECT 198.685 3004.435 198.855 3004.605 ;
        RECT 204.125 3004.435 204.295 3004.605 ;
        RECT 198.685 3003.975 198.855 3004.145 ;
        RECT 204.125 3003.975 204.295 3004.145 ;
        RECT 198.685 3003.515 198.855 3003.685 ;
        RECT 204.125 3003.515 204.295 3003.685 ;
        RECT 198.685 3003.055 198.855 3003.225 ;
        RECT 204.125 3003.055 204.295 3003.225 ;
        RECT 198.685 3002.595 198.855 3002.765 ;
        RECT 204.125 3002.595 204.295 3002.765 ;
        RECT 198.685 3002.135 198.855 3002.305 ;
        RECT 204.125 3002.135 204.295 3002.305 ;
        RECT 198.685 3001.675 198.855 3001.845 ;
        RECT 204.125 3001.675 204.295 3001.845 ;
        RECT 198.685 3001.215 198.855 3001.385 ;
        RECT 204.125 3001.215 204.295 3001.385 ;
        RECT 198.685 3000.755 198.855 3000.925 ;
        RECT 204.125 3000.755 204.295 3000.925 ;
        RECT 198.685 3000.295 198.855 3000.465 ;
        RECT 204.125 3000.295 204.295 3000.465 ;
        RECT 198.685 2999.835 198.855 3000.005 ;
        RECT 204.125 2999.835 204.295 3000.005 ;
        RECT 198.685 2999.375 198.855 2999.545 ;
        RECT 204.125 2999.375 204.295 2999.545 ;
        RECT 198.685 2998.915 198.855 2999.085 ;
        RECT 204.125 2998.915 204.295 2999.085 ;
        RECT 198.685 2998.455 198.855 2998.625 ;
        RECT 204.125 2998.455 204.295 2998.625 ;
        RECT 198.685 2997.995 198.855 2998.165 ;
        RECT 204.125 2997.995 204.295 2998.165 ;
        RECT 198.685 2997.535 198.855 2997.705 ;
        RECT 204.125 2997.535 204.295 2997.705 ;
        RECT 198.685 2997.075 198.855 2997.245 ;
        RECT 204.125 2997.075 204.295 2997.245 ;
        RECT 198.685 2996.615 198.855 2996.785 ;
        RECT 204.125 2996.615 204.295 2996.785 ;
        RECT 198.685 2996.155 198.855 2996.325 ;
        RECT 204.125 2996.155 204.295 2996.325 ;
        RECT 198.685 2995.695 198.855 2995.865 ;
        RECT 204.125 2995.695 204.295 2995.865 ;
        RECT 198.685 2995.235 198.855 2995.405 ;
        RECT 204.125 2995.235 204.295 2995.405 ;
        RECT 198.685 2994.775 198.855 2994.945 ;
        RECT 204.125 2994.775 204.295 2994.945 ;
        RECT 198.685 2994.315 198.855 2994.485 ;
        RECT 204.125 2994.315 204.295 2994.485 ;
        RECT 198.685 2993.855 198.855 2994.025 ;
        RECT 204.125 2993.855 204.295 2994.025 ;
        RECT 198.685 2993.395 198.855 2993.565 ;
        RECT 204.125 2993.395 204.295 2993.565 ;
        RECT 198.685 2992.935 198.855 2993.105 ;
        RECT 204.125 2992.935 204.295 2993.105 ;
        RECT 198.685 2992.475 198.855 2992.645 ;
        RECT 204.125 2992.475 204.295 2992.645 ;
        RECT 198.685 2992.015 198.855 2992.185 ;
        RECT 204.125 2992.015 204.295 2992.185 ;
        RECT 198.685 2991.555 198.855 2991.725 ;
        RECT 204.125 2991.555 204.295 2991.725 ;
        RECT 198.685 2991.095 198.855 2991.265 ;
        RECT 204.125 2991.095 204.295 2991.265 ;
        RECT 198.685 2990.635 198.855 2990.805 ;
        RECT 204.125 2990.635 204.295 2990.805 ;
        RECT 198.685 2990.175 198.855 2990.345 ;
        RECT 204.125 2990.175 204.295 2990.345 ;
        RECT 198.685 2989.715 198.855 2989.885 ;
        RECT 204.125 2989.715 204.295 2989.885 ;
        RECT 198.685 2989.255 198.855 2989.425 ;
        RECT 204.125 2989.255 204.295 2989.425 ;
        RECT 198.685 2988.795 198.855 2988.965 ;
        RECT 204.125 2988.795 204.295 2988.965 ;
        RECT 198.685 2988.335 198.855 2988.505 ;
        RECT 204.125 2988.335 204.295 2988.505 ;
        RECT 198.685 2987.875 198.855 2988.045 ;
        RECT 204.125 2987.875 204.295 2988.045 ;
      LAYER met1 ;
        RECT 198.530 2987.730 199.010 3024.070 ;
        RECT 203.970 2987.730 204.450 3024.070 ;
      LAYER via ;
        RECT 198.655 3020.070 198.955 3021.855 ;
        RECT 204.065 3020.070 204.365 3021.855 ;
      LAYER met2 ;
        RECT 198.570 3020.030 199.000 3021.895 ;
        RECT 203.995 3020.030 204.425 3021.895 ;
      LAYER via2 ;
        RECT 198.655 3020.070 198.955 3021.855 ;
        RECT 204.065 3020.070 204.365 3021.855 ;
      LAYER met3 ;
        RECT 196.915 3020.025 204.440 3021.890 ;
    END
    PORT
      LAYER li1 ;
        RECT 3383.500 2238.065 3383.670 2238.235 ;
        RECT 3388.940 2238.065 3389.110 2238.235 ;
        RECT 3383.500 2237.605 3383.670 2237.775 ;
        RECT 3388.940 2237.605 3389.110 2237.775 ;
        RECT 3383.500 2237.145 3383.670 2237.315 ;
        RECT 3388.940 2237.145 3389.110 2237.315 ;
        RECT 3383.500 2236.685 3383.670 2236.855 ;
        RECT 3388.940 2236.685 3389.110 2236.855 ;
        RECT 3383.500 2236.225 3383.670 2236.395 ;
        RECT 3388.940 2236.225 3389.110 2236.395 ;
        RECT 3383.500 2235.765 3383.670 2235.935 ;
        RECT 3388.940 2235.765 3389.110 2235.935 ;
        RECT 3383.500 2235.305 3383.670 2235.475 ;
        RECT 3388.940 2235.305 3389.110 2235.475 ;
        RECT 3383.500 2234.845 3383.670 2235.015 ;
        RECT 3388.940 2234.845 3389.110 2235.015 ;
        RECT 3383.500 2234.385 3383.670 2234.555 ;
        RECT 3388.940 2234.385 3389.110 2234.555 ;
        RECT 3383.500 2233.925 3383.670 2234.095 ;
        RECT 3388.940 2233.925 3389.110 2234.095 ;
        RECT 3383.500 2233.465 3383.670 2233.635 ;
        RECT 3388.940 2233.465 3389.110 2233.635 ;
        RECT 3383.500 2233.005 3383.670 2233.175 ;
        RECT 3388.940 2233.005 3389.110 2233.175 ;
        RECT 3383.500 2232.545 3383.670 2232.715 ;
        RECT 3388.940 2232.545 3389.110 2232.715 ;
        RECT 3383.500 2232.085 3383.670 2232.255 ;
        RECT 3388.940 2232.085 3389.110 2232.255 ;
        RECT 3383.500 2231.625 3383.670 2231.795 ;
        RECT 3388.940 2231.625 3389.110 2231.795 ;
        RECT 3383.500 2231.165 3383.670 2231.335 ;
        RECT 3388.940 2231.165 3389.110 2231.335 ;
        RECT 3383.500 2230.705 3383.670 2230.875 ;
        RECT 3388.940 2230.705 3389.110 2230.875 ;
        RECT 3383.500 2230.245 3383.670 2230.415 ;
        RECT 3388.940 2230.245 3389.110 2230.415 ;
        RECT 3383.500 2229.785 3383.670 2229.955 ;
        RECT 3388.940 2229.785 3389.110 2229.955 ;
        RECT 3383.500 2229.325 3383.670 2229.495 ;
        RECT 3388.940 2229.325 3389.110 2229.495 ;
        RECT 3383.500 2228.865 3383.670 2229.035 ;
        RECT 3388.940 2228.865 3389.110 2229.035 ;
        RECT 3383.500 2228.405 3383.670 2228.575 ;
        RECT 3388.940 2228.405 3389.110 2228.575 ;
        RECT 3383.500 2227.945 3383.670 2228.115 ;
        RECT 3388.940 2227.945 3389.110 2228.115 ;
        RECT 3383.500 2227.485 3383.670 2227.655 ;
        RECT 3388.940 2227.485 3389.110 2227.655 ;
        RECT 3383.500 2227.025 3383.670 2227.195 ;
        RECT 3388.940 2227.025 3389.110 2227.195 ;
        RECT 3383.500 2226.565 3383.670 2226.735 ;
        RECT 3388.940 2226.565 3389.110 2226.735 ;
        RECT 3383.500 2226.105 3383.670 2226.275 ;
        RECT 3388.940 2226.105 3389.110 2226.275 ;
        RECT 3383.500 2225.645 3383.670 2225.815 ;
        RECT 3388.940 2225.645 3389.110 2225.815 ;
        RECT 3383.500 2225.185 3383.670 2225.355 ;
        RECT 3388.940 2225.185 3389.110 2225.355 ;
        RECT 3383.500 2224.725 3383.670 2224.895 ;
        RECT 3388.940 2224.725 3389.110 2224.895 ;
        RECT 3383.500 2224.265 3383.670 2224.435 ;
        RECT 3388.940 2224.265 3389.110 2224.435 ;
        RECT 3383.500 2223.805 3383.670 2223.975 ;
        RECT 3388.940 2223.805 3389.110 2223.975 ;
        RECT 3383.500 2223.345 3383.670 2223.515 ;
        RECT 3388.940 2223.345 3389.110 2223.515 ;
        RECT 3383.500 2222.885 3383.670 2223.055 ;
        RECT 3388.940 2222.885 3389.110 2223.055 ;
        RECT 3383.500 2222.425 3383.670 2222.595 ;
        RECT 3388.940 2222.425 3389.110 2222.595 ;
        RECT 3383.500 2221.965 3383.670 2222.135 ;
        RECT 3388.940 2221.965 3389.110 2222.135 ;
        RECT 3383.500 2221.505 3383.670 2221.675 ;
        RECT 3388.940 2221.505 3389.110 2221.675 ;
        RECT 3383.500 2221.045 3383.670 2221.215 ;
        RECT 3388.940 2221.045 3389.110 2221.215 ;
        RECT 3383.500 2220.585 3383.670 2220.755 ;
        RECT 3388.940 2220.585 3389.110 2220.755 ;
        RECT 3383.500 2220.125 3383.670 2220.295 ;
        RECT 3388.940 2220.125 3389.110 2220.295 ;
        RECT 3383.500 2219.665 3383.670 2219.835 ;
        RECT 3388.940 2219.665 3389.110 2219.835 ;
        RECT 3383.500 2219.205 3383.670 2219.375 ;
        RECT 3388.940 2219.205 3389.110 2219.375 ;
        RECT 3383.500 2218.745 3383.670 2218.915 ;
        RECT 3388.940 2218.745 3389.110 2218.915 ;
        RECT 3383.500 2218.285 3383.670 2218.455 ;
        RECT 3388.940 2218.285 3389.110 2218.455 ;
        RECT 3383.500 2217.825 3383.670 2217.995 ;
        RECT 3388.940 2217.825 3389.110 2217.995 ;
        RECT 3383.500 2217.365 3383.670 2217.535 ;
        RECT 3388.940 2217.365 3389.110 2217.535 ;
        RECT 3383.500 2216.905 3383.670 2217.075 ;
        RECT 3388.940 2216.905 3389.110 2217.075 ;
        RECT 3383.500 2216.445 3383.670 2216.615 ;
        RECT 3388.940 2216.445 3389.110 2216.615 ;
        RECT 3383.500 2215.985 3383.670 2216.155 ;
        RECT 3388.940 2215.985 3389.110 2216.155 ;
        RECT 3383.500 2215.525 3383.670 2215.695 ;
        RECT 3388.940 2215.525 3389.110 2215.695 ;
        RECT 3383.500 2215.065 3383.670 2215.235 ;
        RECT 3388.940 2215.065 3389.110 2215.235 ;
        RECT 3383.500 2214.605 3383.670 2214.775 ;
        RECT 3388.940 2214.605 3389.110 2214.775 ;
        RECT 3383.500 2214.145 3383.670 2214.315 ;
        RECT 3388.940 2214.145 3389.110 2214.315 ;
        RECT 3383.500 2213.685 3383.670 2213.855 ;
        RECT 3388.940 2213.685 3389.110 2213.855 ;
        RECT 3383.500 2213.225 3383.670 2213.395 ;
        RECT 3388.940 2213.225 3389.110 2213.395 ;
        RECT 3383.500 2212.765 3383.670 2212.935 ;
        RECT 3388.940 2212.765 3389.110 2212.935 ;
        RECT 3383.500 2212.305 3383.670 2212.475 ;
        RECT 3388.940 2212.305 3389.110 2212.475 ;
        RECT 3383.500 2211.845 3383.670 2212.015 ;
        RECT 3388.940 2211.845 3389.110 2212.015 ;
        RECT 3383.500 2211.385 3383.670 2211.555 ;
        RECT 3388.940 2211.385 3389.110 2211.555 ;
        RECT 3383.500 2210.925 3383.670 2211.095 ;
        RECT 3388.940 2210.925 3389.110 2211.095 ;
        RECT 3383.500 2210.465 3383.670 2210.635 ;
        RECT 3388.940 2210.465 3389.110 2210.635 ;
        RECT 3383.500 2210.005 3383.670 2210.175 ;
        RECT 3388.940 2210.005 3389.110 2210.175 ;
        RECT 3383.500 2209.545 3383.670 2209.715 ;
        RECT 3388.940 2209.545 3389.110 2209.715 ;
        RECT 3383.500 2209.085 3383.670 2209.255 ;
        RECT 3388.940 2209.085 3389.110 2209.255 ;
        RECT 3383.500 2208.625 3383.670 2208.795 ;
        RECT 3388.940 2208.625 3389.110 2208.795 ;
        RECT 3383.500 2208.165 3383.670 2208.335 ;
        RECT 3388.940 2208.165 3389.110 2208.335 ;
        RECT 3383.500 2207.705 3383.670 2207.875 ;
        RECT 3388.940 2207.705 3389.110 2207.875 ;
        RECT 3383.500 2207.245 3383.670 2207.415 ;
        RECT 3388.940 2207.245 3389.110 2207.415 ;
        RECT 3383.500 2206.785 3383.670 2206.955 ;
        RECT 3388.940 2206.785 3389.110 2206.955 ;
        RECT 3383.500 2206.325 3383.670 2206.495 ;
        RECT 3388.940 2206.325 3389.110 2206.495 ;
        RECT 3383.500 2205.865 3383.670 2206.035 ;
        RECT 3388.940 2205.865 3389.110 2206.035 ;
        RECT 3383.500 2205.405 3383.670 2205.575 ;
        RECT 3388.940 2205.405 3389.110 2205.575 ;
        RECT 3383.500 2204.945 3383.670 2205.115 ;
        RECT 3388.940 2204.945 3389.110 2205.115 ;
        RECT 3383.500 2204.485 3383.670 2204.655 ;
        RECT 3388.940 2204.485 3389.110 2204.655 ;
        RECT 3383.500 2204.025 3383.670 2204.195 ;
        RECT 3388.940 2204.025 3389.110 2204.195 ;
        RECT 3383.500 2203.565 3383.670 2203.735 ;
        RECT 3388.940 2203.565 3389.110 2203.735 ;
        RECT 3383.500 2203.105 3383.670 2203.275 ;
        RECT 3388.940 2203.105 3389.110 2203.275 ;
        RECT 3383.500 2202.645 3383.670 2202.815 ;
        RECT 3388.940 2202.645 3389.110 2202.815 ;
        RECT 3383.500 2202.185 3383.670 2202.355 ;
        RECT 3388.940 2202.185 3389.110 2202.355 ;
        RECT 3383.500 2201.725 3383.670 2201.895 ;
        RECT 3388.940 2201.725 3389.110 2201.895 ;
        RECT 3383.500 2201.265 3383.670 2201.435 ;
        RECT 3388.940 2201.265 3389.110 2201.435 ;
        RECT 3383.500 2200.805 3383.670 2200.975 ;
        RECT 3388.940 2200.805 3389.110 2200.975 ;
        RECT 3383.500 2200.345 3383.670 2200.515 ;
        RECT 3388.940 2200.345 3389.110 2200.515 ;
        RECT 3383.500 2199.885 3383.670 2200.055 ;
        RECT 3388.940 2199.885 3389.110 2200.055 ;
        RECT 3383.500 2199.425 3383.670 2199.595 ;
        RECT 3388.940 2199.425 3389.110 2199.595 ;
        RECT 3383.500 2198.965 3383.670 2199.135 ;
        RECT 3388.940 2198.965 3389.110 2199.135 ;
        RECT 3383.500 2198.505 3383.670 2198.675 ;
        RECT 3388.940 2198.505 3389.110 2198.675 ;
        RECT 3383.500 2198.045 3383.670 2198.215 ;
        RECT 3388.940 2198.045 3389.110 2198.215 ;
        RECT 3383.500 2197.585 3383.670 2197.755 ;
        RECT 3388.940 2197.585 3389.110 2197.755 ;
        RECT 3383.500 2197.125 3383.670 2197.295 ;
        RECT 3388.940 2197.125 3389.110 2197.295 ;
        RECT 3383.500 2196.665 3383.670 2196.835 ;
        RECT 3388.940 2196.665 3389.110 2196.835 ;
        RECT 3383.500 2196.205 3383.670 2196.375 ;
        RECT 3388.940 2196.205 3389.110 2196.375 ;
      LAYER met1 ;
        RECT 3383.345 2196.060 3383.825 2238.380 ;
        RECT 3388.785 2196.060 3389.265 2238.380 ;
      LAYER via ;
        RECT 3383.425 2228.515 3383.725 2230.300 ;
        RECT 3388.835 2228.515 3389.135 2230.300 ;
      LAYER met2 ;
        RECT 3383.365 2228.475 3383.795 2230.340 ;
        RECT 3388.790 2228.475 3389.220 2230.340 ;
      LAYER via2 ;
        RECT 3383.425 2228.515 3383.725 2230.300 ;
        RECT 3388.835 2228.515 3389.135 2230.300 ;
      LAYER met3 ;
        RECT 3383.350 2228.480 3390.875 2230.345 ;
    END
    PORT
      LAYER li1 ;
        RECT 3383.500 3542.185 3383.670 3542.355 ;
        RECT 3388.940 3542.185 3389.110 3542.355 ;
        RECT 3383.500 3541.725 3383.670 3541.895 ;
        RECT 3388.940 3541.725 3389.110 3541.895 ;
        RECT 3383.500 3541.265 3383.670 3541.435 ;
        RECT 3388.940 3541.265 3389.110 3541.435 ;
        RECT 3383.500 3540.805 3383.670 3540.975 ;
        RECT 3388.940 3540.805 3389.110 3540.975 ;
        RECT 3383.500 3540.345 3383.670 3540.515 ;
        RECT 3388.940 3540.345 3389.110 3540.515 ;
        RECT 3383.500 3539.885 3383.670 3540.055 ;
        RECT 3388.940 3539.885 3389.110 3540.055 ;
        RECT 3383.500 3539.425 3383.670 3539.595 ;
        RECT 3388.940 3539.425 3389.110 3539.595 ;
        RECT 3383.500 3538.965 3383.670 3539.135 ;
        RECT 3388.940 3538.965 3389.110 3539.135 ;
        RECT 3383.500 3538.505 3383.670 3538.675 ;
        RECT 3388.940 3538.505 3389.110 3538.675 ;
        RECT 3383.500 3538.045 3383.670 3538.215 ;
        RECT 3388.940 3538.045 3389.110 3538.215 ;
        RECT 3383.500 3537.585 3383.670 3537.755 ;
        RECT 3388.940 3537.585 3389.110 3537.755 ;
        RECT 3383.500 3537.125 3383.670 3537.295 ;
        RECT 3388.940 3537.125 3389.110 3537.295 ;
        RECT 3383.500 3536.665 3383.670 3536.835 ;
        RECT 3388.940 3536.665 3389.110 3536.835 ;
        RECT 3383.500 3536.205 3383.670 3536.375 ;
        RECT 3388.940 3536.205 3389.110 3536.375 ;
      LAYER met1 ;
        RECT 3383.345 3536.060 3383.825 3542.500 ;
        RECT 3388.785 3536.060 3389.265 3542.500 ;
      LAYER via ;
        RECT 3383.465 3538.540 3383.765 3540.325 ;
        RECT 3388.875 3538.540 3389.175 3540.325 ;
      LAYER met2 ;
        RECT 3383.405 3538.500 3383.835 3540.365 ;
        RECT 3388.830 3538.500 3389.260 3540.365 ;
      LAYER via2 ;
        RECT 3383.465 3538.540 3383.765 3540.325 ;
        RECT 3388.875 3538.540 3389.175 3540.325 ;
      LAYER met3 ;
        RECT 3383.390 3538.505 3390.915 3540.370 ;
    END
  END vssd
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 669.145 1114.320 669.315 1114.490 ;
        RECT 669.605 1114.320 669.775 1114.490 ;
        RECT 670.065 1114.320 670.235 1114.490 ;
        RECT 670.525 1114.320 670.695 1114.490 ;
        RECT 670.985 1114.320 671.155 1114.490 ;
        RECT 671.445 1114.320 671.615 1114.490 ;
        RECT 671.905 1114.320 672.075 1114.490 ;
        RECT 672.365 1114.320 672.535 1114.490 ;
        RECT 672.825 1114.320 672.995 1114.490 ;
        RECT 673.285 1114.320 673.455 1114.490 ;
        RECT 673.745 1114.320 673.915 1114.490 ;
        RECT 674.205 1114.320 674.375 1114.490 ;
        RECT 674.665 1114.320 674.835 1114.490 ;
        RECT 675.125 1114.320 675.295 1114.490 ;
        RECT 675.585 1114.320 675.755 1114.490 ;
        RECT 676.045 1114.320 676.215 1114.490 ;
        RECT 676.505 1114.320 676.675 1114.490 ;
        RECT 676.965 1114.320 677.135 1114.490 ;
        RECT 677.425 1114.320 677.595 1114.490 ;
        RECT 677.885 1114.320 678.055 1114.490 ;
        RECT 678.345 1114.320 678.515 1114.490 ;
        RECT 678.805 1114.320 678.975 1114.490 ;
        RECT 679.265 1114.320 679.435 1114.490 ;
        RECT 679.725 1114.320 679.895 1114.490 ;
        RECT 680.185 1114.320 680.355 1114.490 ;
        RECT 680.645 1114.320 680.815 1114.490 ;
        RECT 681.105 1114.320 681.275 1114.490 ;
        RECT 681.565 1114.320 681.735 1114.490 ;
        RECT 682.025 1114.320 682.195 1114.490 ;
        RECT 682.485 1114.320 682.655 1114.490 ;
        RECT 682.945 1114.320 683.115 1114.490 ;
        RECT 683.405 1114.320 683.575 1114.490 ;
        RECT 683.865 1114.320 684.035 1114.490 ;
        RECT 684.325 1114.320 684.495 1114.490 ;
        RECT 684.785 1114.320 684.955 1114.490 ;
        RECT 685.245 1114.320 685.415 1114.490 ;
        RECT 685.705 1114.320 685.875 1114.490 ;
        RECT 686.165 1114.320 686.335 1114.490 ;
        RECT 686.625 1114.320 686.795 1114.490 ;
        RECT 687.085 1114.320 687.255 1114.490 ;
        RECT 687.545 1114.320 687.715 1114.490 ;
        RECT 688.005 1114.320 688.175 1114.490 ;
        RECT 688.465 1114.320 688.635 1114.490 ;
        RECT 688.925 1114.320 689.095 1114.490 ;
        RECT 689.385 1114.320 689.555 1114.490 ;
        RECT 689.845 1114.320 690.015 1114.490 ;
        RECT 690.305 1114.320 690.475 1114.490 ;
        RECT 690.765 1114.320 690.935 1114.490 ;
        RECT 691.225 1114.320 691.395 1114.490 ;
        RECT 691.685 1114.320 691.855 1114.490 ;
        RECT 692.145 1114.320 692.315 1114.490 ;
        RECT 692.605 1114.320 692.775 1114.490 ;
        RECT 693.065 1114.320 693.235 1114.490 ;
        RECT 693.525 1114.320 693.695 1114.490 ;
        RECT 693.985 1114.320 694.155 1114.490 ;
        RECT 694.445 1114.320 694.615 1114.490 ;
        RECT 694.905 1114.320 695.075 1114.490 ;
        RECT 695.365 1114.320 695.535 1114.490 ;
        RECT 695.825 1114.320 695.995 1114.490 ;
        RECT 696.285 1114.320 696.455 1114.490 ;
        RECT 696.745 1114.320 696.915 1114.490 ;
        RECT 697.205 1114.320 697.375 1114.490 ;
        RECT 697.665 1114.320 697.835 1114.490 ;
        RECT 698.125 1114.320 698.295 1114.490 ;
        RECT 698.585 1114.320 698.755 1114.490 ;
        RECT 699.045 1114.320 699.215 1114.490 ;
        RECT 699.505 1114.320 699.675 1114.490 ;
        RECT 699.965 1114.320 700.135 1114.490 ;
        RECT 700.425 1114.320 700.595 1114.490 ;
        RECT 700.885 1114.320 701.055 1114.490 ;
        RECT 701.345 1114.320 701.515 1114.490 ;
        RECT 701.805 1114.320 701.975 1114.490 ;
        RECT 702.265 1114.320 702.435 1114.490 ;
        RECT 702.725 1114.320 702.895 1114.490 ;
        RECT 703.185 1114.320 703.355 1114.490 ;
        RECT 703.645 1114.320 703.815 1114.490 ;
        RECT 704.105 1114.320 704.275 1114.490 ;
        RECT 704.565 1114.320 704.735 1114.490 ;
        RECT 705.025 1114.320 705.195 1114.490 ;
        RECT 705.485 1114.320 705.655 1114.490 ;
        RECT 705.945 1114.320 706.115 1114.490 ;
        RECT 706.405 1114.320 706.575 1114.490 ;
        RECT 706.865 1114.320 707.035 1114.490 ;
        RECT 707.325 1114.320 707.495 1114.490 ;
        RECT 707.785 1114.320 707.955 1114.490 ;
        RECT 708.245 1114.320 708.415 1114.490 ;
        RECT 708.705 1114.320 708.875 1114.490 ;
        RECT 709.165 1114.320 709.335 1114.490 ;
        RECT 709.625 1114.320 709.795 1114.490 ;
        RECT 710.085 1114.320 710.255 1114.490 ;
        RECT 710.545 1114.320 710.715 1114.490 ;
        RECT 711.005 1114.320 711.175 1114.490 ;
        RECT 711.465 1114.320 711.635 1114.490 ;
        RECT 711.925 1114.320 712.095 1114.490 ;
        RECT 712.385 1114.320 712.555 1114.490 ;
        RECT 712.845 1114.320 713.015 1114.490 ;
        RECT 713.305 1114.320 713.475 1114.490 ;
        RECT 713.765 1114.320 713.935 1114.490 ;
        RECT 714.225 1114.320 714.395 1114.490 ;
        RECT 714.685 1114.320 714.855 1114.490 ;
        RECT 715.145 1114.320 715.315 1114.490 ;
        RECT 715.605 1114.320 715.775 1114.490 ;
        RECT 716.065 1114.320 716.235 1114.490 ;
        RECT 716.525 1114.320 716.695 1114.490 ;
        RECT 716.985 1114.320 717.155 1114.490 ;
        RECT 717.445 1114.320 717.615 1114.490 ;
        RECT 717.905 1114.320 718.075 1114.490 ;
        RECT 718.365 1114.320 718.535 1114.490 ;
        RECT 718.825 1114.320 718.995 1114.490 ;
        RECT 719.285 1114.320 719.455 1114.490 ;
        RECT 719.745 1114.320 719.915 1114.490 ;
        RECT 720.205 1114.320 720.375 1114.490 ;
        RECT 720.665 1114.320 720.835 1114.490 ;
        RECT 721.125 1114.320 721.295 1114.490 ;
        RECT 721.585 1114.320 721.755 1114.490 ;
        RECT 722.045 1114.320 722.215 1114.490 ;
        RECT 722.505 1114.320 722.675 1114.490 ;
        RECT 722.965 1114.320 723.135 1114.490 ;
        RECT 723.425 1114.320 723.595 1114.490 ;
        RECT 723.885 1114.320 724.055 1114.490 ;
        RECT 724.345 1114.320 724.515 1114.490 ;
        RECT 724.805 1114.320 724.975 1114.490 ;
        RECT 725.265 1114.320 725.435 1114.490 ;
        RECT 725.725 1114.320 725.895 1114.490 ;
        RECT 726.185 1114.320 726.355 1114.490 ;
        RECT 726.645 1114.320 726.815 1114.490 ;
        RECT 727.105 1114.320 727.275 1114.490 ;
        RECT 727.565 1114.320 727.735 1114.490 ;
        RECT 728.025 1114.320 728.195 1114.490 ;
        RECT 728.485 1114.320 728.655 1114.490 ;
        RECT 728.945 1114.320 729.115 1114.490 ;
        RECT 729.405 1114.320 729.575 1114.490 ;
        RECT 729.865 1114.320 730.035 1114.490 ;
        RECT 730.325 1114.320 730.495 1114.490 ;
        RECT 730.785 1114.320 730.955 1114.490 ;
        RECT 731.245 1114.320 731.415 1114.490 ;
        RECT 731.705 1114.320 731.875 1114.490 ;
        RECT 732.165 1114.320 732.335 1114.490 ;
        RECT 732.625 1114.320 732.795 1114.490 ;
        RECT 733.085 1114.320 733.255 1114.490 ;
        RECT 733.545 1114.320 733.715 1114.490 ;
        RECT 734.005 1114.320 734.175 1114.490 ;
        RECT 734.465 1114.320 734.635 1114.490 ;
        RECT 734.925 1114.320 735.095 1114.490 ;
        RECT 735.385 1114.320 735.555 1114.490 ;
        RECT 735.845 1114.320 736.015 1114.490 ;
        RECT 736.305 1114.320 736.475 1114.490 ;
        RECT 736.765 1114.320 736.935 1114.490 ;
        RECT 737.225 1114.320 737.395 1114.490 ;
        RECT 737.685 1114.320 737.855 1114.490 ;
        RECT 738.145 1114.320 738.315 1114.490 ;
        RECT 738.605 1114.320 738.775 1114.490 ;
        RECT 739.065 1114.320 739.235 1114.490 ;
        RECT 739.525 1114.320 739.695 1114.490 ;
        RECT 739.985 1114.320 740.155 1114.490 ;
        RECT 740.445 1114.320 740.615 1114.490 ;
        RECT 740.905 1114.320 741.075 1114.490 ;
        RECT 741.365 1114.320 741.535 1114.490 ;
        RECT 741.825 1114.320 741.995 1114.490 ;
        RECT 742.285 1114.320 742.455 1114.490 ;
        RECT 742.745 1114.320 742.915 1114.490 ;
        RECT 743.205 1114.320 743.375 1114.490 ;
        RECT 743.665 1114.320 743.835 1114.490 ;
        RECT 744.125 1114.320 744.295 1114.490 ;
        RECT 744.585 1114.320 744.755 1114.490 ;
        RECT 745.045 1114.320 745.215 1114.490 ;
        RECT 745.505 1114.320 745.675 1114.490 ;
        RECT 745.965 1114.320 746.135 1114.490 ;
        RECT 746.425 1114.320 746.595 1114.490 ;
        RECT 746.885 1114.320 747.055 1114.490 ;
        RECT 747.345 1114.320 747.515 1114.490 ;
        RECT 747.805 1114.320 747.975 1114.490 ;
        RECT 748.265 1114.320 748.435 1114.490 ;
        RECT 748.725 1114.320 748.895 1114.490 ;
        RECT 749.185 1114.320 749.355 1114.490 ;
        RECT 749.645 1114.320 749.815 1114.490 ;
        RECT 750.105 1114.320 750.275 1114.490 ;
        RECT 750.565 1114.320 750.735 1114.490 ;
        RECT 751.025 1114.320 751.195 1114.490 ;
        RECT 751.485 1114.320 751.655 1114.490 ;
        RECT 751.945 1114.320 752.115 1114.490 ;
        RECT 752.405 1114.320 752.575 1114.490 ;
        RECT 752.865 1114.320 753.035 1114.490 ;
        RECT 753.325 1114.320 753.495 1114.490 ;
        RECT 753.785 1114.320 753.955 1114.490 ;
        RECT 754.245 1114.320 754.415 1114.490 ;
        RECT 754.705 1114.320 754.875 1114.490 ;
        RECT 755.165 1114.320 755.335 1114.490 ;
        RECT 755.625 1114.320 755.795 1114.490 ;
        RECT 756.085 1114.320 756.255 1114.490 ;
        RECT 756.545 1114.320 756.715 1114.490 ;
        RECT 757.005 1114.320 757.175 1114.490 ;
        RECT 757.465 1114.320 757.635 1114.490 ;
        RECT 757.925 1114.320 758.095 1114.490 ;
        RECT 758.385 1114.320 758.555 1114.490 ;
        RECT 758.845 1114.320 759.015 1114.490 ;
        RECT 759.305 1114.320 759.475 1114.490 ;
        RECT 759.765 1114.320 759.935 1114.490 ;
        RECT 760.225 1114.320 760.395 1114.490 ;
        RECT 760.685 1114.320 760.855 1114.490 ;
        RECT 761.145 1114.320 761.315 1114.490 ;
        RECT 761.605 1114.320 761.775 1114.490 ;
        RECT 762.065 1114.320 762.235 1114.490 ;
        RECT 762.525 1114.320 762.695 1114.490 ;
        RECT 762.985 1114.320 763.155 1114.490 ;
        RECT 763.445 1114.320 763.615 1114.490 ;
        RECT 763.905 1114.320 764.075 1114.490 ;
        RECT 764.365 1114.320 764.535 1114.490 ;
        RECT 764.825 1114.320 764.995 1114.490 ;
        RECT 765.285 1114.320 765.455 1114.490 ;
        RECT 765.745 1114.320 765.915 1114.490 ;
        RECT 766.205 1114.320 766.375 1114.490 ;
        RECT 766.665 1114.320 766.835 1114.490 ;
        RECT 767.125 1114.320 767.295 1114.490 ;
        RECT 767.585 1114.320 767.755 1114.490 ;
        RECT 768.045 1114.320 768.215 1114.490 ;
        RECT 768.505 1114.320 768.675 1114.490 ;
        RECT 768.965 1114.320 769.135 1114.490 ;
        RECT 769.425 1114.320 769.595 1114.490 ;
        RECT 769.885 1114.320 770.055 1114.490 ;
        RECT 770.345 1114.320 770.515 1114.490 ;
        RECT 770.805 1114.320 770.975 1114.490 ;
      LAYER met1 ;
        RECT 669.000 1114.165 771.120 1114.645 ;
      LAYER via ;
        RECT 730.995 1114.280 732.780 1114.580 ;
      LAYER met2 ;
        RECT 730.955 1114.220 732.820 1114.650 ;
      LAYER via2 ;
        RECT 730.995 1114.280 732.780 1114.580 ;
      LAYER met3 ;
        RECT 730.965 1109.835 732.815 1114.650 ;
    END
    PORT
      LAYER li1 ;
        RECT 1969.145 1114.320 1969.315 1114.490 ;
        RECT 1969.605 1114.320 1969.775 1114.490 ;
        RECT 1970.065 1114.320 1970.235 1114.490 ;
        RECT 1970.525 1114.320 1970.695 1114.490 ;
        RECT 1970.985 1114.320 1971.155 1114.490 ;
        RECT 1971.445 1114.320 1971.615 1114.490 ;
        RECT 1971.905 1114.320 1972.075 1114.490 ;
        RECT 1972.365 1114.320 1972.535 1114.490 ;
        RECT 1972.825 1114.320 1972.995 1114.490 ;
        RECT 1973.285 1114.320 1973.455 1114.490 ;
        RECT 1973.745 1114.320 1973.915 1114.490 ;
        RECT 1974.205 1114.320 1974.375 1114.490 ;
        RECT 1974.665 1114.320 1974.835 1114.490 ;
        RECT 1975.125 1114.320 1975.295 1114.490 ;
        RECT 1975.585 1114.320 1975.755 1114.490 ;
        RECT 1976.045 1114.320 1976.215 1114.490 ;
        RECT 1976.505 1114.320 1976.675 1114.490 ;
        RECT 1976.965 1114.320 1977.135 1114.490 ;
        RECT 1977.425 1114.320 1977.595 1114.490 ;
        RECT 1977.885 1114.320 1978.055 1114.490 ;
        RECT 1978.345 1114.320 1978.515 1114.490 ;
        RECT 1978.805 1114.320 1978.975 1114.490 ;
        RECT 1979.265 1114.320 1979.435 1114.490 ;
        RECT 1979.725 1114.320 1979.895 1114.490 ;
        RECT 1980.185 1114.320 1980.355 1114.490 ;
        RECT 1980.645 1114.320 1980.815 1114.490 ;
        RECT 1981.105 1114.320 1981.275 1114.490 ;
        RECT 1981.565 1114.320 1981.735 1114.490 ;
        RECT 1982.025 1114.320 1982.195 1114.490 ;
        RECT 1982.485 1114.320 1982.655 1114.490 ;
        RECT 1982.945 1114.320 1983.115 1114.490 ;
        RECT 1983.405 1114.320 1983.575 1114.490 ;
        RECT 1983.865 1114.320 1984.035 1114.490 ;
        RECT 1984.325 1114.320 1984.495 1114.490 ;
        RECT 1984.785 1114.320 1984.955 1114.490 ;
        RECT 1985.245 1114.320 1985.415 1114.490 ;
        RECT 1985.705 1114.320 1985.875 1114.490 ;
        RECT 1986.165 1114.320 1986.335 1114.490 ;
        RECT 1986.625 1114.320 1986.795 1114.490 ;
        RECT 1987.085 1114.320 1987.255 1114.490 ;
        RECT 1987.545 1114.320 1987.715 1114.490 ;
        RECT 1988.005 1114.320 1988.175 1114.490 ;
        RECT 1988.465 1114.320 1988.635 1114.490 ;
        RECT 1988.925 1114.320 1989.095 1114.490 ;
        RECT 1989.385 1114.320 1989.555 1114.490 ;
        RECT 1989.845 1114.320 1990.015 1114.490 ;
        RECT 1990.305 1114.320 1990.475 1114.490 ;
        RECT 1990.765 1114.320 1990.935 1114.490 ;
        RECT 1991.225 1114.320 1991.395 1114.490 ;
        RECT 1991.685 1114.320 1991.855 1114.490 ;
        RECT 1992.145 1114.320 1992.315 1114.490 ;
        RECT 1992.605 1114.320 1992.775 1114.490 ;
        RECT 1993.065 1114.320 1993.235 1114.490 ;
        RECT 1993.525 1114.320 1993.695 1114.490 ;
        RECT 1993.985 1114.320 1994.155 1114.490 ;
        RECT 1994.445 1114.320 1994.615 1114.490 ;
        RECT 1994.905 1114.320 1995.075 1114.490 ;
        RECT 1995.365 1114.320 1995.535 1114.490 ;
        RECT 1995.825 1114.320 1995.995 1114.490 ;
        RECT 1996.285 1114.320 1996.455 1114.490 ;
        RECT 1996.745 1114.320 1996.915 1114.490 ;
        RECT 1997.205 1114.320 1997.375 1114.490 ;
        RECT 1997.665 1114.320 1997.835 1114.490 ;
        RECT 1998.125 1114.320 1998.295 1114.490 ;
        RECT 1998.585 1114.320 1998.755 1114.490 ;
        RECT 1999.045 1114.320 1999.215 1114.490 ;
        RECT 1999.505 1114.320 1999.675 1114.490 ;
        RECT 1999.965 1114.320 2000.135 1114.490 ;
        RECT 2000.425 1114.320 2000.595 1114.490 ;
        RECT 2000.885 1114.320 2001.055 1114.490 ;
        RECT 2001.345 1114.320 2001.515 1114.490 ;
        RECT 2001.805 1114.320 2001.975 1114.490 ;
        RECT 2002.265 1114.320 2002.435 1114.490 ;
        RECT 2002.725 1114.320 2002.895 1114.490 ;
        RECT 2003.185 1114.320 2003.355 1114.490 ;
        RECT 2003.645 1114.320 2003.815 1114.490 ;
        RECT 2004.105 1114.320 2004.275 1114.490 ;
        RECT 2004.565 1114.320 2004.735 1114.490 ;
        RECT 2005.025 1114.320 2005.195 1114.490 ;
        RECT 2005.485 1114.320 2005.655 1114.490 ;
        RECT 2005.945 1114.320 2006.115 1114.490 ;
        RECT 2006.405 1114.320 2006.575 1114.490 ;
        RECT 2006.865 1114.320 2007.035 1114.490 ;
        RECT 2007.325 1114.320 2007.495 1114.490 ;
        RECT 2007.785 1114.320 2007.955 1114.490 ;
        RECT 2008.245 1114.320 2008.415 1114.490 ;
        RECT 2008.705 1114.320 2008.875 1114.490 ;
        RECT 2009.165 1114.320 2009.335 1114.490 ;
        RECT 2009.625 1114.320 2009.795 1114.490 ;
        RECT 2010.085 1114.320 2010.255 1114.490 ;
        RECT 2010.545 1114.320 2010.715 1114.490 ;
        RECT 2011.005 1114.320 2011.175 1114.490 ;
        RECT 2011.465 1114.320 2011.635 1114.490 ;
        RECT 2011.925 1114.320 2012.095 1114.490 ;
        RECT 2012.385 1114.320 2012.555 1114.490 ;
        RECT 2012.845 1114.320 2013.015 1114.490 ;
        RECT 2013.305 1114.320 2013.475 1114.490 ;
        RECT 2013.765 1114.320 2013.935 1114.490 ;
        RECT 2014.225 1114.320 2014.395 1114.490 ;
        RECT 2014.685 1114.320 2014.855 1114.490 ;
        RECT 2015.145 1114.320 2015.315 1114.490 ;
        RECT 2015.605 1114.320 2015.775 1114.490 ;
        RECT 2016.065 1114.320 2016.235 1114.490 ;
        RECT 2016.525 1114.320 2016.695 1114.490 ;
        RECT 2016.985 1114.320 2017.155 1114.490 ;
        RECT 2017.445 1114.320 2017.615 1114.490 ;
        RECT 2017.905 1114.320 2018.075 1114.490 ;
        RECT 2018.365 1114.320 2018.535 1114.490 ;
        RECT 2018.825 1114.320 2018.995 1114.490 ;
        RECT 2019.285 1114.320 2019.455 1114.490 ;
        RECT 2019.745 1114.320 2019.915 1114.490 ;
        RECT 2020.205 1114.320 2020.375 1114.490 ;
        RECT 2020.665 1114.320 2020.835 1114.490 ;
        RECT 2021.125 1114.320 2021.295 1114.490 ;
        RECT 2021.585 1114.320 2021.755 1114.490 ;
        RECT 2022.045 1114.320 2022.215 1114.490 ;
        RECT 2022.505 1114.320 2022.675 1114.490 ;
        RECT 2022.965 1114.320 2023.135 1114.490 ;
        RECT 2023.425 1114.320 2023.595 1114.490 ;
        RECT 2023.885 1114.320 2024.055 1114.490 ;
        RECT 2024.345 1114.320 2024.515 1114.490 ;
        RECT 2024.805 1114.320 2024.975 1114.490 ;
        RECT 2025.265 1114.320 2025.435 1114.490 ;
        RECT 2025.725 1114.320 2025.895 1114.490 ;
        RECT 2026.185 1114.320 2026.355 1114.490 ;
        RECT 2026.645 1114.320 2026.815 1114.490 ;
        RECT 2027.105 1114.320 2027.275 1114.490 ;
        RECT 2027.565 1114.320 2027.735 1114.490 ;
        RECT 2028.025 1114.320 2028.195 1114.490 ;
        RECT 2028.485 1114.320 2028.655 1114.490 ;
        RECT 2028.945 1114.320 2029.115 1114.490 ;
        RECT 2029.405 1114.320 2029.575 1114.490 ;
        RECT 2029.865 1114.320 2030.035 1114.490 ;
        RECT 2030.325 1114.320 2030.495 1114.490 ;
        RECT 2030.785 1114.320 2030.955 1114.490 ;
        RECT 2031.245 1114.320 2031.415 1114.490 ;
        RECT 2031.705 1114.320 2031.875 1114.490 ;
        RECT 2032.165 1114.320 2032.335 1114.490 ;
        RECT 2032.625 1114.320 2032.795 1114.490 ;
        RECT 2033.085 1114.320 2033.255 1114.490 ;
        RECT 2033.545 1114.320 2033.715 1114.490 ;
        RECT 2034.005 1114.320 2034.175 1114.490 ;
        RECT 2034.465 1114.320 2034.635 1114.490 ;
        RECT 2034.925 1114.320 2035.095 1114.490 ;
        RECT 2035.385 1114.320 2035.555 1114.490 ;
        RECT 2035.845 1114.320 2036.015 1114.490 ;
        RECT 2036.305 1114.320 2036.475 1114.490 ;
        RECT 2036.765 1114.320 2036.935 1114.490 ;
        RECT 2037.225 1114.320 2037.395 1114.490 ;
        RECT 2037.685 1114.320 2037.855 1114.490 ;
        RECT 2038.145 1114.320 2038.315 1114.490 ;
        RECT 2038.605 1114.320 2038.775 1114.490 ;
        RECT 2039.065 1114.320 2039.235 1114.490 ;
        RECT 2039.525 1114.320 2039.695 1114.490 ;
        RECT 2039.985 1114.320 2040.155 1114.490 ;
        RECT 2040.445 1114.320 2040.615 1114.490 ;
        RECT 2040.905 1114.320 2041.075 1114.490 ;
        RECT 2041.365 1114.320 2041.535 1114.490 ;
        RECT 2041.825 1114.320 2041.995 1114.490 ;
        RECT 2042.285 1114.320 2042.455 1114.490 ;
        RECT 2042.745 1114.320 2042.915 1114.490 ;
        RECT 2043.205 1114.320 2043.375 1114.490 ;
        RECT 2043.665 1114.320 2043.835 1114.490 ;
        RECT 2044.125 1114.320 2044.295 1114.490 ;
        RECT 2044.585 1114.320 2044.755 1114.490 ;
        RECT 2045.045 1114.320 2045.215 1114.490 ;
        RECT 2045.505 1114.320 2045.675 1114.490 ;
        RECT 2045.965 1114.320 2046.135 1114.490 ;
        RECT 2046.425 1114.320 2046.595 1114.490 ;
        RECT 2046.885 1114.320 2047.055 1114.490 ;
        RECT 2047.345 1114.320 2047.515 1114.490 ;
        RECT 2047.805 1114.320 2047.975 1114.490 ;
        RECT 2048.265 1114.320 2048.435 1114.490 ;
        RECT 2048.725 1114.320 2048.895 1114.490 ;
        RECT 2049.185 1114.320 2049.355 1114.490 ;
        RECT 2049.645 1114.320 2049.815 1114.490 ;
        RECT 2050.105 1114.320 2050.275 1114.490 ;
        RECT 2050.565 1114.320 2050.735 1114.490 ;
        RECT 2051.025 1114.320 2051.195 1114.490 ;
        RECT 2051.485 1114.320 2051.655 1114.490 ;
        RECT 2051.945 1114.320 2052.115 1114.490 ;
        RECT 2052.405 1114.320 2052.575 1114.490 ;
        RECT 2052.865 1114.320 2053.035 1114.490 ;
        RECT 2053.325 1114.320 2053.495 1114.490 ;
        RECT 2053.785 1114.320 2053.955 1114.490 ;
        RECT 2054.245 1114.320 2054.415 1114.490 ;
        RECT 2054.705 1114.320 2054.875 1114.490 ;
        RECT 2055.165 1114.320 2055.335 1114.490 ;
        RECT 2055.625 1114.320 2055.795 1114.490 ;
        RECT 2056.085 1114.320 2056.255 1114.490 ;
        RECT 2056.545 1114.320 2056.715 1114.490 ;
        RECT 2057.005 1114.320 2057.175 1114.490 ;
        RECT 2057.465 1114.320 2057.635 1114.490 ;
        RECT 2057.925 1114.320 2058.095 1114.490 ;
        RECT 2058.385 1114.320 2058.555 1114.490 ;
        RECT 2058.845 1114.320 2059.015 1114.490 ;
        RECT 2059.305 1114.320 2059.475 1114.490 ;
        RECT 2059.765 1114.320 2059.935 1114.490 ;
        RECT 2060.225 1114.320 2060.395 1114.490 ;
        RECT 2060.685 1114.320 2060.855 1114.490 ;
        RECT 2061.145 1114.320 2061.315 1114.490 ;
        RECT 2061.605 1114.320 2061.775 1114.490 ;
        RECT 2062.065 1114.320 2062.235 1114.490 ;
        RECT 2062.525 1114.320 2062.695 1114.490 ;
        RECT 2062.985 1114.320 2063.155 1114.490 ;
        RECT 2063.445 1114.320 2063.615 1114.490 ;
        RECT 2063.905 1114.320 2064.075 1114.490 ;
        RECT 2064.365 1114.320 2064.535 1114.490 ;
        RECT 2064.825 1114.320 2064.995 1114.490 ;
        RECT 2065.285 1114.320 2065.455 1114.490 ;
        RECT 2065.745 1114.320 2065.915 1114.490 ;
        RECT 2066.205 1114.320 2066.375 1114.490 ;
        RECT 2066.665 1114.320 2066.835 1114.490 ;
        RECT 2067.125 1114.320 2067.295 1114.490 ;
        RECT 2067.585 1114.320 2067.755 1114.490 ;
        RECT 2068.045 1114.320 2068.215 1114.490 ;
        RECT 2068.505 1114.320 2068.675 1114.490 ;
        RECT 2068.965 1114.320 2069.135 1114.490 ;
        RECT 2069.425 1114.320 2069.595 1114.490 ;
        RECT 2069.885 1114.320 2070.055 1114.490 ;
        RECT 2070.345 1114.320 2070.515 1114.490 ;
        RECT 2070.805 1114.320 2070.975 1114.490 ;
      LAYER met1 ;
        RECT 1969.000 1114.165 2071.120 1114.645 ;
      LAYER via ;
        RECT 2025.150 1114.245 2026.935 1114.545 ;
      LAYER met2 ;
        RECT 2025.110 1114.185 2026.975 1114.615 ;
      LAYER via2 ;
        RECT 2025.150 1114.245 2026.935 1114.545 ;
      LAYER met3 ;
        RECT 2025.120 1109.800 2026.970 1114.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.515 1732.850 201.685 1733.020 ;
        RECT 201.515 1732.390 201.685 1732.560 ;
        RECT 201.515 1731.930 201.685 1732.100 ;
        RECT 201.515 1731.470 201.685 1731.640 ;
        RECT 201.515 1731.010 201.685 1731.180 ;
        RECT 201.515 1730.550 201.685 1730.720 ;
        RECT 201.515 1730.090 201.685 1730.260 ;
        RECT 201.515 1729.630 201.685 1729.800 ;
        RECT 201.515 1729.170 201.685 1729.340 ;
        RECT 201.515 1728.710 201.685 1728.880 ;
        RECT 201.515 1728.250 201.685 1728.420 ;
        RECT 201.515 1727.790 201.685 1727.960 ;
        RECT 201.515 1727.330 201.685 1727.500 ;
        RECT 201.515 1726.870 201.685 1727.040 ;
        RECT 201.515 1726.410 201.685 1726.580 ;
        RECT 201.515 1725.950 201.685 1726.120 ;
        RECT 201.515 1725.490 201.685 1725.660 ;
        RECT 201.515 1725.030 201.685 1725.200 ;
        RECT 201.515 1724.570 201.685 1724.740 ;
        RECT 201.515 1724.110 201.685 1724.280 ;
        RECT 201.515 1723.650 201.685 1723.820 ;
        RECT 201.515 1723.190 201.685 1723.360 ;
        RECT 201.515 1722.730 201.685 1722.900 ;
        RECT 201.515 1722.270 201.685 1722.440 ;
        RECT 201.515 1721.810 201.685 1721.980 ;
        RECT 201.515 1721.350 201.685 1721.520 ;
        RECT 201.515 1720.890 201.685 1721.060 ;
        RECT 201.515 1720.430 201.685 1720.600 ;
        RECT 201.515 1719.970 201.685 1720.140 ;
        RECT 201.515 1719.510 201.685 1719.680 ;
        RECT 201.515 1719.050 201.685 1719.220 ;
        RECT 201.515 1718.590 201.685 1718.760 ;
        RECT 201.515 1718.130 201.685 1718.300 ;
        RECT 201.515 1717.670 201.685 1717.840 ;
        RECT 201.515 1717.210 201.685 1717.380 ;
        RECT 201.515 1716.750 201.685 1716.920 ;
        RECT 201.515 1716.290 201.685 1716.460 ;
        RECT 201.515 1715.830 201.685 1716.000 ;
        RECT 201.515 1715.370 201.685 1715.540 ;
        RECT 201.515 1714.910 201.685 1715.080 ;
        RECT 201.515 1714.450 201.685 1714.620 ;
        RECT 201.515 1713.990 201.685 1714.160 ;
        RECT 201.515 1713.530 201.685 1713.700 ;
        RECT 201.515 1713.070 201.685 1713.240 ;
        RECT 201.515 1712.610 201.685 1712.780 ;
        RECT 201.515 1712.150 201.685 1712.320 ;
        RECT 201.515 1711.690 201.685 1711.860 ;
        RECT 201.515 1711.230 201.685 1711.400 ;
        RECT 201.515 1710.770 201.685 1710.940 ;
        RECT 201.515 1710.310 201.685 1710.480 ;
        RECT 201.515 1709.850 201.685 1710.020 ;
        RECT 201.515 1709.390 201.685 1709.560 ;
        RECT 201.515 1708.930 201.685 1709.100 ;
        RECT 201.515 1708.470 201.685 1708.640 ;
        RECT 201.515 1708.010 201.685 1708.180 ;
        RECT 201.515 1707.550 201.685 1707.720 ;
        RECT 201.515 1707.090 201.685 1707.260 ;
        RECT 201.515 1706.630 201.685 1706.800 ;
        RECT 201.515 1706.170 201.685 1706.340 ;
        RECT 201.515 1705.710 201.685 1705.880 ;
        RECT 201.515 1705.250 201.685 1705.420 ;
        RECT 201.515 1704.790 201.685 1704.960 ;
        RECT 201.515 1704.330 201.685 1704.500 ;
        RECT 201.515 1703.870 201.685 1704.040 ;
        RECT 201.515 1703.410 201.685 1703.580 ;
        RECT 201.515 1702.950 201.685 1703.120 ;
        RECT 201.515 1702.490 201.685 1702.660 ;
        RECT 201.515 1702.030 201.685 1702.200 ;
        RECT 201.515 1701.570 201.685 1701.740 ;
        RECT 201.515 1701.110 201.685 1701.280 ;
        RECT 201.515 1700.650 201.685 1700.820 ;
        RECT 201.515 1700.190 201.685 1700.360 ;
        RECT 201.515 1699.730 201.685 1699.900 ;
        RECT 201.515 1699.270 201.685 1699.440 ;
        RECT 201.515 1698.810 201.685 1698.980 ;
        RECT 201.515 1698.350 201.685 1698.520 ;
        RECT 201.515 1697.890 201.685 1698.060 ;
        RECT 201.515 1697.430 201.685 1697.600 ;
        RECT 201.515 1696.970 201.685 1697.140 ;
        RECT 201.515 1696.510 201.685 1696.680 ;
        RECT 201.515 1696.050 201.685 1696.220 ;
        RECT 201.515 1695.590 201.685 1695.760 ;
        RECT 201.515 1695.130 201.685 1695.300 ;
        RECT 201.515 1694.670 201.685 1694.840 ;
        RECT 201.515 1694.210 201.685 1694.380 ;
        RECT 201.515 1693.750 201.685 1693.920 ;
        RECT 201.515 1693.290 201.685 1693.460 ;
        RECT 201.515 1692.830 201.685 1693.000 ;
        RECT 201.515 1692.370 201.685 1692.540 ;
        RECT 201.515 1691.910 201.685 1692.080 ;
        RECT 201.515 1691.450 201.685 1691.620 ;
        RECT 201.515 1690.990 201.685 1691.160 ;
        RECT 201.515 1690.530 201.685 1690.700 ;
        RECT 201.515 1690.070 201.685 1690.240 ;
        RECT 201.515 1689.610 201.685 1689.780 ;
        RECT 201.515 1689.150 201.685 1689.320 ;
        RECT 201.515 1688.690 201.685 1688.860 ;
        RECT 201.515 1688.230 201.685 1688.400 ;
        RECT 201.515 1687.770 201.685 1687.940 ;
        RECT 201.515 1687.310 201.685 1687.480 ;
        RECT 201.515 1686.850 201.685 1687.020 ;
        RECT 201.515 1686.390 201.685 1686.560 ;
        RECT 201.515 1685.930 201.685 1686.100 ;
        RECT 201.515 1685.470 201.685 1685.640 ;
        RECT 201.515 1685.010 201.685 1685.180 ;
        RECT 201.515 1684.550 201.685 1684.720 ;
        RECT 201.515 1684.090 201.685 1684.260 ;
        RECT 201.515 1683.630 201.685 1683.800 ;
        RECT 201.515 1683.170 201.685 1683.340 ;
        RECT 201.515 1682.710 201.685 1682.880 ;
        RECT 201.515 1682.250 201.685 1682.420 ;
        RECT 201.515 1681.790 201.685 1681.960 ;
        RECT 201.515 1681.330 201.685 1681.500 ;
        RECT 201.515 1680.870 201.685 1681.040 ;
        RECT 201.515 1680.410 201.685 1680.580 ;
        RECT 201.515 1679.950 201.685 1680.120 ;
        RECT 201.515 1679.490 201.685 1679.660 ;
        RECT 201.515 1679.030 201.685 1679.200 ;
        RECT 201.515 1678.570 201.685 1678.740 ;
        RECT 201.515 1678.110 201.685 1678.280 ;
        RECT 201.515 1677.650 201.685 1677.820 ;
        RECT 201.515 1677.190 201.685 1677.360 ;
        RECT 201.515 1676.730 201.685 1676.900 ;
        RECT 201.515 1676.270 201.685 1676.440 ;
        RECT 201.515 1675.810 201.685 1675.980 ;
        RECT 201.515 1675.350 201.685 1675.520 ;
        RECT 201.515 1674.890 201.685 1675.060 ;
        RECT 201.515 1674.430 201.685 1674.600 ;
        RECT 201.515 1673.970 201.685 1674.140 ;
        RECT 201.515 1673.510 201.685 1673.680 ;
        RECT 201.515 1673.050 201.685 1673.220 ;
      LAYER met1 ;
        RECT 201.360 1672.905 201.840 1733.165 ;
      LAYER via ;
        RECT 201.455 1716.855 201.755 1718.640 ;
      LAYER met2 ;
        RECT 201.395 1716.815 201.825 1718.680 ;
      LAYER via2 ;
        RECT 201.455 1716.855 201.755 1718.640 ;
      LAYER met3 ;
        RECT 197.010 1716.820 201.825 1718.670 ;
    END
    PORT
      LAYER li1 ;
        RECT 3386.220 2238.065 3386.390 2238.235 ;
        RECT 3386.220 2237.605 3386.390 2237.775 ;
        RECT 3386.220 2237.145 3386.390 2237.315 ;
        RECT 3386.220 2236.685 3386.390 2236.855 ;
        RECT 3386.220 2236.225 3386.390 2236.395 ;
        RECT 3386.220 2235.765 3386.390 2235.935 ;
        RECT 3386.220 2235.305 3386.390 2235.475 ;
        RECT 3386.220 2234.845 3386.390 2235.015 ;
        RECT 3386.220 2234.385 3386.390 2234.555 ;
        RECT 3386.220 2233.925 3386.390 2234.095 ;
        RECT 3386.220 2233.465 3386.390 2233.635 ;
        RECT 3386.220 2233.005 3386.390 2233.175 ;
        RECT 3386.220 2232.545 3386.390 2232.715 ;
        RECT 3386.220 2232.085 3386.390 2232.255 ;
        RECT 3386.220 2231.625 3386.390 2231.795 ;
        RECT 3386.220 2231.165 3386.390 2231.335 ;
        RECT 3386.220 2230.705 3386.390 2230.875 ;
        RECT 3386.220 2230.245 3386.390 2230.415 ;
        RECT 3386.220 2229.785 3386.390 2229.955 ;
        RECT 3386.220 2229.325 3386.390 2229.495 ;
        RECT 3386.220 2228.865 3386.390 2229.035 ;
        RECT 3386.220 2228.405 3386.390 2228.575 ;
        RECT 3386.220 2227.945 3386.390 2228.115 ;
        RECT 3386.220 2227.485 3386.390 2227.655 ;
        RECT 3386.220 2227.025 3386.390 2227.195 ;
        RECT 3386.220 2226.565 3386.390 2226.735 ;
        RECT 3386.220 2226.105 3386.390 2226.275 ;
        RECT 3386.220 2225.645 3386.390 2225.815 ;
        RECT 3386.220 2225.185 3386.390 2225.355 ;
        RECT 3386.220 2224.725 3386.390 2224.895 ;
        RECT 3386.220 2224.265 3386.390 2224.435 ;
        RECT 3386.220 2223.805 3386.390 2223.975 ;
        RECT 3386.220 2223.345 3386.390 2223.515 ;
        RECT 3386.220 2222.885 3386.390 2223.055 ;
        RECT 3386.220 2222.425 3386.390 2222.595 ;
        RECT 3386.220 2221.965 3386.390 2222.135 ;
        RECT 3386.220 2221.505 3386.390 2221.675 ;
        RECT 3386.220 2221.045 3386.390 2221.215 ;
        RECT 3386.220 2220.585 3386.390 2220.755 ;
        RECT 3386.220 2220.125 3386.390 2220.295 ;
        RECT 3386.220 2219.665 3386.390 2219.835 ;
        RECT 3386.220 2219.205 3386.390 2219.375 ;
        RECT 3386.220 2218.745 3386.390 2218.915 ;
        RECT 3386.220 2218.285 3386.390 2218.455 ;
        RECT 3386.220 2217.825 3386.390 2217.995 ;
        RECT 3386.220 2217.365 3386.390 2217.535 ;
        RECT 3386.220 2216.905 3386.390 2217.075 ;
        RECT 3386.220 2216.445 3386.390 2216.615 ;
        RECT 3386.220 2215.985 3386.390 2216.155 ;
        RECT 3386.220 2215.525 3386.390 2215.695 ;
        RECT 3386.220 2215.065 3386.390 2215.235 ;
        RECT 3386.220 2214.605 3386.390 2214.775 ;
        RECT 3386.220 2214.145 3386.390 2214.315 ;
        RECT 3386.220 2213.685 3386.390 2213.855 ;
        RECT 3386.220 2213.225 3386.390 2213.395 ;
        RECT 3386.220 2212.765 3386.390 2212.935 ;
        RECT 3386.220 2212.305 3386.390 2212.475 ;
        RECT 3386.220 2211.845 3386.390 2212.015 ;
        RECT 3386.220 2211.385 3386.390 2211.555 ;
        RECT 3386.220 2210.925 3386.390 2211.095 ;
        RECT 3386.220 2210.465 3386.390 2210.635 ;
        RECT 3386.220 2210.005 3386.390 2210.175 ;
        RECT 3386.220 2209.545 3386.390 2209.715 ;
        RECT 3386.220 2209.085 3386.390 2209.255 ;
        RECT 3386.220 2208.625 3386.390 2208.795 ;
        RECT 3386.220 2208.165 3386.390 2208.335 ;
        RECT 3386.220 2207.705 3386.390 2207.875 ;
        RECT 3386.220 2207.245 3386.390 2207.415 ;
        RECT 3386.220 2206.785 3386.390 2206.955 ;
        RECT 3386.220 2206.325 3386.390 2206.495 ;
        RECT 3386.220 2205.865 3386.390 2206.035 ;
        RECT 3386.220 2205.405 3386.390 2205.575 ;
        RECT 3386.220 2204.945 3386.390 2205.115 ;
        RECT 3386.220 2204.485 3386.390 2204.655 ;
        RECT 3386.220 2204.025 3386.390 2204.195 ;
        RECT 3386.220 2203.565 3386.390 2203.735 ;
        RECT 3386.220 2203.105 3386.390 2203.275 ;
        RECT 3386.220 2202.645 3386.390 2202.815 ;
        RECT 3386.220 2202.185 3386.390 2202.355 ;
        RECT 3386.220 2201.725 3386.390 2201.895 ;
        RECT 3386.220 2201.265 3386.390 2201.435 ;
        RECT 3386.220 2200.805 3386.390 2200.975 ;
        RECT 3386.220 2200.345 3386.390 2200.515 ;
        RECT 3386.220 2199.885 3386.390 2200.055 ;
        RECT 3386.220 2199.425 3386.390 2199.595 ;
        RECT 3386.220 2198.965 3386.390 2199.135 ;
        RECT 3386.220 2198.505 3386.390 2198.675 ;
        RECT 3386.220 2198.045 3386.390 2198.215 ;
        RECT 3386.220 2197.585 3386.390 2197.755 ;
        RECT 3386.220 2197.125 3386.390 2197.295 ;
        RECT 3386.220 2196.665 3386.390 2196.835 ;
        RECT 3386.220 2196.205 3386.390 2196.375 ;
      LAYER met1 ;
        RECT 3386.065 2196.060 3386.545 2238.380 ;
      LAYER via ;
        RECT 3386.130 2234.495 3386.430 2236.280 ;
      LAYER met2 ;
        RECT 3386.060 2234.455 3386.490 2236.320 ;
      LAYER via2 ;
        RECT 3386.130 2234.495 3386.430 2236.280 ;
      LAYER met3 ;
        RECT 3386.060 2234.465 3390.875 2236.315 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.405 3023.755 201.575 3023.925 ;
        RECT 201.405 3023.295 201.575 3023.465 ;
        RECT 201.405 3022.835 201.575 3023.005 ;
        RECT 201.405 3022.375 201.575 3022.545 ;
        RECT 201.405 3021.915 201.575 3022.085 ;
        RECT 201.405 3021.455 201.575 3021.625 ;
        RECT 201.405 3020.995 201.575 3021.165 ;
        RECT 201.405 3020.535 201.575 3020.705 ;
        RECT 201.405 3020.075 201.575 3020.245 ;
        RECT 201.405 3019.615 201.575 3019.785 ;
        RECT 201.405 3019.155 201.575 3019.325 ;
        RECT 201.405 3018.695 201.575 3018.865 ;
        RECT 201.405 3018.235 201.575 3018.405 ;
        RECT 201.405 3017.775 201.575 3017.945 ;
        RECT 201.405 3017.315 201.575 3017.485 ;
        RECT 201.405 3016.855 201.575 3017.025 ;
        RECT 201.405 3016.395 201.575 3016.565 ;
        RECT 201.405 3015.935 201.575 3016.105 ;
        RECT 201.405 3015.475 201.575 3015.645 ;
        RECT 201.405 3015.015 201.575 3015.185 ;
        RECT 201.405 3014.555 201.575 3014.725 ;
        RECT 201.405 3014.095 201.575 3014.265 ;
        RECT 201.405 3013.635 201.575 3013.805 ;
        RECT 201.405 3013.175 201.575 3013.345 ;
        RECT 201.405 3012.715 201.575 3012.885 ;
        RECT 201.405 3012.255 201.575 3012.425 ;
        RECT 201.405 3011.795 201.575 3011.965 ;
        RECT 201.405 3011.335 201.575 3011.505 ;
        RECT 201.405 3010.875 201.575 3011.045 ;
        RECT 201.405 3010.415 201.575 3010.585 ;
        RECT 201.405 3009.955 201.575 3010.125 ;
        RECT 201.405 3009.495 201.575 3009.665 ;
        RECT 201.405 3009.035 201.575 3009.205 ;
        RECT 201.405 3008.575 201.575 3008.745 ;
        RECT 201.405 3008.115 201.575 3008.285 ;
        RECT 201.405 3007.655 201.575 3007.825 ;
        RECT 201.405 3007.195 201.575 3007.365 ;
        RECT 201.405 3006.735 201.575 3006.905 ;
        RECT 201.405 3006.275 201.575 3006.445 ;
        RECT 201.405 3005.815 201.575 3005.985 ;
        RECT 201.405 3005.355 201.575 3005.525 ;
        RECT 201.405 3004.895 201.575 3005.065 ;
        RECT 201.405 3004.435 201.575 3004.605 ;
        RECT 201.405 3003.975 201.575 3004.145 ;
        RECT 201.405 3003.515 201.575 3003.685 ;
        RECT 201.405 3003.055 201.575 3003.225 ;
        RECT 201.405 3002.595 201.575 3002.765 ;
        RECT 201.405 3002.135 201.575 3002.305 ;
        RECT 201.405 3001.675 201.575 3001.845 ;
        RECT 201.405 3001.215 201.575 3001.385 ;
        RECT 201.405 3000.755 201.575 3000.925 ;
        RECT 201.405 3000.295 201.575 3000.465 ;
        RECT 201.405 2999.835 201.575 3000.005 ;
        RECT 201.405 2999.375 201.575 2999.545 ;
        RECT 201.405 2998.915 201.575 2999.085 ;
        RECT 201.405 2998.455 201.575 2998.625 ;
        RECT 201.405 2997.995 201.575 2998.165 ;
        RECT 201.405 2997.535 201.575 2997.705 ;
        RECT 201.405 2997.075 201.575 2997.245 ;
        RECT 201.405 2996.615 201.575 2996.785 ;
        RECT 201.405 2996.155 201.575 2996.325 ;
        RECT 201.405 2995.695 201.575 2995.865 ;
        RECT 201.405 2995.235 201.575 2995.405 ;
        RECT 201.405 2994.775 201.575 2994.945 ;
        RECT 201.405 2994.315 201.575 2994.485 ;
        RECT 201.405 2993.855 201.575 2994.025 ;
        RECT 201.405 2993.395 201.575 2993.565 ;
        RECT 201.405 2992.935 201.575 2993.105 ;
        RECT 201.405 2992.475 201.575 2992.645 ;
        RECT 201.405 2992.015 201.575 2992.185 ;
        RECT 201.405 2991.555 201.575 2991.725 ;
        RECT 201.405 2991.095 201.575 2991.265 ;
        RECT 201.405 2990.635 201.575 2990.805 ;
        RECT 201.405 2990.175 201.575 2990.345 ;
        RECT 201.405 2989.715 201.575 2989.885 ;
        RECT 201.405 2989.255 201.575 2989.425 ;
        RECT 201.405 2988.795 201.575 2988.965 ;
        RECT 201.405 2988.335 201.575 2988.505 ;
        RECT 201.405 2987.875 201.575 2988.045 ;
      LAYER met1 ;
        RECT 201.250 2987.730 201.730 3024.070 ;
      LAYER via ;
        RECT 201.360 3014.090 201.660 3015.875 ;
      LAYER met2 ;
        RECT 201.300 3014.050 201.730 3015.915 ;
      LAYER via2 ;
        RECT 201.360 3014.090 201.660 3015.875 ;
      LAYER met3 ;
        RECT 196.915 3014.055 201.730 3015.905 ;
    END
    PORT
      LAYER li1 ;
        RECT 3386.220 3542.185 3386.390 3542.355 ;
        RECT 3386.220 3541.725 3386.390 3541.895 ;
        RECT 3386.220 3541.265 3386.390 3541.435 ;
        RECT 3386.220 3540.805 3386.390 3540.975 ;
        RECT 3386.220 3540.345 3386.390 3540.515 ;
        RECT 3386.220 3539.885 3386.390 3540.055 ;
        RECT 3386.220 3539.425 3386.390 3539.595 ;
        RECT 3386.220 3538.965 3386.390 3539.135 ;
        RECT 3386.220 3538.505 3386.390 3538.675 ;
        RECT 3386.220 3538.045 3386.390 3538.215 ;
        RECT 3386.220 3537.585 3386.390 3537.755 ;
        RECT 3386.220 3537.125 3386.390 3537.295 ;
        RECT 3386.220 3536.665 3386.390 3536.835 ;
        RECT 3386.220 3536.205 3386.390 3536.375 ;
      LAYER met1 ;
        RECT 3386.065 3532.490 3386.545 3542.500 ;
      LAYER via ;
        RECT 3386.170 3532.560 3386.470 3534.345 ;
      LAYER met2 ;
        RECT 3386.100 3532.520 3386.530 3534.385 ;
      LAYER via2 ;
        RECT 3386.170 3532.560 3386.470 3534.345 ;
      LAYER met3 ;
        RECT 3386.100 3532.530 3390.915 3534.380 ;
    END
  END vccd
  OBS
      LAYER pwell ;
        RECT 3383.775 3542.055 3384.560 3542.485 ;
        RECT 3383.690 3541.890 3384.600 3542.035 ;
        RECT 3383.500 3541.720 3384.600 3541.890 ;
        RECT 3383.690 3536.905 3384.600 3541.720 ;
        RECT 3383.775 3536.075 3384.560 3536.505 ;
      LAYER nwell ;
        RECT 3384.890 3535.870 3387.720 3542.690 ;
      LAYER pwell ;
        RECT 3388.050 3542.055 3388.835 3542.485 ;
        RECT 3388.010 3536.840 3388.920 3541.655 ;
        RECT 3388.010 3536.670 3389.110 3536.840 ;
        RECT 3388.010 3536.525 3388.920 3536.670 ;
        RECT 3388.050 3536.075 3388.835 3536.505 ;
        RECT 198.960 3023.625 199.745 3024.055 ;
        RECT 198.875 3018.410 199.785 3023.225 ;
        RECT 198.685 3018.240 199.785 3018.410 ;
        RECT 198.875 3018.095 199.785 3018.240 ;
        RECT 198.960 3017.645 199.745 3018.075 ;
        RECT 198.875 3012.430 199.785 3017.245 ;
        RECT 198.685 3012.260 199.785 3012.430 ;
        RECT 198.875 3012.115 199.785 3012.260 ;
        RECT 198.960 3011.665 199.745 3012.095 ;
        RECT 198.875 3006.450 199.785 3011.265 ;
        RECT 198.685 3006.280 199.785 3006.450 ;
        RECT 198.875 3006.135 199.785 3006.280 ;
        RECT 198.960 3005.685 199.745 3006.115 ;
        RECT 198.875 3000.470 199.785 3005.285 ;
        RECT 198.685 3000.300 199.785 3000.470 ;
        RECT 198.875 3000.155 199.785 3000.300 ;
        RECT 198.960 2999.705 199.745 3000.135 ;
        RECT 198.875 2994.490 199.785 2999.305 ;
        RECT 198.685 2994.320 199.785 2994.490 ;
        RECT 198.875 2994.175 199.785 2994.320 ;
        RECT 198.960 2993.725 199.745 2994.155 ;
        RECT 198.875 2988.510 199.785 2993.325 ;
        RECT 198.685 2988.340 199.785 2988.510 ;
        RECT 198.875 2988.195 199.785 2988.340 ;
        RECT 198.960 2987.745 199.745 2988.175 ;
      LAYER nwell ;
        RECT 200.075 2987.540 202.905 3024.260 ;
      LAYER pwell ;
        RECT 203.235 3023.625 204.020 3024.055 ;
        RECT 203.195 3023.460 204.105 3023.605 ;
        RECT 203.195 3023.290 204.295 3023.460 ;
        RECT 203.195 3018.475 204.105 3023.290 ;
        RECT 203.235 3017.645 204.020 3018.075 ;
        RECT 203.195 3017.480 204.105 3017.625 ;
        RECT 203.195 3017.310 204.295 3017.480 ;
        RECT 203.195 3012.495 204.105 3017.310 ;
        RECT 203.235 3011.665 204.020 3012.095 ;
        RECT 203.195 3011.500 204.105 3011.645 ;
        RECT 203.195 3011.330 204.295 3011.500 ;
        RECT 203.195 3006.515 204.105 3011.330 ;
        RECT 203.235 3005.685 204.020 3006.115 ;
        RECT 203.195 3005.520 204.105 3005.665 ;
        RECT 203.195 3005.350 204.295 3005.520 ;
        RECT 203.195 3000.535 204.105 3005.350 ;
        RECT 203.235 2999.705 204.020 3000.135 ;
        RECT 203.195 2999.540 204.105 2999.685 ;
        RECT 203.195 2999.370 204.295 2999.540 ;
        RECT 203.195 2994.555 204.105 2999.370 ;
        RECT 203.235 2993.725 204.020 2994.155 ;
        RECT 203.195 2993.560 204.105 2993.705 ;
        RECT 203.195 2993.390 204.295 2993.560 ;
        RECT 203.195 2988.575 204.105 2993.390 ;
        RECT 203.235 2987.745 204.020 2988.175 ;
        RECT 3383.775 2237.935 3384.560 2238.365 ;
        RECT 3383.690 2237.770 3384.600 2237.915 ;
        RECT 3383.500 2237.600 3384.600 2237.770 ;
        RECT 3383.690 2232.785 3384.600 2237.600 ;
        RECT 3383.775 2231.955 3384.560 2232.385 ;
        RECT 3383.690 2231.790 3384.600 2231.935 ;
        RECT 3383.500 2231.620 3384.600 2231.790 ;
        RECT 3383.690 2226.805 3384.600 2231.620 ;
        RECT 3383.775 2225.975 3384.560 2226.405 ;
        RECT 3383.690 2225.810 3384.600 2225.955 ;
        RECT 3383.500 2225.640 3384.600 2225.810 ;
        RECT 3383.690 2220.825 3384.600 2225.640 ;
        RECT 3383.775 2219.995 3384.560 2220.425 ;
        RECT 3383.690 2219.830 3384.600 2219.975 ;
        RECT 3383.500 2219.660 3384.600 2219.830 ;
        RECT 3383.690 2214.845 3384.600 2219.660 ;
        RECT 3383.775 2214.015 3384.560 2214.445 ;
        RECT 3383.690 2213.850 3384.600 2213.995 ;
        RECT 3383.500 2213.680 3384.600 2213.850 ;
        RECT 3383.690 2208.865 3384.600 2213.680 ;
        RECT 3383.775 2208.035 3384.560 2208.465 ;
        RECT 3383.690 2207.870 3384.600 2208.015 ;
        RECT 3383.500 2207.700 3384.600 2207.870 ;
        RECT 3383.690 2202.885 3384.600 2207.700 ;
        RECT 3383.775 2202.055 3384.560 2202.485 ;
        RECT 3383.690 2201.890 3384.600 2202.035 ;
        RECT 3383.500 2201.720 3384.600 2201.890 ;
        RECT 3383.690 2196.905 3384.600 2201.720 ;
        RECT 3383.775 2196.075 3384.560 2196.505 ;
      LAYER nwell ;
        RECT 3384.890 2195.870 3387.720 2238.570 ;
      LAYER pwell ;
        RECT 3388.050 2237.935 3388.835 2238.365 ;
        RECT 3388.010 2232.720 3388.920 2237.535 ;
        RECT 3388.010 2232.550 3389.110 2232.720 ;
        RECT 3388.010 2232.405 3388.920 2232.550 ;
        RECT 3388.050 2231.955 3388.835 2232.385 ;
        RECT 3388.010 2226.740 3388.920 2231.555 ;
        RECT 3388.010 2226.570 3389.110 2226.740 ;
        RECT 3388.010 2226.425 3388.920 2226.570 ;
        RECT 3388.050 2225.975 3388.835 2226.405 ;
        RECT 3388.010 2220.760 3388.920 2225.575 ;
        RECT 3388.010 2220.590 3389.110 2220.760 ;
        RECT 3388.010 2220.445 3388.920 2220.590 ;
        RECT 3388.050 2219.995 3388.835 2220.425 ;
        RECT 3388.010 2214.780 3388.920 2219.595 ;
        RECT 3388.010 2214.610 3389.110 2214.780 ;
        RECT 3388.010 2214.465 3388.920 2214.610 ;
        RECT 3388.050 2214.015 3388.835 2214.445 ;
        RECT 3388.010 2208.800 3388.920 2213.615 ;
        RECT 3388.010 2208.630 3389.110 2208.800 ;
        RECT 3388.010 2208.485 3388.920 2208.630 ;
        RECT 3388.050 2208.035 3388.835 2208.465 ;
        RECT 3388.010 2202.820 3388.920 2207.635 ;
        RECT 3388.010 2202.650 3389.110 2202.820 ;
        RECT 3388.010 2202.505 3388.920 2202.650 ;
        RECT 3388.050 2202.055 3388.835 2202.485 ;
        RECT 3388.010 2196.840 3388.920 2201.655 ;
        RECT 3388.010 2196.670 3389.110 2196.840 ;
        RECT 3388.010 2196.525 3388.920 2196.670 ;
        RECT 3388.050 2196.075 3388.835 2196.505 ;
        RECT 199.070 1732.720 199.855 1733.150 ;
        RECT 198.985 1727.505 199.895 1732.320 ;
        RECT 198.795 1727.335 199.895 1727.505 ;
        RECT 198.985 1727.190 199.895 1727.335 ;
        RECT 199.070 1726.740 199.855 1727.170 ;
        RECT 198.985 1721.525 199.895 1726.340 ;
        RECT 198.795 1721.355 199.895 1721.525 ;
        RECT 198.985 1721.210 199.895 1721.355 ;
        RECT 199.070 1720.760 199.855 1721.190 ;
        RECT 198.985 1715.545 199.895 1720.360 ;
        RECT 198.795 1715.375 199.895 1715.545 ;
        RECT 198.985 1715.230 199.895 1715.375 ;
        RECT 199.070 1714.780 199.855 1715.210 ;
        RECT 198.985 1709.565 199.895 1714.380 ;
        RECT 198.795 1709.395 199.895 1709.565 ;
        RECT 198.985 1709.250 199.895 1709.395 ;
        RECT 199.070 1708.800 199.855 1709.230 ;
        RECT 198.985 1703.585 199.895 1708.400 ;
        RECT 198.795 1703.415 199.895 1703.585 ;
        RECT 198.985 1703.270 199.895 1703.415 ;
        RECT 199.070 1702.820 199.855 1703.250 ;
        RECT 198.985 1697.605 199.895 1702.420 ;
        RECT 198.795 1697.435 199.895 1697.605 ;
        RECT 198.985 1697.290 199.895 1697.435 ;
        RECT 199.070 1696.840 199.855 1697.270 ;
        RECT 198.985 1691.625 199.895 1696.440 ;
        RECT 198.795 1691.455 199.895 1691.625 ;
        RECT 198.985 1691.310 199.895 1691.455 ;
        RECT 199.070 1690.860 199.855 1691.290 ;
        RECT 198.985 1685.645 199.895 1690.460 ;
        RECT 198.795 1685.475 199.895 1685.645 ;
        RECT 198.985 1685.330 199.895 1685.475 ;
        RECT 199.070 1684.880 199.855 1685.310 ;
        RECT 198.985 1679.665 199.895 1684.480 ;
        RECT 198.795 1679.495 199.895 1679.665 ;
        RECT 198.985 1679.350 199.895 1679.495 ;
        RECT 199.070 1678.900 199.855 1679.330 ;
        RECT 198.985 1673.685 199.895 1678.500 ;
        RECT 198.795 1673.515 199.895 1673.685 ;
        RECT 198.985 1673.370 199.895 1673.515 ;
        RECT 199.070 1672.920 199.855 1673.350 ;
      LAYER nwell ;
        RECT 200.185 1672.715 203.015 1733.355 ;
      LAYER pwell ;
        RECT 203.345 1732.720 204.130 1733.150 ;
        RECT 203.305 1732.555 204.215 1732.700 ;
        RECT 203.305 1732.385 204.405 1732.555 ;
        RECT 203.305 1727.570 204.215 1732.385 ;
        RECT 203.345 1726.740 204.130 1727.170 ;
        RECT 203.305 1726.575 204.215 1726.720 ;
        RECT 203.305 1726.405 204.405 1726.575 ;
        RECT 203.305 1721.590 204.215 1726.405 ;
        RECT 203.345 1720.760 204.130 1721.190 ;
        RECT 203.305 1720.595 204.215 1720.740 ;
        RECT 203.305 1720.425 204.405 1720.595 ;
        RECT 203.305 1715.610 204.215 1720.425 ;
        RECT 203.345 1714.780 204.130 1715.210 ;
        RECT 203.305 1714.615 204.215 1714.760 ;
        RECT 203.305 1714.445 204.405 1714.615 ;
        RECT 203.305 1709.630 204.215 1714.445 ;
        RECT 203.345 1708.800 204.130 1709.230 ;
        RECT 203.305 1708.635 204.215 1708.780 ;
        RECT 203.305 1708.465 204.405 1708.635 ;
        RECT 203.305 1703.650 204.215 1708.465 ;
        RECT 203.345 1702.820 204.130 1703.250 ;
        RECT 203.305 1702.655 204.215 1702.800 ;
        RECT 203.305 1702.485 204.405 1702.655 ;
        RECT 203.305 1697.670 204.215 1702.485 ;
        RECT 203.345 1696.840 204.130 1697.270 ;
        RECT 203.305 1696.675 204.215 1696.820 ;
        RECT 203.305 1696.505 204.405 1696.675 ;
        RECT 203.305 1691.690 204.215 1696.505 ;
        RECT 203.345 1690.860 204.130 1691.290 ;
        RECT 203.305 1690.695 204.215 1690.840 ;
        RECT 203.305 1690.525 204.405 1690.695 ;
        RECT 203.305 1685.710 204.215 1690.525 ;
        RECT 203.345 1684.880 204.130 1685.310 ;
        RECT 203.305 1684.715 204.215 1684.860 ;
        RECT 203.305 1684.545 204.405 1684.715 ;
        RECT 203.305 1679.730 204.215 1684.545 ;
        RECT 203.345 1678.900 204.130 1679.330 ;
        RECT 203.305 1678.735 204.215 1678.880 ;
        RECT 203.305 1678.565 204.405 1678.735 ;
        RECT 203.305 1673.750 204.215 1678.565 ;
        RECT 203.345 1672.920 204.130 1673.350 ;
        RECT 674.660 1117.020 674.830 1117.210 ;
        RECT 680.640 1117.020 680.810 1117.210 ;
        RECT 686.620 1117.020 686.790 1117.210 ;
        RECT 692.600 1117.020 692.770 1117.210 ;
        RECT 698.580 1117.020 698.750 1117.210 ;
        RECT 704.560 1117.020 704.730 1117.210 ;
        RECT 710.540 1117.020 710.710 1117.210 ;
        RECT 716.520 1117.020 716.690 1117.210 ;
        RECT 722.500 1117.020 722.670 1117.210 ;
        RECT 728.480 1117.020 728.650 1117.210 ;
        RECT 734.460 1117.020 734.630 1117.210 ;
        RECT 740.440 1117.020 740.610 1117.210 ;
        RECT 746.420 1117.020 746.590 1117.210 ;
        RECT 752.400 1117.020 752.570 1117.210 ;
        RECT 758.380 1117.020 758.550 1117.210 ;
        RECT 764.360 1117.020 764.530 1117.210 ;
        RECT 770.340 1117.020 770.510 1117.210 ;
        RECT 1974.660 1117.020 1974.830 1117.210 ;
        RECT 1980.640 1117.020 1980.810 1117.210 ;
        RECT 1986.620 1117.020 1986.790 1117.210 ;
        RECT 1992.600 1117.020 1992.770 1117.210 ;
        RECT 1998.580 1117.020 1998.750 1117.210 ;
        RECT 2004.560 1117.020 2004.730 1117.210 ;
        RECT 2010.540 1117.020 2010.710 1117.210 ;
        RECT 2016.520 1117.020 2016.690 1117.210 ;
        RECT 2022.500 1117.020 2022.670 1117.210 ;
        RECT 2028.480 1117.020 2028.650 1117.210 ;
        RECT 2034.460 1117.020 2034.630 1117.210 ;
        RECT 2040.440 1117.020 2040.610 1117.210 ;
        RECT 2046.420 1117.020 2046.590 1117.210 ;
        RECT 2052.400 1117.020 2052.570 1117.210 ;
        RECT 2058.380 1117.020 2058.550 1117.210 ;
        RECT 2064.360 1117.020 2064.530 1117.210 ;
        RECT 2070.340 1117.020 2070.510 1117.210 ;
        RECT 669.015 1116.150 669.445 1116.935 ;
        RECT 669.845 1116.110 674.975 1117.020 ;
        RECT 674.995 1116.150 675.425 1116.935 ;
        RECT 675.825 1116.110 680.955 1117.020 ;
        RECT 680.975 1116.150 681.405 1116.935 ;
        RECT 681.805 1116.110 686.935 1117.020 ;
        RECT 686.955 1116.150 687.385 1116.935 ;
        RECT 687.785 1116.110 692.915 1117.020 ;
        RECT 692.935 1116.150 693.365 1116.935 ;
        RECT 693.765 1116.110 698.895 1117.020 ;
        RECT 698.915 1116.150 699.345 1116.935 ;
        RECT 699.745 1116.110 704.875 1117.020 ;
        RECT 704.895 1116.150 705.325 1116.935 ;
        RECT 705.725 1116.110 710.855 1117.020 ;
        RECT 710.875 1116.150 711.305 1116.935 ;
        RECT 711.705 1116.110 716.835 1117.020 ;
        RECT 716.855 1116.150 717.285 1116.935 ;
        RECT 717.685 1116.110 722.815 1117.020 ;
        RECT 722.835 1116.150 723.265 1116.935 ;
        RECT 723.665 1116.110 728.795 1117.020 ;
        RECT 728.815 1116.150 729.245 1116.935 ;
        RECT 729.645 1116.110 734.775 1117.020 ;
        RECT 734.795 1116.150 735.225 1116.935 ;
        RECT 735.625 1116.110 740.755 1117.020 ;
        RECT 740.775 1116.150 741.205 1116.935 ;
        RECT 741.605 1116.110 746.735 1117.020 ;
        RECT 746.755 1116.150 747.185 1116.935 ;
        RECT 747.585 1116.110 752.715 1117.020 ;
        RECT 752.735 1116.150 753.165 1116.935 ;
        RECT 753.565 1116.110 758.695 1117.020 ;
        RECT 758.715 1116.150 759.145 1116.935 ;
        RECT 759.545 1116.110 764.675 1117.020 ;
        RECT 764.695 1116.150 765.125 1116.935 ;
        RECT 765.525 1116.110 770.655 1117.020 ;
        RECT 770.675 1116.150 771.105 1116.935 ;
        RECT 1969.015 1116.150 1969.445 1116.935 ;
        RECT 1969.845 1116.110 1974.975 1117.020 ;
        RECT 1974.995 1116.150 1975.425 1116.935 ;
        RECT 1975.825 1116.110 1980.955 1117.020 ;
        RECT 1980.975 1116.150 1981.405 1116.935 ;
        RECT 1981.805 1116.110 1986.935 1117.020 ;
        RECT 1986.955 1116.150 1987.385 1116.935 ;
        RECT 1987.785 1116.110 1992.915 1117.020 ;
        RECT 1992.935 1116.150 1993.365 1116.935 ;
        RECT 1993.765 1116.110 1998.895 1117.020 ;
        RECT 1998.915 1116.150 1999.345 1116.935 ;
        RECT 1999.745 1116.110 2004.875 1117.020 ;
        RECT 2004.895 1116.150 2005.325 1116.935 ;
        RECT 2005.725 1116.110 2010.855 1117.020 ;
        RECT 2010.875 1116.150 2011.305 1116.935 ;
        RECT 2011.705 1116.110 2016.835 1117.020 ;
        RECT 2016.855 1116.150 2017.285 1116.935 ;
        RECT 2017.685 1116.110 2022.815 1117.020 ;
        RECT 2022.835 1116.150 2023.265 1116.935 ;
        RECT 2023.665 1116.110 2028.795 1117.020 ;
        RECT 2028.815 1116.150 2029.245 1116.935 ;
        RECT 2029.645 1116.110 2034.775 1117.020 ;
        RECT 2034.795 1116.150 2035.225 1116.935 ;
        RECT 2035.625 1116.110 2040.755 1117.020 ;
        RECT 2040.775 1116.150 2041.205 1116.935 ;
        RECT 2041.605 1116.110 2046.735 1117.020 ;
        RECT 2046.755 1116.150 2047.185 1116.935 ;
        RECT 2047.585 1116.110 2052.715 1117.020 ;
        RECT 2052.735 1116.150 2053.165 1116.935 ;
        RECT 2053.565 1116.110 2058.695 1117.020 ;
        RECT 2058.715 1116.150 2059.145 1116.935 ;
        RECT 2059.545 1116.110 2064.675 1117.020 ;
        RECT 2064.695 1116.150 2065.125 1116.935 ;
        RECT 2065.525 1116.110 2070.655 1117.020 ;
        RECT 2070.675 1116.150 2071.105 1116.935 ;
      LAYER nwell ;
        RECT 668.810 1114.215 771.310 1115.820 ;
        RECT 1968.810 1114.215 2071.310 1115.820 ;
        RECT 674.790 1112.990 771.310 1114.215 ;
        RECT 1974.790 1112.990 2071.310 1114.215 ;
      LAYER pwell ;
        RECT 674.995 1111.875 675.425 1112.660 ;
        RECT 675.445 1111.790 680.575 1112.700 ;
        RECT 680.975 1111.875 681.405 1112.660 ;
        RECT 681.425 1111.790 686.555 1112.700 ;
        RECT 686.955 1111.875 687.385 1112.660 ;
        RECT 687.405 1111.790 692.535 1112.700 ;
        RECT 692.935 1111.875 693.365 1112.660 ;
        RECT 693.385 1111.790 698.515 1112.700 ;
        RECT 698.915 1111.875 699.345 1112.660 ;
        RECT 699.365 1111.790 704.495 1112.700 ;
        RECT 704.895 1111.875 705.325 1112.660 ;
        RECT 705.345 1111.790 710.475 1112.700 ;
        RECT 710.875 1111.875 711.305 1112.660 ;
        RECT 711.325 1111.790 716.455 1112.700 ;
        RECT 716.855 1111.875 717.285 1112.660 ;
        RECT 717.305 1111.790 722.435 1112.700 ;
        RECT 722.835 1111.875 723.265 1112.660 ;
        RECT 723.285 1111.790 728.415 1112.700 ;
        RECT 728.815 1111.875 729.245 1112.660 ;
        RECT 729.265 1111.790 734.395 1112.700 ;
        RECT 734.795 1111.875 735.225 1112.660 ;
        RECT 735.245 1111.790 740.375 1112.700 ;
        RECT 740.775 1111.875 741.205 1112.660 ;
        RECT 741.225 1111.790 746.355 1112.700 ;
        RECT 746.755 1111.875 747.185 1112.660 ;
        RECT 747.205 1111.790 752.335 1112.700 ;
        RECT 752.735 1111.875 753.165 1112.660 ;
        RECT 753.185 1111.790 758.315 1112.700 ;
        RECT 758.715 1111.875 759.145 1112.660 ;
        RECT 759.165 1111.790 764.295 1112.700 ;
        RECT 764.695 1111.875 765.125 1112.660 ;
        RECT 765.525 1111.790 770.655 1112.700 ;
        RECT 770.675 1111.875 771.105 1112.660 ;
        RECT 1974.995 1111.875 1975.425 1112.660 ;
        RECT 1975.445 1111.790 1980.575 1112.700 ;
        RECT 1980.975 1111.875 1981.405 1112.660 ;
        RECT 1981.425 1111.790 1986.555 1112.700 ;
        RECT 1986.955 1111.875 1987.385 1112.660 ;
        RECT 1987.405 1111.790 1992.535 1112.700 ;
        RECT 1992.935 1111.875 1993.365 1112.660 ;
        RECT 1993.385 1111.790 1998.515 1112.700 ;
        RECT 1998.915 1111.875 1999.345 1112.660 ;
        RECT 1999.365 1111.790 2004.495 1112.700 ;
        RECT 2004.895 1111.875 2005.325 1112.660 ;
        RECT 2005.345 1111.790 2010.475 1112.700 ;
        RECT 2010.875 1111.875 2011.305 1112.660 ;
        RECT 2011.325 1111.790 2016.455 1112.700 ;
        RECT 2016.855 1111.875 2017.285 1112.660 ;
        RECT 2017.305 1111.790 2022.435 1112.700 ;
        RECT 2022.835 1111.875 2023.265 1112.660 ;
        RECT 2023.285 1111.790 2028.415 1112.700 ;
        RECT 2028.815 1111.875 2029.245 1112.660 ;
        RECT 2029.265 1111.790 2034.395 1112.700 ;
        RECT 2034.795 1111.875 2035.225 1112.660 ;
        RECT 2035.245 1111.790 2040.375 1112.700 ;
        RECT 2040.775 1111.875 2041.205 1112.660 ;
        RECT 2041.225 1111.790 2046.355 1112.700 ;
        RECT 2046.755 1111.875 2047.185 1112.660 ;
        RECT 2047.205 1111.790 2052.335 1112.700 ;
        RECT 2052.735 1111.875 2053.165 1112.660 ;
        RECT 2053.185 1111.790 2058.315 1112.700 ;
        RECT 2058.715 1111.875 2059.145 1112.660 ;
        RECT 2059.165 1111.790 2064.295 1112.700 ;
        RECT 2064.695 1111.875 2065.125 1112.660 ;
        RECT 2065.525 1111.790 2070.655 1112.700 ;
        RECT 2070.675 1111.875 2071.105 1112.660 ;
        RECT 675.590 1111.600 675.760 1111.790 ;
        RECT 681.570 1111.600 681.740 1111.790 ;
        RECT 687.550 1111.600 687.720 1111.790 ;
        RECT 693.530 1111.600 693.700 1111.790 ;
        RECT 699.510 1111.600 699.680 1111.790 ;
        RECT 705.490 1111.600 705.660 1111.790 ;
        RECT 711.470 1111.600 711.640 1111.790 ;
        RECT 717.450 1111.600 717.620 1111.790 ;
        RECT 723.430 1111.600 723.600 1111.790 ;
        RECT 729.410 1111.600 729.580 1111.790 ;
        RECT 735.390 1111.600 735.560 1111.790 ;
        RECT 741.370 1111.600 741.540 1111.790 ;
        RECT 747.350 1111.600 747.520 1111.790 ;
        RECT 753.330 1111.600 753.500 1111.790 ;
        RECT 759.310 1111.600 759.480 1111.790 ;
        RECT 770.340 1111.600 770.510 1111.790 ;
        RECT 1975.590 1111.600 1975.760 1111.790 ;
        RECT 1981.570 1111.600 1981.740 1111.790 ;
        RECT 1987.550 1111.600 1987.720 1111.790 ;
        RECT 1993.530 1111.600 1993.700 1111.790 ;
        RECT 1999.510 1111.600 1999.680 1111.790 ;
        RECT 2005.490 1111.600 2005.660 1111.790 ;
        RECT 2011.470 1111.600 2011.640 1111.790 ;
        RECT 2017.450 1111.600 2017.620 1111.790 ;
        RECT 2023.430 1111.600 2023.600 1111.790 ;
        RECT 2029.410 1111.600 2029.580 1111.790 ;
        RECT 2035.390 1111.600 2035.560 1111.790 ;
        RECT 2041.370 1111.600 2041.540 1111.790 ;
        RECT 2047.350 1111.600 2047.520 1111.790 ;
        RECT 2053.330 1111.600 2053.500 1111.790 ;
        RECT 2059.310 1111.600 2059.480 1111.790 ;
        RECT 2070.340 1111.600 2070.510 1111.790 ;
      LAYER li1 ;
        RECT 3383.500 3542.415 3383.670 3542.500 ;
        RECT 3386.220 3542.415 3386.390 3542.500 ;
        RECT 3388.940 3542.415 3389.110 3542.500 ;
        RECT 3383.500 3542.355 3384.395 3542.415 ;
        RECT 3383.670 3542.185 3384.395 3542.355 ;
        RECT 3383.500 3542.125 3384.395 3542.185 ;
        RECT 3385.055 3542.355 3387.555 3542.415 ;
        RECT 3385.055 3542.185 3386.220 3542.355 ;
        RECT 3386.390 3542.185 3387.555 3542.355 ;
        RECT 3385.055 3542.125 3387.555 3542.185 ;
        RECT 3388.215 3542.355 3389.110 3542.415 ;
        RECT 3388.215 3542.185 3388.940 3542.355 ;
        RECT 3388.215 3542.125 3389.110 3542.185 ;
        RECT 3383.500 3541.895 3383.670 3542.125 ;
        RECT 3383.500 3541.525 3383.670 3541.725 ;
        RECT 3383.840 3541.695 3384.490 3541.865 ;
        RECT 3383.500 3541.435 3384.150 3541.525 ;
        RECT 3383.670 3541.265 3384.150 3541.435 ;
        RECT 3383.500 3541.195 3384.150 3541.265 ;
        RECT 3383.500 3540.975 3383.670 3541.195 ;
        RECT 3384.320 3541.025 3384.490 3541.695 ;
        RECT 3383.845 3540.855 3384.490 3541.025 ;
        RECT 3383.500 3540.685 3383.670 3540.805 ;
        RECT 3383.500 3540.515 3384.150 3540.685 ;
        RECT 3383.670 3540.355 3384.150 3540.515 ;
        RECT 3384.320 3540.620 3384.490 3540.855 ;
        RECT 3385.030 3541.615 3386.050 3541.945 ;
        RECT 3386.220 3541.895 3386.390 3542.125 ;
        RECT 3388.940 3541.895 3389.110 3542.125 ;
        RECT 3385.030 3541.105 3385.200 3541.615 ;
        RECT 3386.220 3541.565 3386.390 3541.725 ;
        RECT 3388.940 3541.565 3389.110 3541.725 ;
        RECT 3386.220 3541.445 3387.540 3541.565 ;
        RECT 3385.420 3541.435 3387.540 3541.445 ;
        RECT 3385.420 3541.275 3386.220 3541.435 ;
        RECT 3386.390 3541.265 3387.540 3541.435 ;
        RECT 3386.220 3541.235 3387.540 3541.265 ;
        RECT 3388.140 3541.435 3389.110 3541.565 ;
        RECT 3388.140 3541.265 3388.940 3541.435 ;
        RECT 3388.140 3541.235 3389.110 3541.265 ;
        RECT 3385.030 3540.775 3386.050 3541.105 ;
        RECT 3386.220 3540.975 3386.390 3541.235 ;
        RECT 3388.940 3540.975 3389.110 3541.235 ;
        RECT 3385.030 3540.620 3385.200 3540.775 ;
        RECT 3384.320 3540.445 3385.200 3540.620 ;
        RECT 3386.220 3540.725 3386.390 3540.805 ;
        RECT 3388.940 3540.725 3389.110 3540.805 ;
        RECT 3386.220 3540.605 3387.190 3540.725 ;
        RECT 3385.420 3540.515 3387.190 3540.605 ;
        RECT 3383.500 3540.055 3383.670 3540.345 ;
      LAYER li1 ;
        RECT 3383.840 3540.015 3384.490 3540.185 ;
      LAYER li1 ;
        RECT 3383.500 3539.845 3383.670 3539.885 ;
        RECT 3383.500 3539.595 3384.150 3539.845 ;
        RECT 3383.670 3539.515 3384.150 3539.595 ;
        RECT 3383.500 3539.135 3383.670 3539.425 ;
      LAYER li1 ;
        RECT 3384.320 3539.345 3384.490 3540.015 ;
        RECT 3383.840 3539.175 3384.490 3539.345 ;
      LAYER li1 ;
        RECT 3383.670 3538.965 3384.150 3539.005 ;
        RECT 3383.500 3538.675 3384.150 3538.965 ;
      LAYER li1 ;
        RECT 3384.320 3538.505 3384.490 3539.175 ;
      LAYER li1 ;
        RECT 3383.500 3538.215 3383.670 3538.505 ;
      LAYER li1 ;
        RECT 3383.840 3538.335 3384.490 3538.505 ;
      LAYER li1 ;
        RECT 3383.670 3538.045 3384.150 3538.165 ;
        RECT 3383.500 3537.835 3384.150 3538.045 ;
        RECT 3383.500 3537.755 3383.670 3537.835 ;
      LAYER li1 ;
        RECT 3384.320 3537.750 3384.490 3538.335 ;
      LAYER li1 ;
        RECT 3384.660 3537.995 3384.830 3540.445 ;
        RECT 3385.420 3540.435 3386.220 3540.515 ;
        RECT 3386.390 3540.395 3387.190 3540.515 ;
      LAYER li1 ;
        RECT 3385.030 3540.015 3386.050 3540.185 ;
      LAYER li1 ;
        RECT 3386.220 3540.055 3386.390 3540.345 ;
      LAYER li1 ;
        RECT 3385.030 3539.345 3385.200 3540.015 ;
      LAYER li1 ;
        RECT 3386.220 3539.845 3387.190 3539.885 ;
        RECT 3385.420 3539.595 3387.190 3539.845 ;
        RECT 3385.420 3539.515 3386.220 3539.595 ;
        RECT 3386.390 3539.555 3387.190 3539.595 ;
      LAYER li1 ;
        RECT 3385.030 3539.175 3386.050 3539.345 ;
        RECT 3385.030 3538.505 3385.200 3539.175 ;
      LAYER li1 ;
        RECT 3386.220 3539.135 3386.390 3539.425 ;
        RECT 3385.420 3538.965 3386.220 3539.005 ;
        RECT 3386.390 3538.965 3387.190 3539.045 ;
        RECT 3385.420 3538.715 3387.190 3538.965 ;
        RECT 3385.420 3538.675 3386.390 3538.715 ;
      LAYER li1 ;
        RECT 3385.030 3538.335 3386.050 3538.505 ;
        RECT 3385.030 3537.750 3385.200 3538.335 ;
      LAYER li1 ;
        RECT 3386.220 3538.215 3386.390 3538.505 ;
        RECT 3385.420 3538.045 3386.220 3538.165 ;
        RECT 3386.390 3538.045 3387.190 3538.125 ;
        RECT 3387.780 3538.115 3387.950 3540.565 ;
        RECT 3388.460 3540.515 3389.110 3540.725 ;
        RECT 3388.460 3540.395 3388.940 3540.515 ;
        RECT 3388.940 3540.055 3389.110 3540.345 ;
        RECT 3388.460 3539.595 3389.110 3539.885 ;
        RECT 3388.460 3539.555 3388.940 3539.595 ;
        RECT 3388.940 3539.135 3389.110 3539.425 ;
        RECT 3388.460 3538.965 3388.940 3539.045 ;
        RECT 3388.460 3538.715 3389.110 3538.965 ;
        RECT 3388.940 3538.675 3389.110 3538.715 ;
        RECT 3388.940 3538.215 3389.110 3538.505 ;
        RECT 3385.420 3537.955 3387.190 3538.045 ;
        RECT 3385.420 3537.835 3386.390 3537.955 ;
        RECT 3386.220 3537.755 3386.390 3537.835 ;
        RECT 3387.410 3537.940 3388.290 3538.115 ;
        RECT 3387.410 3537.785 3387.580 3537.940 ;
      LAYER li1 ;
        RECT 3384.320 3537.665 3385.200 3537.750 ;
      LAYER li1 ;
        RECT 3383.500 3537.325 3383.670 3537.585 ;
      LAYER li1 ;
        RECT 3383.840 3537.495 3386.050 3537.665 ;
      LAYER li1 ;
        RECT 3386.220 3537.325 3386.390 3537.585 ;
        RECT 3386.560 3537.455 3387.580 3537.785 ;
        RECT 3383.500 3537.295 3384.470 3537.325 ;
        RECT 3383.670 3537.125 3384.470 3537.295 ;
        RECT 3383.500 3536.995 3384.470 3537.125 ;
        RECT 3385.070 3537.295 3386.390 3537.325 ;
        RECT 3385.070 3537.125 3386.220 3537.295 ;
        RECT 3386.390 3537.125 3387.190 3537.285 ;
        RECT 3385.070 3537.115 3387.190 3537.125 ;
        RECT 3385.070 3536.995 3386.390 3537.115 ;
        RECT 3383.500 3536.835 3383.670 3536.995 ;
        RECT 3386.220 3536.835 3386.390 3536.995 ;
        RECT 3387.410 3536.945 3387.580 3537.455 ;
        RECT 3383.500 3536.435 3383.670 3536.665 ;
        RECT 3386.220 3536.435 3386.390 3536.665 ;
        RECT 3386.560 3536.615 3387.580 3536.945 ;
      LAYER li1 ;
        RECT 3387.750 3536.660 3387.950 3537.760 ;
      LAYER li1 ;
        RECT 3388.120 3537.705 3388.290 3537.940 ;
        RECT 3388.460 3538.045 3388.940 3538.205 ;
        RECT 3388.460 3537.875 3389.110 3538.045 ;
        RECT 3388.940 3537.755 3389.110 3537.875 ;
        RECT 3388.120 3537.535 3388.765 3537.705 ;
        RECT 3388.120 3536.865 3388.290 3537.535 ;
        RECT 3388.940 3537.365 3389.110 3537.585 ;
        RECT 3388.460 3537.295 3389.110 3537.365 ;
        RECT 3388.460 3537.125 3388.940 3537.295 ;
        RECT 3388.460 3537.035 3389.110 3537.125 ;
        RECT 3388.120 3536.695 3388.770 3536.865 ;
        RECT 3388.940 3536.835 3389.110 3537.035 ;
        RECT 3388.940 3536.435 3389.110 3536.665 ;
        RECT 3383.500 3536.375 3384.395 3536.435 ;
        RECT 3383.670 3536.205 3384.395 3536.375 ;
        RECT 3383.500 3536.145 3384.395 3536.205 ;
        RECT 3385.055 3536.375 3387.555 3536.435 ;
        RECT 3385.055 3536.205 3386.220 3536.375 ;
        RECT 3386.390 3536.205 3387.555 3536.375 ;
        RECT 3385.055 3536.145 3387.555 3536.205 ;
        RECT 3388.215 3536.375 3389.110 3536.435 ;
        RECT 3388.215 3536.205 3388.940 3536.375 ;
        RECT 3388.215 3536.145 3389.110 3536.205 ;
        RECT 3383.500 3536.060 3383.670 3536.145 ;
        RECT 3386.220 3536.060 3386.390 3536.145 ;
        RECT 3388.940 3536.060 3389.110 3536.145 ;
        RECT 198.685 3023.985 198.855 3024.070 ;
        RECT 201.405 3023.985 201.575 3024.070 ;
        RECT 204.125 3023.985 204.295 3024.070 ;
        RECT 198.685 3023.925 199.580 3023.985 ;
        RECT 198.855 3023.755 199.580 3023.925 ;
        RECT 198.685 3023.695 199.580 3023.755 ;
        RECT 200.240 3023.925 202.740 3023.985 ;
        RECT 200.240 3023.755 201.405 3023.925 ;
        RECT 201.575 3023.755 202.740 3023.925 ;
        RECT 200.240 3023.695 202.740 3023.755 ;
        RECT 203.400 3023.925 204.295 3023.985 ;
        RECT 203.400 3023.755 204.125 3023.925 ;
        RECT 203.400 3023.695 204.295 3023.755 ;
        RECT 198.685 3023.465 198.855 3023.695 ;
        RECT 201.405 3023.465 201.575 3023.695 ;
        RECT 198.685 3023.135 198.855 3023.295 ;
        RECT 201.405 3023.135 201.575 3023.295 ;
        RECT 201.745 3023.185 202.765 3023.515 ;
        RECT 204.125 3023.465 204.295 3023.695 ;
        RECT 198.685 3023.005 199.655 3023.135 ;
        RECT 198.855 3022.835 199.655 3023.005 ;
        RECT 198.685 3022.805 199.655 3022.835 ;
        RECT 200.255 3023.015 201.575 3023.135 ;
        RECT 200.255 3023.005 202.375 3023.015 ;
        RECT 200.255 3022.835 201.405 3023.005 ;
        RECT 201.575 3022.845 202.375 3023.005 ;
        RECT 200.255 3022.805 201.575 3022.835 ;
        RECT 198.685 3022.545 198.855 3022.805 ;
        RECT 201.405 3022.545 201.575 3022.805 ;
        RECT 202.595 3022.675 202.765 3023.185 ;
        RECT 198.685 3022.295 198.855 3022.375 ;
        RECT 201.405 3022.295 201.575 3022.375 ;
        RECT 201.745 3022.345 202.765 3022.675 ;
        RECT 198.685 3022.085 199.335 3022.295 ;
        RECT 200.605 3022.175 201.575 3022.295 ;
        RECT 202.595 3022.190 202.765 3022.345 ;
        RECT 203.305 3023.265 203.955 3023.435 ;
        RECT 203.305 3022.595 203.475 3023.265 ;
        RECT 204.125 3023.095 204.295 3023.295 ;
        RECT 203.645 3023.005 204.295 3023.095 ;
        RECT 203.645 3022.835 204.125 3023.005 ;
        RECT 203.645 3022.765 204.295 3022.835 ;
        RECT 203.305 3022.425 203.950 3022.595 ;
        RECT 204.125 3022.545 204.295 3022.765 ;
        RECT 203.305 3022.190 203.475 3022.425 ;
        RECT 204.125 3022.255 204.295 3022.375 ;
        RECT 198.855 3021.965 199.335 3022.085 ;
        RECT 198.685 3021.625 198.855 3021.915 ;
        RECT 198.685 3021.165 199.335 3021.455 ;
        RECT 198.855 3021.125 199.335 3021.165 ;
        RECT 198.685 3020.705 198.855 3020.995 ;
        RECT 198.855 3020.535 199.335 3020.615 ;
        RECT 198.685 3020.285 199.335 3020.535 ;
        RECT 198.685 3020.245 198.855 3020.285 ;
        RECT 198.685 3019.785 198.855 3020.075 ;
        RECT 198.855 3019.615 199.335 3019.775 ;
        RECT 199.845 3019.685 200.015 3022.135 ;
        RECT 200.605 3022.085 202.375 3022.175 ;
        RECT 200.605 3021.965 201.405 3022.085 ;
        RECT 201.575 3022.005 202.375 3022.085 ;
        RECT 202.595 3022.015 203.475 3022.190 ;
        RECT 203.645 3022.085 204.295 3022.255 ;
        RECT 201.405 3021.625 201.575 3021.915 ;
      LAYER li1 ;
        RECT 201.745 3021.585 202.765 3021.755 ;
      LAYER li1 ;
        RECT 200.605 3021.415 201.575 3021.455 ;
        RECT 200.605 3021.165 202.375 3021.415 ;
        RECT 200.605 3021.125 201.405 3021.165 ;
        RECT 201.575 3021.085 202.375 3021.165 ;
        RECT 201.405 3020.705 201.575 3020.995 ;
      LAYER li1 ;
        RECT 202.595 3020.915 202.765 3021.585 ;
        RECT 201.745 3020.745 202.765 3020.915 ;
      LAYER li1 ;
        RECT 200.605 3020.535 201.405 3020.615 ;
        RECT 201.575 3020.535 202.375 3020.575 ;
        RECT 200.605 3020.285 202.375 3020.535 ;
        RECT 201.405 3020.245 202.375 3020.285 ;
      LAYER li1 ;
        RECT 202.595 3020.075 202.765 3020.745 ;
      LAYER li1 ;
        RECT 201.405 3019.785 201.575 3020.075 ;
      LAYER li1 ;
        RECT 201.745 3019.905 202.765 3020.075 ;
      LAYER li1 ;
        RECT 198.685 3019.445 199.335 3019.615 ;
        RECT 199.505 3019.510 200.385 3019.685 ;
        RECT 200.605 3019.615 201.405 3019.695 ;
        RECT 201.575 3019.615 202.375 3019.735 ;
        RECT 200.605 3019.525 202.375 3019.615 ;
        RECT 198.685 3019.325 198.855 3019.445 ;
        RECT 199.505 3019.275 199.675 3019.510 ;
        RECT 200.215 3019.355 200.385 3019.510 ;
        RECT 201.405 3019.405 202.375 3019.525 ;
        RECT 198.685 3018.935 198.855 3019.155 ;
        RECT 199.030 3019.105 199.675 3019.275 ;
        RECT 198.685 3018.865 199.335 3018.935 ;
        RECT 198.855 3018.695 199.335 3018.865 ;
        RECT 198.685 3018.605 199.335 3018.695 ;
        RECT 198.685 3018.405 198.855 3018.605 ;
        RECT 199.505 3018.435 199.675 3019.105 ;
        RECT 199.025 3018.265 199.675 3018.435 ;
        RECT 198.685 3018.005 198.855 3018.235 ;
      LAYER li1 ;
        RECT 199.845 3018.230 200.045 3019.330 ;
      LAYER li1 ;
        RECT 200.215 3019.025 201.235 3019.355 ;
        RECT 201.405 3019.325 201.575 3019.405 ;
      LAYER li1 ;
        RECT 202.595 3019.320 202.765 3019.905 ;
      LAYER li1 ;
        RECT 202.965 3019.565 203.135 3022.015 ;
        RECT 203.645 3021.925 204.125 3022.085 ;
      LAYER li1 ;
        RECT 203.305 3021.585 203.955 3021.755 ;
      LAYER li1 ;
        RECT 204.125 3021.625 204.295 3021.915 ;
      LAYER li1 ;
        RECT 203.305 3020.915 203.475 3021.585 ;
      LAYER li1 ;
        RECT 204.125 3021.415 204.295 3021.455 ;
        RECT 203.645 3021.165 204.295 3021.415 ;
        RECT 203.645 3021.085 204.125 3021.165 ;
      LAYER li1 ;
        RECT 203.305 3020.745 203.955 3020.915 ;
        RECT 203.305 3020.075 203.475 3020.745 ;
      LAYER li1 ;
        RECT 204.125 3020.705 204.295 3020.995 ;
        RECT 203.645 3020.535 204.125 3020.575 ;
        RECT 203.645 3020.245 204.295 3020.535 ;
      LAYER li1 ;
        RECT 203.305 3019.905 203.955 3020.075 ;
        RECT 203.305 3019.320 203.475 3019.905 ;
      LAYER li1 ;
        RECT 204.125 3019.785 204.295 3020.075 ;
        RECT 203.645 3019.615 204.125 3019.735 ;
        RECT 203.645 3019.405 204.295 3019.615 ;
        RECT 204.125 3019.325 204.295 3019.405 ;
      LAYER li1 ;
        RECT 202.595 3019.235 203.475 3019.320 ;
      LAYER li1 ;
        RECT 200.215 3018.515 200.385 3019.025 ;
        RECT 201.405 3018.895 201.575 3019.155 ;
      LAYER li1 ;
        RECT 201.745 3019.065 203.955 3019.235 ;
      LAYER li1 ;
        RECT 204.125 3018.895 204.295 3019.155 ;
        RECT 201.405 3018.865 202.725 3018.895 ;
        RECT 200.605 3018.695 201.405 3018.855 ;
        RECT 201.575 3018.695 202.725 3018.865 ;
        RECT 200.605 3018.685 202.725 3018.695 ;
        RECT 201.405 3018.565 202.725 3018.685 ;
        RECT 203.325 3018.865 204.295 3018.895 ;
        RECT 203.325 3018.695 204.125 3018.865 ;
        RECT 203.325 3018.565 204.295 3018.695 ;
        RECT 200.215 3018.185 201.235 3018.515 ;
        RECT 201.405 3018.405 201.575 3018.565 ;
        RECT 204.125 3018.405 204.295 3018.565 ;
        RECT 201.405 3018.005 201.575 3018.235 ;
        RECT 204.125 3018.005 204.295 3018.235 ;
        RECT 198.685 3017.945 199.580 3018.005 ;
        RECT 198.855 3017.775 199.580 3017.945 ;
        RECT 198.685 3017.715 199.580 3017.775 ;
        RECT 200.240 3017.945 202.740 3018.005 ;
        RECT 200.240 3017.775 201.405 3017.945 ;
        RECT 201.575 3017.775 202.740 3017.945 ;
        RECT 200.240 3017.715 202.740 3017.775 ;
        RECT 203.400 3017.945 204.295 3018.005 ;
        RECT 203.400 3017.775 204.125 3017.945 ;
        RECT 203.400 3017.715 204.295 3017.775 ;
        RECT 198.685 3017.485 198.855 3017.715 ;
        RECT 201.405 3017.485 201.575 3017.715 ;
        RECT 198.685 3017.155 198.855 3017.315 ;
        RECT 201.405 3017.155 201.575 3017.315 ;
        RECT 201.745 3017.205 202.765 3017.535 ;
        RECT 204.125 3017.485 204.295 3017.715 ;
        RECT 198.685 3017.025 199.655 3017.155 ;
        RECT 198.855 3016.855 199.655 3017.025 ;
        RECT 198.685 3016.825 199.655 3016.855 ;
        RECT 200.255 3017.035 201.575 3017.155 ;
        RECT 200.255 3017.025 202.375 3017.035 ;
        RECT 200.255 3016.855 201.405 3017.025 ;
        RECT 201.575 3016.865 202.375 3017.025 ;
        RECT 200.255 3016.825 201.575 3016.855 ;
        RECT 198.685 3016.565 198.855 3016.825 ;
        RECT 201.405 3016.565 201.575 3016.825 ;
        RECT 202.595 3016.695 202.765 3017.205 ;
        RECT 198.685 3016.315 198.855 3016.395 ;
        RECT 201.405 3016.315 201.575 3016.395 ;
        RECT 201.745 3016.365 202.765 3016.695 ;
        RECT 198.685 3016.105 199.335 3016.315 ;
        RECT 200.605 3016.195 201.575 3016.315 ;
        RECT 202.595 3016.210 202.765 3016.365 ;
        RECT 203.305 3017.285 203.955 3017.455 ;
        RECT 203.305 3016.615 203.475 3017.285 ;
        RECT 204.125 3017.115 204.295 3017.315 ;
        RECT 203.645 3017.025 204.295 3017.115 ;
        RECT 203.645 3016.855 204.125 3017.025 ;
        RECT 203.645 3016.785 204.295 3016.855 ;
        RECT 203.305 3016.445 203.950 3016.615 ;
        RECT 204.125 3016.565 204.295 3016.785 ;
        RECT 203.305 3016.210 203.475 3016.445 ;
        RECT 204.125 3016.275 204.295 3016.395 ;
        RECT 198.855 3015.985 199.335 3016.105 ;
        RECT 198.685 3015.645 198.855 3015.935 ;
        RECT 198.685 3015.185 199.335 3015.475 ;
        RECT 198.855 3015.145 199.335 3015.185 ;
        RECT 198.685 3014.725 198.855 3015.015 ;
        RECT 198.855 3014.555 199.335 3014.635 ;
        RECT 198.685 3014.305 199.335 3014.555 ;
        RECT 198.685 3014.265 198.855 3014.305 ;
        RECT 198.685 3013.805 198.855 3014.095 ;
        RECT 198.855 3013.635 199.335 3013.795 ;
        RECT 199.845 3013.705 200.015 3016.155 ;
        RECT 200.605 3016.105 202.375 3016.195 ;
        RECT 200.605 3015.985 201.405 3016.105 ;
        RECT 201.575 3016.025 202.375 3016.105 ;
        RECT 202.595 3016.035 203.475 3016.210 ;
        RECT 203.645 3016.105 204.295 3016.275 ;
        RECT 201.405 3015.645 201.575 3015.935 ;
      LAYER li1 ;
        RECT 201.745 3015.605 202.765 3015.775 ;
      LAYER li1 ;
        RECT 200.605 3015.435 201.575 3015.475 ;
        RECT 200.605 3015.185 202.375 3015.435 ;
        RECT 200.605 3015.145 201.405 3015.185 ;
        RECT 201.575 3015.105 202.375 3015.185 ;
        RECT 201.405 3014.725 201.575 3015.015 ;
      LAYER li1 ;
        RECT 202.595 3014.935 202.765 3015.605 ;
        RECT 201.745 3014.765 202.765 3014.935 ;
      LAYER li1 ;
        RECT 200.605 3014.555 201.405 3014.635 ;
        RECT 201.575 3014.555 202.375 3014.595 ;
        RECT 200.605 3014.305 202.375 3014.555 ;
        RECT 201.405 3014.265 202.375 3014.305 ;
      LAYER li1 ;
        RECT 202.595 3014.095 202.765 3014.765 ;
      LAYER li1 ;
        RECT 201.405 3013.805 201.575 3014.095 ;
      LAYER li1 ;
        RECT 201.745 3013.925 202.765 3014.095 ;
      LAYER li1 ;
        RECT 198.685 3013.465 199.335 3013.635 ;
        RECT 199.505 3013.530 200.385 3013.705 ;
        RECT 200.605 3013.635 201.405 3013.715 ;
        RECT 201.575 3013.635 202.375 3013.755 ;
        RECT 200.605 3013.545 202.375 3013.635 ;
        RECT 198.685 3013.345 198.855 3013.465 ;
        RECT 199.505 3013.295 199.675 3013.530 ;
        RECT 200.215 3013.375 200.385 3013.530 ;
        RECT 201.405 3013.425 202.375 3013.545 ;
        RECT 198.685 3012.955 198.855 3013.175 ;
        RECT 199.030 3013.125 199.675 3013.295 ;
        RECT 198.685 3012.885 199.335 3012.955 ;
        RECT 198.855 3012.715 199.335 3012.885 ;
        RECT 198.685 3012.625 199.335 3012.715 ;
        RECT 198.685 3012.425 198.855 3012.625 ;
        RECT 199.505 3012.455 199.675 3013.125 ;
        RECT 199.025 3012.285 199.675 3012.455 ;
        RECT 198.685 3012.025 198.855 3012.255 ;
      LAYER li1 ;
        RECT 199.845 3012.250 200.045 3013.350 ;
      LAYER li1 ;
        RECT 200.215 3013.045 201.235 3013.375 ;
        RECT 201.405 3013.345 201.575 3013.425 ;
      LAYER li1 ;
        RECT 202.595 3013.340 202.765 3013.925 ;
      LAYER li1 ;
        RECT 202.965 3013.585 203.135 3016.035 ;
        RECT 203.645 3015.945 204.125 3016.105 ;
      LAYER li1 ;
        RECT 203.305 3015.605 203.955 3015.775 ;
      LAYER li1 ;
        RECT 204.125 3015.645 204.295 3015.935 ;
      LAYER li1 ;
        RECT 203.305 3014.935 203.475 3015.605 ;
      LAYER li1 ;
        RECT 204.125 3015.435 204.295 3015.475 ;
        RECT 203.645 3015.185 204.295 3015.435 ;
        RECT 203.645 3015.105 204.125 3015.185 ;
      LAYER li1 ;
        RECT 203.305 3014.765 203.955 3014.935 ;
        RECT 203.305 3014.095 203.475 3014.765 ;
      LAYER li1 ;
        RECT 204.125 3014.725 204.295 3015.015 ;
        RECT 203.645 3014.555 204.125 3014.595 ;
        RECT 203.645 3014.265 204.295 3014.555 ;
      LAYER li1 ;
        RECT 203.305 3013.925 203.955 3014.095 ;
        RECT 203.305 3013.340 203.475 3013.925 ;
      LAYER li1 ;
        RECT 204.125 3013.805 204.295 3014.095 ;
        RECT 203.645 3013.635 204.125 3013.755 ;
        RECT 203.645 3013.425 204.295 3013.635 ;
        RECT 204.125 3013.345 204.295 3013.425 ;
      LAYER li1 ;
        RECT 202.595 3013.255 203.475 3013.340 ;
      LAYER li1 ;
        RECT 200.215 3012.535 200.385 3013.045 ;
        RECT 201.405 3012.915 201.575 3013.175 ;
      LAYER li1 ;
        RECT 201.745 3013.085 203.955 3013.255 ;
      LAYER li1 ;
        RECT 204.125 3012.915 204.295 3013.175 ;
        RECT 201.405 3012.885 202.725 3012.915 ;
        RECT 200.605 3012.715 201.405 3012.875 ;
        RECT 201.575 3012.715 202.725 3012.885 ;
        RECT 200.605 3012.705 202.725 3012.715 ;
        RECT 201.405 3012.585 202.725 3012.705 ;
        RECT 203.325 3012.885 204.295 3012.915 ;
        RECT 203.325 3012.715 204.125 3012.885 ;
        RECT 203.325 3012.585 204.295 3012.715 ;
        RECT 200.215 3012.205 201.235 3012.535 ;
        RECT 201.405 3012.425 201.575 3012.585 ;
        RECT 204.125 3012.425 204.295 3012.585 ;
        RECT 201.405 3012.025 201.575 3012.255 ;
        RECT 204.125 3012.025 204.295 3012.255 ;
        RECT 198.685 3011.965 199.580 3012.025 ;
        RECT 198.855 3011.795 199.580 3011.965 ;
        RECT 198.685 3011.735 199.580 3011.795 ;
        RECT 200.240 3011.965 202.740 3012.025 ;
        RECT 200.240 3011.795 201.405 3011.965 ;
        RECT 201.575 3011.795 202.740 3011.965 ;
        RECT 200.240 3011.735 202.740 3011.795 ;
        RECT 203.400 3011.965 204.295 3012.025 ;
        RECT 203.400 3011.795 204.125 3011.965 ;
        RECT 203.400 3011.735 204.295 3011.795 ;
        RECT 198.685 3011.505 198.855 3011.735 ;
        RECT 201.405 3011.505 201.575 3011.735 ;
        RECT 198.685 3011.175 198.855 3011.335 ;
        RECT 201.405 3011.175 201.575 3011.335 ;
        RECT 201.745 3011.225 202.765 3011.555 ;
        RECT 204.125 3011.505 204.295 3011.735 ;
        RECT 198.685 3011.045 199.655 3011.175 ;
        RECT 198.855 3010.875 199.655 3011.045 ;
        RECT 198.685 3010.845 199.655 3010.875 ;
        RECT 200.255 3011.055 201.575 3011.175 ;
        RECT 200.255 3011.045 202.375 3011.055 ;
        RECT 200.255 3010.875 201.405 3011.045 ;
        RECT 201.575 3010.885 202.375 3011.045 ;
        RECT 200.255 3010.845 201.575 3010.875 ;
        RECT 198.685 3010.585 198.855 3010.845 ;
        RECT 201.405 3010.585 201.575 3010.845 ;
        RECT 202.595 3010.715 202.765 3011.225 ;
        RECT 198.685 3010.335 198.855 3010.415 ;
        RECT 201.405 3010.335 201.575 3010.415 ;
        RECT 201.745 3010.385 202.765 3010.715 ;
        RECT 198.685 3010.125 199.335 3010.335 ;
        RECT 200.605 3010.215 201.575 3010.335 ;
        RECT 202.595 3010.230 202.765 3010.385 ;
        RECT 203.305 3011.305 203.955 3011.475 ;
        RECT 203.305 3010.635 203.475 3011.305 ;
        RECT 204.125 3011.135 204.295 3011.335 ;
        RECT 203.645 3011.045 204.295 3011.135 ;
        RECT 203.645 3010.875 204.125 3011.045 ;
        RECT 203.645 3010.805 204.295 3010.875 ;
        RECT 203.305 3010.465 203.950 3010.635 ;
        RECT 204.125 3010.585 204.295 3010.805 ;
        RECT 203.305 3010.230 203.475 3010.465 ;
        RECT 204.125 3010.295 204.295 3010.415 ;
        RECT 198.855 3010.005 199.335 3010.125 ;
        RECT 198.685 3009.665 198.855 3009.955 ;
        RECT 198.685 3009.205 199.335 3009.495 ;
        RECT 198.855 3009.165 199.335 3009.205 ;
        RECT 198.685 3008.745 198.855 3009.035 ;
        RECT 198.855 3008.575 199.335 3008.655 ;
        RECT 198.685 3008.325 199.335 3008.575 ;
        RECT 198.685 3008.285 198.855 3008.325 ;
        RECT 198.685 3007.825 198.855 3008.115 ;
        RECT 198.855 3007.655 199.335 3007.815 ;
        RECT 199.845 3007.725 200.015 3010.175 ;
        RECT 200.605 3010.125 202.375 3010.215 ;
        RECT 200.605 3010.005 201.405 3010.125 ;
        RECT 201.575 3010.045 202.375 3010.125 ;
        RECT 202.595 3010.055 203.475 3010.230 ;
        RECT 203.645 3010.125 204.295 3010.295 ;
        RECT 201.405 3009.665 201.575 3009.955 ;
      LAYER li1 ;
        RECT 201.745 3009.625 202.765 3009.795 ;
      LAYER li1 ;
        RECT 200.605 3009.455 201.575 3009.495 ;
        RECT 200.605 3009.205 202.375 3009.455 ;
        RECT 200.605 3009.165 201.405 3009.205 ;
        RECT 201.575 3009.125 202.375 3009.205 ;
        RECT 201.405 3008.745 201.575 3009.035 ;
      LAYER li1 ;
        RECT 202.595 3008.955 202.765 3009.625 ;
        RECT 201.745 3008.785 202.765 3008.955 ;
      LAYER li1 ;
        RECT 200.605 3008.575 201.405 3008.655 ;
        RECT 201.575 3008.575 202.375 3008.615 ;
        RECT 200.605 3008.325 202.375 3008.575 ;
        RECT 201.405 3008.285 202.375 3008.325 ;
      LAYER li1 ;
        RECT 202.595 3008.115 202.765 3008.785 ;
      LAYER li1 ;
        RECT 201.405 3007.825 201.575 3008.115 ;
      LAYER li1 ;
        RECT 201.745 3007.945 202.765 3008.115 ;
      LAYER li1 ;
        RECT 198.685 3007.485 199.335 3007.655 ;
        RECT 199.505 3007.550 200.385 3007.725 ;
        RECT 200.605 3007.655 201.405 3007.735 ;
        RECT 201.575 3007.655 202.375 3007.775 ;
        RECT 200.605 3007.565 202.375 3007.655 ;
        RECT 198.685 3007.365 198.855 3007.485 ;
        RECT 199.505 3007.315 199.675 3007.550 ;
        RECT 200.215 3007.395 200.385 3007.550 ;
        RECT 201.405 3007.445 202.375 3007.565 ;
        RECT 198.685 3006.975 198.855 3007.195 ;
        RECT 199.030 3007.145 199.675 3007.315 ;
        RECT 198.685 3006.905 199.335 3006.975 ;
        RECT 198.855 3006.735 199.335 3006.905 ;
        RECT 198.685 3006.645 199.335 3006.735 ;
        RECT 198.685 3006.445 198.855 3006.645 ;
        RECT 199.505 3006.475 199.675 3007.145 ;
        RECT 199.025 3006.305 199.675 3006.475 ;
        RECT 198.685 3006.045 198.855 3006.275 ;
      LAYER li1 ;
        RECT 199.845 3006.270 200.045 3007.370 ;
      LAYER li1 ;
        RECT 200.215 3007.065 201.235 3007.395 ;
        RECT 201.405 3007.365 201.575 3007.445 ;
      LAYER li1 ;
        RECT 202.595 3007.360 202.765 3007.945 ;
      LAYER li1 ;
        RECT 202.965 3007.605 203.135 3010.055 ;
        RECT 203.645 3009.965 204.125 3010.125 ;
      LAYER li1 ;
        RECT 203.305 3009.625 203.955 3009.795 ;
      LAYER li1 ;
        RECT 204.125 3009.665 204.295 3009.955 ;
      LAYER li1 ;
        RECT 203.305 3008.955 203.475 3009.625 ;
      LAYER li1 ;
        RECT 204.125 3009.455 204.295 3009.495 ;
        RECT 203.645 3009.205 204.295 3009.455 ;
        RECT 203.645 3009.125 204.125 3009.205 ;
      LAYER li1 ;
        RECT 203.305 3008.785 203.955 3008.955 ;
        RECT 203.305 3008.115 203.475 3008.785 ;
      LAYER li1 ;
        RECT 204.125 3008.745 204.295 3009.035 ;
        RECT 203.645 3008.575 204.125 3008.615 ;
        RECT 203.645 3008.285 204.295 3008.575 ;
      LAYER li1 ;
        RECT 203.305 3007.945 203.955 3008.115 ;
        RECT 203.305 3007.360 203.475 3007.945 ;
      LAYER li1 ;
        RECT 204.125 3007.825 204.295 3008.115 ;
        RECT 203.645 3007.655 204.125 3007.775 ;
        RECT 203.645 3007.445 204.295 3007.655 ;
        RECT 204.125 3007.365 204.295 3007.445 ;
      LAYER li1 ;
        RECT 202.595 3007.275 203.475 3007.360 ;
      LAYER li1 ;
        RECT 200.215 3006.555 200.385 3007.065 ;
        RECT 201.405 3006.935 201.575 3007.195 ;
      LAYER li1 ;
        RECT 201.745 3007.105 203.955 3007.275 ;
      LAYER li1 ;
        RECT 204.125 3006.935 204.295 3007.195 ;
        RECT 201.405 3006.905 202.725 3006.935 ;
        RECT 200.605 3006.735 201.405 3006.895 ;
        RECT 201.575 3006.735 202.725 3006.905 ;
        RECT 200.605 3006.725 202.725 3006.735 ;
        RECT 201.405 3006.605 202.725 3006.725 ;
        RECT 203.325 3006.905 204.295 3006.935 ;
        RECT 203.325 3006.735 204.125 3006.905 ;
        RECT 203.325 3006.605 204.295 3006.735 ;
        RECT 200.215 3006.225 201.235 3006.555 ;
        RECT 201.405 3006.445 201.575 3006.605 ;
        RECT 204.125 3006.445 204.295 3006.605 ;
        RECT 201.405 3006.045 201.575 3006.275 ;
        RECT 204.125 3006.045 204.295 3006.275 ;
        RECT 198.685 3005.985 199.580 3006.045 ;
        RECT 198.855 3005.815 199.580 3005.985 ;
        RECT 198.685 3005.755 199.580 3005.815 ;
        RECT 200.240 3005.985 202.740 3006.045 ;
        RECT 200.240 3005.815 201.405 3005.985 ;
        RECT 201.575 3005.815 202.740 3005.985 ;
        RECT 200.240 3005.755 202.740 3005.815 ;
        RECT 203.400 3005.985 204.295 3006.045 ;
        RECT 203.400 3005.815 204.125 3005.985 ;
        RECT 203.400 3005.755 204.295 3005.815 ;
        RECT 198.685 3005.525 198.855 3005.755 ;
        RECT 201.405 3005.525 201.575 3005.755 ;
        RECT 198.685 3005.195 198.855 3005.355 ;
        RECT 201.405 3005.195 201.575 3005.355 ;
        RECT 201.745 3005.245 202.765 3005.575 ;
        RECT 204.125 3005.525 204.295 3005.755 ;
        RECT 198.685 3005.065 199.655 3005.195 ;
        RECT 198.855 3004.895 199.655 3005.065 ;
        RECT 198.685 3004.865 199.655 3004.895 ;
        RECT 200.255 3005.075 201.575 3005.195 ;
        RECT 200.255 3005.065 202.375 3005.075 ;
        RECT 200.255 3004.895 201.405 3005.065 ;
        RECT 201.575 3004.905 202.375 3005.065 ;
        RECT 200.255 3004.865 201.575 3004.895 ;
        RECT 198.685 3004.605 198.855 3004.865 ;
        RECT 201.405 3004.605 201.575 3004.865 ;
        RECT 202.595 3004.735 202.765 3005.245 ;
        RECT 198.685 3004.355 198.855 3004.435 ;
        RECT 201.405 3004.355 201.575 3004.435 ;
        RECT 201.745 3004.405 202.765 3004.735 ;
        RECT 198.685 3004.145 199.335 3004.355 ;
        RECT 200.605 3004.235 201.575 3004.355 ;
        RECT 202.595 3004.250 202.765 3004.405 ;
        RECT 203.305 3005.325 203.955 3005.495 ;
        RECT 203.305 3004.655 203.475 3005.325 ;
        RECT 204.125 3005.155 204.295 3005.355 ;
        RECT 203.645 3005.065 204.295 3005.155 ;
        RECT 203.645 3004.895 204.125 3005.065 ;
        RECT 203.645 3004.825 204.295 3004.895 ;
        RECT 203.305 3004.485 203.950 3004.655 ;
        RECT 204.125 3004.605 204.295 3004.825 ;
        RECT 203.305 3004.250 203.475 3004.485 ;
        RECT 204.125 3004.315 204.295 3004.435 ;
        RECT 198.855 3004.025 199.335 3004.145 ;
        RECT 198.685 3003.685 198.855 3003.975 ;
        RECT 198.685 3003.225 199.335 3003.515 ;
        RECT 198.855 3003.185 199.335 3003.225 ;
        RECT 198.685 3002.765 198.855 3003.055 ;
        RECT 198.855 3002.595 199.335 3002.675 ;
        RECT 198.685 3002.345 199.335 3002.595 ;
        RECT 198.685 3002.305 198.855 3002.345 ;
        RECT 198.685 3001.845 198.855 3002.135 ;
        RECT 198.855 3001.675 199.335 3001.835 ;
        RECT 199.845 3001.745 200.015 3004.195 ;
        RECT 200.605 3004.145 202.375 3004.235 ;
        RECT 200.605 3004.025 201.405 3004.145 ;
        RECT 201.575 3004.065 202.375 3004.145 ;
        RECT 202.595 3004.075 203.475 3004.250 ;
        RECT 203.645 3004.145 204.295 3004.315 ;
        RECT 201.405 3003.685 201.575 3003.975 ;
      LAYER li1 ;
        RECT 201.745 3003.645 202.765 3003.815 ;
      LAYER li1 ;
        RECT 200.605 3003.475 201.575 3003.515 ;
        RECT 200.605 3003.225 202.375 3003.475 ;
        RECT 200.605 3003.185 201.405 3003.225 ;
        RECT 201.575 3003.145 202.375 3003.225 ;
        RECT 201.405 3002.765 201.575 3003.055 ;
      LAYER li1 ;
        RECT 202.595 3002.975 202.765 3003.645 ;
        RECT 201.745 3002.805 202.765 3002.975 ;
      LAYER li1 ;
        RECT 200.605 3002.595 201.405 3002.675 ;
        RECT 201.575 3002.595 202.375 3002.635 ;
        RECT 200.605 3002.345 202.375 3002.595 ;
        RECT 201.405 3002.305 202.375 3002.345 ;
      LAYER li1 ;
        RECT 202.595 3002.135 202.765 3002.805 ;
      LAYER li1 ;
        RECT 201.405 3001.845 201.575 3002.135 ;
      LAYER li1 ;
        RECT 201.745 3001.965 202.765 3002.135 ;
      LAYER li1 ;
        RECT 198.685 3001.505 199.335 3001.675 ;
        RECT 199.505 3001.570 200.385 3001.745 ;
        RECT 200.605 3001.675 201.405 3001.755 ;
        RECT 201.575 3001.675 202.375 3001.795 ;
        RECT 200.605 3001.585 202.375 3001.675 ;
        RECT 198.685 3001.385 198.855 3001.505 ;
        RECT 199.505 3001.335 199.675 3001.570 ;
        RECT 200.215 3001.415 200.385 3001.570 ;
        RECT 201.405 3001.465 202.375 3001.585 ;
        RECT 198.685 3000.995 198.855 3001.215 ;
        RECT 199.030 3001.165 199.675 3001.335 ;
        RECT 198.685 3000.925 199.335 3000.995 ;
        RECT 198.855 3000.755 199.335 3000.925 ;
        RECT 198.685 3000.665 199.335 3000.755 ;
        RECT 198.685 3000.465 198.855 3000.665 ;
        RECT 199.505 3000.495 199.675 3001.165 ;
        RECT 199.025 3000.325 199.675 3000.495 ;
        RECT 198.685 3000.065 198.855 3000.295 ;
      LAYER li1 ;
        RECT 199.845 3000.290 200.045 3001.390 ;
      LAYER li1 ;
        RECT 200.215 3001.085 201.235 3001.415 ;
        RECT 201.405 3001.385 201.575 3001.465 ;
      LAYER li1 ;
        RECT 202.595 3001.380 202.765 3001.965 ;
      LAYER li1 ;
        RECT 202.965 3001.625 203.135 3004.075 ;
        RECT 203.645 3003.985 204.125 3004.145 ;
      LAYER li1 ;
        RECT 203.305 3003.645 203.955 3003.815 ;
      LAYER li1 ;
        RECT 204.125 3003.685 204.295 3003.975 ;
      LAYER li1 ;
        RECT 203.305 3002.975 203.475 3003.645 ;
      LAYER li1 ;
        RECT 204.125 3003.475 204.295 3003.515 ;
        RECT 203.645 3003.225 204.295 3003.475 ;
        RECT 203.645 3003.145 204.125 3003.225 ;
      LAYER li1 ;
        RECT 203.305 3002.805 203.955 3002.975 ;
        RECT 203.305 3002.135 203.475 3002.805 ;
      LAYER li1 ;
        RECT 204.125 3002.765 204.295 3003.055 ;
        RECT 203.645 3002.595 204.125 3002.635 ;
        RECT 203.645 3002.305 204.295 3002.595 ;
      LAYER li1 ;
        RECT 203.305 3001.965 203.955 3002.135 ;
        RECT 203.305 3001.380 203.475 3001.965 ;
      LAYER li1 ;
        RECT 204.125 3001.845 204.295 3002.135 ;
        RECT 203.645 3001.675 204.125 3001.795 ;
        RECT 203.645 3001.465 204.295 3001.675 ;
        RECT 204.125 3001.385 204.295 3001.465 ;
      LAYER li1 ;
        RECT 202.595 3001.295 203.475 3001.380 ;
      LAYER li1 ;
        RECT 200.215 3000.575 200.385 3001.085 ;
        RECT 201.405 3000.955 201.575 3001.215 ;
      LAYER li1 ;
        RECT 201.745 3001.125 203.955 3001.295 ;
      LAYER li1 ;
        RECT 204.125 3000.955 204.295 3001.215 ;
        RECT 201.405 3000.925 202.725 3000.955 ;
        RECT 200.605 3000.755 201.405 3000.915 ;
        RECT 201.575 3000.755 202.725 3000.925 ;
        RECT 200.605 3000.745 202.725 3000.755 ;
        RECT 201.405 3000.625 202.725 3000.745 ;
        RECT 203.325 3000.925 204.295 3000.955 ;
        RECT 203.325 3000.755 204.125 3000.925 ;
        RECT 203.325 3000.625 204.295 3000.755 ;
        RECT 200.215 3000.245 201.235 3000.575 ;
        RECT 201.405 3000.465 201.575 3000.625 ;
        RECT 204.125 3000.465 204.295 3000.625 ;
        RECT 201.405 3000.065 201.575 3000.295 ;
        RECT 204.125 3000.065 204.295 3000.295 ;
        RECT 198.685 3000.005 199.580 3000.065 ;
        RECT 198.855 2999.835 199.580 3000.005 ;
        RECT 198.685 2999.775 199.580 2999.835 ;
        RECT 200.240 3000.005 202.740 3000.065 ;
        RECT 200.240 2999.835 201.405 3000.005 ;
        RECT 201.575 2999.835 202.740 3000.005 ;
        RECT 200.240 2999.775 202.740 2999.835 ;
        RECT 203.400 3000.005 204.295 3000.065 ;
        RECT 203.400 2999.835 204.125 3000.005 ;
        RECT 203.400 2999.775 204.295 2999.835 ;
        RECT 198.685 2999.545 198.855 2999.775 ;
        RECT 201.405 2999.545 201.575 2999.775 ;
        RECT 198.685 2999.215 198.855 2999.375 ;
        RECT 201.405 2999.215 201.575 2999.375 ;
        RECT 201.745 2999.265 202.765 2999.595 ;
        RECT 204.125 2999.545 204.295 2999.775 ;
        RECT 198.685 2999.085 199.655 2999.215 ;
        RECT 198.855 2998.915 199.655 2999.085 ;
        RECT 198.685 2998.885 199.655 2998.915 ;
        RECT 200.255 2999.095 201.575 2999.215 ;
        RECT 200.255 2999.085 202.375 2999.095 ;
        RECT 200.255 2998.915 201.405 2999.085 ;
        RECT 201.575 2998.925 202.375 2999.085 ;
        RECT 200.255 2998.885 201.575 2998.915 ;
        RECT 198.685 2998.625 198.855 2998.885 ;
        RECT 201.405 2998.625 201.575 2998.885 ;
        RECT 202.595 2998.755 202.765 2999.265 ;
        RECT 198.685 2998.375 198.855 2998.455 ;
        RECT 201.405 2998.375 201.575 2998.455 ;
        RECT 201.745 2998.425 202.765 2998.755 ;
        RECT 198.685 2998.165 199.335 2998.375 ;
        RECT 200.605 2998.255 201.575 2998.375 ;
        RECT 202.595 2998.270 202.765 2998.425 ;
        RECT 203.305 2999.345 203.955 2999.515 ;
        RECT 203.305 2998.675 203.475 2999.345 ;
        RECT 204.125 2999.175 204.295 2999.375 ;
        RECT 203.645 2999.085 204.295 2999.175 ;
        RECT 203.645 2998.915 204.125 2999.085 ;
        RECT 203.645 2998.845 204.295 2998.915 ;
        RECT 203.305 2998.505 203.950 2998.675 ;
        RECT 204.125 2998.625 204.295 2998.845 ;
        RECT 203.305 2998.270 203.475 2998.505 ;
        RECT 204.125 2998.335 204.295 2998.455 ;
        RECT 198.855 2998.045 199.335 2998.165 ;
        RECT 198.685 2997.705 198.855 2997.995 ;
        RECT 198.685 2997.245 199.335 2997.535 ;
        RECT 198.855 2997.205 199.335 2997.245 ;
        RECT 198.685 2996.785 198.855 2997.075 ;
        RECT 198.855 2996.615 199.335 2996.695 ;
        RECT 198.685 2996.365 199.335 2996.615 ;
        RECT 198.685 2996.325 198.855 2996.365 ;
        RECT 198.685 2995.865 198.855 2996.155 ;
        RECT 198.855 2995.695 199.335 2995.855 ;
        RECT 199.845 2995.765 200.015 2998.215 ;
        RECT 200.605 2998.165 202.375 2998.255 ;
        RECT 200.605 2998.045 201.405 2998.165 ;
        RECT 201.575 2998.085 202.375 2998.165 ;
        RECT 202.595 2998.095 203.475 2998.270 ;
        RECT 203.645 2998.165 204.295 2998.335 ;
        RECT 201.405 2997.705 201.575 2997.995 ;
      LAYER li1 ;
        RECT 201.745 2997.665 202.765 2997.835 ;
      LAYER li1 ;
        RECT 200.605 2997.495 201.575 2997.535 ;
        RECT 200.605 2997.245 202.375 2997.495 ;
        RECT 200.605 2997.205 201.405 2997.245 ;
        RECT 201.575 2997.165 202.375 2997.245 ;
        RECT 201.405 2996.785 201.575 2997.075 ;
      LAYER li1 ;
        RECT 202.595 2996.995 202.765 2997.665 ;
        RECT 201.745 2996.825 202.765 2996.995 ;
      LAYER li1 ;
        RECT 200.605 2996.615 201.405 2996.695 ;
        RECT 201.575 2996.615 202.375 2996.655 ;
        RECT 200.605 2996.365 202.375 2996.615 ;
        RECT 201.405 2996.325 202.375 2996.365 ;
      LAYER li1 ;
        RECT 202.595 2996.155 202.765 2996.825 ;
      LAYER li1 ;
        RECT 201.405 2995.865 201.575 2996.155 ;
      LAYER li1 ;
        RECT 201.745 2995.985 202.765 2996.155 ;
      LAYER li1 ;
        RECT 198.685 2995.525 199.335 2995.695 ;
        RECT 199.505 2995.590 200.385 2995.765 ;
        RECT 200.605 2995.695 201.405 2995.775 ;
        RECT 201.575 2995.695 202.375 2995.815 ;
        RECT 200.605 2995.605 202.375 2995.695 ;
        RECT 198.685 2995.405 198.855 2995.525 ;
        RECT 199.505 2995.355 199.675 2995.590 ;
        RECT 200.215 2995.435 200.385 2995.590 ;
        RECT 201.405 2995.485 202.375 2995.605 ;
        RECT 198.685 2995.015 198.855 2995.235 ;
        RECT 199.030 2995.185 199.675 2995.355 ;
        RECT 198.685 2994.945 199.335 2995.015 ;
        RECT 198.855 2994.775 199.335 2994.945 ;
        RECT 198.685 2994.685 199.335 2994.775 ;
        RECT 198.685 2994.485 198.855 2994.685 ;
        RECT 199.505 2994.515 199.675 2995.185 ;
        RECT 199.025 2994.345 199.675 2994.515 ;
        RECT 198.685 2994.085 198.855 2994.315 ;
      LAYER li1 ;
        RECT 199.845 2994.310 200.045 2995.410 ;
      LAYER li1 ;
        RECT 200.215 2995.105 201.235 2995.435 ;
        RECT 201.405 2995.405 201.575 2995.485 ;
      LAYER li1 ;
        RECT 202.595 2995.400 202.765 2995.985 ;
      LAYER li1 ;
        RECT 202.965 2995.645 203.135 2998.095 ;
        RECT 203.645 2998.005 204.125 2998.165 ;
      LAYER li1 ;
        RECT 203.305 2997.665 203.955 2997.835 ;
      LAYER li1 ;
        RECT 204.125 2997.705 204.295 2997.995 ;
      LAYER li1 ;
        RECT 203.305 2996.995 203.475 2997.665 ;
      LAYER li1 ;
        RECT 204.125 2997.495 204.295 2997.535 ;
        RECT 203.645 2997.245 204.295 2997.495 ;
        RECT 203.645 2997.165 204.125 2997.245 ;
      LAYER li1 ;
        RECT 203.305 2996.825 203.955 2996.995 ;
        RECT 203.305 2996.155 203.475 2996.825 ;
      LAYER li1 ;
        RECT 204.125 2996.785 204.295 2997.075 ;
        RECT 203.645 2996.615 204.125 2996.655 ;
        RECT 203.645 2996.325 204.295 2996.615 ;
      LAYER li1 ;
        RECT 203.305 2995.985 203.955 2996.155 ;
        RECT 203.305 2995.400 203.475 2995.985 ;
      LAYER li1 ;
        RECT 204.125 2995.865 204.295 2996.155 ;
        RECT 203.645 2995.695 204.125 2995.815 ;
        RECT 203.645 2995.485 204.295 2995.695 ;
        RECT 204.125 2995.405 204.295 2995.485 ;
      LAYER li1 ;
        RECT 202.595 2995.315 203.475 2995.400 ;
      LAYER li1 ;
        RECT 200.215 2994.595 200.385 2995.105 ;
        RECT 201.405 2994.975 201.575 2995.235 ;
      LAYER li1 ;
        RECT 201.745 2995.145 203.955 2995.315 ;
      LAYER li1 ;
        RECT 204.125 2994.975 204.295 2995.235 ;
        RECT 201.405 2994.945 202.725 2994.975 ;
        RECT 200.605 2994.775 201.405 2994.935 ;
        RECT 201.575 2994.775 202.725 2994.945 ;
        RECT 200.605 2994.765 202.725 2994.775 ;
        RECT 201.405 2994.645 202.725 2994.765 ;
        RECT 203.325 2994.945 204.295 2994.975 ;
        RECT 203.325 2994.775 204.125 2994.945 ;
        RECT 203.325 2994.645 204.295 2994.775 ;
        RECT 200.215 2994.265 201.235 2994.595 ;
        RECT 201.405 2994.485 201.575 2994.645 ;
        RECT 204.125 2994.485 204.295 2994.645 ;
        RECT 201.405 2994.085 201.575 2994.315 ;
        RECT 204.125 2994.085 204.295 2994.315 ;
        RECT 198.685 2994.025 199.580 2994.085 ;
        RECT 198.855 2993.855 199.580 2994.025 ;
        RECT 198.685 2993.795 199.580 2993.855 ;
        RECT 200.240 2994.025 202.740 2994.085 ;
        RECT 200.240 2993.855 201.405 2994.025 ;
        RECT 201.575 2993.855 202.740 2994.025 ;
        RECT 200.240 2993.795 202.740 2993.855 ;
        RECT 203.400 2994.025 204.295 2994.085 ;
        RECT 203.400 2993.855 204.125 2994.025 ;
        RECT 203.400 2993.795 204.295 2993.855 ;
        RECT 198.685 2993.565 198.855 2993.795 ;
        RECT 201.405 2993.565 201.575 2993.795 ;
        RECT 198.685 2993.235 198.855 2993.395 ;
        RECT 201.405 2993.235 201.575 2993.395 ;
        RECT 201.745 2993.285 202.765 2993.615 ;
        RECT 204.125 2993.565 204.295 2993.795 ;
        RECT 198.685 2993.105 199.655 2993.235 ;
        RECT 198.855 2992.935 199.655 2993.105 ;
        RECT 198.685 2992.905 199.655 2992.935 ;
        RECT 200.255 2993.115 201.575 2993.235 ;
        RECT 200.255 2993.105 202.375 2993.115 ;
        RECT 200.255 2992.935 201.405 2993.105 ;
        RECT 201.575 2992.945 202.375 2993.105 ;
        RECT 200.255 2992.905 201.575 2992.935 ;
        RECT 198.685 2992.645 198.855 2992.905 ;
        RECT 201.405 2992.645 201.575 2992.905 ;
        RECT 202.595 2992.775 202.765 2993.285 ;
        RECT 198.685 2992.395 198.855 2992.475 ;
        RECT 201.405 2992.395 201.575 2992.475 ;
        RECT 201.745 2992.445 202.765 2992.775 ;
        RECT 198.685 2992.185 199.335 2992.395 ;
        RECT 200.605 2992.275 201.575 2992.395 ;
        RECT 202.595 2992.290 202.765 2992.445 ;
        RECT 203.305 2993.365 203.955 2993.535 ;
        RECT 203.305 2992.695 203.475 2993.365 ;
        RECT 204.125 2993.195 204.295 2993.395 ;
        RECT 203.645 2993.105 204.295 2993.195 ;
        RECT 203.645 2992.935 204.125 2993.105 ;
        RECT 203.645 2992.865 204.295 2992.935 ;
        RECT 203.305 2992.525 203.950 2992.695 ;
        RECT 204.125 2992.645 204.295 2992.865 ;
        RECT 203.305 2992.290 203.475 2992.525 ;
        RECT 204.125 2992.355 204.295 2992.475 ;
        RECT 198.855 2992.065 199.335 2992.185 ;
        RECT 198.685 2991.725 198.855 2992.015 ;
        RECT 198.685 2991.265 199.335 2991.555 ;
        RECT 198.855 2991.225 199.335 2991.265 ;
        RECT 198.685 2990.805 198.855 2991.095 ;
        RECT 198.855 2990.635 199.335 2990.715 ;
        RECT 198.685 2990.385 199.335 2990.635 ;
        RECT 198.685 2990.345 198.855 2990.385 ;
        RECT 198.685 2989.885 198.855 2990.175 ;
        RECT 198.855 2989.715 199.335 2989.875 ;
        RECT 199.845 2989.785 200.015 2992.235 ;
        RECT 200.605 2992.185 202.375 2992.275 ;
        RECT 200.605 2992.065 201.405 2992.185 ;
        RECT 201.575 2992.105 202.375 2992.185 ;
        RECT 202.595 2992.115 203.475 2992.290 ;
        RECT 203.645 2992.185 204.295 2992.355 ;
        RECT 201.405 2991.725 201.575 2992.015 ;
      LAYER li1 ;
        RECT 201.745 2991.685 202.765 2991.855 ;
      LAYER li1 ;
        RECT 200.605 2991.515 201.575 2991.555 ;
        RECT 200.605 2991.265 202.375 2991.515 ;
        RECT 200.605 2991.225 201.405 2991.265 ;
        RECT 201.575 2991.185 202.375 2991.265 ;
        RECT 201.405 2990.805 201.575 2991.095 ;
      LAYER li1 ;
        RECT 202.595 2991.015 202.765 2991.685 ;
        RECT 201.745 2990.845 202.765 2991.015 ;
      LAYER li1 ;
        RECT 200.605 2990.635 201.405 2990.715 ;
        RECT 201.575 2990.635 202.375 2990.675 ;
        RECT 200.605 2990.385 202.375 2990.635 ;
        RECT 201.405 2990.345 202.375 2990.385 ;
      LAYER li1 ;
        RECT 202.595 2990.175 202.765 2990.845 ;
      LAYER li1 ;
        RECT 201.405 2989.885 201.575 2990.175 ;
      LAYER li1 ;
        RECT 201.745 2990.005 202.765 2990.175 ;
      LAYER li1 ;
        RECT 198.685 2989.545 199.335 2989.715 ;
        RECT 199.505 2989.610 200.385 2989.785 ;
        RECT 200.605 2989.715 201.405 2989.795 ;
        RECT 201.575 2989.715 202.375 2989.835 ;
        RECT 200.605 2989.625 202.375 2989.715 ;
        RECT 198.685 2989.425 198.855 2989.545 ;
        RECT 199.505 2989.375 199.675 2989.610 ;
        RECT 200.215 2989.455 200.385 2989.610 ;
        RECT 201.405 2989.505 202.375 2989.625 ;
        RECT 198.685 2989.035 198.855 2989.255 ;
        RECT 199.030 2989.205 199.675 2989.375 ;
        RECT 198.685 2988.965 199.335 2989.035 ;
        RECT 198.855 2988.795 199.335 2988.965 ;
        RECT 198.685 2988.705 199.335 2988.795 ;
        RECT 198.685 2988.505 198.855 2988.705 ;
        RECT 199.505 2988.535 199.675 2989.205 ;
        RECT 199.025 2988.365 199.675 2988.535 ;
        RECT 198.685 2988.105 198.855 2988.335 ;
      LAYER li1 ;
        RECT 199.845 2988.330 200.045 2989.430 ;
      LAYER li1 ;
        RECT 200.215 2989.125 201.235 2989.455 ;
        RECT 201.405 2989.425 201.575 2989.505 ;
      LAYER li1 ;
        RECT 202.595 2989.420 202.765 2990.005 ;
      LAYER li1 ;
        RECT 202.965 2989.665 203.135 2992.115 ;
        RECT 203.645 2992.025 204.125 2992.185 ;
      LAYER li1 ;
        RECT 203.305 2991.685 203.955 2991.855 ;
      LAYER li1 ;
        RECT 204.125 2991.725 204.295 2992.015 ;
      LAYER li1 ;
        RECT 203.305 2991.015 203.475 2991.685 ;
      LAYER li1 ;
        RECT 204.125 2991.515 204.295 2991.555 ;
        RECT 203.645 2991.265 204.295 2991.515 ;
        RECT 203.645 2991.185 204.125 2991.265 ;
      LAYER li1 ;
        RECT 203.305 2990.845 203.955 2991.015 ;
        RECT 203.305 2990.175 203.475 2990.845 ;
      LAYER li1 ;
        RECT 204.125 2990.805 204.295 2991.095 ;
        RECT 203.645 2990.635 204.125 2990.675 ;
        RECT 203.645 2990.345 204.295 2990.635 ;
      LAYER li1 ;
        RECT 203.305 2990.005 203.955 2990.175 ;
        RECT 203.305 2989.420 203.475 2990.005 ;
      LAYER li1 ;
        RECT 204.125 2989.885 204.295 2990.175 ;
        RECT 203.645 2989.715 204.125 2989.835 ;
        RECT 203.645 2989.505 204.295 2989.715 ;
        RECT 204.125 2989.425 204.295 2989.505 ;
      LAYER li1 ;
        RECT 202.595 2989.335 203.475 2989.420 ;
      LAYER li1 ;
        RECT 200.215 2988.615 200.385 2989.125 ;
        RECT 201.405 2988.995 201.575 2989.255 ;
      LAYER li1 ;
        RECT 201.745 2989.165 203.955 2989.335 ;
      LAYER li1 ;
        RECT 204.125 2988.995 204.295 2989.255 ;
        RECT 201.405 2988.965 202.725 2988.995 ;
        RECT 200.605 2988.795 201.405 2988.955 ;
        RECT 201.575 2988.795 202.725 2988.965 ;
        RECT 200.605 2988.785 202.725 2988.795 ;
        RECT 201.405 2988.665 202.725 2988.785 ;
        RECT 203.325 2988.965 204.295 2988.995 ;
        RECT 203.325 2988.795 204.125 2988.965 ;
        RECT 203.325 2988.665 204.295 2988.795 ;
        RECT 200.215 2988.285 201.235 2988.615 ;
        RECT 201.405 2988.505 201.575 2988.665 ;
        RECT 204.125 2988.505 204.295 2988.665 ;
        RECT 201.405 2988.105 201.575 2988.335 ;
        RECT 204.125 2988.105 204.295 2988.335 ;
        RECT 198.685 2988.045 199.580 2988.105 ;
        RECT 198.855 2987.875 199.580 2988.045 ;
        RECT 198.685 2987.815 199.580 2987.875 ;
        RECT 200.240 2988.045 202.740 2988.105 ;
        RECT 200.240 2987.875 201.405 2988.045 ;
        RECT 201.575 2987.875 202.740 2988.045 ;
        RECT 200.240 2987.815 202.740 2987.875 ;
        RECT 203.400 2988.045 204.295 2988.105 ;
        RECT 203.400 2987.875 204.125 2988.045 ;
        RECT 203.400 2987.815 204.295 2987.875 ;
        RECT 198.685 2987.730 198.855 2987.815 ;
        RECT 201.405 2987.730 201.575 2987.815 ;
        RECT 204.125 2987.730 204.295 2987.815 ;
        RECT 3383.500 2238.295 3383.670 2238.380 ;
        RECT 3386.220 2238.295 3386.390 2238.380 ;
        RECT 3388.940 2238.295 3389.110 2238.380 ;
        RECT 3383.500 2238.235 3384.395 2238.295 ;
        RECT 3383.670 2238.065 3384.395 2238.235 ;
        RECT 3383.500 2238.005 3384.395 2238.065 ;
        RECT 3383.500 2237.775 3383.670 2238.005 ;
        RECT 3383.500 2237.405 3383.670 2237.605 ;
        RECT 3383.840 2237.575 3384.490 2237.745 ;
        RECT 3383.500 2237.315 3384.150 2237.405 ;
        RECT 3383.670 2237.145 3384.150 2237.315 ;
        RECT 3383.500 2237.075 3384.150 2237.145 ;
        RECT 3383.500 2236.855 3383.670 2237.075 ;
        RECT 3384.320 2236.905 3384.490 2237.575 ;
        RECT 3383.845 2236.735 3384.490 2236.905 ;
        RECT 3383.500 2236.565 3383.670 2236.685 ;
        RECT 3383.500 2236.395 3384.150 2236.565 ;
        RECT 3383.670 2236.235 3384.150 2236.395 ;
        RECT 3384.320 2236.500 3384.490 2236.735 ;
      LAYER li1 ;
        RECT 3384.660 2236.680 3384.860 2238.270 ;
      LAYER li1 ;
        RECT 3385.055 2238.235 3387.555 2238.295 ;
        RECT 3385.055 2238.065 3386.220 2238.235 ;
        RECT 3386.390 2238.065 3387.555 2238.235 ;
        RECT 3385.055 2238.005 3387.555 2238.065 ;
        RECT 3388.215 2238.235 3389.110 2238.295 ;
        RECT 3388.215 2238.065 3388.940 2238.235 ;
        RECT 3388.215 2238.005 3389.110 2238.065 ;
        RECT 3385.030 2237.495 3386.050 2237.825 ;
        RECT 3386.220 2237.775 3386.390 2238.005 ;
        RECT 3388.940 2237.775 3389.110 2238.005 ;
        RECT 3385.030 2236.985 3385.200 2237.495 ;
        RECT 3386.220 2237.445 3386.390 2237.605 ;
        RECT 3388.940 2237.445 3389.110 2237.605 ;
        RECT 3386.220 2237.325 3387.540 2237.445 ;
        RECT 3385.420 2237.315 3387.540 2237.325 ;
        RECT 3385.420 2237.155 3386.220 2237.315 ;
        RECT 3386.390 2237.145 3387.540 2237.315 ;
        RECT 3386.220 2237.115 3387.540 2237.145 ;
        RECT 3388.140 2237.315 3389.110 2237.445 ;
        RECT 3388.140 2237.145 3388.940 2237.315 ;
        RECT 3388.140 2237.115 3389.110 2237.145 ;
        RECT 3385.030 2236.655 3386.050 2236.985 ;
        RECT 3386.220 2236.855 3386.390 2237.115 ;
      LAYER li1 ;
        RECT 3386.560 2236.775 3388.770 2236.945 ;
      LAYER li1 ;
        RECT 3388.940 2236.855 3389.110 2237.115 ;
      LAYER li1 ;
        RECT 3387.410 2236.690 3388.290 2236.775 ;
      LAYER li1 ;
        RECT 3385.030 2236.500 3385.200 2236.655 ;
        RECT 3384.320 2236.325 3385.200 2236.500 ;
        RECT 3386.220 2236.605 3386.390 2236.685 ;
        RECT 3386.220 2236.485 3387.190 2236.605 ;
        RECT 3385.420 2236.395 3387.190 2236.485 ;
        RECT 3383.500 2235.935 3383.670 2236.225 ;
        RECT 3383.500 2235.725 3383.670 2235.765 ;
        RECT 3383.500 2235.475 3384.150 2235.725 ;
        RECT 3383.670 2235.395 3384.150 2235.475 ;
        RECT 3383.500 2235.015 3383.670 2235.305 ;
        RECT 3383.670 2234.845 3384.150 2234.885 ;
        RECT 3383.500 2234.555 3384.150 2234.845 ;
        RECT 3383.500 2234.095 3383.670 2234.385 ;
        RECT 3383.670 2233.925 3384.150 2234.045 ;
        RECT 3383.500 2233.715 3384.150 2233.925 ;
        RECT 3384.660 2233.875 3384.830 2236.325 ;
        RECT 3385.420 2236.315 3386.220 2236.395 ;
        RECT 3386.390 2236.275 3387.190 2236.395 ;
        RECT 3386.220 2235.935 3386.390 2236.225 ;
      LAYER li1 ;
        RECT 3387.410 2236.105 3387.580 2236.690 ;
        RECT 3386.560 2235.935 3387.580 2236.105 ;
      LAYER li1 ;
        RECT 3386.220 2235.725 3387.190 2235.765 ;
        RECT 3385.420 2235.475 3387.190 2235.725 ;
        RECT 3385.420 2235.395 3386.220 2235.475 ;
        RECT 3386.390 2235.435 3387.190 2235.475 ;
        RECT 3386.220 2235.015 3386.390 2235.305 ;
      LAYER li1 ;
        RECT 3387.410 2235.265 3387.580 2235.935 ;
        RECT 3386.560 2235.095 3387.580 2235.265 ;
      LAYER li1 ;
        RECT 3385.420 2234.845 3386.220 2234.885 ;
        RECT 3386.390 2234.845 3387.190 2234.925 ;
        RECT 3385.420 2234.595 3387.190 2234.845 ;
        RECT 3385.420 2234.555 3386.390 2234.595 ;
      LAYER li1 ;
        RECT 3387.410 2234.425 3387.580 2235.095 ;
      LAYER li1 ;
        RECT 3386.220 2234.095 3386.390 2234.385 ;
      LAYER li1 ;
        RECT 3386.560 2234.255 3387.580 2234.425 ;
      LAYER li1 ;
        RECT 3385.420 2233.925 3386.220 2234.045 ;
        RECT 3386.390 2233.925 3387.190 2234.005 ;
        RECT 3387.780 2233.995 3387.950 2236.445 ;
      LAYER li1 ;
        RECT 3388.120 2236.105 3388.290 2236.690 ;
      LAYER li1 ;
        RECT 3388.940 2236.605 3389.110 2236.685 ;
        RECT 3388.460 2236.395 3389.110 2236.605 ;
        RECT 3388.460 2236.275 3388.940 2236.395 ;
      LAYER li1 ;
        RECT 3388.120 2235.935 3388.770 2236.105 ;
      LAYER li1 ;
        RECT 3388.940 2235.935 3389.110 2236.225 ;
      LAYER li1 ;
        RECT 3388.120 2235.265 3388.290 2235.935 ;
      LAYER li1 ;
        RECT 3388.460 2235.475 3389.110 2235.765 ;
        RECT 3388.460 2235.435 3388.940 2235.475 ;
      LAYER li1 ;
        RECT 3388.120 2235.095 3388.770 2235.265 ;
        RECT 3388.120 2234.425 3388.290 2235.095 ;
      LAYER li1 ;
        RECT 3388.940 2235.015 3389.110 2235.305 ;
        RECT 3388.460 2234.845 3388.940 2234.925 ;
        RECT 3388.460 2234.595 3389.110 2234.845 ;
        RECT 3388.940 2234.555 3389.110 2234.595 ;
      LAYER li1 ;
        RECT 3388.120 2234.255 3388.770 2234.425 ;
      LAYER li1 ;
        RECT 3388.940 2234.095 3389.110 2234.385 ;
        RECT 3385.420 2233.835 3387.190 2233.925 ;
        RECT 3385.420 2233.715 3386.390 2233.835 ;
        RECT 3383.500 2233.635 3383.670 2233.715 ;
        RECT 3386.220 2233.635 3386.390 2233.715 ;
        RECT 3387.410 2233.820 3388.290 2233.995 ;
        RECT 3387.410 2233.665 3387.580 2233.820 ;
        RECT 3383.500 2233.205 3383.670 2233.465 ;
        RECT 3386.220 2233.205 3386.390 2233.465 ;
        RECT 3386.560 2233.335 3387.580 2233.665 ;
        RECT 3383.500 2233.175 3384.470 2233.205 ;
        RECT 3383.670 2233.005 3384.470 2233.175 ;
        RECT 3383.500 2232.875 3384.470 2233.005 ;
        RECT 3385.070 2233.175 3386.390 2233.205 ;
        RECT 3385.070 2233.005 3386.220 2233.175 ;
        RECT 3386.390 2233.005 3387.190 2233.165 ;
        RECT 3385.070 2232.995 3387.190 2233.005 ;
        RECT 3385.070 2232.875 3386.390 2232.995 ;
        RECT 3383.500 2232.715 3383.670 2232.875 ;
        RECT 3386.220 2232.715 3386.390 2232.875 ;
        RECT 3387.410 2232.825 3387.580 2233.335 ;
        RECT 3383.500 2232.315 3383.670 2232.545 ;
        RECT 3386.220 2232.315 3386.390 2232.545 ;
        RECT 3386.560 2232.495 3387.580 2232.825 ;
        RECT 3388.120 2233.585 3388.290 2233.820 ;
        RECT 3388.460 2233.925 3388.940 2234.085 ;
        RECT 3388.460 2233.755 3389.110 2233.925 ;
        RECT 3388.940 2233.635 3389.110 2233.755 ;
        RECT 3388.120 2233.415 3388.765 2233.585 ;
        RECT 3388.120 2232.745 3388.290 2233.415 ;
        RECT 3388.940 2233.245 3389.110 2233.465 ;
        RECT 3388.460 2233.175 3389.110 2233.245 ;
        RECT 3388.460 2233.005 3388.940 2233.175 ;
        RECT 3388.460 2232.915 3389.110 2233.005 ;
        RECT 3388.120 2232.575 3388.770 2232.745 ;
        RECT 3388.940 2232.715 3389.110 2232.915 ;
        RECT 3388.940 2232.315 3389.110 2232.545 ;
        RECT 3383.500 2232.255 3384.395 2232.315 ;
        RECT 3383.670 2232.085 3384.395 2232.255 ;
        RECT 3383.500 2232.025 3384.395 2232.085 ;
        RECT 3385.055 2232.255 3387.555 2232.315 ;
        RECT 3385.055 2232.085 3386.220 2232.255 ;
        RECT 3386.390 2232.085 3387.555 2232.255 ;
        RECT 3385.055 2232.025 3387.555 2232.085 ;
        RECT 3388.215 2232.255 3389.110 2232.315 ;
        RECT 3388.215 2232.085 3388.940 2232.255 ;
        RECT 3388.215 2232.025 3389.110 2232.085 ;
        RECT 3383.500 2231.795 3383.670 2232.025 ;
        RECT 3383.500 2231.425 3383.670 2231.625 ;
        RECT 3383.840 2231.595 3384.490 2231.765 ;
        RECT 3383.500 2231.335 3384.150 2231.425 ;
        RECT 3383.670 2231.165 3384.150 2231.335 ;
        RECT 3383.500 2231.095 3384.150 2231.165 ;
        RECT 3383.500 2230.875 3383.670 2231.095 ;
        RECT 3384.320 2230.925 3384.490 2231.595 ;
        RECT 3383.845 2230.755 3384.490 2230.925 ;
        RECT 3383.500 2230.585 3383.670 2230.705 ;
        RECT 3383.500 2230.415 3384.150 2230.585 ;
        RECT 3383.670 2230.255 3384.150 2230.415 ;
        RECT 3384.320 2230.520 3384.490 2230.755 ;
        RECT 3385.030 2231.515 3386.050 2231.845 ;
        RECT 3386.220 2231.795 3386.390 2232.025 ;
        RECT 3388.940 2231.795 3389.110 2232.025 ;
        RECT 3385.030 2231.005 3385.200 2231.515 ;
        RECT 3386.220 2231.465 3386.390 2231.625 ;
        RECT 3388.940 2231.465 3389.110 2231.625 ;
        RECT 3386.220 2231.345 3387.540 2231.465 ;
        RECT 3385.420 2231.335 3387.540 2231.345 ;
        RECT 3385.420 2231.175 3386.220 2231.335 ;
        RECT 3386.390 2231.165 3387.540 2231.335 ;
        RECT 3386.220 2231.135 3387.540 2231.165 ;
        RECT 3388.140 2231.335 3389.110 2231.465 ;
        RECT 3388.140 2231.165 3388.940 2231.335 ;
        RECT 3388.140 2231.135 3389.110 2231.165 ;
        RECT 3385.030 2230.675 3386.050 2231.005 ;
        RECT 3386.220 2230.875 3386.390 2231.135 ;
        RECT 3388.940 2230.875 3389.110 2231.135 ;
        RECT 3385.030 2230.520 3385.200 2230.675 ;
        RECT 3384.320 2230.345 3385.200 2230.520 ;
        RECT 3386.220 2230.625 3386.390 2230.705 ;
        RECT 3388.940 2230.625 3389.110 2230.705 ;
        RECT 3386.220 2230.505 3387.190 2230.625 ;
        RECT 3385.420 2230.415 3387.190 2230.505 ;
        RECT 3383.500 2229.955 3383.670 2230.245 ;
        RECT 3383.500 2229.745 3383.670 2229.785 ;
        RECT 3383.500 2229.495 3384.150 2229.745 ;
        RECT 3383.670 2229.415 3384.150 2229.495 ;
        RECT 3383.500 2229.035 3383.670 2229.325 ;
        RECT 3383.670 2228.865 3384.150 2228.905 ;
        RECT 3383.500 2228.575 3384.150 2228.865 ;
        RECT 3383.500 2228.115 3383.670 2228.405 ;
        RECT 3383.670 2227.945 3384.150 2228.065 ;
        RECT 3383.500 2227.735 3384.150 2227.945 ;
        RECT 3384.660 2227.895 3384.830 2230.345 ;
        RECT 3385.420 2230.335 3386.220 2230.415 ;
        RECT 3386.390 2230.295 3387.190 2230.415 ;
        RECT 3386.220 2229.955 3386.390 2230.245 ;
        RECT 3386.220 2229.745 3387.190 2229.785 ;
        RECT 3385.420 2229.495 3387.190 2229.745 ;
        RECT 3385.420 2229.415 3386.220 2229.495 ;
        RECT 3386.390 2229.455 3387.190 2229.495 ;
        RECT 3386.220 2229.035 3386.390 2229.325 ;
        RECT 3385.420 2228.865 3386.220 2228.905 ;
        RECT 3386.390 2228.865 3387.190 2228.945 ;
        RECT 3385.420 2228.615 3387.190 2228.865 ;
        RECT 3385.420 2228.575 3386.390 2228.615 ;
        RECT 3386.220 2228.115 3386.390 2228.405 ;
        RECT 3385.420 2227.945 3386.220 2228.065 ;
        RECT 3386.390 2227.945 3387.190 2228.025 ;
        RECT 3387.780 2228.015 3387.950 2230.465 ;
        RECT 3388.460 2230.415 3389.110 2230.625 ;
        RECT 3388.460 2230.295 3388.940 2230.415 ;
        RECT 3388.940 2229.955 3389.110 2230.245 ;
        RECT 3388.460 2229.495 3389.110 2229.785 ;
        RECT 3388.460 2229.455 3388.940 2229.495 ;
        RECT 3388.940 2229.035 3389.110 2229.325 ;
        RECT 3388.460 2228.865 3388.940 2228.945 ;
        RECT 3388.460 2228.615 3389.110 2228.865 ;
        RECT 3388.940 2228.575 3389.110 2228.615 ;
        RECT 3388.940 2228.115 3389.110 2228.405 ;
        RECT 3385.420 2227.855 3387.190 2227.945 ;
        RECT 3385.420 2227.735 3386.390 2227.855 ;
        RECT 3383.500 2227.655 3383.670 2227.735 ;
        RECT 3386.220 2227.655 3386.390 2227.735 ;
        RECT 3387.410 2227.840 3388.290 2228.015 ;
        RECT 3387.410 2227.685 3387.580 2227.840 ;
        RECT 3383.500 2227.225 3383.670 2227.485 ;
        RECT 3386.220 2227.225 3386.390 2227.485 ;
        RECT 3386.560 2227.355 3387.580 2227.685 ;
        RECT 3383.500 2227.195 3384.470 2227.225 ;
        RECT 3383.670 2227.025 3384.470 2227.195 ;
        RECT 3383.500 2226.895 3384.470 2227.025 ;
        RECT 3385.070 2227.195 3386.390 2227.225 ;
        RECT 3385.070 2227.025 3386.220 2227.195 ;
        RECT 3386.390 2227.025 3387.190 2227.185 ;
        RECT 3385.070 2227.015 3387.190 2227.025 ;
        RECT 3385.070 2226.895 3386.390 2227.015 ;
        RECT 3383.500 2226.735 3383.670 2226.895 ;
        RECT 3386.220 2226.735 3386.390 2226.895 ;
        RECT 3387.410 2226.845 3387.580 2227.355 ;
        RECT 3383.500 2226.335 3383.670 2226.565 ;
        RECT 3386.220 2226.335 3386.390 2226.565 ;
        RECT 3386.560 2226.515 3387.580 2226.845 ;
        RECT 3388.120 2227.605 3388.290 2227.840 ;
        RECT 3388.460 2227.945 3388.940 2228.105 ;
        RECT 3388.460 2227.775 3389.110 2227.945 ;
        RECT 3388.940 2227.655 3389.110 2227.775 ;
        RECT 3388.120 2227.435 3388.765 2227.605 ;
        RECT 3388.120 2226.765 3388.290 2227.435 ;
        RECT 3388.940 2227.265 3389.110 2227.485 ;
        RECT 3388.460 2227.195 3389.110 2227.265 ;
        RECT 3388.460 2227.025 3388.940 2227.195 ;
        RECT 3388.460 2226.935 3389.110 2227.025 ;
        RECT 3388.120 2226.595 3388.770 2226.765 ;
        RECT 3388.940 2226.735 3389.110 2226.935 ;
        RECT 3388.940 2226.335 3389.110 2226.565 ;
        RECT 3383.500 2226.275 3384.395 2226.335 ;
        RECT 3383.670 2226.105 3384.395 2226.275 ;
        RECT 3383.500 2226.045 3384.395 2226.105 ;
        RECT 3385.055 2226.275 3387.555 2226.335 ;
        RECT 3385.055 2226.105 3386.220 2226.275 ;
        RECT 3386.390 2226.105 3387.555 2226.275 ;
        RECT 3385.055 2226.045 3387.555 2226.105 ;
        RECT 3388.215 2226.275 3389.110 2226.335 ;
        RECT 3388.215 2226.105 3388.940 2226.275 ;
        RECT 3388.215 2226.045 3389.110 2226.105 ;
        RECT 3383.500 2225.815 3383.670 2226.045 ;
        RECT 3383.500 2225.445 3383.670 2225.645 ;
        RECT 3383.840 2225.615 3384.490 2225.785 ;
        RECT 3383.500 2225.355 3384.150 2225.445 ;
        RECT 3383.670 2225.185 3384.150 2225.355 ;
        RECT 3383.500 2225.115 3384.150 2225.185 ;
        RECT 3383.500 2224.895 3383.670 2225.115 ;
        RECT 3384.320 2224.945 3384.490 2225.615 ;
        RECT 3383.845 2224.775 3384.490 2224.945 ;
        RECT 3383.500 2224.605 3383.670 2224.725 ;
        RECT 3383.500 2224.435 3384.150 2224.605 ;
        RECT 3383.670 2224.275 3384.150 2224.435 ;
        RECT 3384.320 2224.540 3384.490 2224.775 ;
        RECT 3385.030 2225.535 3386.050 2225.865 ;
        RECT 3386.220 2225.815 3386.390 2226.045 ;
        RECT 3388.940 2225.815 3389.110 2226.045 ;
        RECT 3385.030 2225.025 3385.200 2225.535 ;
        RECT 3386.220 2225.485 3386.390 2225.645 ;
        RECT 3388.940 2225.485 3389.110 2225.645 ;
        RECT 3386.220 2225.365 3387.540 2225.485 ;
        RECT 3385.420 2225.355 3387.540 2225.365 ;
        RECT 3385.420 2225.195 3386.220 2225.355 ;
        RECT 3386.390 2225.185 3387.540 2225.355 ;
        RECT 3386.220 2225.155 3387.540 2225.185 ;
        RECT 3388.140 2225.355 3389.110 2225.485 ;
        RECT 3388.140 2225.185 3388.940 2225.355 ;
        RECT 3388.140 2225.155 3389.110 2225.185 ;
        RECT 3385.030 2224.695 3386.050 2225.025 ;
        RECT 3386.220 2224.895 3386.390 2225.155 ;
        RECT 3388.940 2224.895 3389.110 2225.155 ;
        RECT 3385.030 2224.540 3385.200 2224.695 ;
        RECT 3384.320 2224.365 3385.200 2224.540 ;
        RECT 3386.220 2224.645 3386.390 2224.725 ;
        RECT 3388.940 2224.645 3389.110 2224.725 ;
        RECT 3386.220 2224.525 3387.190 2224.645 ;
        RECT 3385.420 2224.435 3387.190 2224.525 ;
        RECT 3383.500 2223.975 3383.670 2224.265 ;
        RECT 3383.500 2223.765 3383.670 2223.805 ;
        RECT 3383.500 2223.515 3384.150 2223.765 ;
        RECT 3383.670 2223.435 3384.150 2223.515 ;
        RECT 3383.500 2223.055 3383.670 2223.345 ;
        RECT 3383.670 2222.885 3384.150 2222.925 ;
        RECT 3383.500 2222.595 3384.150 2222.885 ;
        RECT 3383.500 2222.135 3383.670 2222.425 ;
        RECT 3383.670 2221.965 3384.150 2222.085 ;
        RECT 3383.500 2221.755 3384.150 2221.965 ;
        RECT 3384.660 2221.915 3384.830 2224.365 ;
        RECT 3385.420 2224.355 3386.220 2224.435 ;
        RECT 3386.390 2224.315 3387.190 2224.435 ;
        RECT 3386.220 2223.975 3386.390 2224.265 ;
        RECT 3386.220 2223.765 3387.190 2223.805 ;
        RECT 3385.420 2223.515 3387.190 2223.765 ;
        RECT 3385.420 2223.435 3386.220 2223.515 ;
        RECT 3386.390 2223.475 3387.190 2223.515 ;
        RECT 3386.220 2223.055 3386.390 2223.345 ;
        RECT 3385.420 2222.885 3386.220 2222.925 ;
        RECT 3386.390 2222.885 3387.190 2222.965 ;
        RECT 3385.420 2222.635 3387.190 2222.885 ;
        RECT 3385.420 2222.595 3386.390 2222.635 ;
        RECT 3386.220 2222.135 3386.390 2222.425 ;
        RECT 3385.420 2221.965 3386.220 2222.085 ;
        RECT 3386.390 2221.965 3387.190 2222.045 ;
        RECT 3387.780 2222.035 3387.950 2224.485 ;
        RECT 3388.460 2224.435 3389.110 2224.645 ;
        RECT 3388.460 2224.315 3388.940 2224.435 ;
        RECT 3388.940 2223.975 3389.110 2224.265 ;
        RECT 3388.460 2223.515 3389.110 2223.805 ;
        RECT 3388.460 2223.475 3388.940 2223.515 ;
        RECT 3388.940 2223.055 3389.110 2223.345 ;
        RECT 3388.460 2222.885 3388.940 2222.965 ;
        RECT 3388.460 2222.635 3389.110 2222.885 ;
        RECT 3388.940 2222.595 3389.110 2222.635 ;
        RECT 3388.940 2222.135 3389.110 2222.425 ;
        RECT 3385.420 2221.875 3387.190 2221.965 ;
        RECT 3385.420 2221.755 3386.390 2221.875 ;
        RECT 3383.500 2221.675 3383.670 2221.755 ;
        RECT 3386.220 2221.675 3386.390 2221.755 ;
        RECT 3387.410 2221.860 3388.290 2222.035 ;
        RECT 3387.410 2221.705 3387.580 2221.860 ;
        RECT 3383.500 2221.245 3383.670 2221.505 ;
        RECT 3386.220 2221.245 3386.390 2221.505 ;
        RECT 3386.560 2221.375 3387.580 2221.705 ;
        RECT 3383.500 2221.215 3384.470 2221.245 ;
        RECT 3383.670 2221.045 3384.470 2221.215 ;
        RECT 3383.500 2220.915 3384.470 2221.045 ;
        RECT 3385.070 2221.215 3386.390 2221.245 ;
        RECT 3385.070 2221.045 3386.220 2221.215 ;
        RECT 3386.390 2221.045 3387.190 2221.205 ;
        RECT 3385.070 2221.035 3387.190 2221.045 ;
        RECT 3385.070 2220.915 3386.390 2221.035 ;
        RECT 3383.500 2220.755 3383.670 2220.915 ;
        RECT 3386.220 2220.755 3386.390 2220.915 ;
        RECT 3387.410 2220.865 3387.580 2221.375 ;
        RECT 3383.500 2220.355 3383.670 2220.585 ;
        RECT 3386.220 2220.355 3386.390 2220.585 ;
        RECT 3386.560 2220.535 3387.580 2220.865 ;
        RECT 3388.120 2221.625 3388.290 2221.860 ;
        RECT 3388.460 2221.965 3388.940 2222.125 ;
        RECT 3388.460 2221.795 3389.110 2221.965 ;
        RECT 3388.940 2221.675 3389.110 2221.795 ;
        RECT 3388.120 2221.455 3388.765 2221.625 ;
        RECT 3388.120 2220.785 3388.290 2221.455 ;
        RECT 3388.940 2221.285 3389.110 2221.505 ;
        RECT 3388.460 2221.215 3389.110 2221.285 ;
        RECT 3388.460 2221.045 3388.940 2221.215 ;
        RECT 3388.460 2220.955 3389.110 2221.045 ;
        RECT 3388.120 2220.615 3388.770 2220.785 ;
        RECT 3388.940 2220.755 3389.110 2220.955 ;
        RECT 3388.940 2220.355 3389.110 2220.585 ;
        RECT 3383.500 2220.295 3384.395 2220.355 ;
        RECT 3383.670 2220.125 3384.395 2220.295 ;
        RECT 3383.500 2220.065 3384.395 2220.125 ;
        RECT 3385.055 2220.295 3387.555 2220.355 ;
        RECT 3385.055 2220.125 3386.220 2220.295 ;
        RECT 3386.390 2220.125 3387.555 2220.295 ;
        RECT 3385.055 2220.065 3387.555 2220.125 ;
        RECT 3388.215 2220.295 3389.110 2220.355 ;
        RECT 3388.215 2220.125 3388.940 2220.295 ;
        RECT 3388.215 2220.065 3389.110 2220.125 ;
        RECT 3383.500 2219.835 3383.670 2220.065 ;
        RECT 3383.500 2219.465 3383.670 2219.665 ;
        RECT 3383.840 2219.635 3384.490 2219.805 ;
        RECT 3383.500 2219.375 3384.150 2219.465 ;
        RECT 3383.670 2219.205 3384.150 2219.375 ;
        RECT 3383.500 2219.135 3384.150 2219.205 ;
        RECT 3383.500 2218.915 3383.670 2219.135 ;
        RECT 3384.320 2218.965 3384.490 2219.635 ;
        RECT 3383.845 2218.795 3384.490 2218.965 ;
        RECT 3383.500 2218.625 3383.670 2218.745 ;
        RECT 3383.500 2218.455 3384.150 2218.625 ;
        RECT 3383.670 2218.295 3384.150 2218.455 ;
        RECT 3384.320 2218.560 3384.490 2218.795 ;
        RECT 3385.030 2219.555 3386.050 2219.885 ;
        RECT 3386.220 2219.835 3386.390 2220.065 ;
        RECT 3388.940 2219.835 3389.110 2220.065 ;
        RECT 3385.030 2219.045 3385.200 2219.555 ;
        RECT 3386.220 2219.505 3386.390 2219.665 ;
        RECT 3388.940 2219.505 3389.110 2219.665 ;
        RECT 3386.220 2219.385 3387.540 2219.505 ;
        RECT 3385.420 2219.375 3387.540 2219.385 ;
        RECT 3385.420 2219.215 3386.220 2219.375 ;
        RECT 3386.390 2219.205 3387.540 2219.375 ;
        RECT 3386.220 2219.175 3387.540 2219.205 ;
        RECT 3388.140 2219.375 3389.110 2219.505 ;
        RECT 3388.140 2219.205 3388.940 2219.375 ;
        RECT 3388.140 2219.175 3389.110 2219.205 ;
        RECT 3385.030 2218.715 3386.050 2219.045 ;
        RECT 3386.220 2218.915 3386.390 2219.175 ;
        RECT 3388.940 2218.915 3389.110 2219.175 ;
        RECT 3385.030 2218.560 3385.200 2218.715 ;
        RECT 3384.320 2218.385 3385.200 2218.560 ;
        RECT 3386.220 2218.665 3386.390 2218.745 ;
        RECT 3388.940 2218.665 3389.110 2218.745 ;
        RECT 3386.220 2218.545 3387.190 2218.665 ;
        RECT 3385.420 2218.455 3387.190 2218.545 ;
        RECT 3383.500 2217.995 3383.670 2218.285 ;
        RECT 3383.500 2217.785 3383.670 2217.825 ;
        RECT 3383.500 2217.535 3384.150 2217.785 ;
        RECT 3383.670 2217.455 3384.150 2217.535 ;
        RECT 3383.500 2217.075 3383.670 2217.365 ;
        RECT 3383.670 2216.905 3384.150 2216.945 ;
        RECT 3383.500 2216.615 3384.150 2216.905 ;
        RECT 3383.500 2216.155 3383.670 2216.445 ;
        RECT 3383.670 2215.985 3384.150 2216.105 ;
        RECT 3383.500 2215.775 3384.150 2215.985 ;
        RECT 3384.660 2215.935 3384.830 2218.385 ;
        RECT 3385.420 2218.375 3386.220 2218.455 ;
        RECT 3386.390 2218.335 3387.190 2218.455 ;
        RECT 3386.220 2217.995 3386.390 2218.285 ;
        RECT 3386.220 2217.785 3387.190 2217.825 ;
        RECT 3385.420 2217.535 3387.190 2217.785 ;
        RECT 3385.420 2217.455 3386.220 2217.535 ;
        RECT 3386.390 2217.495 3387.190 2217.535 ;
        RECT 3386.220 2217.075 3386.390 2217.365 ;
        RECT 3385.420 2216.905 3386.220 2216.945 ;
        RECT 3386.390 2216.905 3387.190 2216.985 ;
        RECT 3385.420 2216.655 3387.190 2216.905 ;
        RECT 3385.420 2216.615 3386.390 2216.655 ;
        RECT 3386.220 2216.155 3386.390 2216.445 ;
        RECT 3385.420 2215.985 3386.220 2216.105 ;
        RECT 3386.390 2215.985 3387.190 2216.065 ;
        RECT 3387.780 2216.055 3387.950 2218.505 ;
        RECT 3388.460 2218.455 3389.110 2218.665 ;
        RECT 3388.460 2218.335 3388.940 2218.455 ;
        RECT 3388.940 2217.995 3389.110 2218.285 ;
        RECT 3388.460 2217.535 3389.110 2217.825 ;
        RECT 3388.460 2217.495 3388.940 2217.535 ;
        RECT 3388.940 2217.075 3389.110 2217.365 ;
        RECT 3388.460 2216.905 3388.940 2216.985 ;
        RECT 3388.460 2216.655 3389.110 2216.905 ;
        RECT 3388.940 2216.615 3389.110 2216.655 ;
        RECT 3388.940 2216.155 3389.110 2216.445 ;
        RECT 3385.420 2215.895 3387.190 2215.985 ;
        RECT 3385.420 2215.775 3386.390 2215.895 ;
        RECT 3383.500 2215.695 3383.670 2215.775 ;
        RECT 3386.220 2215.695 3386.390 2215.775 ;
        RECT 3387.410 2215.880 3388.290 2216.055 ;
        RECT 3387.410 2215.725 3387.580 2215.880 ;
        RECT 3383.500 2215.265 3383.670 2215.525 ;
        RECT 3386.220 2215.265 3386.390 2215.525 ;
        RECT 3386.560 2215.395 3387.580 2215.725 ;
        RECT 3383.500 2215.235 3384.470 2215.265 ;
        RECT 3383.670 2215.065 3384.470 2215.235 ;
        RECT 3383.500 2214.935 3384.470 2215.065 ;
        RECT 3385.070 2215.235 3386.390 2215.265 ;
        RECT 3385.070 2215.065 3386.220 2215.235 ;
        RECT 3386.390 2215.065 3387.190 2215.225 ;
        RECT 3385.070 2215.055 3387.190 2215.065 ;
        RECT 3385.070 2214.935 3386.390 2215.055 ;
        RECT 3383.500 2214.775 3383.670 2214.935 ;
        RECT 3386.220 2214.775 3386.390 2214.935 ;
        RECT 3387.410 2214.885 3387.580 2215.395 ;
        RECT 3383.500 2214.375 3383.670 2214.605 ;
        RECT 3386.220 2214.375 3386.390 2214.605 ;
        RECT 3386.560 2214.555 3387.580 2214.885 ;
        RECT 3388.120 2215.645 3388.290 2215.880 ;
        RECT 3388.460 2215.985 3388.940 2216.145 ;
        RECT 3388.460 2215.815 3389.110 2215.985 ;
        RECT 3388.940 2215.695 3389.110 2215.815 ;
        RECT 3388.120 2215.475 3388.765 2215.645 ;
        RECT 3388.120 2214.805 3388.290 2215.475 ;
        RECT 3388.940 2215.305 3389.110 2215.525 ;
        RECT 3388.460 2215.235 3389.110 2215.305 ;
        RECT 3388.460 2215.065 3388.940 2215.235 ;
        RECT 3388.460 2214.975 3389.110 2215.065 ;
        RECT 3388.120 2214.635 3388.770 2214.805 ;
        RECT 3388.940 2214.775 3389.110 2214.975 ;
        RECT 3388.940 2214.375 3389.110 2214.605 ;
        RECT 3383.500 2214.315 3384.395 2214.375 ;
        RECT 3383.670 2214.145 3384.395 2214.315 ;
        RECT 3383.500 2214.085 3384.395 2214.145 ;
        RECT 3385.055 2214.315 3387.555 2214.375 ;
        RECT 3385.055 2214.145 3386.220 2214.315 ;
        RECT 3386.390 2214.145 3387.555 2214.315 ;
        RECT 3385.055 2214.085 3387.555 2214.145 ;
        RECT 3388.215 2214.315 3389.110 2214.375 ;
        RECT 3388.215 2214.145 3388.940 2214.315 ;
        RECT 3388.215 2214.085 3389.110 2214.145 ;
        RECT 3383.500 2213.855 3383.670 2214.085 ;
        RECT 3383.500 2213.485 3383.670 2213.685 ;
        RECT 3383.840 2213.655 3384.490 2213.825 ;
        RECT 3383.500 2213.395 3384.150 2213.485 ;
        RECT 3383.670 2213.225 3384.150 2213.395 ;
        RECT 3383.500 2213.155 3384.150 2213.225 ;
        RECT 3383.500 2212.935 3383.670 2213.155 ;
        RECT 3384.320 2212.985 3384.490 2213.655 ;
        RECT 3383.845 2212.815 3384.490 2212.985 ;
        RECT 3383.500 2212.645 3383.670 2212.765 ;
        RECT 3383.500 2212.475 3384.150 2212.645 ;
        RECT 3383.670 2212.315 3384.150 2212.475 ;
        RECT 3384.320 2212.580 3384.490 2212.815 ;
        RECT 3385.030 2213.575 3386.050 2213.905 ;
        RECT 3386.220 2213.855 3386.390 2214.085 ;
        RECT 3388.940 2213.855 3389.110 2214.085 ;
        RECT 3385.030 2213.065 3385.200 2213.575 ;
        RECT 3386.220 2213.525 3386.390 2213.685 ;
        RECT 3388.940 2213.525 3389.110 2213.685 ;
        RECT 3386.220 2213.405 3387.540 2213.525 ;
        RECT 3385.420 2213.395 3387.540 2213.405 ;
        RECT 3385.420 2213.235 3386.220 2213.395 ;
        RECT 3386.390 2213.225 3387.540 2213.395 ;
        RECT 3386.220 2213.195 3387.540 2213.225 ;
        RECT 3388.140 2213.395 3389.110 2213.525 ;
        RECT 3388.140 2213.225 3388.940 2213.395 ;
        RECT 3388.140 2213.195 3389.110 2213.225 ;
        RECT 3385.030 2212.735 3386.050 2213.065 ;
        RECT 3386.220 2212.935 3386.390 2213.195 ;
        RECT 3388.940 2212.935 3389.110 2213.195 ;
        RECT 3385.030 2212.580 3385.200 2212.735 ;
        RECT 3384.320 2212.405 3385.200 2212.580 ;
        RECT 3386.220 2212.685 3386.390 2212.765 ;
        RECT 3388.940 2212.685 3389.110 2212.765 ;
        RECT 3386.220 2212.565 3387.190 2212.685 ;
        RECT 3385.420 2212.475 3387.190 2212.565 ;
        RECT 3383.500 2212.015 3383.670 2212.305 ;
        RECT 3383.500 2211.805 3383.670 2211.845 ;
        RECT 3383.500 2211.555 3384.150 2211.805 ;
        RECT 3383.670 2211.475 3384.150 2211.555 ;
        RECT 3383.500 2211.095 3383.670 2211.385 ;
        RECT 3383.670 2210.925 3384.150 2210.965 ;
        RECT 3383.500 2210.635 3384.150 2210.925 ;
        RECT 3383.500 2210.175 3383.670 2210.465 ;
        RECT 3383.670 2210.005 3384.150 2210.125 ;
        RECT 3383.500 2209.795 3384.150 2210.005 ;
        RECT 3384.660 2209.955 3384.830 2212.405 ;
        RECT 3385.420 2212.395 3386.220 2212.475 ;
        RECT 3386.390 2212.355 3387.190 2212.475 ;
        RECT 3386.220 2212.015 3386.390 2212.305 ;
        RECT 3386.220 2211.805 3387.190 2211.845 ;
        RECT 3385.420 2211.555 3387.190 2211.805 ;
        RECT 3385.420 2211.475 3386.220 2211.555 ;
        RECT 3386.390 2211.515 3387.190 2211.555 ;
        RECT 3386.220 2211.095 3386.390 2211.385 ;
        RECT 3385.420 2210.925 3386.220 2210.965 ;
        RECT 3386.390 2210.925 3387.190 2211.005 ;
        RECT 3385.420 2210.675 3387.190 2210.925 ;
        RECT 3385.420 2210.635 3386.390 2210.675 ;
        RECT 3386.220 2210.175 3386.390 2210.465 ;
        RECT 3385.420 2210.005 3386.220 2210.125 ;
        RECT 3386.390 2210.005 3387.190 2210.085 ;
        RECT 3387.780 2210.075 3387.950 2212.525 ;
        RECT 3388.460 2212.475 3389.110 2212.685 ;
        RECT 3388.460 2212.355 3388.940 2212.475 ;
        RECT 3388.940 2212.015 3389.110 2212.305 ;
        RECT 3388.460 2211.555 3389.110 2211.845 ;
        RECT 3388.460 2211.515 3388.940 2211.555 ;
        RECT 3388.940 2211.095 3389.110 2211.385 ;
        RECT 3388.460 2210.925 3388.940 2211.005 ;
        RECT 3388.460 2210.675 3389.110 2210.925 ;
        RECT 3388.940 2210.635 3389.110 2210.675 ;
        RECT 3388.940 2210.175 3389.110 2210.465 ;
        RECT 3385.420 2209.915 3387.190 2210.005 ;
        RECT 3385.420 2209.795 3386.390 2209.915 ;
        RECT 3383.500 2209.715 3383.670 2209.795 ;
        RECT 3386.220 2209.715 3386.390 2209.795 ;
        RECT 3387.410 2209.900 3388.290 2210.075 ;
        RECT 3387.410 2209.745 3387.580 2209.900 ;
        RECT 3383.500 2209.285 3383.670 2209.545 ;
        RECT 3386.220 2209.285 3386.390 2209.545 ;
        RECT 3386.560 2209.415 3387.580 2209.745 ;
        RECT 3383.500 2209.255 3384.470 2209.285 ;
        RECT 3383.670 2209.085 3384.470 2209.255 ;
        RECT 3383.500 2208.955 3384.470 2209.085 ;
        RECT 3385.070 2209.255 3386.390 2209.285 ;
        RECT 3385.070 2209.085 3386.220 2209.255 ;
        RECT 3386.390 2209.085 3387.190 2209.245 ;
        RECT 3385.070 2209.075 3387.190 2209.085 ;
        RECT 3385.070 2208.955 3386.390 2209.075 ;
        RECT 3383.500 2208.795 3383.670 2208.955 ;
        RECT 3386.220 2208.795 3386.390 2208.955 ;
        RECT 3387.410 2208.905 3387.580 2209.415 ;
        RECT 3383.500 2208.395 3383.670 2208.625 ;
        RECT 3386.220 2208.395 3386.390 2208.625 ;
        RECT 3386.560 2208.575 3387.580 2208.905 ;
        RECT 3388.120 2209.665 3388.290 2209.900 ;
        RECT 3388.460 2210.005 3388.940 2210.165 ;
        RECT 3388.460 2209.835 3389.110 2210.005 ;
        RECT 3388.940 2209.715 3389.110 2209.835 ;
        RECT 3388.120 2209.495 3388.765 2209.665 ;
        RECT 3388.120 2208.825 3388.290 2209.495 ;
        RECT 3388.940 2209.325 3389.110 2209.545 ;
        RECT 3388.460 2209.255 3389.110 2209.325 ;
        RECT 3388.460 2209.085 3388.940 2209.255 ;
        RECT 3388.460 2208.995 3389.110 2209.085 ;
        RECT 3388.120 2208.655 3388.770 2208.825 ;
        RECT 3388.940 2208.795 3389.110 2208.995 ;
        RECT 3388.940 2208.395 3389.110 2208.625 ;
        RECT 3383.500 2208.335 3384.395 2208.395 ;
        RECT 3383.670 2208.165 3384.395 2208.335 ;
        RECT 3383.500 2208.105 3384.395 2208.165 ;
        RECT 3385.055 2208.335 3387.555 2208.395 ;
        RECT 3385.055 2208.165 3386.220 2208.335 ;
        RECT 3386.390 2208.165 3387.555 2208.335 ;
        RECT 3385.055 2208.105 3387.555 2208.165 ;
        RECT 3388.215 2208.335 3389.110 2208.395 ;
        RECT 3388.215 2208.165 3388.940 2208.335 ;
        RECT 3388.215 2208.105 3389.110 2208.165 ;
        RECT 3383.500 2207.875 3383.670 2208.105 ;
        RECT 3383.500 2207.505 3383.670 2207.705 ;
        RECT 3383.840 2207.675 3384.490 2207.845 ;
        RECT 3383.500 2207.415 3384.150 2207.505 ;
        RECT 3383.670 2207.245 3384.150 2207.415 ;
        RECT 3383.500 2207.175 3384.150 2207.245 ;
        RECT 3383.500 2206.955 3383.670 2207.175 ;
        RECT 3384.320 2207.005 3384.490 2207.675 ;
        RECT 3383.845 2206.835 3384.490 2207.005 ;
        RECT 3383.500 2206.665 3383.670 2206.785 ;
        RECT 3383.500 2206.495 3384.150 2206.665 ;
        RECT 3383.670 2206.335 3384.150 2206.495 ;
        RECT 3384.320 2206.600 3384.490 2206.835 ;
        RECT 3385.030 2207.595 3386.050 2207.925 ;
        RECT 3386.220 2207.875 3386.390 2208.105 ;
        RECT 3388.940 2207.875 3389.110 2208.105 ;
        RECT 3385.030 2207.085 3385.200 2207.595 ;
        RECT 3386.220 2207.545 3386.390 2207.705 ;
        RECT 3388.940 2207.545 3389.110 2207.705 ;
        RECT 3386.220 2207.425 3387.540 2207.545 ;
        RECT 3385.420 2207.415 3387.540 2207.425 ;
        RECT 3385.420 2207.255 3386.220 2207.415 ;
        RECT 3386.390 2207.245 3387.540 2207.415 ;
        RECT 3386.220 2207.215 3387.540 2207.245 ;
        RECT 3388.140 2207.415 3389.110 2207.545 ;
        RECT 3388.140 2207.245 3388.940 2207.415 ;
        RECT 3388.140 2207.215 3389.110 2207.245 ;
        RECT 3385.030 2206.755 3386.050 2207.085 ;
        RECT 3386.220 2206.955 3386.390 2207.215 ;
        RECT 3388.940 2206.955 3389.110 2207.215 ;
        RECT 3385.030 2206.600 3385.200 2206.755 ;
        RECT 3384.320 2206.425 3385.200 2206.600 ;
        RECT 3386.220 2206.705 3386.390 2206.785 ;
        RECT 3388.940 2206.705 3389.110 2206.785 ;
        RECT 3386.220 2206.585 3387.190 2206.705 ;
        RECT 3385.420 2206.495 3387.190 2206.585 ;
        RECT 3383.500 2206.035 3383.670 2206.325 ;
        RECT 3383.500 2205.825 3383.670 2205.865 ;
        RECT 3383.500 2205.575 3384.150 2205.825 ;
        RECT 3383.670 2205.495 3384.150 2205.575 ;
        RECT 3383.500 2205.115 3383.670 2205.405 ;
        RECT 3383.670 2204.945 3384.150 2204.985 ;
        RECT 3383.500 2204.655 3384.150 2204.945 ;
        RECT 3383.500 2204.195 3383.670 2204.485 ;
        RECT 3383.670 2204.025 3384.150 2204.145 ;
        RECT 3383.500 2203.815 3384.150 2204.025 ;
        RECT 3384.660 2203.975 3384.830 2206.425 ;
        RECT 3385.420 2206.415 3386.220 2206.495 ;
        RECT 3386.390 2206.375 3387.190 2206.495 ;
        RECT 3386.220 2206.035 3386.390 2206.325 ;
        RECT 3386.220 2205.825 3387.190 2205.865 ;
        RECT 3385.420 2205.575 3387.190 2205.825 ;
        RECT 3385.420 2205.495 3386.220 2205.575 ;
        RECT 3386.390 2205.535 3387.190 2205.575 ;
        RECT 3386.220 2205.115 3386.390 2205.405 ;
        RECT 3385.420 2204.945 3386.220 2204.985 ;
        RECT 3386.390 2204.945 3387.190 2205.025 ;
        RECT 3385.420 2204.695 3387.190 2204.945 ;
        RECT 3385.420 2204.655 3386.390 2204.695 ;
        RECT 3386.220 2204.195 3386.390 2204.485 ;
        RECT 3385.420 2204.025 3386.220 2204.145 ;
        RECT 3386.390 2204.025 3387.190 2204.105 ;
        RECT 3387.780 2204.095 3387.950 2206.545 ;
        RECT 3388.460 2206.495 3389.110 2206.705 ;
        RECT 3388.460 2206.375 3388.940 2206.495 ;
        RECT 3388.940 2206.035 3389.110 2206.325 ;
        RECT 3388.460 2205.575 3389.110 2205.865 ;
        RECT 3388.460 2205.535 3388.940 2205.575 ;
        RECT 3388.940 2205.115 3389.110 2205.405 ;
        RECT 3388.460 2204.945 3388.940 2205.025 ;
        RECT 3388.460 2204.695 3389.110 2204.945 ;
        RECT 3388.940 2204.655 3389.110 2204.695 ;
        RECT 3388.940 2204.195 3389.110 2204.485 ;
        RECT 3385.420 2203.935 3387.190 2204.025 ;
        RECT 3385.420 2203.815 3386.390 2203.935 ;
        RECT 3383.500 2203.735 3383.670 2203.815 ;
        RECT 3386.220 2203.735 3386.390 2203.815 ;
        RECT 3387.410 2203.920 3388.290 2204.095 ;
        RECT 3387.410 2203.765 3387.580 2203.920 ;
        RECT 3383.500 2203.305 3383.670 2203.565 ;
        RECT 3386.220 2203.305 3386.390 2203.565 ;
        RECT 3386.560 2203.435 3387.580 2203.765 ;
        RECT 3383.500 2203.275 3384.470 2203.305 ;
        RECT 3383.670 2203.105 3384.470 2203.275 ;
        RECT 3383.500 2202.975 3384.470 2203.105 ;
        RECT 3385.070 2203.275 3386.390 2203.305 ;
        RECT 3385.070 2203.105 3386.220 2203.275 ;
        RECT 3386.390 2203.105 3387.190 2203.265 ;
        RECT 3385.070 2203.095 3387.190 2203.105 ;
        RECT 3385.070 2202.975 3386.390 2203.095 ;
        RECT 3383.500 2202.815 3383.670 2202.975 ;
        RECT 3386.220 2202.815 3386.390 2202.975 ;
        RECT 3387.410 2202.925 3387.580 2203.435 ;
        RECT 3383.500 2202.415 3383.670 2202.645 ;
        RECT 3386.220 2202.415 3386.390 2202.645 ;
        RECT 3386.560 2202.595 3387.580 2202.925 ;
        RECT 3388.120 2203.685 3388.290 2203.920 ;
        RECT 3388.460 2204.025 3388.940 2204.185 ;
        RECT 3388.460 2203.855 3389.110 2204.025 ;
        RECT 3388.940 2203.735 3389.110 2203.855 ;
        RECT 3388.120 2203.515 3388.765 2203.685 ;
        RECT 3388.120 2202.845 3388.290 2203.515 ;
        RECT 3388.940 2203.345 3389.110 2203.565 ;
        RECT 3388.460 2203.275 3389.110 2203.345 ;
        RECT 3388.460 2203.105 3388.940 2203.275 ;
        RECT 3388.460 2203.015 3389.110 2203.105 ;
        RECT 3388.120 2202.675 3388.770 2202.845 ;
        RECT 3388.940 2202.815 3389.110 2203.015 ;
        RECT 3388.940 2202.415 3389.110 2202.645 ;
        RECT 3383.500 2202.355 3384.395 2202.415 ;
        RECT 3383.670 2202.185 3384.395 2202.355 ;
        RECT 3383.500 2202.125 3384.395 2202.185 ;
        RECT 3385.055 2202.355 3387.555 2202.415 ;
        RECT 3385.055 2202.185 3386.220 2202.355 ;
        RECT 3386.390 2202.185 3387.555 2202.355 ;
        RECT 3385.055 2202.125 3387.555 2202.185 ;
        RECT 3388.215 2202.355 3389.110 2202.415 ;
        RECT 3388.215 2202.185 3388.940 2202.355 ;
        RECT 3388.215 2202.125 3389.110 2202.185 ;
        RECT 3383.500 2201.895 3383.670 2202.125 ;
        RECT 3383.500 2201.525 3383.670 2201.725 ;
        RECT 3383.840 2201.695 3384.490 2201.865 ;
        RECT 3383.500 2201.435 3384.150 2201.525 ;
        RECT 3383.670 2201.265 3384.150 2201.435 ;
        RECT 3383.500 2201.195 3384.150 2201.265 ;
        RECT 3383.500 2200.975 3383.670 2201.195 ;
        RECT 3384.320 2201.025 3384.490 2201.695 ;
        RECT 3383.845 2200.855 3384.490 2201.025 ;
        RECT 3383.500 2200.685 3383.670 2200.805 ;
        RECT 3383.500 2200.515 3384.150 2200.685 ;
        RECT 3383.670 2200.355 3384.150 2200.515 ;
        RECT 3384.320 2200.620 3384.490 2200.855 ;
        RECT 3385.030 2201.615 3386.050 2201.945 ;
        RECT 3386.220 2201.895 3386.390 2202.125 ;
        RECT 3388.940 2201.895 3389.110 2202.125 ;
        RECT 3385.030 2201.105 3385.200 2201.615 ;
        RECT 3386.220 2201.565 3386.390 2201.725 ;
        RECT 3388.940 2201.565 3389.110 2201.725 ;
        RECT 3386.220 2201.445 3387.540 2201.565 ;
        RECT 3385.420 2201.435 3387.540 2201.445 ;
        RECT 3385.420 2201.275 3386.220 2201.435 ;
        RECT 3386.390 2201.265 3387.540 2201.435 ;
        RECT 3386.220 2201.235 3387.540 2201.265 ;
        RECT 3388.140 2201.435 3389.110 2201.565 ;
        RECT 3388.140 2201.265 3388.940 2201.435 ;
        RECT 3388.140 2201.235 3389.110 2201.265 ;
        RECT 3385.030 2200.775 3386.050 2201.105 ;
        RECT 3386.220 2200.975 3386.390 2201.235 ;
        RECT 3388.940 2200.975 3389.110 2201.235 ;
        RECT 3385.030 2200.620 3385.200 2200.775 ;
        RECT 3384.320 2200.445 3385.200 2200.620 ;
        RECT 3386.220 2200.725 3386.390 2200.805 ;
        RECT 3388.940 2200.725 3389.110 2200.805 ;
        RECT 3386.220 2200.605 3387.190 2200.725 ;
        RECT 3385.420 2200.515 3387.190 2200.605 ;
        RECT 3383.500 2200.055 3383.670 2200.345 ;
        RECT 3383.500 2199.845 3383.670 2199.885 ;
        RECT 3383.500 2199.595 3384.150 2199.845 ;
        RECT 3383.670 2199.515 3384.150 2199.595 ;
        RECT 3383.500 2199.135 3383.670 2199.425 ;
        RECT 3383.670 2198.965 3384.150 2199.005 ;
        RECT 3383.500 2198.675 3384.150 2198.965 ;
        RECT 3383.500 2198.215 3383.670 2198.505 ;
        RECT 3383.670 2198.045 3384.150 2198.165 ;
        RECT 3383.500 2197.835 3384.150 2198.045 ;
        RECT 3384.660 2197.995 3384.830 2200.445 ;
        RECT 3385.420 2200.435 3386.220 2200.515 ;
        RECT 3386.390 2200.395 3387.190 2200.515 ;
        RECT 3386.220 2200.055 3386.390 2200.345 ;
        RECT 3386.220 2199.845 3387.190 2199.885 ;
        RECT 3385.420 2199.595 3387.190 2199.845 ;
        RECT 3385.420 2199.515 3386.220 2199.595 ;
        RECT 3386.390 2199.555 3387.190 2199.595 ;
        RECT 3386.220 2199.135 3386.390 2199.425 ;
        RECT 3385.420 2198.965 3386.220 2199.005 ;
        RECT 3386.390 2198.965 3387.190 2199.045 ;
        RECT 3385.420 2198.715 3387.190 2198.965 ;
        RECT 3385.420 2198.675 3386.390 2198.715 ;
        RECT 3386.220 2198.215 3386.390 2198.505 ;
        RECT 3385.420 2198.045 3386.220 2198.165 ;
        RECT 3386.390 2198.045 3387.190 2198.125 ;
        RECT 3387.780 2198.115 3387.950 2200.565 ;
        RECT 3388.460 2200.515 3389.110 2200.725 ;
        RECT 3388.460 2200.395 3388.940 2200.515 ;
        RECT 3388.940 2200.055 3389.110 2200.345 ;
        RECT 3388.460 2199.595 3389.110 2199.885 ;
        RECT 3388.460 2199.555 3388.940 2199.595 ;
        RECT 3388.940 2199.135 3389.110 2199.425 ;
        RECT 3388.460 2198.965 3388.940 2199.045 ;
        RECT 3388.460 2198.715 3389.110 2198.965 ;
        RECT 3388.940 2198.675 3389.110 2198.715 ;
        RECT 3388.940 2198.215 3389.110 2198.505 ;
        RECT 3385.420 2197.955 3387.190 2198.045 ;
        RECT 3385.420 2197.835 3386.390 2197.955 ;
        RECT 3383.500 2197.755 3383.670 2197.835 ;
        RECT 3386.220 2197.755 3386.390 2197.835 ;
        RECT 3387.410 2197.940 3388.290 2198.115 ;
        RECT 3387.410 2197.785 3387.580 2197.940 ;
        RECT 3383.500 2197.325 3383.670 2197.585 ;
        RECT 3386.220 2197.325 3386.390 2197.585 ;
        RECT 3386.560 2197.455 3387.580 2197.785 ;
        RECT 3383.500 2197.295 3384.470 2197.325 ;
        RECT 3383.670 2197.125 3384.470 2197.295 ;
        RECT 3383.500 2196.995 3384.470 2197.125 ;
        RECT 3385.070 2197.295 3386.390 2197.325 ;
        RECT 3385.070 2197.125 3386.220 2197.295 ;
        RECT 3386.390 2197.125 3387.190 2197.285 ;
        RECT 3385.070 2197.115 3387.190 2197.125 ;
        RECT 3385.070 2196.995 3386.390 2197.115 ;
        RECT 3383.500 2196.835 3383.670 2196.995 ;
        RECT 3386.220 2196.835 3386.390 2196.995 ;
        RECT 3387.410 2196.945 3387.580 2197.455 ;
        RECT 3383.500 2196.435 3383.670 2196.665 ;
        RECT 3386.220 2196.435 3386.390 2196.665 ;
        RECT 3386.560 2196.615 3387.580 2196.945 ;
        RECT 3388.120 2197.705 3388.290 2197.940 ;
        RECT 3388.460 2198.045 3388.940 2198.205 ;
        RECT 3388.460 2197.875 3389.110 2198.045 ;
        RECT 3388.940 2197.755 3389.110 2197.875 ;
        RECT 3388.120 2197.535 3388.765 2197.705 ;
        RECT 3388.120 2196.865 3388.290 2197.535 ;
        RECT 3388.940 2197.365 3389.110 2197.585 ;
        RECT 3388.460 2197.295 3389.110 2197.365 ;
        RECT 3388.460 2197.125 3388.940 2197.295 ;
        RECT 3388.460 2197.035 3389.110 2197.125 ;
        RECT 3388.120 2196.695 3388.770 2196.865 ;
        RECT 3388.940 2196.835 3389.110 2197.035 ;
        RECT 3388.940 2196.435 3389.110 2196.665 ;
        RECT 3383.500 2196.375 3384.395 2196.435 ;
        RECT 3383.670 2196.205 3384.395 2196.375 ;
        RECT 3383.500 2196.145 3384.395 2196.205 ;
        RECT 3385.055 2196.375 3387.555 2196.435 ;
        RECT 3385.055 2196.205 3386.220 2196.375 ;
        RECT 3386.390 2196.205 3387.555 2196.375 ;
        RECT 3385.055 2196.145 3387.555 2196.205 ;
        RECT 3388.215 2196.375 3389.110 2196.435 ;
        RECT 3388.215 2196.205 3388.940 2196.375 ;
        RECT 3388.215 2196.145 3389.110 2196.205 ;
        RECT 3383.500 2196.060 3383.670 2196.145 ;
        RECT 3386.220 2196.060 3386.390 2196.145 ;
        RECT 3388.940 2196.060 3389.110 2196.145 ;
        RECT 198.795 1733.080 198.965 1733.165 ;
        RECT 201.515 1733.080 201.685 1733.165 ;
        RECT 204.235 1733.080 204.405 1733.165 ;
        RECT 198.795 1733.020 199.690 1733.080 ;
        RECT 198.965 1732.850 199.690 1733.020 ;
        RECT 198.795 1732.790 199.690 1732.850 ;
        RECT 200.350 1733.020 202.850 1733.080 ;
        RECT 200.350 1732.850 201.515 1733.020 ;
        RECT 201.685 1732.850 202.850 1733.020 ;
        RECT 200.350 1732.790 202.850 1732.850 ;
        RECT 198.795 1732.560 198.965 1732.790 ;
        RECT 201.515 1732.560 201.685 1732.790 ;
        RECT 198.795 1732.230 198.965 1732.390 ;
        RECT 201.515 1732.230 201.685 1732.390 ;
        RECT 201.855 1732.280 202.875 1732.610 ;
        RECT 198.795 1732.100 199.765 1732.230 ;
        RECT 198.965 1731.930 199.765 1732.100 ;
        RECT 198.795 1731.900 199.765 1731.930 ;
        RECT 200.365 1732.110 201.685 1732.230 ;
        RECT 200.365 1732.100 202.485 1732.110 ;
        RECT 200.365 1731.930 201.515 1732.100 ;
        RECT 201.685 1731.940 202.485 1732.100 ;
        RECT 200.365 1731.900 201.685 1731.930 ;
        RECT 198.795 1731.640 198.965 1731.900 ;
      LAYER li1 ;
        RECT 199.135 1731.560 201.345 1731.730 ;
      LAYER li1 ;
        RECT 201.515 1731.640 201.685 1731.900 ;
        RECT 202.705 1731.770 202.875 1732.280 ;
      LAYER li1 ;
        RECT 199.615 1731.475 200.495 1731.560 ;
      LAYER li1 ;
        RECT 198.795 1731.390 198.965 1731.470 ;
        RECT 198.795 1731.180 199.445 1731.390 ;
        RECT 198.965 1731.060 199.445 1731.180 ;
        RECT 198.795 1730.720 198.965 1731.010 ;
      LAYER li1 ;
        RECT 199.615 1730.890 199.785 1731.475 ;
        RECT 199.135 1730.720 199.785 1730.890 ;
      LAYER li1 ;
        RECT 198.795 1730.260 199.445 1730.550 ;
        RECT 198.965 1730.220 199.445 1730.260 ;
        RECT 198.795 1729.800 198.965 1730.090 ;
      LAYER li1 ;
        RECT 199.615 1730.050 199.785 1730.720 ;
        RECT 199.135 1729.880 199.785 1730.050 ;
      LAYER li1 ;
        RECT 198.965 1729.630 199.445 1729.710 ;
        RECT 198.795 1729.380 199.445 1729.630 ;
        RECT 198.795 1729.340 198.965 1729.380 ;
      LAYER li1 ;
        RECT 199.615 1729.210 199.785 1729.880 ;
      LAYER li1 ;
        RECT 198.795 1728.880 198.965 1729.170 ;
      LAYER li1 ;
        RECT 199.135 1729.040 199.785 1729.210 ;
      LAYER li1 ;
        RECT 198.965 1728.710 199.445 1728.870 ;
        RECT 199.955 1728.780 200.125 1731.230 ;
      LAYER li1 ;
        RECT 200.325 1730.890 200.495 1731.475 ;
      LAYER li1 ;
        RECT 201.515 1731.390 201.685 1731.470 ;
        RECT 201.855 1731.440 202.875 1731.770 ;
      LAYER li1 ;
        RECT 203.045 1731.465 203.245 1733.055 ;
      LAYER li1 ;
        RECT 203.510 1733.020 204.405 1733.080 ;
        RECT 203.510 1732.850 204.235 1733.020 ;
        RECT 203.510 1732.790 204.405 1732.850 ;
        RECT 204.235 1732.560 204.405 1732.790 ;
        RECT 203.415 1732.360 204.065 1732.530 ;
        RECT 203.415 1731.690 203.585 1732.360 ;
        RECT 204.235 1732.190 204.405 1732.390 ;
        RECT 203.755 1732.100 204.405 1732.190 ;
        RECT 203.755 1731.930 204.235 1732.100 ;
        RECT 203.755 1731.860 204.405 1731.930 ;
        RECT 203.415 1731.520 204.060 1731.690 ;
        RECT 204.235 1731.640 204.405 1731.860 ;
        RECT 200.715 1731.270 201.685 1731.390 ;
        RECT 202.705 1731.285 202.875 1731.440 ;
        RECT 203.415 1731.285 203.585 1731.520 ;
        RECT 204.235 1731.350 204.405 1731.470 ;
        RECT 200.715 1731.180 202.485 1731.270 ;
        RECT 200.715 1731.060 201.515 1731.180 ;
        RECT 201.685 1731.100 202.485 1731.180 ;
        RECT 202.705 1731.110 203.585 1731.285 ;
        RECT 203.755 1731.180 204.405 1731.350 ;
      LAYER li1 ;
        RECT 200.325 1730.720 201.345 1730.890 ;
      LAYER li1 ;
        RECT 201.515 1730.720 201.685 1731.010 ;
      LAYER li1 ;
        RECT 200.325 1730.050 200.495 1730.720 ;
        RECT 201.855 1730.680 202.875 1730.850 ;
      LAYER li1 ;
        RECT 200.715 1730.510 201.685 1730.550 ;
        RECT 200.715 1730.260 202.485 1730.510 ;
        RECT 200.715 1730.220 201.515 1730.260 ;
        RECT 201.685 1730.180 202.485 1730.260 ;
      LAYER li1 ;
        RECT 200.325 1729.880 201.345 1730.050 ;
        RECT 200.325 1729.210 200.495 1729.880 ;
      LAYER li1 ;
        RECT 201.515 1729.800 201.685 1730.090 ;
      LAYER li1 ;
        RECT 202.705 1730.010 202.875 1730.680 ;
        RECT 201.855 1729.840 202.875 1730.010 ;
      LAYER li1 ;
        RECT 200.715 1729.630 201.515 1729.710 ;
        RECT 201.685 1729.630 202.485 1729.670 ;
        RECT 200.715 1729.380 202.485 1729.630 ;
        RECT 201.515 1729.340 202.485 1729.380 ;
      LAYER li1 ;
        RECT 200.325 1729.040 201.345 1729.210 ;
        RECT 202.705 1729.170 202.875 1729.840 ;
      LAYER li1 ;
        RECT 201.515 1728.880 201.685 1729.170 ;
      LAYER li1 ;
        RECT 201.855 1729.000 202.875 1729.170 ;
      LAYER li1 ;
        RECT 198.795 1728.540 199.445 1728.710 ;
        RECT 199.615 1728.605 200.495 1728.780 ;
        RECT 200.715 1728.710 201.515 1728.790 ;
        RECT 201.685 1728.710 202.485 1728.830 ;
        RECT 200.715 1728.620 202.485 1728.710 ;
        RECT 198.795 1728.420 198.965 1728.540 ;
        RECT 199.615 1728.370 199.785 1728.605 ;
        RECT 200.325 1728.450 200.495 1728.605 ;
        RECT 201.515 1728.500 202.485 1728.620 ;
        RECT 198.795 1728.030 198.965 1728.250 ;
        RECT 199.140 1728.200 199.785 1728.370 ;
        RECT 198.795 1727.960 199.445 1728.030 ;
        RECT 198.965 1727.790 199.445 1727.960 ;
        RECT 198.795 1727.700 199.445 1727.790 ;
        RECT 198.795 1727.500 198.965 1727.700 ;
        RECT 199.615 1727.530 199.785 1728.200 ;
        RECT 199.135 1727.360 199.785 1727.530 ;
        RECT 198.795 1727.100 198.965 1727.330 ;
      LAYER li1 ;
        RECT 199.955 1727.325 200.155 1728.425 ;
      LAYER li1 ;
        RECT 200.325 1728.120 201.345 1728.450 ;
        RECT 201.515 1728.420 201.685 1728.500 ;
      LAYER li1 ;
        RECT 202.705 1728.415 202.875 1729.000 ;
      LAYER li1 ;
        RECT 203.075 1728.660 203.245 1731.110 ;
        RECT 203.755 1731.020 204.235 1731.180 ;
      LAYER li1 ;
        RECT 203.415 1730.680 204.065 1730.850 ;
      LAYER li1 ;
        RECT 204.235 1730.720 204.405 1731.010 ;
      LAYER li1 ;
        RECT 203.415 1730.010 203.585 1730.680 ;
      LAYER li1 ;
        RECT 204.235 1730.510 204.405 1730.550 ;
        RECT 203.755 1730.260 204.405 1730.510 ;
        RECT 203.755 1730.180 204.235 1730.260 ;
      LAYER li1 ;
        RECT 203.415 1729.840 204.065 1730.010 ;
        RECT 203.415 1729.170 203.585 1729.840 ;
      LAYER li1 ;
        RECT 204.235 1729.800 204.405 1730.090 ;
        RECT 203.755 1729.630 204.235 1729.670 ;
        RECT 203.755 1729.340 204.405 1729.630 ;
      LAYER li1 ;
        RECT 203.415 1729.000 204.065 1729.170 ;
        RECT 203.415 1728.415 203.585 1729.000 ;
      LAYER li1 ;
        RECT 204.235 1728.880 204.405 1729.170 ;
        RECT 203.755 1728.710 204.235 1728.830 ;
        RECT 203.755 1728.500 204.405 1728.710 ;
        RECT 204.235 1728.420 204.405 1728.500 ;
      LAYER li1 ;
        RECT 202.705 1728.330 203.585 1728.415 ;
      LAYER li1 ;
        RECT 200.325 1727.610 200.495 1728.120 ;
        RECT 201.515 1727.990 201.685 1728.250 ;
      LAYER li1 ;
        RECT 201.855 1728.160 204.065 1728.330 ;
      LAYER li1 ;
        RECT 204.235 1727.990 204.405 1728.250 ;
        RECT 201.515 1727.960 202.835 1727.990 ;
        RECT 200.715 1727.790 201.515 1727.950 ;
        RECT 201.685 1727.790 202.835 1727.960 ;
        RECT 200.715 1727.780 202.835 1727.790 ;
        RECT 201.515 1727.660 202.835 1727.780 ;
        RECT 203.435 1727.960 204.405 1727.990 ;
        RECT 203.435 1727.790 204.235 1727.960 ;
        RECT 203.435 1727.660 204.405 1727.790 ;
        RECT 200.325 1727.280 201.345 1727.610 ;
        RECT 201.515 1727.500 201.685 1727.660 ;
        RECT 204.235 1727.500 204.405 1727.660 ;
        RECT 201.515 1727.100 201.685 1727.330 ;
        RECT 204.235 1727.100 204.405 1727.330 ;
        RECT 198.795 1727.040 199.690 1727.100 ;
        RECT 198.965 1726.870 199.690 1727.040 ;
        RECT 198.795 1726.810 199.690 1726.870 ;
        RECT 200.350 1727.040 202.850 1727.100 ;
        RECT 200.350 1726.870 201.515 1727.040 ;
        RECT 201.685 1726.870 202.850 1727.040 ;
        RECT 200.350 1726.810 202.850 1726.870 ;
        RECT 198.795 1726.580 198.965 1726.810 ;
        RECT 201.515 1726.580 201.685 1726.810 ;
        RECT 198.795 1726.250 198.965 1726.410 ;
        RECT 201.515 1726.250 201.685 1726.410 ;
        RECT 201.855 1726.300 202.875 1726.630 ;
        RECT 198.795 1726.120 199.765 1726.250 ;
        RECT 198.965 1725.950 199.765 1726.120 ;
        RECT 198.795 1725.920 199.765 1725.950 ;
        RECT 200.365 1726.130 201.685 1726.250 ;
        RECT 200.365 1726.120 202.485 1726.130 ;
        RECT 200.365 1725.950 201.515 1726.120 ;
        RECT 201.685 1725.960 202.485 1726.120 ;
        RECT 200.365 1725.920 201.685 1725.950 ;
        RECT 198.795 1725.660 198.965 1725.920 ;
      LAYER li1 ;
        RECT 199.135 1725.580 201.345 1725.750 ;
      LAYER li1 ;
        RECT 201.515 1725.660 201.685 1725.920 ;
        RECT 202.705 1725.790 202.875 1726.300 ;
      LAYER li1 ;
        RECT 199.615 1725.495 200.495 1725.580 ;
      LAYER li1 ;
        RECT 198.795 1725.410 198.965 1725.490 ;
        RECT 198.795 1725.200 199.445 1725.410 ;
        RECT 198.965 1725.080 199.445 1725.200 ;
        RECT 198.795 1724.740 198.965 1725.030 ;
      LAYER li1 ;
        RECT 199.615 1724.910 199.785 1725.495 ;
        RECT 199.135 1724.740 199.785 1724.910 ;
      LAYER li1 ;
        RECT 198.795 1724.280 199.445 1724.570 ;
        RECT 198.965 1724.240 199.445 1724.280 ;
        RECT 198.795 1723.820 198.965 1724.110 ;
      LAYER li1 ;
        RECT 199.615 1724.070 199.785 1724.740 ;
        RECT 199.135 1723.900 199.785 1724.070 ;
      LAYER li1 ;
        RECT 198.965 1723.650 199.445 1723.730 ;
        RECT 198.795 1723.400 199.445 1723.650 ;
        RECT 198.795 1723.360 198.965 1723.400 ;
      LAYER li1 ;
        RECT 199.615 1723.230 199.785 1723.900 ;
      LAYER li1 ;
        RECT 198.795 1722.900 198.965 1723.190 ;
      LAYER li1 ;
        RECT 199.135 1723.060 199.785 1723.230 ;
      LAYER li1 ;
        RECT 198.965 1722.730 199.445 1722.890 ;
        RECT 199.955 1722.800 200.125 1725.250 ;
      LAYER li1 ;
        RECT 200.325 1724.910 200.495 1725.495 ;
      LAYER li1 ;
        RECT 201.515 1725.410 201.685 1725.490 ;
        RECT 201.855 1725.460 202.875 1725.790 ;
      LAYER li1 ;
        RECT 203.045 1725.485 203.245 1727.075 ;
      LAYER li1 ;
        RECT 203.510 1727.040 204.405 1727.100 ;
        RECT 203.510 1726.870 204.235 1727.040 ;
        RECT 203.510 1726.810 204.405 1726.870 ;
        RECT 204.235 1726.580 204.405 1726.810 ;
        RECT 203.415 1726.380 204.065 1726.550 ;
        RECT 203.415 1725.710 203.585 1726.380 ;
        RECT 204.235 1726.210 204.405 1726.410 ;
        RECT 203.755 1726.120 204.405 1726.210 ;
        RECT 203.755 1725.950 204.235 1726.120 ;
        RECT 203.755 1725.880 204.405 1725.950 ;
        RECT 203.415 1725.540 204.060 1725.710 ;
        RECT 204.235 1725.660 204.405 1725.880 ;
        RECT 200.715 1725.290 201.685 1725.410 ;
        RECT 202.705 1725.305 202.875 1725.460 ;
        RECT 203.415 1725.305 203.585 1725.540 ;
        RECT 204.235 1725.370 204.405 1725.490 ;
        RECT 200.715 1725.200 202.485 1725.290 ;
        RECT 200.715 1725.080 201.515 1725.200 ;
        RECT 201.685 1725.120 202.485 1725.200 ;
        RECT 202.705 1725.130 203.585 1725.305 ;
        RECT 203.755 1725.200 204.405 1725.370 ;
      LAYER li1 ;
        RECT 200.325 1724.740 201.345 1724.910 ;
      LAYER li1 ;
        RECT 201.515 1724.740 201.685 1725.030 ;
      LAYER li1 ;
        RECT 200.325 1724.070 200.495 1724.740 ;
        RECT 201.855 1724.700 202.875 1724.870 ;
      LAYER li1 ;
        RECT 200.715 1724.530 201.685 1724.570 ;
        RECT 200.715 1724.280 202.485 1724.530 ;
        RECT 200.715 1724.240 201.515 1724.280 ;
        RECT 201.685 1724.200 202.485 1724.280 ;
      LAYER li1 ;
        RECT 200.325 1723.900 201.345 1724.070 ;
        RECT 200.325 1723.230 200.495 1723.900 ;
      LAYER li1 ;
        RECT 201.515 1723.820 201.685 1724.110 ;
      LAYER li1 ;
        RECT 202.705 1724.030 202.875 1724.700 ;
        RECT 201.855 1723.860 202.875 1724.030 ;
      LAYER li1 ;
        RECT 200.715 1723.650 201.515 1723.730 ;
        RECT 201.685 1723.650 202.485 1723.690 ;
        RECT 200.715 1723.400 202.485 1723.650 ;
        RECT 201.515 1723.360 202.485 1723.400 ;
      LAYER li1 ;
        RECT 200.325 1723.060 201.345 1723.230 ;
        RECT 202.705 1723.190 202.875 1723.860 ;
      LAYER li1 ;
        RECT 201.515 1722.900 201.685 1723.190 ;
      LAYER li1 ;
        RECT 201.855 1723.020 202.875 1723.190 ;
      LAYER li1 ;
        RECT 198.795 1722.560 199.445 1722.730 ;
        RECT 199.615 1722.625 200.495 1722.800 ;
        RECT 200.715 1722.730 201.515 1722.810 ;
        RECT 201.685 1722.730 202.485 1722.850 ;
        RECT 200.715 1722.640 202.485 1722.730 ;
        RECT 198.795 1722.440 198.965 1722.560 ;
        RECT 199.615 1722.390 199.785 1722.625 ;
        RECT 200.325 1722.470 200.495 1722.625 ;
        RECT 201.515 1722.520 202.485 1722.640 ;
        RECT 198.795 1722.050 198.965 1722.270 ;
        RECT 199.140 1722.220 199.785 1722.390 ;
        RECT 198.795 1721.980 199.445 1722.050 ;
        RECT 198.965 1721.810 199.445 1721.980 ;
        RECT 198.795 1721.720 199.445 1721.810 ;
        RECT 198.795 1721.520 198.965 1721.720 ;
        RECT 199.615 1721.550 199.785 1722.220 ;
        RECT 199.135 1721.380 199.785 1721.550 ;
        RECT 198.795 1721.120 198.965 1721.350 ;
      LAYER li1 ;
        RECT 199.955 1721.345 200.155 1722.445 ;
      LAYER li1 ;
        RECT 200.325 1722.140 201.345 1722.470 ;
        RECT 201.515 1722.440 201.685 1722.520 ;
      LAYER li1 ;
        RECT 202.705 1722.435 202.875 1723.020 ;
      LAYER li1 ;
        RECT 203.075 1722.680 203.245 1725.130 ;
        RECT 203.755 1725.040 204.235 1725.200 ;
      LAYER li1 ;
        RECT 203.415 1724.700 204.065 1724.870 ;
      LAYER li1 ;
        RECT 204.235 1724.740 204.405 1725.030 ;
      LAYER li1 ;
        RECT 203.415 1724.030 203.585 1724.700 ;
      LAYER li1 ;
        RECT 204.235 1724.530 204.405 1724.570 ;
        RECT 203.755 1724.280 204.405 1724.530 ;
        RECT 203.755 1724.200 204.235 1724.280 ;
      LAYER li1 ;
        RECT 203.415 1723.860 204.065 1724.030 ;
        RECT 203.415 1723.190 203.585 1723.860 ;
      LAYER li1 ;
        RECT 204.235 1723.820 204.405 1724.110 ;
        RECT 203.755 1723.650 204.235 1723.690 ;
        RECT 203.755 1723.360 204.405 1723.650 ;
      LAYER li1 ;
        RECT 203.415 1723.020 204.065 1723.190 ;
        RECT 203.415 1722.435 203.585 1723.020 ;
      LAYER li1 ;
        RECT 204.235 1722.900 204.405 1723.190 ;
        RECT 203.755 1722.730 204.235 1722.850 ;
        RECT 203.755 1722.520 204.405 1722.730 ;
        RECT 204.235 1722.440 204.405 1722.520 ;
      LAYER li1 ;
        RECT 202.705 1722.350 203.585 1722.435 ;
      LAYER li1 ;
        RECT 200.325 1721.630 200.495 1722.140 ;
        RECT 201.515 1722.010 201.685 1722.270 ;
      LAYER li1 ;
        RECT 201.855 1722.180 204.065 1722.350 ;
      LAYER li1 ;
        RECT 204.235 1722.010 204.405 1722.270 ;
        RECT 201.515 1721.980 202.835 1722.010 ;
        RECT 200.715 1721.810 201.515 1721.970 ;
        RECT 201.685 1721.810 202.835 1721.980 ;
        RECT 200.715 1721.800 202.835 1721.810 ;
        RECT 201.515 1721.680 202.835 1721.800 ;
        RECT 203.435 1721.980 204.405 1722.010 ;
        RECT 203.435 1721.810 204.235 1721.980 ;
        RECT 203.435 1721.680 204.405 1721.810 ;
        RECT 200.325 1721.300 201.345 1721.630 ;
        RECT 201.515 1721.520 201.685 1721.680 ;
        RECT 204.235 1721.520 204.405 1721.680 ;
        RECT 201.515 1721.120 201.685 1721.350 ;
        RECT 204.235 1721.120 204.405 1721.350 ;
        RECT 198.795 1721.060 199.690 1721.120 ;
        RECT 198.965 1720.890 199.690 1721.060 ;
        RECT 198.795 1720.830 199.690 1720.890 ;
        RECT 200.350 1721.060 202.850 1721.120 ;
        RECT 200.350 1720.890 201.515 1721.060 ;
        RECT 201.685 1720.890 202.850 1721.060 ;
        RECT 200.350 1720.830 202.850 1720.890 ;
        RECT 198.795 1720.600 198.965 1720.830 ;
        RECT 201.515 1720.600 201.685 1720.830 ;
        RECT 198.795 1720.270 198.965 1720.430 ;
        RECT 201.515 1720.270 201.685 1720.430 ;
        RECT 201.855 1720.320 202.875 1720.650 ;
        RECT 198.795 1720.140 199.765 1720.270 ;
        RECT 198.965 1719.970 199.765 1720.140 ;
        RECT 198.795 1719.940 199.765 1719.970 ;
        RECT 200.365 1720.150 201.685 1720.270 ;
        RECT 200.365 1720.140 202.485 1720.150 ;
        RECT 200.365 1719.970 201.515 1720.140 ;
        RECT 201.685 1719.980 202.485 1720.140 ;
        RECT 200.365 1719.940 201.685 1719.970 ;
        RECT 198.795 1719.680 198.965 1719.940 ;
      LAYER li1 ;
        RECT 199.135 1719.600 201.345 1719.770 ;
      LAYER li1 ;
        RECT 201.515 1719.680 201.685 1719.940 ;
        RECT 202.705 1719.810 202.875 1720.320 ;
      LAYER li1 ;
        RECT 199.615 1719.515 200.495 1719.600 ;
      LAYER li1 ;
        RECT 198.795 1719.430 198.965 1719.510 ;
        RECT 198.795 1719.220 199.445 1719.430 ;
        RECT 198.965 1719.100 199.445 1719.220 ;
        RECT 198.795 1718.760 198.965 1719.050 ;
      LAYER li1 ;
        RECT 199.615 1718.930 199.785 1719.515 ;
        RECT 199.135 1718.760 199.785 1718.930 ;
      LAYER li1 ;
        RECT 198.795 1718.300 199.445 1718.590 ;
        RECT 198.965 1718.260 199.445 1718.300 ;
        RECT 198.795 1717.840 198.965 1718.130 ;
      LAYER li1 ;
        RECT 199.615 1718.090 199.785 1718.760 ;
        RECT 199.135 1717.920 199.785 1718.090 ;
      LAYER li1 ;
        RECT 198.965 1717.670 199.445 1717.750 ;
        RECT 198.795 1717.420 199.445 1717.670 ;
        RECT 198.795 1717.380 198.965 1717.420 ;
      LAYER li1 ;
        RECT 199.615 1717.250 199.785 1717.920 ;
      LAYER li1 ;
        RECT 198.795 1716.920 198.965 1717.210 ;
      LAYER li1 ;
        RECT 199.135 1717.080 199.785 1717.250 ;
      LAYER li1 ;
        RECT 198.965 1716.750 199.445 1716.910 ;
        RECT 199.955 1716.820 200.125 1719.270 ;
      LAYER li1 ;
        RECT 200.325 1718.930 200.495 1719.515 ;
      LAYER li1 ;
        RECT 201.515 1719.430 201.685 1719.510 ;
        RECT 201.855 1719.480 202.875 1719.810 ;
      LAYER li1 ;
        RECT 203.045 1719.505 203.245 1721.095 ;
      LAYER li1 ;
        RECT 203.510 1721.060 204.405 1721.120 ;
        RECT 203.510 1720.890 204.235 1721.060 ;
        RECT 203.510 1720.830 204.405 1720.890 ;
        RECT 204.235 1720.600 204.405 1720.830 ;
        RECT 203.415 1720.400 204.065 1720.570 ;
        RECT 203.415 1719.730 203.585 1720.400 ;
        RECT 204.235 1720.230 204.405 1720.430 ;
        RECT 203.755 1720.140 204.405 1720.230 ;
        RECT 203.755 1719.970 204.235 1720.140 ;
        RECT 203.755 1719.900 204.405 1719.970 ;
        RECT 203.415 1719.560 204.060 1719.730 ;
        RECT 204.235 1719.680 204.405 1719.900 ;
        RECT 200.715 1719.310 201.685 1719.430 ;
        RECT 202.705 1719.325 202.875 1719.480 ;
        RECT 203.415 1719.325 203.585 1719.560 ;
        RECT 204.235 1719.390 204.405 1719.510 ;
        RECT 200.715 1719.220 202.485 1719.310 ;
        RECT 200.715 1719.100 201.515 1719.220 ;
        RECT 201.685 1719.140 202.485 1719.220 ;
        RECT 202.705 1719.150 203.585 1719.325 ;
        RECT 203.755 1719.220 204.405 1719.390 ;
      LAYER li1 ;
        RECT 200.325 1718.760 201.345 1718.930 ;
      LAYER li1 ;
        RECT 201.515 1718.760 201.685 1719.050 ;
      LAYER li1 ;
        RECT 200.325 1718.090 200.495 1718.760 ;
        RECT 201.855 1718.720 202.875 1718.890 ;
      LAYER li1 ;
        RECT 200.715 1718.550 201.685 1718.590 ;
        RECT 200.715 1718.300 202.485 1718.550 ;
        RECT 200.715 1718.260 201.515 1718.300 ;
        RECT 201.685 1718.220 202.485 1718.300 ;
      LAYER li1 ;
        RECT 200.325 1717.920 201.345 1718.090 ;
        RECT 200.325 1717.250 200.495 1717.920 ;
      LAYER li1 ;
        RECT 201.515 1717.840 201.685 1718.130 ;
      LAYER li1 ;
        RECT 202.705 1718.050 202.875 1718.720 ;
        RECT 201.855 1717.880 202.875 1718.050 ;
      LAYER li1 ;
        RECT 200.715 1717.670 201.515 1717.750 ;
        RECT 201.685 1717.670 202.485 1717.710 ;
        RECT 200.715 1717.420 202.485 1717.670 ;
        RECT 201.515 1717.380 202.485 1717.420 ;
      LAYER li1 ;
        RECT 200.325 1717.080 201.345 1717.250 ;
        RECT 202.705 1717.210 202.875 1717.880 ;
      LAYER li1 ;
        RECT 201.515 1716.920 201.685 1717.210 ;
      LAYER li1 ;
        RECT 201.855 1717.040 202.875 1717.210 ;
      LAYER li1 ;
        RECT 198.795 1716.580 199.445 1716.750 ;
        RECT 199.615 1716.645 200.495 1716.820 ;
        RECT 200.715 1716.750 201.515 1716.830 ;
        RECT 201.685 1716.750 202.485 1716.870 ;
        RECT 200.715 1716.660 202.485 1716.750 ;
        RECT 198.795 1716.460 198.965 1716.580 ;
        RECT 199.615 1716.410 199.785 1716.645 ;
        RECT 200.325 1716.490 200.495 1716.645 ;
        RECT 201.515 1716.540 202.485 1716.660 ;
        RECT 198.795 1716.070 198.965 1716.290 ;
        RECT 199.140 1716.240 199.785 1716.410 ;
        RECT 198.795 1716.000 199.445 1716.070 ;
        RECT 198.965 1715.830 199.445 1716.000 ;
        RECT 198.795 1715.740 199.445 1715.830 ;
        RECT 198.795 1715.540 198.965 1715.740 ;
        RECT 199.615 1715.570 199.785 1716.240 ;
        RECT 199.135 1715.400 199.785 1715.570 ;
        RECT 198.795 1715.140 198.965 1715.370 ;
      LAYER li1 ;
        RECT 199.955 1715.365 200.155 1716.465 ;
      LAYER li1 ;
        RECT 200.325 1716.160 201.345 1716.490 ;
        RECT 201.515 1716.460 201.685 1716.540 ;
      LAYER li1 ;
        RECT 202.705 1716.455 202.875 1717.040 ;
      LAYER li1 ;
        RECT 203.075 1716.700 203.245 1719.150 ;
        RECT 203.755 1719.060 204.235 1719.220 ;
      LAYER li1 ;
        RECT 203.415 1718.720 204.065 1718.890 ;
      LAYER li1 ;
        RECT 204.235 1718.760 204.405 1719.050 ;
      LAYER li1 ;
        RECT 203.415 1718.050 203.585 1718.720 ;
      LAYER li1 ;
        RECT 204.235 1718.550 204.405 1718.590 ;
        RECT 203.755 1718.300 204.405 1718.550 ;
        RECT 203.755 1718.220 204.235 1718.300 ;
      LAYER li1 ;
        RECT 203.415 1717.880 204.065 1718.050 ;
        RECT 203.415 1717.210 203.585 1717.880 ;
      LAYER li1 ;
        RECT 204.235 1717.840 204.405 1718.130 ;
        RECT 203.755 1717.670 204.235 1717.710 ;
        RECT 203.755 1717.380 204.405 1717.670 ;
      LAYER li1 ;
        RECT 203.415 1717.040 204.065 1717.210 ;
        RECT 203.415 1716.455 203.585 1717.040 ;
      LAYER li1 ;
        RECT 204.235 1716.920 204.405 1717.210 ;
        RECT 203.755 1716.750 204.235 1716.870 ;
        RECT 203.755 1716.540 204.405 1716.750 ;
        RECT 204.235 1716.460 204.405 1716.540 ;
      LAYER li1 ;
        RECT 202.705 1716.370 203.585 1716.455 ;
      LAYER li1 ;
        RECT 200.325 1715.650 200.495 1716.160 ;
        RECT 201.515 1716.030 201.685 1716.290 ;
      LAYER li1 ;
        RECT 201.855 1716.200 204.065 1716.370 ;
      LAYER li1 ;
        RECT 204.235 1716.030 204.405 1716.290 ;
        RECT 201.515 1716.000 202.835 1716.030 ;
        RECT 200.715 1715.830 201.515 1715.990 ;
        RECT 201.685 1715.830 202.835 1716.000 ;
        RECT 200.715 1715.820 202.835 1715.830 ;
        RECT 201.515 1715.700 202.835 1715.820 ;
        RECT 203.435 1716.000 204.405 1716.030 ;
        RECT 203.435 1715.830 204.235 1716.000 ;
        RECT 203.435 1715.700 204.405 1715.830 ;
        RECT 200.325 1715.320 201.345 1715.650 ;
        RECT 201.515 1715.540 201.685 1715.700 ;
        RECT 204.235 1715.540 204.405 1715.700 ;
        RECT 201.515 1715.140 201.685 1715.370 ;
        RECT 204.235 1715.140 204.405 1715.370 ;
        RECT 198.795 1715.080 199.690 1715.140 ;
        RECT 198.965 1714.910 199.690 1715.080 ;
        RECT 198.795 1714.850 199.690 1714.910 ;
        RECT 200.350 1715.080 202.850 1715.140 ;
        RECT 200.350 1714.910 201.515 1715.080 ;
        RECT 201.685 1714.910 202.850 1715.080 ;
        RECT 200.350 1714.850 202.850 1714.910 ;
        RECT 198.795 1714.620 198.965 1714.850 ;
        RECT 201.515 1714.620 201.685 1714.850 ;
        RECT 198.795 1714.290 198.965 1714.450 ;
        RECT 201.515 1714.290 201.685 1714.450 ;
        RECT 201.855 1714.340 202.875 1714.670 ;
        RECT 198.795 1714.160 199.765 1714.290 ;
        RECT 198.965 1713.990 199.765 1714.160 ;
        RECT 198.795 1713.960 199.765 1713.990 ;
        RECT 200.365 1714.170 201.685 1714.290 ;
        RECT 200.365 1714.160 202.485 1714.170 ;
        RECT 200.365 1713.990 201.515 1714.160 ;
        RECT 201.685 1714.000 202.485 1714.160 ;
        RECT 200.365 1713.960 201.685 1713.990 ;
        RECT 198.795 1713.700 198.965 1713.960 ;
      LAYER li1 ;
        RECT 199.135 1713.620 201.345 1713.790 ;
      LAYER li1 ;
        RECT 201.515 1713.700 201.685 1713.960 ;
        RECT 202.705 1713.830 202.875 1714.340 ;
      LAYER li1 ;
        RECT 199.615 1713.535 200.495 1713.620 ;
      LAYER li1 ;
        RECT 198.795 1713.450 198.965 1713.530 ;
        RECT 198.795 1713.240 199.445 1713.450 ;
        RECT 198.965 1713.120 199.445 1713.240 ;
        RECT 198.795 1712.780 198.965 1713.070 ;
      LAYER li1 ;
        RECT 199.615 1712.950 199.785 1713.535 ;
        RECT 199.135 1712.780 199.785 1712.950 ;
      LAYER li1 ;
        RECT 198.795 1712.320 199.445 1712.610 ;
        RECT 198.965 1712.280 199.445 1712.320 ;
        RECT 198.795 1711.860 198.965 1712.150 ;
      LAYER li1 ;
        RECT 199.615 1712.110 199.785 1712.780 ;
        RECT 199.135 1711.940 199.785 1712.110 ;
      LAYER li1 ;
        RECT 198.965 1711.690 199.445 1711.770 ;
        RECT 198.795 1711.440 199.445 1711.690 ;
        RECT 198.795 1711.400 198.965 1711.440 ;
      LAYER li1 ;
        RECT 199.615 1711.270 199.785 1711.940 ;
      LAYER li1 ;
        RECT 198.795 1710.940 198.965 1711.230 ;
      LAYER li1 ;
        RECT 199.135 1711.100 199.785 1711.270 ;
      LAYER li1 ;
        RECT 198.965 1710.770 199.445 1710.930 ;
        RECT 199.955 1710.840 200.125 1713.290 ;
      LAYER li1 ;
        RECT 200.325 1712.950 200.495 1713.535 ;
      LAYER li1 ;
        RECT 201.515 1713.450 201.685 1713.530 ;
        RECT 201.855 1713.500 202.875 1713.830 ;
      LAYER li1 ;
        RECT 203.045 1713.525 203.245 1715.115 ;
      LAYER li1 ;
        RECT 203.510 1715.080 204.405 1715.140 ;
        RECT 203.510 1714.910 204.235 1715.080 ;
        RECT 203.510 1714.850 204.405 1714.910 ;
        RECT 204.235 1714.620 204.405 1714.850 ;
        RECT 203.415 1714.420 204.065 1714.590 ;
        RECT 203.415 1713.750 203.585 1714.420 ;
        RECT 204.235 1714.250 204.405 1714.450 ;
        RECT 203.755 1714.160 204.405 1714.250 ;
        RECT 203.755 1713.990 204.235 1714.160 ;
        RECT 203.755 1713.920 204.405 1713.990 ;
        RECT 203.415 1713.580 204.060 1713.750 ;
        RECT 204.235 1713.700 204.405 1713.920 ;
        RECT 200.715 1713.330 201.685 1713.450 ;
        RECT 202.705 1713.345 202.875 1713.500 ;
        RECT 203.415 1713.345 203.585 1713.580 ;
        RECT 204.235 1713.410 204.405 1713.530 ;
        RECT 200.715 1713.240 202.485 1713.330 ;
        RECT 200.715 1713.120 201.515 1713.240 ;
        RECT 201.685 1713.160 202.485 1713.240 ;
        RECT 202.705 1713.170 203.585 1713.345 ;
        RECT 203.755 1713.240 204.405 1713.410 ;
      LAYER li1 ;
        RECT 200.325 1712.780 201.345 1712.950 ;
      LAYER li1 ;
        RECT 201.515 1712.780 201.685 1713.070 ;
      LAYER li1 ;
        RECT 200.325 1712.110 200.495 1712.780 ;
        RECT 201.855 1712.740 202.875 1712.910 ;
      LAYER li1 ;
        RECT 200.715 1712.570 201.685 1712.610 ;
        RECT 200.715 1712.320 202.485 1712.570 ;
        RECT 200.715 1712.280 201.515 1712.320 ;
        RECT 201.685 1712.240 202.485 1712.320 ;
      LAYER li1 ;
        RECT 200.325 1711.940 201.345 1712.110 ;
        RECT 200.325 1711.270 200.495 1711.940 ;
      LAYER li1 ;
        RECT 201.515 1711.860 201.685 1712.150 ;
      LAYER li1 ;
        RECT 202.705 1712.070 202.875 1712.740 ;
        RECT 201.855 1711.900 202.875 1712.070 ;
      LAYER li1 ;
        RECT 200.715 1711.690 201.515 1711.770 ;
        RECT 201.685 1711.690 202.485 1711.730 ;
        RECT 200.715 1711.440 202.485 1711.690 ;
        RECT 201.515 1711.400 202.485 1711.440 ;
      LAYER li1 ;
        RECT 200.325 1711.100 201.345 1711.270 ;
        RECT 202.705 1711.230 202.875 1711.900 ;
      LAYER li1 ;
        RECT 201.515 1710.940 201.685 1711.230 ;
      LAYER li1 ;
        RECT 201.855 1711.060 202.875 1711.230 ;
      LAYER li1 ;
        RECT 198.795 1710.600 199.445 1710.770 ;
        RECT 199.615 1710.665 200.495 1710.840 ;
        RECT 200.715 1710.770 201.515 1710.850 ;
        RECT 201.685 1710.770 202.485 1710.890 ;
        RECT 200.715 1710.680 202.485 1710.770 ;
        RECT 198.795 1710.480 198.965 1710.600 ;
        RECT 199.615 1710.430 199.785 1710.665 ;
        RECT 200.325 1710.510 200.495 1710.665 ;
        RECT 201.515 1710.560 202.485 1710.680 ;
        RECT 198.795 1710.090 198.965 1710.310 ;
        RECT 199.140 1710.260 199.785 1710.430 ;
        RECT 198.795 1710.020 199.445 1710.090 ;
        RECT 198.965 1709.850 199.445 1710.020 ;
        RECT 198.795 1709.760 199.445 1709.850 ;
        RECT 198.795 1709.560 198.965 1709.760 ;
        RECT 199.615 1709.590 199.785 1710.260 ;
        RECT 199.135 1709.420 199.785 1709.590 ;
        RECT 198.795 1709.160 198.965 1709.390 ;
      LAYER li1 ;
        RECT 199.955 1709.385 200.155 1710.485 ;
      LAYER li1 ;
        RECT 200.325 1710.180 201.345 1710.510 ;
        RECT 201.515 1710.480 201.685 1710.560 ;
      LAYER li1 ;
        RECT 202.705 1710.475 202.875 1711.060 ;
      LAYER li1 ;
        RECT 203.075 1710.720 203.245 1713.170 ;
        RECT 203.755 1713.080 204.235 1713.240 ;
      LAYER li1 ;
        RECT 203.415 1712.740 204.065 1712.910 ;
      LAYER li1 ;
        RECT 204.235 1712.780 204.405 1713.070 ;
      LAYER li1 ;
        RECT 203.415 1712.070 203.585 1712.740 ;
      LAYER li1 ;
        RECT 204.235 1712.570 204.405 1712.610 ;
        RECT 203.755 1712.320 204.405 1712.570 ;
        RECT 203.755 1712.240 204.235 1712.320 ;
      LAYER li1 ;
        RECT 203.415 1711.900 204.065 1712.070 ;
        RECT 203.415 1711.230 203.585 1711.900 ;
      LAYER li1 ;
        RECT 204.235 1711.860 204.405 1712.150 ;
        RECT 203.755 1711.690 204.235 1711.730 ;
        RECT 203.755 1711.400 204.405 1711.690 ;
      LAYER li1 ;
        RECT 203.415 1711.060 204.065 1711.230 ;
        RECT 203.415 1710.475 203.585 1711.060 ;
      LAYER li1 ;
        RECT 204.235 1710.940 204.405 1711.230 ;
        RECT 203.755 1710.770 204.235 1710.890 ;
        RECT 203.755 1710.560 204.405 1710.770 ;
        RECT 204.235 1710.480 204.405 1710.560 ;
      LAYER li1 ;
        RECT 202.705 1710.390 203.585 1710.475 ;
      LAYER li1 ;
        RECT 200.325 1709.670 200.495 1710.180 ;
        RECT 201.515 1710.050 201.685 1710.310 ;
      LAYER li1 ;
        RECT 201.855 1710.220 204.065 1710.390 ;
      LAYER li1 ;
        RECT 204.235 1710.050 204.405 1710.310 ;
        RECT 201.515 1710.020 202.835 1710.050 ;
        RECT 200.715 1709.850 201.515 1710.010 ;
        RECT 201.685 1709.850 202.835 1710.020 ;
        RECT 200.715 1709.840 202.835 1709.850 ;
        RECT 201.515 1709.720 202.835 1709.840 ;
        RECT 203.435 1710.020 204.405 1710.050 ;
        RECT 203.435 1709.850 204.235 1710.020 ;
        RECT 203.435 1709.720 204.405 1709.850 ;
        RECT 200.325 1709.340 201.345 1709.670 ;
        RECT 201.515 1709.560 201.685 1709.720 ;
        RECT 204.235 1709.560 204.405 1709.720 ;
        RECT 201.515 1709.160 201.685 1709.390 ;
        RECT 204.235 1709.160 204.405 1709.390 ;
        RECT 198.795 1709.100 199.690 1709.160 ;
        RECT 198.965 1708.930 199.690 1709.100 ;
        RECT 198.795 1708.870 199.690 1708.930 ;
        RECT 200.350 1709.100 202.850 1709.160 ;
        RECT 200.350 1708.930 201.515 1709.100 ;
        RECT 201.685 1708.930 202.850 1709.100 ;
        RECT 200.350 1708.870 202.850 1708.930 ;
        RECT 198.795 1708.640 198.965 1708.870 ;
        RECT 201.515 1708.640 201.685 1708.870 ;
        RECT 198.795 1708.310 198.965 1708.470 ;
        RECT 201.515 1708.310 201.685 1708.470 ;
        RECT 201.855 1708.360 202.875 1708.690 ;
        RECT 198.795 1708.180 199.765 1708.310 ;
        RECT 198.965 1708.010 199.765 1708.180 ;
        RECT 198.795 1707.980 199.765 1708.010 ;
        RECT 200.365 1708.190 201.685 1708.310 ;
        RECT 200.365 1708.180 202.485 1708.190 ;
        RECT 200.365 1708.010 201.515 1708.180 ;
        RECT 201.685 1708.020 202.485 1708.180 ;
        RECT 200.365 1707.980 201.685 1708.010 ;
        RECT 198.795 1707.720 198.965 1707.980 ;
      LAYER li1 ;
        RECT 199.135 1707.640 201.345 1707.810 ;
      LAYER li1 ;
        RECT 201.515 1707.720 201.685 1707.980 ;
        RECT 202.705 1707.850 202.875 1708.360 ;
      LAYER li1 ;
        RECT 199.615 1707.555 200.495 1707.640 ;
      LAYER li1 ;
        RECT 198.795 1707.470 198.965 1707.550 ;
        RECT 198.795 1707.260 199.445 1707.470 ;
        RECT 198.965 1707.140 199.445 1707.260 ;
        RECT 198.795 1706.800 198.965 1707.090 ;
      LAYER li1 ;
        RECT 199.615 1706.970 199.785 1707.555 ;
        RECT 199.135 1706.800 199.785 1706.970 ;
      LAYER li1 ;
        RECT 198.795 1706.340 199.445 1706.630 ;
        RECT 198.965 1706.300 199.445 1706.340 ;
        RECT 198.795 1705.880 198.965 1706.170 ;
      LAYER li1 ;
        RECT 199.615 1706.130 199.785 1706.800 ;
        RECT 199.135 1705.960 199.785 1706.130 ;
      LAYER li1 ;
        RECT 198.965 1705.710 199.445 1705.790 ;
        RECT 198.795 1705.460 199.445 1705.710 ;
        RECT 198.795 1705.420 198.965 1705.460 ;
      LAYER li1 ;
        RECT 199.615 1705.290 199.785 1705.960 ;
      LAYER li1 ;
        RECT 198.795 1704.960 198.965 1705.250 ;
      LAYER li1 ;
        RECT 199.135 1705.120 199.785 1705.290 ;
      LAYER li1 ;
        RECT 198.965 1704.790 199.445 1704.950 ;
        RECT 199.955 1704.860 200.125 1707.310 ;
      LAYER li1 ;
        RECT 200.325 1706.970 200.495 1707.555 ;
      LAYER li1 ;
        RECT 201.515 1707.470 201.685 1707.550 ;
        RECT 201.855 1707.520 202.875 1707.850 ;
      LAYER li1 ;
        RECT 203.045 1707.545 203.245 1709.135 ;
      LAYER li1 ;
        RECT 203.510 1709.100 204.405 1709.160 ;
        RECT 203.510 1708.930 204.235 1709.100 ;
        RECT 203.510 1708.870 204.405 1708.930 ;
        RECT 204.235 1708.640 204.405 1708.870 ;
        RECT 203.415 1708.440 204.065 1708.610 ;
        RECT 203.415 1707.770 203.585 1708.440 ;
        RECT 204.235 1708.270 204.405 1708.470 ;
        RECT 203.755 1708.180 204.405 1708.270 ;
        RECT 203.755 1708.010 204.235 1708.180 ;
        RECT 203.755 1707.940 204.405 1708.010 ;
        RECT 203.415 1707.600 204.060 1707.770 ;
        RECT 204.235 1707.720 204.405 1707.940 ;
        RECT 200.715 1707.350 201.685 1707.470 ;
        RECT 202.705 1707.365 202.875 1707.520 ;
        RECT 203.415 1707.365 203.585 1707.600 ;
        RECT 204.235 1707.430 204.405 1707.550 ;
        RECT 200.715 1707.260 202.485 1707.350 ;
        RECT 200.715 1707.140 201.515 1707.260 ;
        RECT 201.685 1707.180 202.485 1707.260 ;
        RECT 202.705 1707.190 203.585 1707.365 ;
        RECT 203.755 1707.260 204.405 1707.430 ;
      LAYER li1 ;
        RECT 200.325 1706.800 201.345 1706.970 ;
      LAYER li1 ;
        RECT 201.515 1706.800 201.685 1707.090 ;
      LAYER li1 ;
        RECT 200.325 1706.130 200.495 1706.800 ;
        RECT 201.855 1706.760 202.875 1706.930 ;
      LAYER li1 ;
        RECT 200.715 1706.590 201.685 1706.630 ;
        RECT 200.715 1706.340 202.485 1706.590 ;
        RECT 200.715 1706.300 201.515 1706.340 ;
        RECT 201.685 1706.260 202.485 1706.340 ;
      LAYER li1 ;
        RECT 200.325 1705.960 201.345 1706.130 ;
        RECT 200.325 1705.290 200.495 1705.960 ;
      LAYER li1 ;
        RECT 201.515 1705.880 201.685 1706.170 ;
      LAYER li1 ;
        RECT 202.705 1706.090 202.875 1706.760 ;
        RECT 201.855 1705.920 202.875 1706.090 ;
      LAYER li1 ;
        RECT 200.715 1705.710 201.515 1705.790 ;
        RECT 201.685 1705.710 202.485 1705.750 ;
        RECT 200.715 1705.460 202.485 1705.710 ;
        RECT 201.515 1705.420 202.485 1705.460 ;
      LAYER li1 ;
        RECT 200.325 1705.120 201.345 1705.290 ;
        RECT 202.705 1705.250 202.875 1705.920 ;
      LAYER li1 ;
        RECT 201.515 1704.960 201.685 1705.250 ;
      LAYER li1 ;
        RECT 201.855 1705.080 202.875 1705.250 ;
      LAYER li1 ;
        RECT 198.795 1704.620 199.445 1704.790 ;
        RECT 199.615 1704.685 200.495 1704.860 ;
        RECT 200.715 1704.790 201.515 1704.870 ;
        RECT 201.685 1704.790 202.485 1704.910 ;
        RECT 200.715 1704.700 202.485 1704.790 ;
        RECT 198.795 1704.500 198.965 1704.620 ;
        RECT 199.615 1704.450 199.785 1704.685 ;
        RECT 200.325 1704.530 200.495 1704.685 ;
        RECT 201.515 1704.580 202.485 1704.700 ;
        RECT 198.795 1704.110 198.965 1704.330 ;
        RECT 199.140 1704.280 199.785 1704.450 ;
        RECT 198.795 1704.040 199.445 1704.110 ;
        RECT 198.965 1703.870 199.445 1704.040 ;
        RECT 198.795 1703.780 199.445 1703.870 ;
        RECT 198.795 1703.580 198.965 1703.780 ;
        RECT 199.615 1703.610 199.785 1704.280 ;
        RECT 199.135 1703.440 199.785 1703.610 ;
        RECT 198.795 1703.180 198.965 1703.410 ;
      LAYER li1 ;
        RECT 199.955 1703.405 200.155 1704.505 ;
      LAYER li1 ;
        RECT 200.325 1704.200 201.345 1704.530 ;
        RECT 201.515 1704.500 201.685 1704.580 ;
      LAYER li1 ;
        RECT 202.705 1704.495 202.875 1705.080 ;
      LAYER li1 ;
        RECT 203.075 1704.740 203.245 1707.190 ;
        RECT 203.755 1707.100 204.235 1707.260 ;
      LAYER li1 ;
        RECT 203.415 1706.760 204.065 1706.930 ;
      LAYER li1 ;
        RECT 204.235 1706.800 204.405 1707.090 ;
      LAYER li1 ;
        RECT 203.415 1706.090 203.585 1706.760 ;
      LAYER li1 ;
        RECT 204.235 1706.590 204.405 1706.630 ;
        RECT 203.755 1706.340 204.405 1706.590 ;
        RECT 203.755 1706.260 204.235 1706.340 ;
      LAYER li1 ;
        RECT 203.415 1705.920 204.065 1706.090 ;
        RECT 203.415 1705.250 203.585 1705.920 ;
      LAYER li1 ;
        RECT 204.235 1705.880 204.405 1706.170 ;
        RECT 203.755 1705.710 204.235 1705.750 ;
        RECT 203.755 1705.420 204.405 1705.710 ;
      LAYER li1 ;
        RECT 203.415 1705.080 204.065 1705.250 ;
        RECT 203.415 1704.495 203.585 1705.080 ;
      LAYER li1 ;
        RECT 204.235 1704.960 204.405 1705.250 ;
        RECT 203.755 1704.790 204.235 1704.910 ;
        RECT 203.755 1704.580 204.405 1704.790 ;
        RECT 204.235 1704.500 204.405 1704.580 ;
      LAYER li1 ;
        RECT 202.705 1704.410 203.585 1704.495 ;
      LAYER li1 ;
        RECT 200.325 1703.690 200.495 1704.200 ;
        RECT 201.515 1704.070 201.685 1704.330 ;
      LAYER li1 ;
        RECT 201.855 1704.240 204.065 1704.410 ;
      LAYER li1 ;
        RECT 204.235 1704.070 204.405 1704.330 ;
        RECT 201.515 1704.040 202.835 1704.070 ;
        RECT 200.715 1703.870 201.515 1704.030 ;
        RECT 201.685 1703.870 202.835 1704.040 ;
        RECT 200.715 1703.860 202.835 1703.870 ;
        RECT 201.515 1703.740 202.835 1703.860 ;
        RECT 203.435 1704.040 204.405 1704.070 ;
        RECT 203.435 1703.870 204.235 1704.040 ;
        RECT 203.435 1703.740 204.405 1703.870 ;
        RECT 200.325 1703.360 201.345 1703.690 ;
        RECT 201.515 1703.580 201.685 1703.740 ;
        RECT 204.235 1703.580 204.405 1703.740 ;
        RECT 201.515 1703.180 201.685 1703.410 ;
        RECT 204.235 1703.180 204.405 1703.410 ;
        RECT 198.795 1703.120 199.690 1703.180 ;
        RECT 198.965 1702.950 199.690 1703.120 ;
        RECT 198.795 1702.890 199.690 1702.950 ;
        RECT 200.350 1703.120 202.850 1703.180 ;
        RECT 200.350 1702.950 201.515 1703.120 ;
        RECT 201.685 1702.950 202.850 1703.120 ;
        RECT 200.350 1702.890 202.850 1702.950 ;
        RECT 198.795 1702.660 198.965 1702.890 ;
        RECT 201.515 1702.660 201.685 1702.890 ;
        RECT 198.795 1702.330 198.965 1702.490 ;
        RECT 201.515 1702.330 201.685 1702.490 ;
        RECT 201.855 1702.380 202.875 1702.710 ;
        RECT 198.795 1702.200 199.765 1702.330 ;
        RECT 198.965 1702.030 199.765 1702.200 ;
        RECT 198.795 1702.000 199.765 1702.030 ;
        RECT 200.365 1702.210 201.685 1702.330 ;
        RECT 200.365 1702.200 202.485 1702.210 ;
        RECT 200.365 1702.030 201.515 1702.200 ;
        RECT 201.685 1702.040 202.485 1702.200 ;
        RECT 200.365 1702.000 201.685 1702.030 ;
        RECT 198.795 1701.740 198.965 1702.000 ;
      LAYER li1 ;
        RECT 199.135 1701.660 201.345 1701.830 ;
      LAYER li1 ;
        RECT 201.515 1701.740 201.685 1702.000 ;
        RECT 202.705 1701.870 202.875 1702.380 ;
      LAYER li1 ;
        RECT 199.615 1701.575 200.495 1701.660 ;
      LAYER li1 ;
        RECT 198.795 1701.490 198.965 1701.570 ;
        RECT 198.795 1701.280 199.445 1701.490 ;
        RECT 198.965 1701.160 199.445 1701.280 ;
        RECT 198.795 1700.820 198.965 1701.110 ;
      LAYER li1 ;
        RECT 199.615 1700.990 199.785 1701.575 ;
        RECT 199.135 1700.820 199.785 1700.990 ;
      LAYER li1 ;
        RECT 198.795 1700.360 199.445 1700.650 ;
        RECT 198.965 1700.320 199.445 1700.360 ;
        RECT 198.795 1699.900 198.965 1700.190 ;
      LAYER li1 ;
        RECT 199.615 1700.150 199.785 1700.820 ;
        RECT 199.135 1699.980 199.785 1700.150 ;
      LAYER li1 ;
        RECT 198.965 1699.730 199.445 1699.810 ;
        RECT 198.795 1699.480 199.445 1699.730 ;
        RECT 198.795 1699.440 198.965 1699.480 ;
      LAYER li1 ;
        RECT 199.615 1699.310 199.785 1699.980 ;
      LAYER li1 ;
        RECT 198.795 1698.980 198.965 1699.270 ;
      LAYER li1 ;
        RECT 199.135 1699.140 199.785 1699.310 ;
      LAYER li1 ;
        RECT 198.965 1698.810 199.445 1698.970 ;
        RECT 199.955 1698.880 200.125 1701.330 ;
      LAYER li1 ;
        RECT 200.325 1700.990 200.495 1701.575 ;
      LAYER li1 ;
        RECT 201.515 1701.490 201.685 1701.570 ;
        RECT 201.855 1701.540 202.875 1701.870 ;
      LAYER li1 ;
        RECT 203.045 1701.565 203.245 1703.155 ;
      LAYER li1 ;
        RECT 203.510 1703.120 204.405 1703.180 ;
        RECT 203.510 1702.950 204.235 1703.120 ;
        RECT 203.510 1702.890 204.405 1702.950 ;
        RECT 204.235 1702.660 204.405 1702.890 ;
        RECT 203.415 1702.460 204.065 1702.630 ;
        RECT 203.415 1701.790 203.585 1702.460 ;
        RECT 204.235 1702.290 204.405 1702.490 ;
        RECT 203.755 1702.200 204.405 1702.290 ;
        RECT 203.755 1702.030 204.235 1702.200 ;
        RECT 203.755 1701.960 204.405 1702.030 ;
        RECT 203.415 1701.620 204.060 1701.790 ;
        RECT 204.235 1701.740 204.405 1701.960 ;
        RECT 200.715 1701.370 201.685 1701.490 ;
        RECT 202.705 1701.385 202.875 1701.540 ;
        RECT 203.415 1701.385 203.585 1701.620 ;
        RECT 204.235 1701.450 204.405 1701.570 ;
        RECT 200.715 1701.280 202.485 1701.370 ;
        RECT 200.715 1701.160 201.515 1701.280 ;
        RECT 201.685 1701.200 202.485 1701.280 ;
        RECT 202.705 1701.210 203.585 1701.385 ;
        RECT 203.755 1701.280 204.405 1701.450 ;
      LAYER li1 ;
        RECT 200.325 1700.820 201.345 1700.990 ;
      LAYER li1 ;
        RECT 201.515 1700.820 201.685 1701.110 ;
      LAYER li1 ;
        RECT 200.325 1700.150 200.495 1700.820 ;
        RECT 201.855 1700.780 202.875 1700.950 ;
      LAYER li1 ;
        RECT 200.715 1700.610 201.685 1700.650 ;
        RECT 200.715 1700.360 202.485 1700.610 ;
        RECT 200.715 1700.320 201.515 1700.360 ;
        RECT 201.685 1700.280 202.485 1700.360 ;
      LAYER li1 ;
        RECT 200.325 1699.980 201.345 1700.150 ;
        RECT 200.325 1699.310 200.495 1699.980 ;
      LAYER li1 ;
        RECT 201.515 1699.900 201.685 1700.190 ;
      LAYER li1 ;
        RECT 202.705 1700.110 202.875 1700.780 ;
        RECT 201.855 1699.940 202.875 1700.110 ;
      LAYER li1 ;
        RECT 200.715 1699.730 201.515 1699.810 ;
        RECT 201.685 1699.730 202.485 1699.770 ;
        RECT 200.715 1699.480 202.485 1699.730 ;
        RECT 201.515 1699.440 202.485 1699.480 ;
      LAYER li1 ;
        RECT 200.325 1699.140 201.345 1699.310 ;
        RECT 202.705 1699.270 202.875 1699.940 ;
      LAYER li1 ;
        RECT 201.515 1698.980 201.685 1699.270 ;
      LAYER li1 ;
        RECT 201.855 1699.100 202.875 1699.270 ;
      LAYER li1 ;
        RECT 198.795 1698.640 199.445 1698.810 ;
        RECT 199.615 1698.705 200.495 1698.880 ;
        RECT 200.715 1698.810 201.515 1698.890 ;
        RECT 201.685 1698.810 202.485 1698.930 ;
        RECT 200.715 1698.720 202.485 1698.810 ;
        RECT 198.795 1698.520 198.965 1698.640 ;
        RECT 199.615 1698.470 199.785 1698.705 ;
        RECT 200.325 1698.550 200.495 1698.705 ;
        RECT 201.515 1698.600 202.485 1698.720 ;
        RECT 198.795 1698.130 198.965 1698.350 ;
        RECT 199.140 1698.300 199.785 1698.470 ;
        RECT 198.795 1698.060 199.445 1698.130 ;
        RECT 198.965 1697.890 199.445 1698.060 ;
        RECT 198.795 1697.800 199.445 1697.890 ;
        RECT 198.795 1697.600 198.965 1697.800 ;
        RECT 199.615 1697.630 199.785 1698.300 ;
        RECT 199.135 1697.460 199.785 1697.630 ;
        RECT 198.795 1697.200 198.965 1697.430 ;
      LAYER li1 ;
        RECT 199.955 1697.425 200.155 1698.525 ;
      LAYER li1 ;
        RECT 200.325 1698.220 201.345 1698.550 ;
        RECT 201.515 1698.520 201.685 1698.600 ;
      LAYER li1 ;
        RECT 202.705 1698.515 202.875 1699.100 ;
      LAYER li1 ;
        RECT 203.075 1698.760 203.245 1701.210 ;
        RECT 203.755 1701.120 204.235 1701.280 ;
      LAYER li1 ;
        RECT 203.415 1700.780 204.065 1700.950 ;
      LAYER li1 ;
        RECT 204.235 1700.820 204.405 1701.110 ;
      LAYER li1 ;
        RECT 203.415 1700.110 203.585 1700.780 ;
      LAYER li1 ;
        RECT 204.235 1700.610 204.405 1700.650 ;
        RECT 203.755 1700.360 204.405 1700.610 ;
        RECT 203.755 1700.280 204.235 1700.360 ;
      LAYER li1 ;
        RECT 203.415 1699.940 204.065 1700.110 ;
        RECT 203.415 1699.270 203.585 1699.940 ;
      LAYER li1 ;
        RECT 204.235 1699.900 204.405 1700.190 ;
        RECT 203.755 1699.730 204.235 1699.770 ;
        RECT 203.755 1699.440 204.405 1699.730 ;
      LAYER li1 ;
        RECT 203.415 1699.100 204.065 1699.270 ;
        RECT 203.415 1698.515 203.585 1699.100 ;
      LAYER li1 ;
        RECT 204.235 1698.980 204.405 1699.270 ;
        RECT 203.755 1698.810 204.235 1698.930 ;
        RECT 203.755 1698.600 204.405 1698.810 ;
        RECT 204.235 1698.520 204.405 1698.600 ;
      LAYER li1 ;
        RECT 202.705 1698.430 203.585 1698.515 ;
      LAYER li1 ;
        RECT 200.325 1697.710 200.495 1698.220 ;
        RECT 201.515 1698.090 201.685 1698.350 ;
      LAYER li1 ;
        RECT 201.855 1698.260 204.065 1698.430 ;
      LAYER li1 ;
        RECT 204.235 1698.090 204.405 1698.350 ;
        RECT 201.515 1698.060 202.835 1698.090 ;
        RECT 200.715 1697.890 201.515 1698.050 ;
        RECT 201.685 1697.890 202.835 1698.060 ;
        RECT 200.715 1697.880 202.835 1697.890 ;
        RECT 201.515 1697.760 202.835 1697.880 ;
        RECT 203.435 1698.060 204.405 1698.090 ;
        RECT 203.435 1697.890 204.235 1698.060 ;
        RECT 203.435 1697.760 204.405 1697.890 ;
        RECT 200.325 1697.380 201.345 1697.710 ;
        RECT 201.515 1697.600 201.685 1697.760 ;
        RECT 204.235 1697.600 204.405 1697.760 ;
        RECT 201.515 1697.200 201.685 1697.430 ;
        RECT 204.235 1697.200 204.405 1697.430 ;
        RECT 198.795 1697.140 199.690 1697.200 ;
        RECT 198.965 1696.970 199.690 1697.140 ;
        RECT 198.795 1696.910 199.690 1696.970 ;
        RECT 200.350 1697.140 202.850 1697.200 ;
        RECT 200.350 1696.970 201.515 1697.140 ;
        RECT 201.685 1696.970 202.850 1697.140 ;
        RECT 200.350 1696.910 202.850 1696.970 ;
        RECT 203.510 1697.140 204.405 1697.200 ;
        RECT 203.510 1696.970 204.235 1697.140 ;
        RECT 203.510 1696.910 204.405 1696.970 ;
        RECT 198.795 1696.680 198.965 1696.910 ;
        RECT 201.515 1696.680 201.685 1696.910 ;
        RECT 198.795 1696.350 198.965 1696.510 ;
        RECT 201.515 1696.350 201.685 1696.510 ;
        RECT 201.855 1696.400 202.875 1696.730 ;
        RECT 204.235 1696.680 204.405 1696.910 ;
        RECT 198.795 1696.220 199.765 1696.350 ;
        RECT 198.965 1696.050 199.765 1696.220 ;
        RECT 198.795 1696.020 199.765 1696.050 ;
        RECT 200.365 1696.230 201.685 1696.350 ;
        RECT 200.365 1696.220 202.485 1696.230 ;
        RECT 200.365 1696.050 201.515 1696.220 ;
        RECT 201.685 1696.060 202.485 1696.220 ;
        RECT 200.365 1696.020 201.685 1696.050 ;
        RECT 198.795 1695.760 198.965 1696.020 ;
        RECT 201.515 1695.760 201.685 1696.020 ;
        RECT 202.705 1695.890 202.875 1696.400 ;
        RECT 198.795 1695.510 198.965 1695.590 ;
        RECT 201.515 1695.510 201.685 1695.590 ;
        RECT 201.855 1695.560 202.875 1695.890 ;
        RECT 198.795 1695.300 199.445 1695.510 ;
        RECT 200.715 1695.390 201.685 1695.510 ;
        RECT 202.705 1695.405 202.875 1695.560 ;
        RECT 203.415 1696.480 204.065 1696.650 ;
        RECT 203.415 1695.810 203.585 1696.480 ;
        RECT 204.235 1696.310 204.405 1696.510 ;
        RECT 203.755 1696.220 204.405 1696.310 ;
        RECT 203.755 1696.050 204.235 1696.220 ;
        RECT 203.755 1695.980 204.405 1696.050 ;
        RECT 203.415 1695.640 204.060 1695.810 ;
        RECT 204.235 1695.760 204.405 1695.980 ;
        RECT 203.415 1695.405 203.585 1695.640 ;
        RECT 204.235 1695.470 204.405 1695.590 ;
        RECT 198.965 1695.180 199.445 1695.300 ;
        RECT 198.795 1694.840 198.965 1695.130 ;
        RECT 198.795 1694.380 199.445 1694.670 ;
        RECT 198.965 1694.340 199.445 1694.380 ;
        RECT 198.795 1693.920 198.965 1694.210 ;
        RECT 198.965 1693.750 199.445 1693.830 ;
        RECT 198.795 1693.500 199.445 1693.750 ;
        RECT 198.795 1693.460 198.965 1693.500 ;
        RECT 198.795 1693.000 198.965 1693.290 ;
        RECT 198.965 1692.830 199.445 1692.990 ;
        RECT 199.955 1692.900 200.125 1695.350 ;
        RECT 200.715 1695.300 202.485 1695.390 ;
        RECT 200.715 1695.180 201.515 1695.300 ;
        RECT 201.685 1695.220 202.485 1695.300 ;
        RECT 202.705 1695.230 203.585 1695.405 ;
        RECT 203.755 1695.300 204.405 1695.470 ;
        RECT 201.515 1694.840 201.685 1695.130 ;
      LAYER li1 ;
        RECT 201.855 1694.800 202.875 1694.970 ;
      LAYER li1 ;
        RECT 200.715 1694.630 201.685 1694.670 ;
        RECT 200.715 1694.380 202.485 1694.630 ;
        RECT 200.715 1694.340 201.515 1694.380 ;
        RECT 201.685 1694.300 202.485 1694.380 ;
        RECT 201.515 1693.920 201.685 1694.210 ;
      LAYER li1 ;
        RECT 202.705 1694.130 202.875 1694.800 ;
        RECT 201.855 1693.960 202.875 1694.130 ;
      LAYER li1 ;
        RECT 200.715 1693.750 201.515 1693.830 ;
        RECT 201.685 1693.750 202.485 1693.790 ;
        RECT 200.715 1693.500 202.485 1693.750 ;
        RECT 201.515 1693.460 202.485 1693.500 ;
      LAYER li1 ;
        RECT 202.705 1693.290 202.875 1693.960 ;
      LAYER li1 ;
        RECT 201.515 1693.000 201.685 1693.290 ;
      LAYER li1 ;
        RECT 201.855 1693.120 202.875 1693.290 ;
      LAYER li1 ;
        RECT 198.795 1692.660 199.445 1692.830 ;
        RECT 199.615 1692.725 200.495 1692.900 ;
        RECT 200.715 1692.830 201.515 1692.910 ;
        RECT 201.685 1692.830 202.485 1692.950 ;
        RECT 200.715 1692.740 202.485 1692.830 ;
        RECT 198.795 1692.540 198.965 1692.660 ;
        RECT 199.615 1692.490 199.785 1692.725 ;
        RECT 200.325 1692.570 200.495 1692.725 ;
        RECT 201.515 1692.620 202.485 1692.740 ;
        RECT 198.795 1692.150 198.965 1692.370 ;
        RECT 199.140 1692.320 199.785 1692.490 ;
        RECT 198.795 1692.080 199.445 1692.150 ;
        RECT 198.965 1691.910 199.445 1692.080 ;
        RECT 198.795 1691.820 199.445 1691.910 ;
        RECT 198.795 1691.620 198.965 1691.820 ;
        RECT 199.615 1691.650 199.785 1692.320 ;
        RECT 199.135 1691.480 199.785 1691.650 ;
        RECT 198.795 1691.220 198.965 1691.450 ;
      LAYER li1 ;
        RECT 199.955 1691.445 200.155 1692.545 ;
      LAYER li1 ;
        RECT 200.325 1692.240 201.345 1692.570 ;
        RECT 201.515 1692.540 201.685 1692.620 ;
      LAYER li1 ;
        RECT 202.705 1692.535 202.875 1693.120 ;
      LAYER li1 ;
        RECT 203.075 1692.780 203.245 1695.230 ;
        RECT 203.755 1695.140 204.235 1695.300 ;
      LAYER li1 ;
        RECT 203.415 1694.800 204.065 1694.970 ;
      LAYER li1 ;
        RECT 204.235 1694.840 204.405 1695.130 ;
      LAYER li1 ;
        RECT 203.415 1694.130 203.585 1694.800 ;
      LAYER li1 ;
        RECT 204.235 1694.630 204.405 1694.670 ;
        RECT 203.755 1694.380 204.405 1694.630 ;
        RECT 203.755 1694.300 204.235 1694.380 ;
      LAYER li1 ;
        RECT 203.415 1693.960 204.065 1694.130 ;
        RECT 203.415 1693.290 203.585 1693.960 ;
      LAYER li1 ;
        RECT 204.235 1693.920 204.405 1694.210 ;
        RECT 203.755 1693.750 204.235 1693.790 ;
        RECT 203.755 1693.460 204.405 1693.750 ;
      LAYER li1 ;
        RECT 203.415 1693.120 204.065 1693.290 ;
        RECT 203.415 1692.535 203.585 1693.120 ;
      LAYER li1 ;
        RECT 204.235 1693.000 204.405 1693.290 ;
        RECT 203.755 1692.830 204.235 1692.950 ;
        RECT 203.755 1692.620 204.405 1692.830 ;
        RECT 204.235 1692.540 204.405 1692.620 ;
      LAYER li1 ;
        RECT 202.705 1692.450 203.585 1692.535 ;
      LAYER li1 ;
        RECT 200.325 1691.730 200.495 1692.240 ;
        RECT 201.515 1692.110 201.685 1692.370 ;
      LAYER li1 ;
        RECT 201.855 1692.280 204.065 1692.450 ;
      LAYER li1 ;
        RECT 204.235 1692.110 204.405 1692.370 ;
        RECT 201.515 1692.080 202.835 1692.110 ;
        RECT 200.715 1691.910 201.515 1692.070 ;
        RECT 201.685 1691.910 202.835 1692.080 ;
        RECT 200.715 1691.900 202.835 1691.910 ;
        RECT 201.515 1691.780 202.835 1691.900 ;
        RECT 203.435 1692.080 204.405 1692.110 ;
        RECT 203.435 1691.910 204.235 1692.080 ;
        RECT 203.435 1691.780 204.405 1691.910 ;
        RECT 200.325 1691.400 201.345 1691.730 ;
        RECT 201.515 1691.620 201.685 1691.780 ;
        RECT 204.235 1691.620 204.405 1691.780 ;
        RECT 201.515 1691.220 201.685 1691.450 ;
        RECT 204.235 1691.220 204.405 1691.450 ;
        RECT 198.795 1691.160 199.690 1691.220 ;
        RECT 198.965 1690.990 199.690 1691.160 ;
        RECT 198.795 1690.930 199.690 1690.990 ;
        RECT 200.350 1691.160 202.850 1691.220 ;
        RECT 200.350 1690.990 201.515 1691.160 ;
        RECT 201.685 1690.990 202.850 1691.160 ;
        RECT 200.350 1690.930 202.850 1690.990 ;
        RECT 203.510 1691.160 204.405 1691.220 ;
        RECT 203.510 1690.990 204.235 1691.160 ;
        RECT 203.510 1690.930 204.405 1690.990 ;
        RECT 198.795 1690.700 198.965 1690.930 ;
        RECT 201.515 1690.700 201.685 1690.930 ;
        RECT 198.795 1690.370 198.965 1690.530 ;
        RECT 201.515 1690.370 201.685 1690.530 ;
        RECT 201.855 1690.420 202.875 1690.750 ;
        RECT 204.235 1690.700 204.405 1690.930 ;
        RECT 198.795 1690.240 199.765 1690.370 ;
        RECT 198.965 1690.070 199.765 1690.240 ;
        RECT 198.795 1690.040 199.765 1690.070 ;
        RECT 200.365 1690.250 201.685 1690.370 ;
        RECT 200.365 1690.240 202.485 1690.250 ;
        RECT 200.365 1690.070 201.515 1690.240 ;
        RECT 201.685 1690.080 202.485 1690.240 ;
        RECT 200.365 1690.040 201.685 1690.070 ;
        RECT 198.795 1689.780 198.965 1690.040 ;
        RECT 201.515 1689.780 201.685 1690.040 ;
        RECT 202.705 1689.910 202.875 1690.420 ;
        RECT 198.795 1689.530 198.965 1689.610 ;
        RECT 201.515 1689.530 201.685 1689.610 ;
        RECT 201.855 1689.580 202.875 1689.910 ;
        RECT 198.795 1689.320 199.445 1689.530 ;
        RECT 200.715 1689.410 201.685 1689.530 ;
        RECT 202.705 1689.425 202.875 1689.580 ;
        RECT 203.415 1690.500 204.065 1690.670 ;
        RECT 203.415 1689.830 203.585 1690.500 ;
        RECT 204.235 1690.330 204.405 1690.530 ;
        RECT 203.755 1690.240 204.405 1690.330 ;
        RECT 203.755 1690.070 204.235 1690.240 ;
        RECT 203.755 1690.000 204.405 1690.070 ;
        RECT 203.415 1689.660 204.060 1689.830 ;
        RECT 204.235 1689.780 204.405 1690.000 ;
        RECT 203.415 1689.425 203.585 1689.660 ;
        RECT 204.235 1689.490 204.405 1689.610 ;
        RECT 198.965 1689.200 199.445 1689.320 ;
        RECT 198.795 1688.860 198.965 1689.150 ;
        RECT 198.795 1688.400 199.445 1688.690 ;
        RECT 198.965 1688.360 199.445 1688.400 ;
        RECT 198.795 1687.940 198.965 1688.230 ;
        RECT 198.965 1687.770 199.445 1687.850 ;
        RECT 198.795 1687.520 199.445 1687.770 ;
        RECT 198.795 1687.480 198.965 1687.520 ;
        RECT 198.795 1687.020 198.965 1687.310 ;
        RECT 198.965 1686.850 199.445 1687.010 ;
        RECT 199.955 1686.920 200.125 1689.370 ;
        RECT 200.715 1689.320 202.485 1689.410 ;
        RECT 200.715 1689.200 201.515 1689.320 ;
        RECT 201.685 1689.240 202.485 1689.320 ;
        RECT 202.705 1689.250 203.585 1689.425 ;
        RECT 203.755 1689.320 204.405 1689.490 ;
        RECT 201.515 1688.860 201.685 1689.150 ;
      LAYER li1 ;
        RECT 201.855 1688.820 202.875 1688.990 ;
      LAYER li1 ;
        RECT 200.715 1688.650 201.685 1688.690 ;
        RECT 200.715 1688.400 202.485 1688.650 ;
        RECT 200.715 1688.360 201.515 1688.400 ;
        RECT 201.685 1688.320 202.485 1688.400 ;
        RECT 201.515 1687.940 201.685 1688.230 ;
      LAYER li1 ;
        RECT 202.705 1688.150 202.875 1688.820 ;
        RECT 201.855 1687.980 202.875 1688.150 ;
      LAYER li1 ;
        RECT 200.715 1687.770 201.515 1687.850 ;
        RECT 201.685 1687.770 202.485 1687.810 ;
        RECT 200.715 1687.520 202.485 1687.770 ;
        RECT 201.515 1687.480 202.485 1687.520 ;
      LAYER li1 ;
        RECT 202.705 1687.310 202.875 1687.980 ;
      LAYER li1 ;
        RECT 201.515 1687.020 201.685 1687.310 ;
      LAYER li1 ;
        RECT 201.855 1687.140 202.875 1687.310 ;
      LAYER li1 ;
        RECT 198.795 1686.680 199.445 1686.850 ;
        RECT 199.615 1686.745 200.495 1686.920 ;
        RECT 200.715 1686.850 201.515 1686.930 ;
        RECT 201.685 1686.850 202.485 1686.970 ;
        RECT 200.715 1686.760 202.485 1686.850 ;
        RECT 198.795 1686.560 198.965 1686.680 ;
        RECT 199.615 1686.510 199.785 1686.745 ;
        RECT 200.325 1686.590 200.495 1686.745 ;
        RECT 201.515 1686.640 202.485 1686.760 ;
        RECT 198.795 1686.170 198.965 1686.390 ;
        RECT 199.140 1686.340 199.785 1686.510 ;
        RECT 198.795 1686.100 199.445 1686.170 ;
        RECT 198.965 1685.930 199.445 1686.100 ;
        RECT 198.795 1685.840 199.445 1685.930 ;
        RECT 198.795 1685.640 198.965 1685.840 ;
        RECT 199.615 1685.670 199.785 1686.340 ;
        RECT 199.135 1685.500 199.785 1685.670 ;
        RECT 198.795 1685.240 198.965 1685.470 ;
      LAYER li1 ;
        RECT 199.955 1685.465 200.155 1686.565 ;
      LAYER li1 ;
        RECT 200.325 1686.260 201.345 1686.590 ;
        RECT 201.515 1686.560 201.685 1686.640 ;
      LAYER li1 ;
        RECT 202.705 1686.555 202.875 1687.140 ;
      LAYER li1 ;
        RECT 203.075 1686.800 203.245 1689.250 ;
        RECT 203.755 1689.160 204.235 1689.320 ;
      LAYER li1 ;
        RECT 203.415 1688.820 204.065 1688.990 ;
      LAYER li1 ;
        RECT 204.235 1688.860 204.405 1689.150 ;
      LAYER li1 ;
        RECT 203.415 1688.150 203.585 1688.820 ;
      LAYER li1 ;
        RECT 204.235 1688.650 204.405 1688.690 ;
        RECT 203.755 1688.400 204.405 1688.650 ;
        RECT 203.755 1688.320 204.235 1688.400 ;
      LAYER li1 ;
        RECT 203.415 1687.980 204.065 1688.150 ;
        RECT 203.415 1687.310 203.585 1687.980 ;
      LAYER li1 ;
        RECT 204.235 1687.940 204.405 1688.230 ;
        RECT 203.755 1687.770 204.235 1687.810 ;
        RECT 203.755 1687.480 204.405 1687.770 ;
      LAYER li1 ;
        RECT 203.415 1687.140 204.065 1687.310 ;
        RECT 203.415 1686.555 203.585 1687.140 ;
      LAYER li1 ;
        RECT 204.235 1687.020 204.405 1687.310 ;
        RECT 203.755 1686.850 204.235 1686.970 ;
        RECT 203.755 1686.640 204.405 1686.850 ;
        RECT 204.235 1686.560 204.405 1686.640 ;
      LAYER li1 ;
        RECT 202.705 1686.470 203.585 1686.555 ;
      LAYER li1 ;
        RECT 200.325 1685.750 200.495 1686.260 ;
        RECT 201.515 1686.130 201.685 1686.390 ;
      LAYER li1 ;
        RECT 201.855 1686.300 204.065 1686.470 ;
      LAYER li1 ;
        RECT 204.235 1686.130 204.405 1686.390 ;
        RECT 201.515 1686.100 202.835 1686.130 ;
        RECT 200.715 1685.930 201.515 1686.090 ;
        RECT 201.685 1685.930 202.835 1686.100 ;
        RECT 200.715 1685.920 202.835 1685.930 ;
        RECT 201.515 1685.800 202.835 1685.920 ;
        RECT 203.435 1686.100 204.405 1686.130 ;
        RECT 203.435 1685.930 204.235 1686.100 ;
        RECT 203.435 1685.800 204.405 1685.930 ;
        RECT 200.325 1685.420 201.345 1685.750 ;
        RECT 201.515 1685.640 201.685 1685.800 ;
        RECT 204.235 1685.640 204.405 1685.800 ;
        RECT 201.515 1685.240 201.685 1685.470 ;
        RECT 204.235 1685.240 204.405 1685.470 ;
        RECT 198.795 1685.180 199.690 1685.240 ;
        RECT 198.965 1685.010 199.690 1685.180 ;
        RECT 198.795 1684.950 199.690 1685.010 ;
        RECT 200.350 1685.180 202.850 1685.240 ;
        RECT 200.350 1685.010 201.515 1685.180 ;
        RECT 201.685 1685.010 202.850 1685.180 ;
        RECT 200.350 1684.950 202.850 1685.010 ;
        RECT 203.510 1685.180 204.405 1685.240 ;
        RECT 203.510 1685.010 204.235 1685.180 ;
        RECT 203.510 1684.950 204.405 1685.010 ;
        RECT 198.795 1684.720 198.965 1684.950 ;
        RECT 201.515 1684.720 201.685 1684.950 ;
        RECT 198.795 1684.390 198.965 1684.550 ;
        RECT 201.515 1684.390 201.685 1684.550 ;
        RECT 201.855 1684.440 202.875 1684.770 ;
        RECT 204.235 1684.720 204.405 1684.950 ;
        RECT 198.795 1684.260 199.765 1684.390 ;
        RECT 198.965 1684.090 199.765 1684.260 ;
        RECT 198.795 1684.060 199.765 1684.090 ;
        RECT 200.365 1684.270 201.685 1684.390 ;
        RECT 200.365 1684.260 202.485 1684.270 ;
        RECT 200.365 1684.090 201.515 1684.260 ;
        RECT 201.685 1684.100 202.485 1684.260 ;
        RECT 200.365 1684.060 201.685 1684.090 ;
        RECT 198.795 1683.800 198.965 1684.060 ;
        RECT 201.515 1683.800 201.685 1684.060 ;
        RECT 202.705 1683.930 202.875 1684.440 ;
        RECT 198.795 1683.550 198.965 1683.630 ;
        RECT 201.515 1683.550 201.685 1683.630 ;
        RECT 201.855 1683.600 202.875 1683.930 ;
        RECT 198.795 1683.340 199.445 1683.550 ;
        RECT 200.715 1683.430 201.685 1683.550 ;
        RECT 202.705 1683.445 202.875 1683.600 ;
        RECT 203.415 1684.520 204.065 1684.690 ;
        RECT 203.415 1683.850 203.585 1684.520 ;
        RECT 204.235 1684.350 204.405 1684.550 ;
        RECT 203.755 1684.260 204.405 1684.350 ;
        RECT 203.755 1684.090 204.235 1684.260 ;
        RECT 203.755 1684.020 204.405 1684.090 ;
        RECT 203.415 1683.680 204.060 1683.850 ;
        RECT 204.235 1683.800 204.405 1684.020 ;
        RECT 203.415 1683.445 203.585 1683.680 ;
        RECT 204.235 1683.510 204.405 1683.630 ;
        RECT 198.965 1683.220 199.445 1683.340 ;
        RECT 198.795 1682.880 198.965 1683.170 ;
        RECT 198.795 1682.420 199.445 1682.710 ;
        RECT 198.965 1682.380 199.445 1682.420 ;
        RECT 198.795 1681.960 198.965 1682.250 ;
        RECT 198.965 1681.790 199.445 1681.870 ;
        RECT 198.795 1681.540 199.445 1681.790 ;
        RECT 198.795 1681.500 198.965 1681.540 ;
        RECT 198.795 1681.040 198.965 1681.330 ;
        RECT 198.965 1680.870 199.445 1681.030 ;
        RECT 199.955 1680.940 200.125 1683.390 ;
        RECT 200.715 1683.340 202.485 1683.430 ;
        RECT 200.715 1683.220 201.515 1683.340 ;
        RECT 201.685 1683.260 202.485 1683.340 ;
        RECT 202.705 1683.270 203.585 1683.445 ;
        RECT 203.755 1683.340 204.405 1683.510 ;
        RECT 201.515 1682.880 201.685 1683.170 ;
      LAYER li1 ;
        RECT 201.855 1682.840 202.875 1683.010 ;
      LAYER li1 ;
        RECT 200.715 1682.670 201.685 1682.710 ;
        RECT 200.715 1682.420 202.485 1682.670 ;
        RECT 200.715 1682.380 201.515 1682.420 ;
        RECT 201.685 1682.340 202.485 1682.420 ;
        RECT 201.515 1681.960 201.685 1682.250 ;
      LAYER li1 ;
        RECT 202.705 1682.170 202.875 1682.840 ;
        RECT 201.855 1682.000 202.875 1682.170 ;
      LAYER li1 ;
        RECT 200.715 1681.790 201.515 1681.870 ;
        RECT 201.685 1681.790 202.485 1681.830 ;
        RECT 200.715 1681.540 202.485 1681.790 ;
        RECT 201.515 1681.500 202.485 1681.540 ;
      LAYER li1 ;
        RECT 202.705 1681.330 202.875 1682.000 ;
      LAYER li1 ;
        RECT 201.515 1681.040 201.685 1681.330 ;
      LAYER li1 ;
        RECT 201.855 1681.160 202.875 1681.330 ;
      LAYER li1 ;
        RECT 198.795 1680.700 199.445 1680.870 ;
        RECT 199.615 1680.765 200.495 1680.940 ;
        RECT 200.715 1680.870 201.515 1680.950 ;
        RECT 201.685 1680.870 202.485 1680.990 ;
        RECT 200.715 1680.780 202.485 1680.870 ;
        RECT 198.795 1680.580 198.965 1680.700 ;
        RECT 199.615 1680.530 199.785 1680.765 ;
        RECT 200.325 1680.610 200.495 1680.765 ;
        RECT 201.515 1680.660 202.485 1680.780 ;
        RECT 198.795 1680.190 198.965 1680.410 ;
        RECT 199.140 1680.360 199.785 1680.530 ;
        RECT 198.795 1680.120 199.445 1680.190 ;
        RECT 198.965 1679.950 199.445 1680.120 ;
        RECT 198.795 1679.860 199.445 1679.950 ;
        RECT 198.795 1679.660 198.965 1679.860 ;
        RECT 199.615 1679.690 199.785 1680.360 ;
        RECT 199.135 1679.520 199.785 1679.690 ;
        RECT 198.795 1679.260 198.965 1679.490 ;
      LAYER li1 ;
        RECT 199.955 1679.485 200.155 1680.585 ;
      LAYER li1 ;
        RECT 200.325 1680.280 201.345 1680.610 ;
        RECT 201.515 1680.580 201.685 1680.660 ;
      LAYER li1 ;
        RECT 202.705 1680.575 202.875 1681.160 ;
      LAYER li1 ;
        RECT 203.075 1680.820 203.245 1683.270 ;
        RECT 203.755 1683.180 204.235 1683.340 ;
      LAYER li1 ;
        RECT 203.415 1682.840 204.065 1683.010 ;
      LAYER li1 ;
        RECT 204.235 1682.880 204.405 1683.170 ;
      LAYER li1 ;
        RECT 203.415 1682.170 203.585 1682.840 ;
      LAYER li1 ;
        RECT 204.235 1682.670 204.405 1682.710 ;
        RECT 203.755 1682.420 204.405 1682.670 ;
        RECT 203.755 1682.340 204.235 1682.420 ;
      LAYER li1 ;
        RECT 203.415 1682.000 204.065 1682.170 ;
        RECT 203.415 1681.330 203.585 1682.000 ;
      LAYER li1 ;
        RECT 204.235 1681.960 204.405 1682.250 ;
        RECT 203.755 1681.790 204.235 1681.830 ;
        RECT 203.755 1681.500 204.405 1681.790 ;
      LAYER li1 ;
        RECT 203.415 1681.160 204.065 1681.330 ;
        RECT 203.415 1680.575 203.585 1681.160 ;
      LAYER li1 ;
        RECT 204.235 1681.040 204.405 1681.330 ;
        RECT 203.755 1680.870 204.235 1680.990 ;
        RECT 203.755 1680.660 204.405 1680.870 ;
        RECT 204.235 1680.580 204.405 1680.660 ;
      LAYER li1 ;
        RECT 202.705 1680.490 203.585 1680.575 ;
      LAYER li1 ;
        RECT 200.325 1679.770 200.495 1680.280 ;
        RECT 201.515 1680.150 201.685 1680.410 ;
      LAYER li1 ;
        RECT 201.855 1680.320 204.065 1680.490 ;
      LAYER li1 ;
        RECT 204.235 1680.150 204.405 1680.410 ;
        RECT 201.515 1680.120 202.835 1680.150 ;
        RECT 200.715 1679.950 201.515 1680.110 ;
        RECT 201.685 1679.950 202.835 1680.120 ;
        RECT 200.715 1679.940 202.835 1679.950 ;
        RECT 201.515 1679.820 202.835 1679.940 ;
        RECT 203.435 1680.120 204.405 1680.150 ;
        RECT 203.435 1679.950 204.235 1680.120 ;
        RECT 203.435 1679.820 204.405 1679.950 ;
        RECT 200.325 1679.440 201.345 1679.770 ;
        RECT 201.515 1679.660 201.685 1679.820 ;
        RECT 204.235 1679.660 204.405 1679.820 ;
        RECT 201.515 1679.260 201.685 1679.490 ;
        RECT 204.235 1679.260 204.405 1679.490 ;
        RECT 198.795 1679.200 199.690 1679.260 ;
        RECT 198.965 1679.030 199.690 1679.200 ;
        RECT 198.795 1678.970 199.690 1679.030 ;
        RECT 200.350 1679.200 202.850 1679.260 ;
        RECT 200.350 1679.030 201.515 1679.200 ;
        RECT 201.685 1679.030 202.850 1679.200 ;
        RECT 200.350 1678.970 202.850 1679.030 ;
        RECT 203.510 1679.200 204.405 1679.260 ;
        RECT 203.510 1679.030 204.235 1679.200 ;
        RECT 203.510 1678.970 204.405 1679.030 ;
        RECT 198.795 1678.740 198.965 1678.970 ;
        RECT 201.515 1678.740 201.685 1678.970 ;
        RECT 198.795 1678.410 198.965 1678.570 ;
        RECT 201.515 1678.410 201.685 1678.570 ;
        RECT 201.855 1678.460 202.875 1678.790 ;
        RECT 204.235 1678.740 204.405 1678.970 ;
        RECT 198.795 1678.280 199.765 1678.410 ;
        RECT 198.965 1678.110 199.765 1678.280 ;
        RECT 198.795 1678.080 199.765 1678.110 ;
        RECT 200.365 1678.290 201.685 1678.410 ;
        RECT 200.365 1678.280 202.485 1678.290 ;
        RECT 200.365 1678.110 201.515 1678.280 ;
        RECT 201.685 1678.120 202.485 1678.280 ;
        RECT 200.365 1678.080 201.685 1678.110 ;
        RECT 198.795 1677.820 198.965 1678.080 ;
        RECT 201.515 1677.820 201.685 1678.080 ;
        RECT 202.705 1677.950 202.875 1678.460 ;
        RECT 198.795 1677.570 198.965 1677.650 ;
        RECT 201.515 1677.570 201.685 1677.650 ;
        RECT 201.855 1677.620 202.875 1677.950 ;
        RECT 198.795 1677.360 199.445 1677.570 ;
        RECT 200.715 1677.450 201.685 1677.570 ;
        RECT 202.705 1677.465 202.875 1677.620 ;
        RECT 203.415 1678.540 204.065 1678.710 ;
        RECT 203.415 1677.870 203.585 1678.540 ;
        RECT 204.235 1678.370 204.405 1678.570 ;
        RECT 203.755 1678.280 204.405 1678.370 ;
        RECT 203.755 1678.110 204.235 1678.280 ;
        RECT 203.755 1678.040 204.405 1678.110 ;
        RECT 203.415 1677.700 204.060 1677.870 ;
        RECT 204.235 1677.820 204.405 1678.040 ;
        RECT 203.415 1677.465 203.585 1677.700 ;
        RECT 204.235 1677.530 204.405 1677.650 ;
        RECT 198.965 1677.240 199.445 1677.360 ;
        RECT 198.795 1676.900 198.965 1677.190 ;
        RECT 198.795 1676.440 199.445 1676.730 ;
        RECT 198.965 1676.400 199.445 1676.440 ;
        RECT 198.795 1675.980 198.965 1676.270 ;
        RECT 198.965 1675.810 199.445 1675.890 ;
        RECT 198.795 1675.560 199.445 1675.810 ;
        RECT 198.795 1675.520 198.965 1675.560 ;
        RECT 198.795 1675.060 198.965 1675.350 ;
        RECT 198.965 1674.890 199.445 1675.050 ;
        RECT 199.955 1674.960 200.125 1677.410 ;
        RECT 200.715 1677.360 202.485 1677.450 ;
        RECT 200.715 1677.240 201.515 1677.360 ;
        RECT 201.685 1677.280 202.485 1677.360 ;
        RECT 202.705 1677.290 203.585 1677.465 ;
        RECT 203.755 1677.360 204.405 1677.530 ;
        RECT 201.515 1676.900 201.685 1677.190 ;
      LAYER li1 ;
        RECT 201.855 1676.860 202.875 1677.030 ;
      LAYER li1 ;
        RECT 200.715 1676.690 201.685 1676.730 ;
        RECT 200.715 1676.440 202.485 1676.690 ;
        RECT 200.715 1676.400 201.515 1676.440 ;
        RECT 201.685 1676.360 202.485 1676.440 ;
        RECT 201.515 1675.980 201.685 1676.270 ;
      LAYER li1 ;
        RECT 202.705 1676.190 202.875 1676.860 ;
        RECT 201.855 1676.020 202.875 1676.190 ;
      LAYER li1 ;
        RECT 200.715 1675.810 201.515 1675.890 ;
        RECT 201.685 1675.810 202.485 1675.850 ;
        RECT 200.715 1675.560 202.485 1675.810 ;
        RECT 201.515 1675.520 202.485 1675.560 ;
      LAYER li1 ;
        RECT 202.705 1675.350 202.875 1676.020 ;
      LAYER li1 ;
        RECT 201.515 1675.060 201.685 1675.350 ;
      LAYER li1 ;
        RECT 201.855 1675.180 202.875 1675.350 ;
      LAYER li1 ;
        RECT 198.795 1674.720 199.445 1674.890 ;
        RECT 199.615 1674.785 200.495 1674.960 ;
        RECT 200.715 1674.890 201.515 1674.970 ;
        RECT 201.685 1674.890 202.485 1675.010 ;
        RECT 200.715 1674.800 202.485 1674.890 ;
        RECT 198.795 1674.600 198.965 1674.720 ;
        RECT 199.615 1674.550 199.785 1674.785 ;
        RECT 200.325 1674.630 200.495 1674.785 ;
        RECT 201.515 1674.680 202.485 1674.800 ;
        RECT 198.795 1674.210 198.965 1674.430 ;
        RECT 199.140 1674.380 199.785 1674.550 ;
        RECT 198.795 1674.140 199.445 1674.210 ;
        RECT 198.965 1673.970 199.445 1674.140 ;
        RECT 198.795 1673.880 199.445 1673.970 ;
        RECT 198.795 1673.680 198.965 1673.880 ;
        RECT 199.615 1673.710 199.785 1674.380 ;
        RECT 199.135 1673.540 199.785 1673.710 ;
        RECT 198.795 1673.280 198.965 1673.510 ;
      LAYER li1 ;
        RECT 199.955 1673.505 200.155 1674.605 ;
      LAYER li1 ;
        RECT 200.325 1674.300 201.345 1674.630 ;
        RECT 201.515 1674.600 201.685 1674.680 ;
      LAYER li1 ;
        RECT 202.705 1674.595 202.875 1675.180 ;
      LAYER li1 ;
        RECT 203.075 1674.840 203.245 1677.290 ;
        RECT 203.755 1677.200 204.235 1677.360 ;
      LAYER li1 ;
        RECT 203.415 1676.860 204.065 1677.030 ;
      LAYER li1 ;
        RECT 204.235 1676.900 204.405 1677.190 ;
      LAYER li1 ;
        RECT 203.415 1676.190 203.585 1676.860 ;
      LAYER li1 ;
        RECT 204.235 1676.690 204.405 1676.730 ;
        RECT 203.755 1676.440 204.405 1676.690 ;
        RECT 203.755 1676.360 204.235 1676.440 ;
      LAYER li1 ;
        RECT 203.415 1676.020 204.065 1676.190 ;
        RECT 203.415 1675.350 203.585 1676.020 ;
      LAYER li1 ;
        RECT 204.235 1675.980 204.405 1676.270 ;
        RECT 203.755 1675.810 204.235 1675.850 ;
        RECT 203.755 1675.520 204.405 1675.810 ;
      LAYER li1 ;
        RECT 203.415 1675.180 204.065 1675.350 ;
        RECT 203.415 1674.595 203.585 1675.180 ;
      LAYER li1 ;
        RECT 204.235 1675.060 204.405 1675.350 ;
        RECT 203.755 1674.890 204.235 1675.010 ;
        RECT 203.755 1674.680 204.405 1674.890 ;
        RECT 204.235 1674.600 204.405 1674.680 ;
      LAYER li1 ;
        RECT 202.705 1674.510 203.585 1674.595 ;
      LAYER li1 ;
        RECT 200.325 1673.790 200.495 1674.300 ;
        RECT 201.515 1674.170 201.685 1674.430 ;
      LAYER li1 ;
        RECT 201.855 1674.340 204.065 1674.510 ;
      LAYER li1 ;
        RECT 204.235 1674.170 204.405 1674.430 ;
        RECT 201.515 1674.140 202.835 1674.170 ;
        RECT 200.715 1673.970 201.515 1674.130 ;
        RECT 201.685 1673.970 202.835 1674.140 ;
        RECT 200.715 1673.960 202.835 1673.970 ;
        RECT 201.515 1673.840 202.835 1673.960 ;
        RECT 203.435 1674.140 204.405 1674.170 ;
        RECT 203.435 1673.970 204.235 1674.140 ;
        RECT 203.435 1673.840 204.405 1673.970 ;
        RECT 200.325 1673.460 201.345 1673.790 ;
        RECT 201.515 1673.680 201.685 1673.840 ;
        RECT 204.235 1673.680 204.405 1673.840 ;
        RECT 201.515 1673.280 201.685 1673.510 ;
        RECT 204.235 1673.280 204.405 1673.510 ;
        RECT 198.795 1673.220 199.690 1673.280 ;
        RECT 198.965 1673.050 199.690 1673.220 ;
        RECT 198.795 1672.990 199.690 1673.050 ;
        RECT 200.350 1673.220 202.850 1673.280 ;
        RECT 200.350 1673.050 201.515 1673.220 ;
        RECT 201.685 1673.050 202.850 1673.220 ;
        RECT 200.350 1672.990 202.850 1673.050 ;
        RECT 203.510 1673.220 204.405 1673.280 ;
        RECT 203.510 1673.050 204.235 1673.220 ;
        RECT 203.510 1672.990 204.405 1673.050 ;
        RECT 198.795 1672.905 198.965 1672.990 ;
        RECT 201.515 1672.905 201.685 1672.990 ;
        RECT 204.235 1672.905 204.405 1672.990 ;
        RECT 669.000 1117.040 669.145 1117.210 ;
        RECT 669.315 1117.040 669.605 1117.210 ;
        RECT 669.775 1117.040 670.065 1117.210 ;
        RECT 670.235 1117.040 670.525 1117.210 ;
        RECT 670.695 1117.040 670.985 1117.210 ;
        RECT 671.155 1117.040 671.445 1117.210 ;
        RECT 671.615 1117.040 671.905 1117.210 ;
        RECT 672.075 1117.040 672.365 1117.210 ;
        RECT 672.535 1117.040 672.825 1117.210 ;
        RECT 672.995 1117.040 673.285 1117.210 ;
        RECT 673.455 1117.040 673.745 1117.210 ;
        RECT 673.915 1117.040 674.205 1117.210 ;
        RECT 674.375 1117.040 674.665 1117.210 ;
        RECT 674.835 1117.040 675.125 1117.210 ;
        RECT 675.295 1117.040 675.585 1117.210 ;
        RECT 675.755 1117.040 676.045 1117.210 ;
        RECT 676.215 1117.040 676.505 1117.210 ;
        RECT 676.675 1117.040 676.965 1117.210 ;
        RECT 677.135 1117.040 677.425 1117.210 ;
        RECT 677.595 1117.040 677.885 1117.210 ;
        RECT 678.055 1117.040 678.345 1117.210 ;
        RECT 678.515 1117.040 678.805 1117.210 ;
        RECT 678.975 1117.040 679.265 1117.210 ;
        RECT 679.435 1117.040 679.725 1117.210 ;
        RECT 679.895 1117.040 680.185 1117.210 ;
        RECT 680.355 1117.040 680.645 1117.210 ;
        RECT 680.815 1117.040 681.105 1117.210 ;
        RECT 681.275 1117.040 681.565 1117.210 ;
        RECT 681.735 1117.040 682.025 1117.210 ;
        RECT 682.195 1117.040 682.485 1117.210 ;
        RECT 682.655 1117.040 682.945 1117.210 ;
        RECT 683.115 1117.040 683.405 1117.210 ;
        RECT 683.575 1117.040 683.865 1117.210 ;
        RECT 684.035 1117.040 684.325 1117.210 ;
        RECT 684.495 1117.040 684.785 1117.210 ;
        RECT 684.955 1117.040 685.245 1117.210 ;
        RECT 685.415 1117.040 685.705 1117.210 ;
        RECT 685.875 1117.040 686.165 1117.210 ;
        RECT 686.335 1117.040 686.625 1117.210 ;
        RECT 686.795 1117.040 687.085 1117.210 ;
        RECT 687.255 1117.040 687.545 1117.210 ;
        RECT 687.715 1117.040 688.005 1117.210 ;
        RECT 688.175 1117.040 688.465 1117.210 ;
        RECT 688.635 1117.040 688.925 1117.210 ;
        RECT 689.095 1117.040 689.385 1117.210 ;
        RECT 689.555 1117.040 689.845 1117.210 ;
        RECT 690.015 1117.040 690.305 1117.210 ;
        RECT 690.475 1117.040 690.765 1117.210 ;
        RECT 690.935 1117.040 691.225 1117.210 ;
        RECT 691.395 1117.040 691.685 1117.210 ;
        RECT 691.855 1117.040 692.145 1117.210 ;
        RECT 692.315 1117.040 692.605 1117.210 ;
        RECT 692.775 1117.040 693.065 1117.210 ;
        RECT 693.235 1117.040 693.525 1117.210 ;
        RECT 693.695 1117.040 693.985 1117.210 ;
        RECT 694.155 1117.040 694.445 1117.210 ;
        RECT 694.615 1117.040 694.905 1117.210 ;
        RECT 695.075 1117.040 695.365 1117.210 ;
        RECT 695.535 1117.040 695.825 1117.210 ;
        RECT 695.995 1117.040 696.285 1117.210 ;
        RECT 696.455 1117.040 696.745 1117.210 ;
        RECT 696.915 1117.040 697.205 1117.210 ;
        RECT 697.375 1117.040 697.665 1117.210 ;
        RECT 697.835 1117.040 698.125 1117.210 ;
        RECT 698.295 1117.040 698.585 1117.210 ;
        RECT 698.755 1117.040 699.045 1117.210 ;
        RECT 699.215 1117.040 699.505 1117.210 ;
        RECT 699.675 1117.040 699.965 1117.210 ;
        RECT 700.135 1117.040 700.425 1117.210 ;
        RECT 700.595 1117.040 700.885 1117.210 ;
        RECT 701.055 1117.040 701.345 1117.210 ;
        RECT 701.515 1117.040 701.805 1117.210 ;
        RECT 701.975 1117.040 702.265 1117.210 ;
        RECT 702.435 1117.040 702.725 1117.210 ;
        RECT 702.895 1117.040 703.185 1117.210 ;
        RECT 703.355 1117.040 703.645 1117.210 ;
        RECT 703.815 1117.040 704.105 1117.210 ;
        RECT 704.275 1117.040 704.565 1117.210 ;
        RECT 704.735 1117.040 705.025 1117.210 ;
        RECT 705.195 1117.040 705.485 1117.210 ;
        RECT 705.655 1117.040 705.945 1117.210 ;
        RECT 706.115 1117.040 706.405 1117.210 ;
        RECT 706.575 1117.040 706.865 1117.210 ;
        RECT 707.035 1117.040 707.325 1117.210 ;
        RECT 707.495 1117.040 707.785 1117.210 ;
        RECT 707.955 1117.040 708.245 1117.210 ;
        RECT 708.415 1117.040 708.705 1117.210 ;
        RECT 708.875 1117.040 709.165 1117.210 ;
        RECT 709.335 1117.040 709.625 1117.210 ;
        RECT 709.795 1117.040 710.085 1117.210 ;
        RECT 710.255 1117.040 710.545 1117.210 ;
        RECT 710.715 1117.040 711.005 1117.210 ;
        RECT 711.175 1117.040 711.465 1117.210 ;
        RECT 711.635 1117.040 711.925 1117.210 ;
        RECT 712.095 1117.040 712.385 1117.210 ;
        RECT 712.555 1117.040 712.845 1117.210 ;
        RECT 713.015 1117.040 713.305 1117.210 ;
        RECT 713.475 1117.040 713.765 1117.210 ;
        RECT 713.935 1117.040 714.225 1117.210 ;
        RECT 714.395 1117.040 714.685 1117.210 ;
        RECT 714.855 1117.040 715.145 1117.210 ;
        RECT 715.315 1117.040 715.605 1117.210 ;
        RECT 715.775 1117.040 716.065 1117.210 ;
        RECT 716.235 1117.040 716.525 1117.210 ;
        RECT 716.695 1117.040 716.985 1117.210 ;
        RECT 717.155 1117.040 717.445 1117.210 ;
        RECT 717.615 1117.040 717.905 1117.210 ;
        RECT 718.075 1117.040 718.365 1117.210 ;
        RECT 718.535 1117.040 718.825 1117.210 ;
        RECT 718.995 1117.040 719.285 1117.210 ;
        RECT 719.455 1117.040 719.745 1117.210 ;
        RECT 719.915 1117.040 720.205 1117.210 ;
        RECT 720.375 1117.040 720.665 1117.210 ;
        RECT 720.835 1117.040 721.125 1117.210 ;
        RECT 721.295 1117.040 721.585 1117.210 ;
        RECT 721.755 1117.040 722.045 1117.210 ;
        RECT 722.215 1117.040 722.505 1117.210 ;
        RECT 722.675 1117.040 722.965 1117.210 ;
        RECT 723.135 1117.040 723.425 1117.210 ;
        RECT 723.595 1117.040 723.885 1117.210 ;
        RECT 724.055 1117.040 724.345 1117.210 ;
        RECT 724.515 1117.040 724.805 1117.210 ;
        RECT 724.975 1117.040 725.265 1117.210 ;
        RECT 725.435 1117.040 725.725 1117.210 ;
        RECT 725.895 1117.040 726.185 1117.210 ;
        RECT 726.355 1117.040 726.645 1117.210 ;
        RECT 726.815 1117.040 727.105 1117.210 ;
        RECT 727.275 1117.040 727.565 1117.210 ;
        RECT 727.735 1117.040 728.025 1117.210 ;
        RECT 728.195 1117.040 728.485 1117.210 ;
        RECT 728.655 1117.040 728.945 1117.210 ;
        RECT 729.115 1117.040 729.405 1117.210 ;
        RECT 729.575 1117.040 729.865 1117.210 ;
        RECT 730.035 1117.040 730.325 1117.210 ;
        RECT 730.495 1117.040 730.785 1117.210 ;
        RECT 730.955 1117.040 731.245 1117.210 ;
        RECT 731.415 1117.040 731.705 1117.210 ;
        RECT 731.875 1117.040 732.165 1117.210 ;
        RECT 732.335 1117.040 732.625 1117.210 ;
        RECT 732.795 1117.040 733.085 1117.210 ;
        RECT 733.255 1117.040 733.545 1117.210 ;
        RECT 733.715 1117.040 734.005 1117.210 ;
        RECT 734.175 1117.040 734.465 1117.210 ;
        RECT 734.635 1117.040 734.925 1117.210 ;
        RECT 735.095 1117.040 735.385 1117.210 ;
        RECT 735.555 1117.040 735.845 1117.210 ;
        RECT 736.015 1117.040 736.305 1117.210 ;
        RECT 736.475 1117.040 736.765 1117.210 ;
        RECT 736.935 1117.040 737.225 1117.210 ;
        RECT 737.395 1117.040 737.685 1117.210 ;
        RECT 737.855 1117.040 738.145 1117.210 ;
        RECT 738.315 1117.040 738.605 1117.210 ;
        RECT 738.775 1117.040 739.065 1117.210 ;
        RECT 739.235 1117.040 739.525 1117.210 ;
        RECT 739.695 1117.040 739.985 1117.210 ;
        RECT 740.155 1117.040 740.445 1117.210 ;
        RECT 740.615 1117.040 740.905 1117.210 ;
        RECT 741.075 1117.040 741.365 1117.210 ;
        RECT 741.535 1117.040 741.825 1117.210 ;
        RECT 741.995 1117.040 742.285 1117.210 ;
        RECT 742.455 1117.040 742.745 1117.210 ;
        RECT 742.915 1117.040 743.205 1117.210 ;
        RECT 743.375 1117.040 743.665 1117.210 ;
        RECT 743.835 1117.040 744.125 1117.210 ;
        RECT 744.295 1117.040 744.585 1117.210 ;
        RECT 744.755 1117.040 745.045 1117.210 ;
        RECT 745.215 1117.040 745.505 1117.210 ;
        RECT 745.675 1117.040 745.965 1117.210 ;
        RECT 746.135 1117.040 746.425 1117.210 ;
        RECT 746.595 1117.040 746.885 1117.210 ;
        RECT 747.055 1117.040 747.345 1117.210 ;
        RECT 747.515 1117.040 747.805 1117.210 ;
        RECT 747.975 1117.040 748.265 1117.210 ;
        RECT 748.435 1117.040 748.725 1117.210 ;
        RECT 748.895 1117.040 749.185 1117.210 ;
        RECT 749.355 1117.040 749.645 1117.210 ;
        RECT 749.815 1117.040 750.105 1117.210 ;
        RECT 750.275 1117.040 750.565 1117.210 ;
        RECT 750.735 1117.040 751.025 1117.210 ;
        RECT 751.195 1117.040 751.485 1117.210 ;
        RECT 751.655 1117.040 751.945 1117.210 ;
        RECT 752.115 1117.040 752.405 1117.210 ;
        RECT 752.575 1117.040 752.865 1117.210 ;
        RECT 753.035 1117.040 753.325 1117.210 ;
        RECT 753.495 1117.040 753.785 1117.210 ;
        RECT 753.955 1117.040 754.245 1117.210 ;
        RECT 754.415 1117.040 754.705 1117.210 ;
        RECT 754.875 1117.040 755.165 1117.210 ;
        RECT 755.335 1117.040 755.625 1117.210 ;
        RECT 755.795 1117.040 756.085 1117.210 ;
        RECT 756.255 1117.040 756.545 1117.210 ;
        RECT 756.715 1117.040 757.005 1117.210 ;
        RECT 757.175 1117.040 757.465 1117.210 ;
        RECT 757.635 1117.040 757.925 1117.210 ;
        RECT 758.095 1117.040 758.385 1117.210 ;
        RECT 758.555 1117.040 758.845 1117.210 ;
        RECT 759.015 1117.040 759.305 1117.210 ;
        RECT 759.475 1117.040 759.765 1117.210 ;
        RECT 759.935 1117.040 760.225 1117.210 ;
        RECT 760.395 1117.040 760.685 1117.210 ;
        RECT 760.855 1117.040 761.145 1117.210 ;
        RECT 761.315 1117.040 761.605 1117.210 ;
        RECT 761.775 1117.040 762.065 1117.210 ;
        RECT 762.235 1117.040 762.525 1117.210 ;
        RECT 762.695 1117.040 762.985 1117.210 ;
        RECT 763.155 1117.040 763.445 1117.210 ;
        RECT 763.615 1117.040 763.905 1117.210 ;
        RECT 764.075 1117.040 764.365 1117.210 ;
        RECT 764.535 1117.040 764.825 1117.210 ;
        RECT 764.995 1117.040 765.285 1117.210 ;
        RECT 765.455 1117.040 765.745 1117.210 ;
        RECT 765.915 1117.040 766.205 1117.210 ;
        RECT 766.375 1117.040 766.665 1117.210 ;
        RECT 766.835 1117.040 767.125 1117.210 ;
        RECT 767.295 1117.040 767.585 1117.210 ;
        RECT 767.755 1117.040 768.045 1117.210 ;
        RECT 768.215 1117.040 768.505 1117.210 ;
        RECT 768.675 1117.040 768.965 1117.210 ;
        RECT 769.135 1117.040 769.425 1117.210 ;
        RECT 769.595 1117.040 769.885 1117.210 ;
        RECT 770.055 1117.040 770.345 1117.210 ;
        RECT 770.515 1117.040 770.805 1117.210 ;
        RECT 770.975 1117.040 771.120 1117.210 ;
        RECT 1969.000 1117.040 1969.145 1117.210 ;
        RECT 1969.315 1117.040 1969.605 1117.210 ;
        RECT 1969.775 1117.040 1970.065 1117.210 ;
        RECT 1970.235 1117.040 1970.525 1117.210 ;
        RECT 1970.695 1117.040 1970.985 1117.210 ;
        RECT 1971.155 1117.040 1971.445 1117.210 ;
        RECT 1971.615 1117.040 1971.905 1117.210 ;
        RECT 1972.075 1117.040 1972.365 1117.210 ;
        RECT 1972.535 1117.040 1972.825 1117.210 ;
        RECT 1972.995 1117.040 1973.285 1117.210 ;
        RECT 1973.455 1117.040 1973.745 1117.210 ;
        RECT 1973.915 1117.040 1974.205 1117.210 ;
        RECT 1974.375 1117.040 1974.665 1117.210 ;
        RECT 1974.835 1117.040 1975.125 1117.210 ;
        RECT 1975.295 1117.040 1975.585 1117.210 ;
        RECT 1975.755 1117.040 1976.045 1117.210 ;
        RECT 1976.215 1117.040 1976.505 1117.210 ;
        RECT 1976.675 1117.040 1976.965 1117.210 ;
        RECT 1977.135 1117.040 1977.425 1117.210 ;
        RECT 1977.595 1117.040 1977.885 1117.210 ;
        RECT 1978.055 1117.040 1978.345 1117.210 ;
        RECT 1978.515 1117.040 1978.805 1117.210 ;
        RECT 1978.975 1117.040 1979.265 1117.210 ;
        RECT 1979.435 1117.040 1979.725 1117.210 ;
        RECT 1979.895 1117.040 1980.185 1117.210 ;
        RECT 1980.355 1117.040 1980.645 1117.210 ;
        RECT 1980.815 1117.040 1981.105 1117.210 ;
        RECT 1981.275 1117.040 1981.565 1117.210 ;
        RECT 1981.735 1117.040 1982.025 1117.210 ;
        RECT 1982.195 1117.040 1982.485 1117.210 ;
        RECT 1982.655 1117.040 1982.945 1117.210 ;
        RECT 1983.115 1117.040 1983.405 1117.210 ;
        RECT 1983.575 1117.040 1983.865 1117.210 ;
        RECT 1984.035 1117.040 1984.325 1117.210 ;
        RECT 1984.495 1117.040 1984.785 1117.210 ;
        RECT 1984.955 1117.040 1985.245 1117.210 ;
        RECT 1985.415 1117.040 1985.705 1117.210 ;
        RECT 1985.875 1117.040 1986.165 1117.210 ;
        RECT 1986.335 1117.040 1986.625 1117.210 ;
        RECT 1986.795 1117.040 1987.085 1117.210 ;
        RECT 1987.255 1117.040 1987.545 1117.210 ;
        RECT 1987.715 1117.040 1988.005 1117.210 ;
        RECT 1988.175 1117.040 1988.465 1117.210 ;
        RECT 1988.635 1117.040 1988.925 1117.210 ;
        RECT 1989.095 1117.040 1989.385 1117.210 ;
        RECT 1989.555 1117.040 1989.845 1117.210 ;
        RECT 1990.015 1117.040 1990.305 1117.210 ;
        RECT 1990.475 1117.040 1990.765 1117.210 ;
        RECT 1990.935 1117.040 1991.225 1117.210 ;
        RECT 1991.395 1117.040 1991.685 1117.210 ;
        RECT 1991.855 1117.040 1992.145 1117.210 ;
        RECT 1992.315 1117.040 1992.605 1117.210 ;
        RECT 1992.775 1117.040 1993.065 1117.210 ;
        RECT 1993.235 1117.040 1993.525 1117.210 ;
        RECT 1993.695 1117.040 1993.985 1117.210 ;
        RECT 1994.155 1117.040 1994.445 1117.210 ;
        RECT 1994.615 1117.040 1994.905 1117.210 ;
        RECT 1995.075 1117.040 1995.365 1117.210 ;
        RECT 1995.535 1117.040 1995.825 1117.210 ;
        RECT 1995.995 1117.040 1996.285 1117.210 ;
        RECT 1996.455 1117.040 1996.745 1117.210 ;
        RECT 1996.915 1117.040 1997.205 1117.210 ;
        RECT 1997.375 1117.040 1997.665 1117.210 ;
        RECT 1997.835 1117.040 1998.125 1117.210 ;
        RECT 1998.295 1117.040 1998.585 1117.210 ;
        RECT 1998.755 1117.040 1999.045 1117.210 ;
        RECT 1999.215 1117.040 1999.505 1117.210 ;
        RECT 1999.675 1117.040 1999.965 1117.210 ;
        RECT 2000.135 1117.040 2000.425 1117.210 ;
        RECT 2000.595 1117.040 2000.885 1117.210 ;
        RECT 2001.055 1117.040 2001.345 1117.210 ;
        RECT 2001.515 1117.040 2001.805 1117.210 ;
        RECT 2001.975 1117.040 2002.265 1117.210 ;
        RECT 2002.435 1117.040 2002.725 1117.210 ;
        RECT 2002.895 1117.040 2003.185 1117.210 ;
        RECT 2003.355 1117.040 2003.645 1117.210 ;
        RECT 2003.815 1117.040 2004.105 1117.210 ;
        RECT 2004.275 1117.040 2004.565 1117.210 ;
        RECT 2004.735 1117.040 2005.025 1117.210 ;
        RECT 2005.195 1117.040 2005.485 1117.210 ;
        RECT 2005.655 1117.040 2005.945 1117.210 ;
        RECT 2006.115 1117.040 2006.405 1117.210 ;
        RECT 2006.575 1117.040 2006.865 1117.210 ;
        RECT 2007.035 1117.040 2007.325 1117.210 ;
        RECT 2007.495 1117.040 2007.785 1117.210 ;
        RECT 2007.955 1117.040 2008.245 1117.210 ;
        RECT 2008.415 1117.040 2008.705 1117.210 ;
        RECT 2008.875 1117.040 2009.165 1117.210 ;
        RECT 2009.335 1117.040 2009.625 1117.210 ;
        RECT 2009.795 1117.040 2010.085 1117.210 ;
        RECT 2010.255 1117.040 2010.545 1117.210 ;
        RECT 2010.715 1117.040 2011.005 1117.210 ;
        RECT 2011.175 1117.040 2011.465 1117.210 ;
        RECT 2011.635 1117.040 2011.925 1117.210 ;
        RECT 2012.095 1117.040 2012.385 1117.210 ;
        RECT 2012.555 1117.040 2012.845 1117.210 ;
        RECT 2013.015 1117.040 2013.305 1117.210 ;
        RECT 2013.475 1117.040 2013.765 1117.210 ;
        RECT 2013.935 1117.040 2014.225 1117.210 ;
        RECT 2014.395 1117.040 2014.685 1117.210 ;
        RECT 2014.855 1117.040 2015.145 1117.210 ;
        RECT 2015.315 1117.040 2015.605 1117.210 ;
        RECT 2015.775 1117.040 2016.065 1117.210 ;
        RECT 2016.235 1117.040 2016.525 1117.210 ;
        RECT 2016.695 1117.040 2016.985 1117.210 ;
        RECT 2017.155 1117.040 2017.445 1117.210 ;
        RECT 2017.615 1117.040 2017.905 1117.210 ;
        RECT 2018.075 1117.040 2018.365 1117.210 ;
        RECT 2018.535 1117.040 2018.825 1117.210 ;
        RECT 2018.995 1117.040 2019.285 1117.210 ;
        RECT 2019.455 1117.040 2019.745 1117.210 ;
        RECT 2019.915 1117.040 2020.205 1117.210 ;
        RECT 2020.375 1117.040 2020.665 1117.210 ;
        RECT 2020.835 1117.040 2021.125 1117.210 ;
        RECT 2021.295 1117.040 2021.585 1117.210 ;
        RECT 2021.755 1117.040 2022.045 1117.210 ;
        RECT 2022.215 1117.040 2022.505 1117.210 ;
        RECT 2022.675 1117.040 2022.965 1117.210 ;
        RECT 2023.135 1117.040 2023.425 1117.210 ;
        RECT 2023.595 1117.040 2023.885 1117.210 ;
        RECT 2024.055 1117.040 2024.345 1117.210 ;
        RECT 2024.515 1117.040 2024.805 1117.210 ;
        RECT 2024.975 1117.040 2025.265 1117.210 ;
        RECT 2025.435 1117.040 2025.725 1117.210 ;
        RECT 2025.895 1117.040 2026.185 1117.210 ;
        RECT 2026.355 1117.040 2026.645 1117.210 ;
        RECT 2026.815 1117.040 2027.105 1117.210 ;
        RECT 2027.275 1117.040 2027.565 1117.210 ;
        RECT 2027.735 1117.040 2028.025 1117.210 ;
        RECT 2028.195 1117.040 2028.485 1117.210 ;
        RECT 2028.655 1117.040 2028.945 1117.210 ;
        RECT 2029.115 1117.040 2029.405 1117.210 ;
        RECT 2029.575 1117.040 2029.865 1117.210 ;
        RECT 2030.035 1117.040 2030.325 1117.210 ;
        RECT 2030.495 1117.040 2030.785 1117.210 ;
        RECT 2030.955 1117.040 2031.245 1117.210 ;
        RECT 2031.415 1117.040 2031.705 1117.210 ;
        RECT 2031.875 1117.040 2032.165 1117.210 ;
        RECT 2032.335 1117.040 2032.625 1117.210 ;
        RECT 2032.795 1117.040 2033.085 1117.210 ;
        RECT 2033.255 1117.040 2033.545 1117.210 ;
        RECT 2033.715 1117.040 2034.005 1117.210 ;
        RECT 2034.175 1117.040 2034.465 1117.210 ;
        RECT 2034.635 1117.040 2034.925 1117.210 ;
        RECT 2035.095 1117.040 2035.385 1117.210 ;
        RECT 2035.555 1117.040 2035.845 1117.210 ;
        RECT 2036.015 1117.040 2036.305 1117.210 ;
        RECT 2036.475 1117.040 2036.765 1117.210 ;
        RECT 2036.935 1117.040 2037.225 1117.210 ;
        RECT 2037.395 1117.040 2037.685 1117.210 ;
        RECT 2037.855 1117.040 2038.145 1117.210 ;
        RECT 2038.315 1117.040 2038.605 1117.210 ;
        RECT 2038.775 1117.040 2039.065 1117.210 ;
        RECT 2039.235 1117.040 2039.525 1117.210 ;
        RECT 2039.695 1117.040 2039.985 1117.210 ;
        RECT 2040.155 1117.040 2040.445 1117.210 ;
        RECT 2040.615 1117.040 2040.905 1117.210 ;
        RECT 2041.075 1117.040 2041.365 1117.210 ;
        RECT 2041.535 1117.040 2041.825 1117.210 ;
        RECT 2041.995 1117.040 2042.285 1117.210 ;
        RECT 2042.455 1117.040 2042.745 1117.210 ;
        RECT 2042.915 1117.040 2043.205 1117.210 ;
        RECT 2043.375 1117.040 2043.665 1117.210 ;
        RECT 2043.835 1117.040 2044.125 1117.210 ;
        RECT 2044.295 1117.040 2044.585 1117.210 ;
        RECT 2044.755 1117.040 2045.045 1117.210 ;
        RECT 2045.215 1117.040 2045.505 1117.210 ;
        RECT 2045.675 1117.040 2045.965 1117.210 ;
        RECT 2046.135 1117.040 2046.425 1117.210 ;
        RECT 2046.595 1117.040 2046.885 1117.210 ;
        RECT 2047.055 1117.040 2047.345 1117.210 ;
        RECT 2047.515 1117.040 2047.805 1117.210 ;
        RECT 2047.975 1117.040 2048.265 1117.210 ;
        RECT 2048.435 1117.040 2048.725 1117.210 ;
        RECT 2048.895 1117.040 2049.185 1117.210 ;
        RECT 2049.355 1117.040 2049.645 1117.210 ;
        RECT 2049.815 1117.040 2050.105 1117.210 ;
        RECT 2050.275 1117.040 2050.565 1117.210 ;
        RECT 2050.735 1117.040 2051.025 1117.210 ;
        RECT 2051.195 1117.040 2051.485 1117.210 ;
        RECT 2051.655 1117.040 2051.945 1117.210 ;
        RECT 2052.115 1117.040 2052.405 1117.210 ;
        RECT 2052.575 1117.040 2052.865 1117.210 ;
        RECT 2053.035 1117.040 2053.325 1117.210 ;
        RECT 2053.495 1117.040 2053.785 1117.210 ;
        RECT 2053.955 1117.040 2054.245 1117.210 ;
        RECT 2054.415 1117.040 2054.705 1117.210 ;
        RECT 2054.875 1117.040 2055.165 1117.210 ;
        RECT 2055.335 1117.040 2055.625 1117.210 ;
        RECT 2055.795 1117.040 2056.085 1117.210 ;
        RECT 2056.255 1117.040 2056.545 1117.210 ;
        RECT 2056.715 1117.040 2057.005 1117.210 ;
        RECT 2057.175 1117.040 2057.465 1117.210 ;
        RECT 2057.635 1117.040 2057.925 1117.210 ;
        RECT 2058.095 1117.040 2058.385 1117.210 ;
        RECT 2058.555 1117.040 2058.845 1117.210 ;
        RECT 2059.015 1117.040 2059.305 1117.210 ;
        RECT 2059.475 1117.040 2059.765 1117.210 ;
        RECT 2059.935 1117.040 2060.225 1117.210 ;
        RECT 2060.395 1117.040 2060.685 1117.210 ;
        RECT 2060.855 1117.040 2061.145 1117.210 ;
        RECT 2061.315 1117.040 2061.605 1117.210 ;
        RECT 2061.775 1117.040 2062.065 1117.210 ;
        RECT 2062.235 1117.040 2062.525 1117.210 ;
        RECT 2062.695 1117.040 2062.985 1117.210 ;
        RECT 2063.155 1117.040 2063.445 1117.210 ;
        RECT 2063.615 1117.040 2063.905 1117.210 ;
        RECT 2064.075 1117.040 2064.365 1117.210 ;
        RECT 2064.535 1117.040 2064.825 1117.210 ;
        RECT 2064.995 1117.040 2065.285 1117.210 ;
        RECT 2065.455 1117.040 2065.745 1117.210 ;
        RECT 2065.915 1117.040 2066.205 1117.210 ;
        RECT 2066.375 1117.040 2066.665 1117.210 ;
        RECT 2066.835 1117.040 2067.125 1117.210 ;
        RECT 2067.295 1117.040 2067.585 1117.210 ;
        RECT 2067.755 1117.040 2068.045 1117.210 ;
        RECT 2068.215 1117.040 2068.505 1117.210 ;
        RECT 2068.675 1117.040 2068.965 1117.210 ;
        RECT 2069.135 1117.040 2069.425 1117.210 ;
        RECT 2069.595 1117.040 2069.885 1117.210 ;
        RECT 2070.055 1117.040 2070.345 1117.210 ;
        RECT 2070.515 1117.040 2070.805 1117.210 ;
        RECT 2070.975 1117.040 2071.120 1117.210 ;
        RECT 669.085 1116.315 669.375 1117.040 ;
        RECT 669.935 1116.240 670.265 1117.040 ;
      LAYER li1 ;
        RECT 670.435 1116.390 670.605 1116.870 ;
      LAYER li1 ;
        RECT 670.775 1116.560 671.105 1117.040 ;
      LAYER li1 ;
        RECT 671.275 1116.390 671.445 1116.870 ;
      LAYER li1 ;
        RECT 671.615 1116.560 671.945 1117.040 ;
      LAYER li1 ;
        RECT 672.115 1116.390 672.285 1116.870 ;
      LAYER li1 ;
        RECT 672.455 1116.560 672.785 1117.040 ;
      LAYER li1 ;
        RECT 672.955 1116.390 673.125 1116.870 ;
      LAYER li1 ;
        RECT 673.295 1116.560 673.625 1117.040 ;
        RECT 673.795 1116.390 673.965 1116.865 ;
        RECT 674.135 1116.560 674.465 1117.040 ;
        RECT 674.635 1116.390 674.805 1116.870 ;
      LAYER li1 ;
        RECT 670.435 1116.220 673.125 1116.390 ;
      LAYER li1 ;
        RECT 673.385 1116.220 674.805 1116.390 ;
        RECT 675.065 1116.315 675.355 1117.040 ;
        RECT 675.915 1116.240 676.245 1117.040 ;
      LAYER li1 ;
        RECT 676.415 1116.390 676.585 1116.870 ;
      LAYER li1 ;
        RECT 676.755 1116.560 677.085 1117.040 ;
      LAYER li1 ;
        RECT 677.255 1116.390 677.425 1116.870 ;
      LAYER li1 ;
        RECT 677.595 1116.560 677.925 1117.040 ;
      LAYER li1 ;
        RECT 678.095 1116.390 678.265 1116.870 ;
      LAYER li1 ;
        RECT 678.435 1116.560 678.765 1117.040 ;
      LAYER li1 ;
        RECT 678.935 1116.390 679.105 1116.870 ;
      LAYER li1 ;
        RECT 679.275 1116.560 679.605 1117.040 ;
        RECT 679.775 1116.390 679.945 1116.865 ;
        RECT 680.115 1116.560 680.445 1117.040 ;
        RECT 680.615 1116.390 680.785 1116.870 ;
      LAYER li1 ;
        RECT 676.415 1116.220 679.105 1116.390 ;
      LAYER li1 ;
        RECT 679.365 1116.220 680.785 1116.390 ;
        RECT 681.045 1116.315 681.335 1117.040 ;
        RECT 681.895 1116.240 682.225 1117.040 ;
      LAYER li1 ;
        RECT 682.395 1116.390 682.565 1116.870 ;
      LAYER li1 ;
        RECT 682.735 1116.560 683.065 1117.040 ;
      LAYER li1 ;
        RECT 683.235 1116.390 683.405 1116.870 ;
      LAYER li1 ;
        RECT 683.575 1116.560 683.905 1117.040 ;
      LAYER li1 ;
        RECT 684.075 1116.390 684.245 1116.870 ;
      LAYER li1 ;
        RECT 684.415 1116.560 684.745 1117.040 ;
      LAYER li1 ;
        RECT 684.915 1116.390 685.085 1116.870 ;
      LAYER li1 ;
        RECT 685.255 1116.560 685.585 1117.040 ;
        RECT 685.755 1116.390 685.925 1116.865 ;
        RECT 686.095 1116.560 686.425 1117.040 ;
        RECT 686.595 1116.390 686.765 1116.870 ;
      LAYER li1 ;
        RECT 682.395 1116.220 685.085 1116.390 ;
      LAYER li1 ;
        RECT 685.345 1116.220 686.765 1116.390 ;
        RECT 687.025 1116.315 687.315 1117.040 ;
        RECT 687.875 1116.240 688.205 1117.040 ;
      LAYER li1 ;
        RECT 688.375 1116.390 688.545 1116.870 ;
      LAYER li1 ;
        RECT 688.715 1116.560 689.045 1117.040 ;
      LAYER li1 ;
        RECT 689.215 1116.390 689.385 1116.870 ;
      LAYER li1 ;
        RECT 689.555 1116.560 689.885 1117.040 ;
      LAYER li1 ;
        RECT 690.055 1116.390 690.225 1116.870 ;
      LAYER li1 ;
        RECT 690.395 1116.560 690.725 1117.040 ;
      LAYER li1 ;
        RECT 690.895 1116.390 691.065 1116.870 ;
      LAYER li1 ;
        RECT 691.235 1116.560 691.565 1117.040 ;
        RECT 691.735 1116.390 691.905 1116.865 ;
        RECT 692.075 1116.560 692.405 1117.040 ;
        RECT 692.575 1116.390 692.745 1116.870 ;
      LAYER li1 ;
        RECT 688.375 1116.220 691.065 1116.390 ;
      LAYER li1 ;
        RECT 691.325 1116.220 692.745 1116.390 ;
        RECT 693.005 1116.315 693.295 1117.040 ;
        RECT 693.855 1116.240 694.185 1117.040 ;
      LAYER li1 ;
        RECT 694.355 1116.390 694.525 1116.870 ;
      LAYER li1 ;
        RECT 694.695 1116.560 695.025 1117.040 ;
      LAYER li1 ;
        RECT 695.195 1116.390 695.365 1116.870 ;
      LAYER li1 ;
        RECT 695.535 1116.560 695.865 1117.040 ;
      LAYER li1 ;
        RECT 696.035 1116.390 696.205 1116.870 ;
      LAYER li1 ;
        RECT 696.375 1116.560 696.705 1117.040 ;
      LAYER li1 ;
        RECT 696.875 1116.390 697.045 1116.870 ;
      LAYER li1 ;
        RECT 697.215 1116.560 697.545 1117.040 ;
        RECT 697.715 1116.390 697.885 1116.865 ;
        RECT 698.055 1116.560 698.385 1117.040 ;
        RECT 698.555 1116.390 698.725 1116.870 ;
      LAYER li1 ;
        RECT 694.355 1116.220 697.045 1116.390 ;
      LAYER li1 ;
        RECT 697.305 1116.220 698.725 1116.390 ;
        RECT 698.985 1116.315 699.275 1117.040 ;
        RECT 699.835 1116.240 700.165 1117.040 ;
      LAYER li1 ;
        RECT 700.335 1116.390 700.505 1116.870 ;
      LAYER li1 ;
        RECT 700.675 1116.560 701.005 1117.040 ;
      LAYER li1 ;
        RECT 701.175 1116.390 701.345 1116.870 ;
      LAYER li1 ;
        RECT 701.515 1116.560 701.845 1117.040 ;
      LAYER li1 ;
        RECT 702.015 1116.390 702.185 1116.870 ;
      LAYER li1 ;
        RECT 702.355 1116.560 702.685 1117.040 ;
      LAYER li1 ;
        RECT 702.855 1116.390 703.025 1116.870 ;
      LAYER li1 ;
        RECT 703.195 1116.560 703.525 1117.040 ;
        RECT 703.695 1116.390 703.865 1116.865 ;
        RECT 704.035 1116.560 704.365 1117.040 ;
        RECT 704.535 1116.390 704.705 1116.870 ;
      LAYER li1 ;
        RECT 700.335 1116.220 703.025 1116.390 ;
      LAYER li1 ;
        RECT 703.285 1116.220 704.705 1116.390 ;
        RECT 704.965 1116.315 705.255 1117.040 ;
        RECT 705.815 1116.240 706.145 1117.040 ;
      LAYER li1 ;
        RECT 706.315 1116.390 706.485 1116.870 ;
      LAYER li1 ;
        RECT 706.655 1116.560 706.985 1117.040 ;
      LAYER li1 ;
        RECT 707.155 1116.390 707.325 1116.870 ;
      LAYER li1 ;
        RECT 707.495 1116.560 707.825 1117.040 ;
      LAYER li1 ;
        RECT 707.995 1116.390 708.165 1116.870 ;
      LAYER li1 ;
        RECT 708.335 1116.560 708.665 1117.040 ;
      LAYER li1 ;
        RECT 708.835 1116.390 709.005 1116.870 ;
      LAYER li1 ;
        RECT 709.175 1116.560 709.505 1117.040 ;
        RECT 709.675 1116.390 709.845 1116.865 ;
        RECT 710.015 1116.560 710.345 1117.040 ;
        RECT 710.515 1116.390 710.685 1116.870 ;
      LAYER li1 ;
        RECT 706.315 1116.220 709.005 1116.390 ;
      LAYER li1 ;
        RECT 709.265 1116.220 710.685 1116.390 ;
        RECT 710.945 1116.315 711.235 1117.040 ;
        RECT 711.795 1116.240 712.125 1117.040 ;
      LAYER li1 ;
        RECT 712.295 1116.390 712.465 1116.870 ;
      LAYER li1 ;
        RECT 712.635 1116.560 712.965 1117.040 ;
      LAYER li1 ;
        RECT 713.135 1116.390 713.305 1116.870 ;
      LAYER li1 ;
        RECT 713.475 1116.560 713.805 1117.040 ;
      LAYER li1 ;
        RECT 713.975 1116.390 714.145 1116.870 ;
      LAYER li1 ;
        RECT 714.315 1116.560 714.645 1117.040 ;
      LAYER li1 ;
        RECT 714.815 1116.390 714.985 1116.870 ;
      LAYER li1 ;
        RECT 715.155 1116.560 715.485 1117.040 ;
        RECT 715.655 1116.390 715.825 1116.865 ;
        RECT 715.995 1116.560 716.325 1117.040 ;
        RECT 716.495 1116.390 716.665 1116.870 ;
      LAYER li1 ;
        RECT 712.295 1116.220 714.985 1116.390 ;
      LAYER li1 ;
        RECT 715.245 1116.220 716.665 1116.390 ;
        RECT 716.925 1116.315 717.215 1117.040 ;
        RECT 717.775 1116.240 718.105 1117.040 ;
      LAYER li1 ;
        RECT 718.275 1116.390 718.445 1116.870 ;
      LAYER li1 ;
        RECT 718.615 1116.560 718.945 1117.040 ;
      LAYER li1 ;
        RECT 719.115 1116.390 719.285 1116.870 ;
      LAYER li1 ;
        RECT 719.455 1116.560 719.785 1117.040 ;
      LAYER li1 ;
        RECT 719.955 1116.390 720.125 1116.870 ;
      LAYER li1 ;
        RECT 720.295 1116.560 720.625 1117.040 ;
      LAYER li1 ;
        RECT 720.795 1116.390 720.965 1116.870 ;
      LAYER li1 ;
        RECT 721.135 1116.560 721.465 1117.040 ;
        RECT 721.635 1116.390 721.805 1116.865 ;
        RECT 721.975 1116.560 722.305 1117.040 ;
        RECT 722.475 1116.390 722.645 1116.870 ;
      LAYER li1 ;
        RECT 718.275 1116.220 720.965 1116.390 ;
      LAYER li1 ;
        RECT 721.225 1116.220 722.645 1116.390 ;
        RECT 722.905 1116.315 723.195 1117.040 ;
        RECT 723.755 1116.240 724.085 1117.040 ;
      LAYER li1 ;
        RECT 724.255 1116.390 724.425 1116.870 ;
      LAYER li1 ;
        RECT 724.595 1116.560 724.925 1117.040 ;
      LAYER li1 ;
        RECT 725.095 1116.390 725.265 1116.870 ;
      LAYER li1 ;
        RECT 725.435 1116.560 725.765 1117.040 ;
      LAYER li1 ;
        RECT 725.935 1116.390 726.105 1116.870 ;
      LAYER li1 ;
        RECT 726.275 1116.560 726.605 1117.040 ;
      LAYER li1 ;
        RECT 726.775 1116.390 726.945 1116.870 ;
      LAYER li1 ;
        RECT 727.115 1116.560 727.445 1117.040 ;
        RECT 727.615 1116.390 727.785 1116.865 ;
        RECT 727.955 1116.560 728.285 1117.040 ;
        RECT 728.455 1116.390 728.625 1116.870 ;
      LAYER li1 ;
        RECT 724.255 1116.220 726.945 1116.390 ;
      LAYER li1 ;
        RECT 727.205 1116.220 728.625 1116.390 ;
        RECT 728.885 1116.315 729.175 1117.040 ;
        RECT 729.735 1116.240 730.065 1117.040 ;
      LAYER li1 ;
        RECT 730.235 1116.390 730.405 1116.870 ;
      LAYER li1 ;
        RECT 730.575 1116.560 730.905 1117.040 ;
      LAYER li1 ;
        RECT 731.075 1116.390 731.245 1116.870 ;
      LAYER li1 ;
        RECT 731.415 1116.560 731.745 1117.040 ;
      LAYER li1 ;
        RECT 731.915 1116.390 732.085 1116.870 ;
      LAYER li1 ;
        RECT 732.255 1116.560 732.585 1117.040 ;
      LAYER li1 ;
        RECT 732.755 1116.390 732.925 1116.870 ;
      LAYER li1 ;
        RECT 733.095 1116.560 733.425 1117.040 ;
        RECT 733.595 1116.390 733.765 1116.865 ;
        RECT 733.935 1116.560 734.265 1117.040 ;
        RECT 734.435 1116.390 734.605 1116.870 ;
      LAYER li1 ;
        RECT 730.235 1116.220 732.925 1116.390 ;
      LAYER li1 ;
        RECT 733.185 1116.220 734.605 1116.390 ;
        RECT 734.865 1116.315 735.155 1117.040 ;
        RECT 735.715 1116.240 736.045 1117.040 ;
        RECT 736.555 1116.560 736.885 1117.040 ;
        RECT 737.395 1116.560 737.725 1117.040 ;
        RECT 738.235 1116.560 738.565 1117.040 ;
        RECT 739.075 1116.560 739.405 1117.040 ;
        RECT 739.575 1116.390 739.745 1116.865 ;
        RECT 739.915 1116.560 740.245 1117.040 ;
        RECT 740.415 1116.390 740.585 1116.870 ;
        RECT 739.165 1116.220 740.585 1116.390 ;
        RECT 740.845 1116.315 741.135 1117.040 ;
        RECT 741.695 1116.240 742.025 1117.040 ;
        RECT 742.535 1116.560 742.865 1117.040 ;
        RECT 743.375 1116.560 743.705 1117.040 ;
        RECT 744.215 1116.560 744.545 1117.040 ;
        RECT 745.055 1116.560 745.385 1117.040 ;
        RECT 745.555 1116.390 745.725 1116.865 ;
        RECT 745.895 1116.560 746.225 1117.040 ;
        RECT 746.395 1116.390 746.565 1116.870 ;
        RECT 745.145 1116.220 746.565 1116.390 ;
        RECT 746.825 1116.315 747.115 1117.040 ;
        RECT 747.675 1116.240 748.005 1117.040 ;
        RECT 748.515 1116.560 748.845 1117.040 ;
        RECT 749.355 1116.560 749.685 1117.040 ;
        RECT 750.195 1116.560 750.525 1117.040 ;
        RECT 751.035 1116.560 751.365 1117.040 ;
        RECT 751.535 1116.390 751.705 1116.865 ;
        RECT 751.875 1116.560 752.205 1117.040 ;
        RECT 752.375 1116.390 752.545 1116.870 ;
        RECT 751.125 1116.220 752.545 1116.390 ;
        RECT 752.805 1116.315 753.095 1117.040 ;
        RECT 753.655 1116.240 753.985 1117.040 ;
        RECT 754.495 1116.560 754.825 1117.040 ;
        RECT 755.335 1116.560 755.665 1117.040 ;
        RECT 756.175 1116.560 756.505 1117.040 ;
        RECT 757.015 1116.560 757.345 1117.040 ;
        RECT 757.515 1116.390 757.685 1116.865 ;
        RECT 757.855 1116.560 758.185 1117.040 ;
        RECT 758.355 1116.390 758.525 1116.870 ;
        RECT 757.105 1116.220 758.525 1116.390 ;
        RECT 758.785 1116.315 759.075 1117.040 ;
        RECT 759.635 1116.240 759.965 1117.040 ;
        RECT 760.475 1116.560 760.805 1117.040 ;
        RECT 761.315 1116.560 761.645 1117.040 ;
        RECT 762.155 1116.560 762.485 1117.040 ;
        RECT 762.995 1116.560 763.325 1117.040 ;
        RECT 763.495 1116.390 763.665 1116.865 ;
        RECT 763.835 1116.560 764.165 1117.040 ;
        RECT 764.335 1116.390 764.505 1116.870 ;
        RECT 763.085 1116.220 764.505 1116.390 ;
        RECT 764.765 1116.315 765.055 1117.040 ;
        RECT 765.615 1116.240 765.945 1117.040 ;
        RECT 766.455 1116.560 766.785 1117.040 ;
        RECT 767.295 1116.560 767.625 1117.040 ;
        RECT 768.135 1116.560 768.465 1117.040 ;
        RECT 768.975 1116.560 769.305 1117.040 ;
        RECT 769.475 1116.390 769.645 1116.865 ;
        RECT 769.815 1116.560 770.145 1117.040 ;
        RECT 770.315 1116.390 770.485 1116.870 ;
        RECT 769.065 1116.220 770.485 1116.390 ;
        RECT 770.745 1116.315 771.035 1117.040 ;
        RECT 1969.085 1116.315 1969.375 1117.040 ;
        RECT 1969.935 1116.240 1970.265 1117.040 ;
      LAYER li1 ;
        RECT 1970.435 1116.390 1970.605 1116.870 ;
      LAYER li1 ;
        RECT 1970.775 1116.560 1971.105 1117.040 ;
      LAYER li1 ;
        RECT 1971.275 1116.390 1971.445 1116.870 ;
      LAYER li1 ;
        RECT 1971.615 1116.560 1971.945 1117.040 ;
      LAYER li1 ;
        RECT 1972.115 1116.390 1972.285 1116.870 ;
      LAYER li1 ;
        RECT 1972.455 1116.560 1972.785 1117.040 ;
      LAYER li1 ;
        RECT 1972.955 1116.390 1973.125 1116.870 ;
      LAYER li1 ;
        RECT 1973.295 1116.560 1973.625 1117.040 ;
        RECT 1973.795 1116.390 1973.965 1116.865 ;
        RECT 1974.135 1116.560 1974.465 1117.040 ;
        RECT 1974.635 1116.390 1974.805 1116.870 ;
      LAYER li1 ;
        RECT 1970.435 1116.220 1973.125 1116.390 ;
      LAYER li1 ;
        RECT 1973.385 1116.220 1974.805 1116.390 ;
        RECT 1975.065 1116.315 1975.355 1117.040 ;
        RECT 1975.915 1116.240 1976.245 1117.040 ;
      LAYER li1 ;
        RECT 1976.415 1116.390 1976.585 1116.870 ;
      LAYER li1 ;
        RECT 1976.755 1116.560 1977.085 1117.040 ;
      LAYER li1 ;
        RECT 1977.255 1116.390 1977.425 1116.870 ;
      LAYER li1 ;
        RECT 1977.595 1116.560 1977.925 1117.040 ;
      LAYER li1 ;
        RECT 1978.095 1116.390 1978.265 1116.870 ;
      LAYER li1 ;
        RECT 1978.435 1116.560 1978.765 1117.040 ;
      LAYER li1 ;
        RECT 1978.935 1116.390 1979.105 1116.870 ;
      LAYER li1 ;
        RECT 1979.275 1116.560 1979.605 1117.040 ;
        RECT 1979.775 1116.390 1979.945 1116.865 ;
        RECT 1980.115 1116.560 1980.445 1117.040 ;
        RECT 1980.615 1116.390 1980.785 1116.870 ;
      LAYER li1 ;
        RECT 1976.415 1116.220 1979.105 1116.390 ;
      LAYER li1 ;
        RECT 1979.365 1116.220 1980.785 1116.390 ;
        RECT 1981.045 1116.315 1981.335 1117.040 ;
        RECT 1981.895 1116.240 1982.225 1117.040 ;
      LAYER li1 ;
        RECT 1982.395 1116.390 1982.565 1116.870 ;
      LAYER li1 ;
        RECT 1982.735 1116.560 1983.065 1117.040 ;
      LAYER li1 ;
        RECT 1983.235 1116.390 1983.405 1116.870 ;
      LAYER li1 ;
        RECT 1983.575 1116.560 1983.905 1117.040 ;
      LAYER li1 ;
        RECT 1984.075 1116.390 1984.245 1116.870 ;
      LAYER li1 ;
        RECT 1984.415 1116.560 1984.745 1117.040 ;
      LAYER li1 ;
        RECT 1984.915 1116.390 1985.085 1116.870 ;
      LAYER li1 ;
        RECT 1985.255 1116.560 1985.585 1117.040 ;
        RECT 1985.755 1116.390 1985.925 1116.865 ;
        RECT 1986.095 1116.560 1986.425 1117.040 ;
        RECT 1986.595 1116.390 1986.765 1116.870 ;
      LAYER li1 ;
        RECT 1982.395 1116.220 1985.085 1116.390 ;
      LAYER li1 ;
        RECT 1985.345 1116.220 1986.765 1116.390 ;
        RECT 1987.025 1116.315 1987.315 1117.040 ;
        RECT 1987.875 1116.240 1988.205 1117.040 ;
      LAYER li1 ;
        RECT 1988.375 1116.390 1988.545 1116.870 ;
      LAYER li1 ;
        RECT 1988.715 1116.560 1989.045 1117.040 ;
      LAYER li1 ;
        RECT 1989.215 1116.390 1989.385 1116.870 ;
      LAYER li1 ;
        RECT 1989.555 1116.560 1989.885 1117.040 ;
      LAYER li1 ;
        RECT 1990.055 1116.390 1990.225 1116.870 ;
      LAYER li1 ;
        RECT 1990.395 1116.560 1990.725 1117.040 ;
      LAYER li1 ;
        RECT 1990.895 1116.390 1991.065 1116.870 ;
      LAYER li1 ;
        RECT 1991.235 1116.560 1991.565 1117.040 ;
        RECT 1991.735 1116.390 1991.905 1116.865 ;
        RECT 1992.075 1116.560 1992.405 1117.040 ;
        RECT 1992.575 1116.390 1992.745 1116.870 ;
      LAYER li1 ;
        RECT 1988.375 1116.220 1991.065 1116.390 ;
      LAYER li1 ;
        RECT 1991.325 1116.220 1992.745 1116.390 ;
        RECT 1993.005 1116.315 1993.295 1117.040 ;
        RECT 1993.855 1116.240 1994.185 1117.040 ;
      LAYER li1 ;
        RECT 1994.355 1116.390 1994.525 1116.870 ;
      LAYER li1 ;
        RECT 1994.695 1116.560 1995.025 1117.040 ;
      LAYER li1 ;
        RECT 1995.195 1116.390 1995.365 1116.870 ;
      LAYER li1 ;
        RECT 1995.535 1116.560 1995.865 1117.040 ;
      LAYER li1 ;
        RECT 1996.035 1116.390 1996.205 1116.870 ;
      LAYER li1 ;
        RECT 1996.375 1116.560 1996.705 1117.040 ;
      LAYER li1 ;
        RECT 1996.875 1116.390 1997.045 1116.870 ;
      LAYER li1 ;
        RECT 1997.215 1116.560 1997.545 1117.040 ;
        RECT 1997.715 1116.390 1997.885 1116.865 ;
        RECT 1998.055 1116.560 1998.385 1117.040 ;
        RECT 1998.555 1116.390 1998.725 1116.870 ;
      LAYER li1 ;
        RECT 1994.355 1116.220 1997.045 1116.390 ;
      LAYER li1 ;
        RECT 1997.305 1116.220 1998.725 1116.390 ;
        RECT 1998.985 1116.315 1999.275 1117.040 ;
        RECT 1999.835 1116.240 2000.165 1117.040 ;
      LAYER li1 ;
        RECT 2000.335 1116.390 2000.505 1116.870 ;
      LAYER li1 ;
        RECT 2000.675 1116.560 2001.005 1117.040 ;
      LAYER li1 ;
        RECT 2001.175 1116.390 2001.345 1116.870 ;
      LAYER li1 ;
        RECT 2001.515 1116.560 2001.845 1117.040 ;
      LAYER li1 ;
        RECT 2002.015 1116.390 2002.185 1116.870 ;
      LAYER li1 ;
        RECT 2002.355 1116.560 2002.685 1117.040 ;
      LAYER li1 ;
        RECT 2002.855 1116.390 2003.025 1116.870 ;
      LAYER li1 ;
        RECT 2003.195 1116.560 2003.525 1117.040 ;
        RECT 2003.695 1116.390 2003.865 1116.865 ;
        RECT 2004.035 1116.560 2004.365 1117.040 ;
        RECT 2004.535 1116.390 2004.705 1116.870 ;
      LAYER li1 ;
        RECT 2000.335 1116.220 2003.025 1116.390 ;
      LAYER li1 ;
        RECT 2003.285 1116.220 2004.705 1116.390 ;
        RECT 2004.965 1116.315 2005.255 1117.040 ;
        RECT 2005.815 1116.240 2006.145 1117.040 ;
      LAYER li1 ;
        RECT 2006.315 1116.390 2006.485 1116.870 ;
      LAYER li1 ;
        RECT 2006.655 1116.560 2006.985 1117.040 ;
      LAYER li1 ;
        RECT 2007.155 1116.390 2007.325 1116.870 ;
      LAYER li1 ;
        RECT 2007.495 1116.560 2007.825 1117.040 ;
      LAYER li1 ;
        RECT 2007.995 1116.390 2008.165 1116.870 ;
      LAYER li1 ;
        RECT 2008.335 1116.560 2008.665 1117.040 ;
      LAYER li1 ;
        RECT 2008.835 1116.390 2009.005 1116.870 ;
      LAYER li1 ;
        RECT 2009.175 1116.560 2009.505 1117.040 ;
        RECT 2009.675 1116.390 2009.845 1116.865 ;
        RECT 2010.015 1116.560 2010.345 1117.040 ;
        RECT 2010.515 1116.390 2010.685 1116.870 ;
      LAYER li1 ;
        RECT 2006.315 1116.220 2009.005 1116.390 ;
      LAYER li1 ;
        RECT 2009.265 1116.220 2010.685 1116.390 ;
        RECT 2010.945 1116.315 2011.235 1117.040 ;
        RECT 2011.795 1116.240 2012.125 1117.040 ;
      LAYER li1 ;
        RECT 2012.295 1116.390 2012.465 1116.870 ;
      LAYER li1 ;
        RECT 2012.635 1116.560 2012.965 1117.040 ;
      LAYER li1 ;
        RECT 2013.135 1116.390 2013.305 1116.870 ;
      LAYER li1 ;
        RECT 2013.475 1116.560 2013.805 1117.040 ;
      LAYER li1 ;
        RECT 2013.975 1116.390 2014.145 1116.870 ;
      LAYER li1 ;
        RECT 2014.315 1116.560 2014.645 1117.040 ;
      LAYER li1 ;
        RECT 2014.815 1116.390 2014.985 1116.870 ;
      LAYER li1 ;
        RECT 2015.155 1116.560 2015.485 1117.040 ;
        RECT 2015.655 1116.390 2015.825 1116.865 ;
        RECT 2015.995 1116.560 2016.325 1117.040 ;
        RECT 2016.495 1116.390 2016.665 1116.870 ;
      LAYER li1 ;
        RECT 2012.295 1116.220 2014.985 1116.390 ;
      LAYER li1 ;
        RECT 2015.245 1116.220 2016.665 1116.390 ;
        RECT 2016.925 1116.315 2017.215 1117.040 ;
        RECT 2017.775 1116.240 2018.105 1117.040 ;
      LAYER li1 ;
        RECT 2018.275 1116.390 2018.445 1116.870 ;
      LAYER li1 ;
        RECT 2018.615 1116.560 2018.945 1117.040 ;
      LAYER li1 ;
        RECT 2019.115 1116.390 2019.285 1116.870 ;
      LAYER li1 ;
        RECT 2019.455 1116.560 2019.785 1117.040 ;
      LAYER li1 ;
        RECT 2019.955 1116.390 2020.125 1116.870 ;
      LAYER li1 ;
        RECT 2020.295 1116.560 2020.625 1117.040 ;
      LAYER li1 ;
        RECT 2020.795 1116.390 2020.965 1116.870 ;
      LAYER li1 ;
        RECT 2021.135 1116.560 2021.465 1117.040 ;
        RECT 2021.635 1116.390 2021.805 1116.865 ;
        RECT 2021.975 1116.560 2022.305 1117.040 ;
        RECT 2022.475 1116.390 2022.645 1116.870 ;
      LAYER li1 ;
        RECT 2018.275 1116.220 2020.965 1116.390 ;
      LAYER li1 ;
        RECT 2021.225 1116.220 2022.645 1116.390 ;
        RECT 2022.905 1116.315 2023.195 1117.040 ;
        RECT 2023.755 1116.240 2024.085 1117.040 ;
      LAYER li1 ;
        RECT 2024.255 1116.390 2024.425 1116.870 ;
      LAYER li1 ;
        RECT 2024.595 1116.560 2024.925 1117.040 ;
      LAYER li1 ;
        RECT 2025.095 1116.390 2025.265 1116.870 ;
      LAYER li1 ;
        RECT 2025.435 1116.560 2025.765 1117.040 ;
      LAYER li1 ;
        RECT 2025.935 1116.390 2026.105 1116.870 ;
      LAYER li1 ;
        RECT 2026.275 1116.560 2026.605 1117.040 ;
      LAYER li1 ;
        RECT 2026.775 1116.390 2026.945 1116.870 ;
      LAYER li1 ;
        RECT 2027.115 1116.560 2027.445 1117.040 ;
        RECT 2027.615 1116.390 2027.785 1116.865 ;
        RECT 2027.955 1116.560 2028.285 1117.040 ;
        RECT 2028.455 1116.390 2028.625 1116.870 ;
      LAYER li1 ;
        RECT 2024.255 1116.220 2026.945 1116.390 ;
      LAYER li1 ;
        RECT 2027.205 1116.220 2028.625 1116.390 ;
        RECT 2028.885 1116.315 2029.175 1117.040 ;
        RECT 2029.735 1116.240 2030.065 1117.040 ;
      LAYER li1 ;
        RECT 2030.235 1116.390 2030.405 1116.870 ;
      LAYER li1 ;
        RECT 2030.575 1116.560 2030.905 1117.040 ;
      LAYER li1 ;
        RECT 2031.075 1116.390 2031.245 1116.870 ;
      LAYER li1 ;
        RECT 2031.415 1116.560 2031.745 1117.040 ;
      LAYER li1 ;
        RECT 2031.915 1116.390 2032.085 1116.870 ;
      LAYER li1 ;
        RECT 2032.255 1116.560 2032.585 1117.040 ;
      LAYER li1 ;
        RECT 2032.755 1116.390 2032.925 1116.870 ;
      LAYER li1 ;
        RECT 2033.095 1116.560 2033.425 1117.040 ;
        RECT 2033.595 1116.390 2033.765 1116.865 ;
        RECT 2033.935 1116.560 2034.265 1117.040 ;
        RECT 2034.435 1116.390 2034.605 1116.870 ;
      LAYER li1 ;
        RECT 2030.235 1116.220 2032.925 1116.390 ;
      LAYER li1 ;
        RECT 2033.185 1116.220 2034.605 1116.390 ;
        RECT 2034.865 1116.315 2035.155 1117.040 ;
        RECT 2035.715 1116.240 2036.045 1117.040 ;
      LAYER li1 ;
        RECT 2036.215 1116.390 2036.385 1116.870 ;
      LAYER li1 ;
        RECT 2036.555 1116.560 2036.885 1117.040 ;
      LAYER li1 ;
        RECT 2037.055 1116.390 2037.225 1116.870 ;
      LAYER li1 ;
        RECT 2037.395 1116.560 2037.725 1117.040 ;
      LAYER li1 ;
        RECT 2037.895 1116.390 2038.065 1116.870 ;
      LAYER li1 ;
        RECT 2038.235 1116.560 2038.565 1117.040 ;
      LAYER li1 ;
        RECT 2038.735 1116.390 2038.905 1116.870 ;
      LAYER li1 ;
        RECT 2039.075 1116.560 2039.405 1117.040 ;
        RECT 2039.575 1116.390 2039.745 1116.865 ;
        RECT 2039.915 1116.560 2040.245 1117.040 ;
        RECT 2040.415 1116.390 2040.585 1116.870 ;
      LAYER li1 ;
        RECT 2036.215 1116.220 2038.905 1116.390 ;
      LAYER li1 ;
        RECT 2039.165 1116.220 2040.585 1116.390 ;
        RECT 2040.845 1116.315 2041.135 1117.040 ;
        RECT 2041.695 1116.240 2042.025 1117.040 ;
      LAYER li1 ;
        RECT 2042.195 1116.390 2042.365 1116.870 ;
      LAYER li1 ;
        RECT 2042.535 1116.560 2042.865 1117.040 ;
      LAYER li1 ;
        RECT 2043.035 1116.390 2043.205 1116.870 ;
      LAYER li1 ;
        RECT 2043.375 1116.560 2043.705 1117.040 ;
      LAYER li1 ;
        RECT 2043.875 1116.390 2044.045 1116.870 ;
      LAYER li1 ;
        RECT 2044.215 1116.560 2044.545 1117.040 ;
      LAYER li1 ;
        RECT 2044.715 1116.390 2044.885 1116.870 ;
      LAYER li1 ;
        RECT 2045.055 1116.560 2045.385 1117.040 ;
        RECT 2045.555 1116.390 2045.725 1116.865 ;
        RECT 2045.895 1116.560 2046.225 1117.040 ;
        RECT 2046.395 1116.390 2046.565 1116.870 ;
      LAYER li1 ;
        RECT 2042.195 1116.220 2044.885 1116.390 ;
      LAYER li1 ;
        RECT 2045.145 1116.220 2046.565 1116.390 ;
        RECT 2046.825 1116.315 2047.115 1117.040 ;
        RECT 2047.675 1116.240 2048.005 1117.040 ;
      LAYER li1 ;
        RECT 2048.175 1116.390 2048.345 1116.870 ;
      LAYER li1 ;
        RECT 2048.515 1116.560 2048.845 1117.040 ;
      LAYER li1 ;
        RECT 2049.015 1116.390 2049.185 1116.870 ;
      LAYER li1 ;
        RECT 2049.355 1116.560 2049.685 1117.040 ;
      LAYER li1 ;
        RECT 2049.855 1116.390 2050.025 1116.870 ;
      LAYER li1 ;
        RECT 2050.195 1116.560 2050.525 1117.040 ;
      LAYER li1 ;
        RECT 2050.695 1116.390 2050.865 1116.870 ;
      LAYER li1 ;
        RECT 2051.035 1116.560 2051.365 1117.040 ;
        RECT 2051.535 1116.390 2051.705 1116.865 ;
        RECT 2051.875 1116.560 2052.205 1117.040 ;
        RECT 2052.375 1116.390 2052.545 1116.870 ;
      LAYER li1 ;
        RECT 2048.175 1116.220 2050.865 1116.390 ;
      LAYER li1 ;
        RECT 2051.125 1116.220 2052.545 1116.390 ;
        RECT 2052.805 1116.315 2053.095 1117.040 ;
        RECT 2053.655 1116.240 2053.985 1117.040 ;
      LAYER li1 ;
        RECT 2054.155 1116.390 2054.325 1116.870 ;
      LAYER li1 ;
        RECT 2054.495 1116.560 2054.825 1117.040 ;
      LAYER li1 ;
        RECT 2054.995 1116.390 2055.165 1116.870 ;
      LAYER li1 ;
        RECT 2055.335 1116.560 2055.665 1117.040 ;
      LAYER li1 ;
        RECT 2055.835 1116.390 2056.005 1116.870 ;
      LAYER li1 ;
        RECT 2056.175 1116.560 2056.505 1117.040 ;
      LAYER li1 ;
        RECT 2056.675 1116.390 2056.845 1116.870 ;
      LAYER li1 ;
        RECT 2057.015 1116.560 2057.345 1117.040 ;
        RECT 2057.515 1116.390 2057.685 1116.865 ;
        RECT 2057.855 1116.560 2058.185 1117.040 ;
        RECT 2058.355 1116.390 2058.525 1116.870 ;
      LAYER li1 ;
        RECT 2054.155 1116.220 2056.845 1116.390 ;
      LAYER li1 ;
        RECT 2057.105 1116.220 2058.525 1116.390 ;
        RECT 2058.785 1116.315 2059.075 1117.040 ;
        RECT 2059.635 1116.240 2059.965 1117.040 ;
      LAYER li1 ;
        RECT 2060.135 1116.390 2060.305 1116.870 ;
      LAYER li1 ;
        RECT 2060.475 1116.560 2060.805 1117.040 ;
      LAYER li1 ;
        RECT 2060.975 1116.390 2061.145 1116.870 ;
      LAYER li1 ;
        RECT 2061.315 1116.560 2061.645 1117.040 ;
      LAYER li1 ;
        RECT 2061.815 1116.390 2061.985 1116.870 ;
      LAYER li1 ;
        RECT 2062.155 1116.560 2062.485 1117.040 ;
      LAYER li1 ;
        RECT 2062.655 1116.390 2062.825 1116.870 ;
      LAYER li1 ;
        RECT 2062.995 1116.560 2063.325 1117.040 ;
        RECT 2063.495 1116.390 2063.665 1116.865 ;
        RECT 2063.835 1116.560 2064.165 1117.040 ;
        RECT 2064.335 1116.390 2064.505 1116.870 ;
      LAYER li1 ;
        RECT 2060.135 1116.220 2062.825 1116.390 ;
      LAYER li1 ;
        RECT 2063.085 1116.220 2064.505 1116.390 ;
        RECT 2064.765 1116.315 2065.055 1117.040 ;
        RECT 2065.615 1116.240 2065.945 1117.040 ;
      LAYER li1 ;
        RECT 2066.115 1116.390 2066.285 1116.870 ;
      LAYER li1 ;
        RECT 2066.455 1116.560 2066.785 1117.040 ;
      LAYER li1 ;
        RECT 2066.955 1116.390 2067.125 1116.870 ;
      LAYER li1 ;
        RECT 2067.295 1116.560 2067.625 1117.040 ;
      LAYER li1 ;
        RECT 2067.795 1116.390 2067.965 1116.870 ;
      LAYER li1 ;
        RECT 2068.135 1116.560 2068.465 1117.040 ;
      LAYER li1 ;
        RECT 2068.635 1116.390 2068.805 1116.870 ;
      LAYER li1 ;
        RECT 2068.975 1116.560 2069.305 1117.040 ;
        RECT 2069.475 1116.390 2069.645 1116.865 ;
        RECT 2069.815 1116.560 2070.145 1117.040 ;
        RECT 2070.315 1116.390 2070.485 1116.870 ;
      LAYER li1 ;
        RECT 2066.115 1116.220 2068.805 1116.390 ;
      LAYER li1 ;
        RECT 2069.065 1116.220 2070.485 1116.390 ;
        RECT 2070.745 1116.315 2071.035 1117.040 ;
      LAYER li1 ;
        RECT 670.435 1115.680 670.690 1116.220 ;
      LAYER li1 ;
        RECT 673.385 1116.050 673.560 1116.220 ;
        RECT 670.935 1115.880 673.560 1116.050 ;
        RECT 673.385 1115.680 673.560 1115.880 ;
      LAYER li1 ;
        RECT 673.740 1115.850 675.330 1116.050 ;
        RECT 676.415 1115.680 676.670 1116.220 ;
      LAYER li1 ;
        RECT 679.365 1116.050 679.540 1116.220 ;
        RECT 676.915 1115.880 679.540 1116.050 ;
        RECT 679.365 1115.680 679.540 1115.880 ;
      LAYER li1 ;
        RECT 679.720 1115.850 681.310 1116.050 ;
        RECT 682.395 1115.680 682.650 1116.220 ;
      LAYER li1 ;
        RECT 685.345 1116.050 685.520 1116.220 ;
        RECT 682.895 1115.880 685.520 1116.050 ;
        RECT 685.345 1115.680 685.520 1115.880 ;
      LAYER li1 ;
        RECT 685.700 1115.850 687.290 1116.050 ;
        RECT 688.375 1115.680 688.630 1116.220 ;
      LAYER li1 ;
        RECT 691.325 1116.050 691.500 1116.220 ;
        RECT 688.875 1115.880 691.500 1116.050 ;
        RECT 691.325 1115.680 691.500 1115.880 ;
      LAYER li1 ;
        RECT 691.680 1115.850 693.270 1116.050 ;
        RECT 694.355 1115.680 694.610 1116.220 ;
      LAYER li1 ;
        RECT 697.305 1116.050 697.480 1116.220 ;
        RECT 694.855 1115.880 697.480 1116.050 ;
        RECT 697.305 1115.680 697.480 1115.880 ;
      LAYER li1 ;
        RECT 697.660 1115.850 699.250 1116.050 ;
        RECT 700.335 1115.680 700.590 1116.220 ;
      LAYER li1 ;
        RECT 703.285 1116.050 703.460 1116.220 ;
        RECT 700.835 1115.880 703.460 1116.050 ;
        RECT 703.285 1115.680 703.460 1115.880 ;
      LAYER li1 ;
        RECT 703.640 1115.850 705.230 1116.050 ;
        RECT 706.315 1115.680 706.570 1116.220 ;
      LAYER li1 ;
        RECT 709.265 1116.050 709.440 1116.220 ;
        RECT 706.815 1115.880 709.440 1116.050 ;
        RECT 709.265 1115.680 709.440 1115.880 ;
      LAYER li1 ;
        RECT 709.620 1115.850 711.210 1116.050 ;
        RECT 712.295 1115.680 712.550 1116.220 ;
      LAYER li1 ;
        RECT 715.245 1116.050 715.420 1116.220 ;
        RECT 712.795 1115.880 715.420 1116.050 ;
        RECT 715.245 1115.680 715.420 1115.880 ;
      LAYER li1 ;
        RECT 715.600 1115.850 717.190 1116.050 ;
        RECT 718.275 1115.680 718.530 1116.220 ;
      LAYER li1 ;
        RECT 721.225 1116.050 721.400 1116.220 ;
        RECT 718.775 1115.880 721.400 1116.050 ;
        RECT 721.225 1115.680 721.400 1115.880 ;
      LAYER li1 ;
        RECT 721.580 1115.850 723.170 1116.050 ;
        RECT 724.255 1115.680 724.510 1116.220 ;
      LAYER li1 ;
        RECT 727.205 1116.050 727.380 1116.220 ;
        RECT 724.755 1115.880 727.380 1116.050 ;
        RECT 727.205 1115.680 727.380 1115.880 ;
      LAYER li1 ;
        RECT 727.560 1115.850 729.150 1116.050 ;
        RECT 730.235 1115.680 730.490 1116.220 ;
      LAYER li1 ;
        RECT 733.185 1116.050 733.360 1116.220 ;
        RECT 739.165 1116.050 739.340 1116.220 ;
        RECT 745.145 1116.050 745.320 1116.220 ;
        RECT 751.125 1116.050 751.300 1116.220 ;
        RECT 757.105 1116.050 757.280 1116.220 ;
        RECT 763.085 1116.050 763.260 1116.220 ;
        RECT 769.065 1116.050 769.240 1116.220 ;
        RECT 730.735 1115.880 733.360 1116.050 ;
        RECT 733.185 1115.680 733.360 1115.880 ;
      LAYER li1 ;
        RECT 733.540 1115.850 734.640 1116.050 ;
      LAYER li1 ;
        RECT 736.715 1115.880 739.340 1116.050 ;
        RECT 739.165 1115.680 739.340 1115.880 ;
      LAYER li1 ;
        RECT 739.520 1115.850 741.110 1116.050 ;
      LAYER li1 ;
        RECT 742.695 1115.880 745.320 1116.050 ;
        RECT 745.145 1115.680 745.320 1115.880 ;
      LAYER li1 ;
        RECT 745.500 1115.850 747.090 1116.050 ;
      LAYER li1 ;
        RECT 748.675 1115.880 751.300 1116.050 ;
        RECT 751.125 1115.680 751.300 1115.880 ;
      LAYER li1 ;
        RECT 751.480 1115.850 753.070 1116.050 ;
      LAYER li1 ;
        RECT 754.655 1115.880 757.280 1116.050 ;
        RECT 757.105 1115.680 757.280 1115.880 ;
      LAYER li1 ;
        RECT 757.460 1115.850 759.050 1116.050 ;
      LAYER li1 ;
        RECT 760.635 1115.880 763.260 1116.050 ;
        RECT 763.085 1115.680 763.260 1115.880 ;
      LAYER li1 ;
        RECT 763.440 1115.850 765.030 1116.050 ;
      LAYER li1 ;
        RECT 766.615 1115.880 769.240 1116.050 ;
        RECT 769.065 1115.680 769.240 1115.880 ;
      LAYER li1 ;
        RECT 769.420 1115.850 771.010 1116.050 ;
        RECT 1970.435 1115.680 1970.690 1116.220 ;
      LAYER li1 ;
        RECT 1973.385 1116.050 1973.560 1116.220 ;
        RECT 1970.935 1115.880 1973.560 1116.050 ;
        RECT 1973.385 1115.680 1973.560 1115.880 ;
      LAYER li1 ;
        RECT 1976.415 1115.680 1976.670 1116.220 ;
      LAYER li1 ;
        RECT 1979.365 1116.050 1979.540 1116.220 ;
        RECT 1976.915 1115.880 1979.540 1116.050 ;
        RECT 1979.365 1115.680 1979.540 1115.880 ;
      LAYER li1 ;
        RECT 1982.395 1115.680 1982.650 1116.220 ;
      LAYER li1 ;
        RECT 1985.345 1116.050 1985.520 1116.220 ;
        RECT 1982.895 1115.880 1985.520 1116.050 ;
        RECT 1985.345 1115.680 1985.520 1115.880 ;
      LAYER li1 ;
        RECT 1988.375 1115.680 1988.630 1116.220 ;
      LAYER li1 ;
        RECT 1991.325 1116.050 1991.500 1116.220 ;
        RECT 1988.875 1115.880 1991.500 1116.050 ;
        RECT 1991.325 1115.680 1991.500 1115.880 ;
      LAYER li1 ;
        RECT 1994.355 1115.680 1994.610 1116.220 ;
      LAYER li1 ;
        RECT 1997.305 1116.050 1997.480 1116.220 ;
        RECT 1994.855 1115.880 1997.480 1116.050 ;
        RECT 1997.305 1115.680 1997.480 1115.880 ;
      LAYER li1 ;
        RECT 2000.335 1115.680 2000.590 1116.220 ;
      LAYER li1 ;
        RECT 2003.285 1116.050 2003.460 1116.220 ;
        RECT 2000.835 1115.880 2003.460 1116.050 ;
        RECT 2003.285 1115.680 2003.460 1115.880 ;
      LAYER li1 ;
        RECT 2006.315 1115.680 2006.570 1116.220 ;
      LAYER li1 ;
        RECT 2009.265 1116.050 2009.440 1116.220 ;
        RECT 2006.815 1115.880 2009.440 1116.050 ;
        RECT 2009.265 1115.680 2009.440 1115.880 ;
      LAYER li1 ;
        RECT 2012.295 1115.680 2012.550 1116.220 ;
      LAYER li1 ;
        RECT 2015.245 1116.050 2015.420 1116.220 ;
        RECT 2012.795 1115.880 2015.420 1116.050 ;
        RECT 2015.245 1115.680 2015.420 1115.880 ;
      LAYER li1 ;
        RECT 2018.275 1115.680 2018.530 1116.220 ;
      LAYER li1 ;
        RECT 2021.225 1116.050 2021.400 1116.220 ;
        RECT 2018.775 1115.880 2021.400 1116.050 ;
        RECT 2021.225 1115.680 2021.400 1115.880 ;
      LAYER li1 ;
        RECT 2024.255 1115.680 2024.510 1116.220 ;
      LAYER li1 ;
        RECT 2027.205 1116.050 2027.380 1116.220 ;
        RECT 2024.755 1115.880 2027.380 1116.050 ;
        RECT 2027.205 1115.680 2027.380 1115.880 ;
      LAYER li1 ;
        RECT 2030.235 1115.680 2030.490 1116.220 ;
      LAYER li1 ;
        RECT 2033.185 1116.050 2033.360 1116.220 ;
        RECT 2030.735 1115.880 2033.360 1116.050 ;
        RECT 2033.185 1115.680 2033.360 1115.880 ;
      LAYER li1 ;
        RECT 2033.540 1115.850 2034.640 1116.050 ;
        RECT 2036.215 1115.680 2036.470 1116.220 ;
      LAYER li1 ;
        RECT 2039.165 1116.050 2039.340 1116.220 ;
        RECT 2036.715 1115.880 2039.340 1116.050 ;
        RECT 2039.165 1115.680 2039.340 1115.880 ;
      LAYER li1 ;
        RECT 2042.195 1115.680 2042.450 1116.220 ;
      LAYER li1 ;
        RECT 2045.145 1116.050 2045.320 1116.220 ;
        RECT 2042.695 1115.880 2045.320 1116.050 ;
        RECT 2045.145 1115.680 2045.320 1115.880 ;
      LAYER li1 ;
        RECT 2048.175 1115.680 2048.430 1116.220 ;
      LAYER li1 ;
        RECT 2051.125 1116.050 2051.300 1116.220 ;
        RECT 2048.675 1115.880 2051.300 1116.050 ;
        RECT 2051.125 1115.680 2051.300 1115.880 ;
      LAYER li1 ;
        RECT 2054.155 1115.680 2054.410 1116.220 ;
      LAYER li1 ;
        RECT 2057.105 1116.050 2057.280 1116.220 ;
        RECT 2054.655 1115.880 2057.280 1116.050 ;
        RECT 2057.105 1115.680 2057.280 1115.880 ;
      LAYER li1 ;
        RECT 2060.135 1115.680 2060.390 1116.220 ;
      LAYER li1 ;
        RECT 2063.085 1116.050 2063.260 1116.220 ;
        RECT 2060.635 1115.880 2063.260 1116.050 ;
        RECT 2063.085 1115.680 2063.260 1115.880 ;
      LAYER li1 ;
        RECT 2066.115 1115.680 2066.370 1116.220 ;
      LAYER li1 ;
        RECT 2069.065 1116.050 2069.240 1116.220 ;
        RECT 2066.615 1115.880 2069.240 1116.050 ;
        RECT 2069.065 1115.680 2069.240 1115.880 ;
        RECT 669.085 1114.490 669.375 1115.655 ;
        RECT 669.935 1114.490 670.265 1115.640 ;
      LAYER li1 ;
        RECT 670.435 1115.510 673.125 1115.680 ;
      LAYER li1 ;
        RECT 673.385 1115.510 674.885 1115.680 ;
      LAYER li1 ;
        RECT 670.435 1114.660 670.605 1115.510 ;
      LAYER li1 ;
        RECT 670.775 1114.490 671.105 1115.290 ;
      LAYER li1 ;
        RECT 671.275 1114.660 671.445 1115.510 ;
      LAYER li1 ;
        RECT 671.615 1114.490 671.945 1115.290 ;
      LAYER li1 ;
        RECT 672.115 1114.660 672.285 1115.510 ;
      LAYER li1 ;
        RECT 672.455 1114.490 672.785 1115.290 ;
      LAYER li1 ;
        RECT 672.955 1114.660 673.125 1115.510 ;
      LAYER li1 ;
        RECT 673.375 1114.490 673.545 1115.290 ;
        RECT 673.715 1114.660 674.045 1115.510 ;
        RECT 674.215 1114.490 674.385 1115.290 ;
        RECT 674.555 1114.660 674.885 1115.510 ;
        RECT 675.065 1114.490 675.355 1115.655 ;
        RECT 675.915 1114.490 676.245 1115.640 ;
      LAYER li1 ;
        RECT 676.415 1115.510 679.105 1115.680 ;
      LAYER li1 ;
        RECT 679.365 1115.510 680.865 1115.680 ;
      LAYER li1 ;
        RECT 676.415 1114.660 676.585 1115.510 ;
      LAYER li1 ;
        RECT 676.755 1114.490 677.085 1115.290 ;
      LAYER li1 ;
        RECT 677.255 1114.660 677.425 1115.510 ;
      LAYER li1 ;
        RECT 677.595 1114.490 677.925 1115.290 ;
      LAYER li1 ;
        RECT 678.095 1114.660 678.265 1115.510 ;
      LAYER li1 ;
        RECT 678.435 1114.490 678.765 1115.290 ;
      LAYER li1 ;
        RECT 678.935 1114.660 679.105 1115.510 ;
      LAYER li1 ;
        RECT 679.355 1114.490 679.525 1115.290 ;
        RECT 679.695 1114.660 680.025 1115.510 ;
        RECT 680.195 1114.490 680.365 1115.290 ;
        RECT 680.535 1114.660 680.865 1115.510 ;
        RECT 681.045 1114.490 681.335 1115.655 ;
        RECT 681.895 1114.490 682.225 1115.640 ;
      LAYER li1 ;
        RECT 682.395 1115.510 685.085 1115.680 ;
      LAYER li1 ;
        RECT 685.345 1115.510 686.845 1115.680 ;
      LAYER li1 ;
        RECT 682.395 1114.660 682.565 1115.510 ;
      LAYER li1 ;
        RECT 682.735 1114.490 683.065 1115.290 ;
      LAYER li1 ;
        RECT 683.235 1114.660 683.405 1115.510 ;
      LAYER li1 ;
        RECT 683.575 1114.490 683.905 1115.290 ;
      LAYER li1 ;
        RECT 684.075 1114.660 684.245 1115.510 ;
      LAYER li1 ;
        RECT 684.415 1114.490 684.745 1115.290 ;
      LAYER li1 ;
        RECT 684.915 1114.660 685.085 1115.510 ;
      LAYER li1 ;
        RECT 685.335 1114.490 685.505 1115.290 ;
        RECT 685.675 1114.660 686.005 1115.510 ;
        RECT 686.175 1114.490 686.345 1115.290 ;
        RECT 686.515 1114.660 686.845 1115.510 ;
        RECT 687.025 1114.490 687.315 1115.655 ;
        RECT 687.875 1114.490 688.205 1115.640 ;
      LAYER li1 ;
        RECT 688.375 1115.510 691.065 1115.680 ;
      LAYER li1 ;
        RECT 691.325 1115.510 692.825 1115.680 ;
      LAYER li1 ;
        RECT 688.375 1114.660 688.545 1115.510 ;
      LAYER li1 ;
        RECT 688.715 1114.490 689.045 1115.290 ;
      LAYER li1 ;
        RECT 689.215 1114.660 689.385 1115.510 ;
      LAYER li1 ;
        RECT 689.555 1114.490 689.885 1115.290 ;
      LAYER li1 ;
        RECT 690.055 1114.660 690.225 1115.510 ;
      LAYER li1 ;
        RECT 690.395 1114.490 690.725 1115.290 ;
      LAYER li1 ;
        RECT 690.895 1114.660 691.065 1115.510 ;
      LAYER li1 ;
        RECT 691.315 1114.490 691.485 1115.290 ;
        RECT 691.655 1114.660 691.985 1115.510 ;
        RECT 692.155 1114.490 692.325 1115.290 ;
        RECT 692.495 1114.660 692.825 1115.510 ;
        RECT 693.005 1114.490 693.295 1115.655 ;
        RECT 693.855 1114.490 694.185 1115.640 ;
      LAYER li1 ;
        RECT 694.355 1115.510 697.045 1115.680 ;
      LAYER li1 ;
        RECT 697.305 1115.510 698.805 1115.680 ;
      LAYER li1 ;
        RECT 694.355 1114.660 694.525 1115.510 ;
      LAYER li1 ;
        RECT 694.695 1114.490 695.025 1115.290 ;
      LAYER li1 ;
        RECT 695.195 1114.660 695.365 1115.510 ;
      LAYER li1 ;
        RECT 695.535 1114.490 695.865 1115.290 ;
      LAYER li1 ;
        RECT 696.035 1114.660 696.205 1115.510 ;
      LAYER li1 ;
        RECT 696.375 1114.490 696.705 1115.290 ;
      LAYER li1 ;
        RECT 696.875 1114.660 697.045 1115.510 ;
      LAYER li1 ;
        RECT 697.295 1114.490 697.465 1115.290 ;
        RECT 697.635 1114.660 697.965 1115.510 ;
        RECT 698.135 1114.490 698.305 1115.290 ;
        RECT 698.475 1114.660 698.805 1115.510 ;
        RECT 698.985 1114.490 699.275 1115.655 ;
        RECT 699.835 1114.490 700.165 1115.640 ;
      LAYER li1 ;
        RECT 700.335 1115.510 703.025 1115.680 ;
      LAYER li1 ;
        RECT 703.285 1115.510 704.785 1115.680 ;
      LAYER li1 ;
        RECT 700.335 1114.660 700.505 1115.510 ;
      LAYER li1 ;
        RECT 700.675 1114.490 701.005 1115.290 ;
      LAYER li1 ;
        RECT 701.175 1114.660 701.345 1115.510 ;
      LAYER li1 ;
        RECT 701.515 1114.490 701.845 1115.290 ;
      LAYER li1 ;
        RECT 702.015 1114.660 702.185 1115.510 ;
      LAYER li1 ;
        RECT 702.355 1114.490 702.685 1115.290 ;
      LAYER li1 ;
        RECT 702.855 1114.660 703.025 1115.510 ;
      LAYER li1 ;
        RECT 703.275 1114.490 703.445 1115.290 ;
        RECT 703.615 1114.660 703.945 1115.510 ;
        RECT 704.115 1114.490 704.285 1115.290 ;
        RECT 704.455 1114.660 704.785 1115.510 ;
        RECT 704.965 1114.490 705.255 1115.655 ;
        RECT 705.815 1114.490 706.145 1115.640 ;
      LAYER li1 ;
        RECT 706.315 1115.510 709.005 1115.680 ;
      LAYER li1 ;
        RECT 709.265 1115.510 710.765 1115.680 ;
      LAYER li1 ;
        RECT 706.315 1114.660 706.485 1115.510 ;
      LAYER li1 ;
        RECT 706.655 1114.490 706.985 1115.290 ;
      LAYER li1 ;
        RECT 707.155 1114.660 707.325 1115.510 ;
      LAYER li1 ;
        RECT 707.495 1114.490 707.825 1115.290 ;
      LAYER li1 ;
        RECT 707.995 1114.660 708.165 1115.510 ;
      LAYER li1 ;
        RECT 708.335 1114.490 708.665 1115.290 ;
      LAYER li1 ;
        RECT 708.835 1114.660 709.005 1115.510 ;
      LAYER li1 ;
        RECT 709.255 1114.490 709.425 1115.290 ;
        RECT 709.595 1114.660 709.925 1115.510 ;
        RECT 710.095 1114.490 710.265 1115.290 ;
        RECT 710.435 1114.660 710.765 1115.510 ;
        RECT 710.945 1114.490 711.235 1115.655 ;
        RECT 711.795 1114.490 712.125 1115.640 ;
      LAYER li1 ;
        RECT 712.295 1115.510 714.985 1115.680 ;
      LAYER li1 ;
        RECT 715.245 1115.510 716.745 1115.680 ;
      LAYER li1 ;
        RECT 712.295 1114.660 712.465 1115.510 ;
      LAYER li1 ;
        RECT 712.635 1114.490 712.965 1115.290 ;
      LAYER li1 ;
        RECT 713.135 1114.660 713.305 1115.510 ;
      LAYER li1 ;
        RECT 713.475 1114.490 713.805 1115.290 ;
      LAYER li1 ;
        RECT 713.975 1114.660 714.145 1115.510 ;
      LAYER li1 ;
        RECT 714.315 1114.490 714.645 1115.290 ;
      LAYER li1 ;
        RECT 714.815 1114.660 714.985 1115.510 ;
      LAYER li1 ;
        RECT 715.235 1114.490 715.405 1115.290 ;
        RECT 715.575 1114.660 715.905 1115.510 ;
        RECT 716.075 1114.490 716.245 1115.290 ;
        RECT 716.415 1114.660 716.745 1115.510 ;
        RECT 716.925 1114.490 717.215 1115.655 ;
        RECT 717.775 1114.490 718.105 1115.640 ;
      LAYER li1 ;
        RECT 718.275 1115.510 720.965 1115.680 ;
      LAYER li1 ;
        RECT 721.225 1115.510 722.725 1115.680 ;
      LAYER li1 ;
        RECT 718.275 1114.660 718.445 1115.510 ;
      LAYER li1 ;
        RECT 718.615 1114.490 718.945 1115.290 ;
      LAYER li1 ;
        RECT 719.115 1114.660 719.285 1115.510 ;
      LAYER li1 ;
        RECT 719.455 1114.490 719.785 1115.290 ;
      LAYER li1 ;
        RECT 719.955 1114.660 720.125 1115.510 ;
      LAYER li1 ;
        RECT 720.295 1114.490 720.625 1115.290 ;
      LAYER li1 ;
        RECT 720.795 1114.660 720.965 1115.510 ;
      LAYER li1 ;
        RECT 721.215 1114.490 721.385 1115.290 ;
        RECT 721.555 1114.660 721.885 1115.510 ;
        RECT 722.055 1114.490 722.225 1115.290 ;
        RECT 722.395 1114.660 722.725 1115.510 ;
        RECT 722.905 1114.490 723.195 1115.655 ;
        RECT 723.755 1114.490 724.085 1115.640 ;
      LAYER li1 ;
        RECT 724.255 1115.510 726.945 1115.680 ;
      LAYER li1 ;
        RECT 727.205 1115.510 728.705 1115.680 ;
      LAYER li1 ;
        RECT 724.255 1114.660 724.425 1115.510 ;
      LAYER li1 ;
        RECT 724.595 1114.490 724.925 1115.290 ;
      LAYER li1 ;
        RECT 725.095 1114.660 725.265 1115.510 ;
      LAYER li1 ;
        RECT 725.435 1114.490 725.765 1115.290 ;
      LAYER li1 ;
        RECT 725.935 1114.660 726.105 1115.510 ;
      LAYER li1 ;
        RECT 726.275 1114.490 726.605 1115.290 ;
      LAYER li1 ;
        RECT 726.775 1114.660 726.945 1115.510 ;
      LAYER li1 ;
        RECT 727.195 1114.490 727.365 1115.290 ;
        RECT 727.535 1114.660 727.865 1115.510 ;
        RECT 728.035 1114.490 728.205 1115.290 ;
        RECT 728.375 1114.660 728.705 1115.510 ;
        RECT 728.885 1114.490 729.175 1115.655 ;
        RECT 729.735 1114.490 730.065 1115.640 ;
      LAYER li1 ;
        RECT 730.235 1115.510 732.925 1115.680 ;
      LAYER li1 ;
        RECT 733.185 1115.510 734.685 1115.680 ;
      LAYER li1 ;
        RECT 730.235 1114.660 730.405 1115.510 ;
      LAYER li1 ;
        RECT 730.575 1114.490 730.905 1115.290 ;
      LAYER li1 ;
        RECT 731.075 1114.660 731.245 1115.510 ;
      LAYER li1 ;
        RECT 731.415 1114.490 731.745 1115.290 ;
      LAYER li1 ;
        RECT 731.915 1114.660 732.085 1115.510 ;
      LAYER li1 ;
        RECT 732.255 1114.490 732.585 1115.290 ;
      LAYER li1 ;
        RECT 732.755 1114.660 732.925 1115.510 ;
      LAYER li1 ;
        RECT 733.175 1114.490 733.345 1115.290 ;
        RECT 733.515 1114.660 733.845 1115.510 ;
        RECT 734.015 1114.490 734.185 1115.290 ;
        RECT 734.355 1114.660 734.685 1115.510 ;
        RECT 734.865 1114.490 735.155 1115.655 ;
        RECT 735.715 1114.490 736.045 1115.640 ;
        RECT 739.165 1115.510 740.665 1115.680 ;
        RECT 736.555 1114.490 736.885 1115.290 ;
        RECT 737.395 1114.490 737.725 1115.290 ;
        RECT 738.235 1114.490 738.565 1115.290 ;
        RECT 739.155 1114.490 739.325 1115.290 ;
        RECT 739.495 1114.660 739.825 1115.510 ;
        RECT 739.995 1114.490 740.165 1115.290 ;
        RECT 740.335 1114.660 740.665 1115.510 ;
        RECT 740.845 1114.490 741.135 1115.655 ;
        RECT 741.695 1114.490 742.025 1115.640 ;
        RECT 745.145 1115.510 746.645 1115.680 ;
        RECT 742.535 1114.490 742.865 1115.290 ;
        RECT 743.375 1114.490 743.705 1115.290 ;
        RECT 744.215 1114.490 744.545 1115.290 ;
        RECT 745.135 1114.490 745.305 1115.290 ;
        RECT 745.475 1114.660 745.805 1115.510 ;
        RECT 745.975 1114.490 746.145 1115.290 ;
        RECT 746.315 1114.660 746.645 1115.510 ;
        RECT 746.825 1114.490 747.115 1115.655 ;
        RECT 747.675 1114.490 748.005 1115.640 ;
        RECT 751.125 1115.510 752.625 1115.680 ;
        RECT 748.515 1114.490 748.845 1115.290 ;
        RECT 749.355 1114.490 749.685 1115.290 ;
        RECT 750.195 1114.490 750.525 1115.290 ;
        RECT 751.115 1114.490 751.285 1115.290 ;
        RECT 751.455 1114.660 751.785 1115.510 ;
        RECT 751.955 1114.490 752.125 1115.290 ;
        RECT 752.295 1114.660 752.625 1115.510 ;
        RECT 752.805 1114.490 753.095 1115.655 ;
        RECT 753.655 1114.490 753.985 1115.640 ;
        RECT 757.105 1115.510 758.605 1115.680 ;
        RECT 754.495 1114.490 754.825 1115.290 ;
        RECT 755.335 1114.490 755.665 1115.290 ;
        RECT 756.175 1114.490 756.505 1115.290 ;
        RECT 757.095 1114.490 757.265 1115.290 ;
        RECT 757.435 1114.660 757.765 1115.510 ;
        RECT 757.935 1114.490 758.105 1115.290 ;
        RECT 758.275 1114.660 758.605 1115.510 ;
        RECT 758.785 1114.490 759.075 1115.655 ;
        RECT 759.635 1114.490 759.965 1115.640 ;
        RECT 763.085 1115.510 764.585 1115.680 ;
        RECT 760.475 1114.490 760.805 1115.290 ;
        RECT 761.315 1114.490 761.645 1115.290 ;
        RECT 762.155 1114.490 762.485 1115.290 ;
        RECT 763.075 1114.490 763.245 1115.290 ;
        RECT 763.415 1114.660 763.745 1115.510 ;
        RECT 763.915 1114.490 764.085 1115.290 ;
        RECT 764.255 1114.660 764.585 1115.510 ;
        RECT 764.765 1114.490 765.055 1115.655 ;
        RECT 765.615 1114.490 765.945 1115.640 ;
        RECT 769.065 1115.510 770.565 1115.680 ;
        RECT 766.455 1114.490 766.785 1115.290 ;
        RECT 767.295 1114.490 767.625 1115.290 ;
        RECT 768.135 1114.490 768.465 1115.290 ;
        RECT 769.055 1114.490 769.225 1115.290 ;
        RECT 769.395 1114.660 769.725 1115.510 ;
        RECT 769.895 1114.490 770.065 1115.290 ;
        RECT 770.235 1114.660 770.565 1115.510 ;
        RECT 770.745 1114.490 771.035 1115.655 ;
        RECT 1969.085 1114.490 1969.375 1115.655 ;
        RECT 1969.935 1114.490 1970.265 1115.640 ;
      LAYER li1 ;
        RECT 1970.435 1115.510 1973.125 1115.680 ;
      LAYER li1 ;
        RECT 1973.385 1115.510 1974.885 1115.680 ;
      LAYER li1 ;
        RECT 1970.435 1114.660 1970.605 1115.510 ;
      LAYER li1 ;
        RECT 1970.775 1114.490 1971.105 1115.290 ;
      LAYER li1 ;
        RECT 1971.275 1114.660 1971.445 1115.510 ;
      LAYER li1 ;
        RECT 1971.615 1114.490 1971.945 1115.290 ;
      LAYER li1 ;
        RECT 1972.115 1114.660 1972.285 1115.510 ;
      LAYER li1 ;
        RECT 1972.455 1114.490 1972.785 1115.290 ;
      LAYER li1 ;
        RECT 1972.955 1114.660 1973.125 1115.510 ;
      LAYER li1 ;
        RECT 1973.375 1114.490 1973.545 1115.290 ;
        RECT 1973.715 1114.660 1974.045 1115.510 ;
        RECT 1974.215 1114.490 1974.385 1115.290 ;
        RECT 1974.555 1114.660 1974.885 1115.510 ;
        RECT 1975.065 1114.490 1975.355 1115.655 ;
        RECT 1975.915 1114.490 1976.245 1115.640 ;
      LAYER li1 ;
        RECT 1976.415 1115.510 1979.105 1115.680 ;
      LAYER li1 ;
        RECT 1979.365 1115.510 1980.865 1115.680 ;
      LAYER li1 ;
        RECT 1976.415 1114.660 1976.585 1115.510 ;
      LAYER li1 ;
        RECT 1976.755 1114.490 1977.085 1115.290 ;
      LAYER li1 ;
        RECT 1977.255 1114.660 1977.425 1115.510 ;
      LAYER li1 ;
        RECT 1977.595 1114.490 1977.925 1115.290 ;
      LAYER li1 ;
        RECT 1978.095 1114.660 1978.265 1115.510 ;
      LAYER li1 ;
        RECT 1978.435 1114.490 1978.765 1115.290 ;
      LAYER li1 ;
        RECT 1978.935 1114.660 1979.105 1115.510 ;
      LAYER li1 ;
        RECT 1979.355 1114.490 1979.525 1115.290 ;
        RECT 1979.695 1114.660 1980.025 1115.510 ;
        RECT 1980.195 1114.490 1980.365 1115.290 ;
        RECT 1980.535 1114.660 1980.865 1115.510 ;
        RECT 1981.045 1114.490 1981.335 1115.655 ;
        RECT 1981.895 1114.490 1982.225 1115.640 ;
      LAYER li1 ;
        RECT 1982.395 1115.510 1985.085 1115.680 ;
      LAYER li1 ;
        RECT 1985.345 1115.510 1986.845 1115.680 ;
      LAYER li1 ;
        RECT 1982.395 1114.660 1982.565 1115.510 ;
      LAYER li1 ;
        RECT 1982.735 1114.490 1983.065 1115.290 ;
      LAYER li1 ;
        RECT 1983.235 1114.660 1983.405 1115.510 ;
      LAYER li1 ;
        RECT 1983.575 1114.490 1983.905 1115.290 ;
      LAYER li1 ;
        RECT 1984.075 1114.660 1984.245 1115.510 ;
      LAYER li1 ;
        RECT 1984.415 1114.490 1984.745 1115.290 ;
      LAYER li1 ;
        RECT 1984.915 1114.660 1985.085 1115.510 ;
      LAYER li1 ;
        RECT 1985.335 1114.490 1985.505 1115.290 ;
        RECT 1985.675 1114.660 1986.005 1115.510 ;
        RECT 1986.175 1114.490 1986.345 1115.290 ;
        RECT 1986.515 1114.660 1986.845 1115.510 ;
        RECT 1987.025 1114.490 1987.315 1115.655 ;
        RECT 1987.875 1114.490 1988.205 1115.640 ;
      LAYER li1 ;
        RECT 1988.375 1115.510 1991.065 1115.680 ;
      LAYER li1 ;
        RECT 1991.325 1115.510 1992.825 1115.680 ;
      LAYER li1 ;
        RECT 1988.375 1114.660 1988.545 1115.510 ;
      LAYER li1 ;
        RECT 1988.715 1114.490 1989.045 1115.290 ;
      LAYER li1 ;
        RECT 1989.215 1114.660 1989.385 1115.510 ;
      LAYER li1 ;
        RECT 1989.555 1114.490 1989.885 1115.290 ;
      LAYER li1 ;
        RECT 1990.055 1114.660 1990.225 1115.510 ;
      LAYER li1 ;
        RECT 1990.395 1114.490 1990.725 1115.290 ;
      LAYER li1 ;
        RECT 1990.895 1114.660 1991.065 1115.510 ;
      LAYER li1 ;
        RECT 1991.315 1114.490 1991.485 1115.290 ;
        RECT 1991.655 1114.660 1991.985 1115.510 ;
        RECT 1992.155 1114.490 1992.325 1115.290 ;
        RECT 1992.495 1114.660 1992.825 1115.510 ;
        RECT 1993.005 1114.490 1993.295 1115.655 ;
        RECT 1993.855 1114.490 1994.185 1115.640 ;
      LAYER li1 ;
        RECT 1994.355 1115.510 1997.045 1115.680 ;
      LAYER li1 ;
        RECT 1997.305 1115.510 1998.805 1115.680 ;
      LAYER li1 ;
        RECT 1994.355 1114.660 1994.525 1115.510 ;
      LAYER li1 ;
        RECT 1994.695 1114.490 1995.025 1115.290 ;
      LAYER li1 ;
        RECT 1995.195 1114.660 1995.365 1115.510 ;
      LAYER li1 ;
        RECT 1995.535 1114.490 1995.865 1115.290 ;
      LAYER li1 ;
        RECT 1996.035 1114.660 1996.205 1115.510 ;
      LAYER li1 ;
        RECT 1996.375 1114.490 1996.705 1115.290 ;
      LAYER li1 ;
        RECT 1996.875 1114.660 1997.045 1115.510 ;
      LAYER li1 ;
        RECT 1997.295 1114.490 1997.465 1115.290 ;
        RECT 1997.635 1114.660 1997.965 1115.510 ;
        RECT 1998.135 1114.490 1998.305 1115.290 ;
        RECT 1998.475 1114.660 1998.805 1115.510 ;
        RECT 1998.985 1114.490 1999.275 1115.655 ;
        RECT 1999.835 1114.490 2000.165 1115.640 ;
      LAYER li1 ;
        RECT 2000.335 1115.510 2003.025 1115.680 ;
      LAYER li1 ;
        RECT 2003.285 1115.510 2004.785 1115.680 ;
      LAYER li1 ;
        RECT 2000.335 1114.660 2000.505 1115.510 ;
      LAYER li1 ;
        RECT 2000.675 1114.490 2001.005 1115.290 ;
      LAYER li1 ;
        RECT 2001.175 1114.660 2001.345 1115.510 ;
      LAYER li1 ;
        RECT 2001.515 1114.490 2001.845 1115.290 ;
      LAYER li1 ;
        RECT 2002.015 1114.660 2002.185 1115.510 ;
      LAYER li1 ;
        RECT 2002.355 1114.490 2002.685 1115.290 ;
      LAYER li1 ;
        RECT 2002.855 1114.660 2003.025 1115.510 ;
      LAYER li1 ;
        RECT 2003.275 1114.490 2003.445 1115.290 ;
        RECT 2003.615 1114.660 2003.945 1115.510 ;
        RECT 2004.115 1114.490 2004.285 1115.290 ;
        RECT 2004.455 1114.660 2004.785 1115.510 ;
        RECT 2004.965 1114.490 2005.255 1115.655 ;
        RECT 2005.815 1114.490 2006.145 1115.640 ;
      LAYER li1 ;
        RECT 2006.315 1115.510 2009.005 1115.680 ;
      LAYER li1 ;
        RECT 2009.265 1115.510 2010.765 1115.680 ;
      LAYER li1 ;
        RECT 2006.315 1114.660 2006.485 1115.510 ;
      LAYER li1 ;
        RECT 2006.655 1114.490 2006.985 1115.290 ;
      LAYER li1 ;
        RECT 2007.155 1114.660 2007.325 1115.510 ;
      LAYER li1 ;
        RECT 2007.495 1114.490 2007.825 1115.290 ;
      LAYER li1 ;
        RECT 2007.995 1114.660 2008.165 1115.510 ;
      LAYER li1 ;
        RECT 2008.335 1114.490 2008.665 1115.290 ;
      LAYER li1 ;
        RECT 2008.835 1114.660 2009.005 1115.510 ;
      LAYER li1 ;
        RECT 2009.255 1114.490 2009.425 1115.290 ;
        RECT 2009.595 1114.660 2009.925 1115.510 ;
        RECT 2010.095 1114.490 2010.265 1115.290 ;
        RECT 2010.435 1114.660 2010.765 1115.510 ;
        RECT 2010.945 1114.490 2011.235 1115.655 ;
        RECT 2011.795 1114.490 2012.125 1115.640 ;
      LAYER li1 ;
        RECT 2012.295 1115.510 2014.985 1115.680 ;
      LAYER li1 ;
        RECT 2015.245 1115.510 2016.745 1115.680 ;
      LAYER li1 ;
        RECT 2012.295 1114.660 2012.465 1115.510 ;
      LAYER li1 ;
        RECT 2012.635 1114.490 2012.965 1115.290 ;
      LAYER li1 ;
        RECT 2013.135 1114.660 2013.305 1115.510 ;
      LAYER li1 ;
        RECT 2013.475 1114.490 2013.805 1115.290 ;
      LAYER li1 ;
        RECT 2013.975 1114.660 2014.145 1115.510 ;
      LAYER li1 ;
        RECT 2014.315 1114.490 2014.645 1115.290 ;
      LAYER li1 ;
        RECT 2014.815 1114.660 2014.985 1115.510 ;
      LAYER li1 ;
        RECT 2015.235 1114.490 2015.405 1115.290 ;
        RECT 2015.575 1114.660 2015.905 1115.510 ;
        RECT 2016.075 1114.490 2016.245 1115.290 ;
        RECT 2016.415 1114.660 2016.745 1115.510 ;
        RECT 2016.925 1114.490 2017.215 1115.655 ;
        RECT 2017.775 1114.490 2018.105 1115.640 ;
      LAYER li1 ;
        RECT 2018.275 1115.510 2020.965 1115.680 ;
      LAYER li1 ;
        RECT 2021.225 1115.510 2022.725 1115.680 ;
      LAYER li1 ;
        RECT 2018.275 1114.660 2018.445 1115.510 ;
      LAYER li1 ;
        RECT 2018.615 1114.490 2018.945 1115.290 ;
      LAYER li1 ;
        RECT 2019.115 1114.660 2019.285 1115.510 ;
      LAYER li1 ;
        RECT 2019.455 1114.490 2019.785 1115.290 ;
      LAYER li1 ;
        RECT 2019.955 1114.660 2020.125 1115.510 ;
      LAYER li1 ;
        RECT 2020.295 1114.490 2020.625 1115.290 ;
      LAYER li1 ;
        RECT 2020.795 1114.660 2020.965 1115.510 ;
      LAYER li1 ;
        RECT 2021.215 1114.490 2021.385 1115.290 ;
        RECT 2021.555 1114.660 2021.885 1115.510 ;
        RECT 2022.055 1114.490 2022.225 1115.290 ;
        RECT 2022.395 1114.660 2022.725 1115.510 ;
        RECT 2022.905 1114.490 2023.195 1115.655 ;
        RECT 2023.755 1114.490 2024.085 1115.640 ;
      LAYER li1 ;
        RECT 2024.255 1115.510 2026.945 1115.680 ;
      LAYER li1 ;
        RECT 2027.205 1115.510 2028.705 1115.680 ;
      LAYER li1 ;
        RECT 2024.255 1114.660 2024.425 1115.510 ;
      LAYER li1 ;
        RECT 2024.595 1114.490 2024.925 1115.290 ;
      LAYER li1 ;
        RECT 2025.095 1114.660 2025.265 1115.510 ;
      LAYER li1 ;
        RECT 2025.435 1114.490 2025.765 1115.290 ;
      LAYER li1 ;
        RECT 2025.935 1114.660 2026.105 1115.510 ;
      LAYER li1 ;
        RECT 2026.275 1114.490 2026.605 1115.290 ;
      LAYER li1 ;
        RECT 2026.775 1114.660 2026.945 1115.510 ;
      LAYER li1 ;
        RECT 2027.195 1114.490 2027.365 1115.290 ;
        RECT 2027.535 1114.660 2027.865 1115.510 ;
        RECT 2028.035 1114.490 2028.205 1115.290 ;
        RECT 2028.375 1114.660 2028.705 1115.510 ;
        RECT 2028.885 1114.490 2029.175 1115.655 ;
        RECT 2029.735 1114.490 2030.065 1115.640 ;
      LAYER li1 ;
        RECT 2030.235 1115.510 2032.925 1115.680 ;
      LAYER li1 ;
        RECT 2033.185 1115.510 2034.685 1115.680 ;
      LAYER li1 ;
        RECT 2030.235 1114.660 2030.405 1115.510 ;
      LAYER li1 ;
        RECT 2030.575 1114.490 2030.905 1115.290 ;
      LAYER li1 ;
        RECT 2031.075 1114.660 2031.245 1115.510 ;
      LAYER li1 ;
        RECT 2031.415 1114.490 2031.745 1115.290 ;
      LAYER li1 ;
        RECT 2031.915 1114.660 2032.085 1115.510 ;
      LAYER li1 ;
        RECT 2032.255 1114.490 2032.585 1115.290 ;
      LAYER li1 ;
        RECT 2032.755 1114.660 2032.925 1115.510 ;
      LAYER li1 ;
        RECT 2033.175 1114.490 2033.345 1115.290 ;
        RECT 2033.515 1114.660 2033.845 1115.510 ;
        RECT 2034.015 1114.490 2034.185 1115.290 ;
        RECT 2034.355 1114.660 2034.685 1115.510 ;
        RECT 2034.865 1114.490 2035.155 1115.655 ;
        RECT 2035.715 1114.490 2036.045 1115.640 ;
      LAYER li1 ;
        RECT 2036.215 1115.510 2038.905 1115.680 ;
      LAYER li1 ;
        RECT 2039.165 1115.510 2040.665 1115.680 ;
      LAYER li1 ;
        RECT 2036.215 1114.660 2036.385 1115.510 ;
      LAYER li1 ;
        RECT 2036.555 1114.490 2036.885 1115.290 ;
      LAYER li1 ;
        RECT 2037.055 1114.660 2037.225 1115.510 ;
      LAYER li1 ;
        RECT 2037.395 1114.490 2037.725 1115.290 ;
      LAYER li1 ;
        RECT 2037.895 1114.660 2038.065 1115.510 ;
      LAYER li1 ;
        RECT 2038.235 1114.490 2038.565 1115.290 ;
      LAYER li1 ;
        RECT 2038.735 1114.660 2038.905 1115.510 ;
      LAYER li1 ;
        RECT 2039.155 1114.490 2039.325 1115.290 ;
        RECT 2039.495 1114.660 2039.825 1115.510 ;
        RECT 2039.995 1114.490 2040.165 1115.290 ;
        RECT 2040.335 1114.660 2040.665 1115.510 ;
        RECT 2040.845 1114.490 2041.135 1115.655 ;
        RECT 2041.695 1114.490 2042.025 1115.640 ;
      LAYER li1 ;
        RECT 2042.195 1115.510 2044.885 1115.680 ;
      LAYER li1 ;
        RECT 2045.145 1115.510 2046.645 1115.680 ;
      LAYER li1 ;
        RECT 2042.195 1114.660 2042.365 1115.510 ;
      LAYER li1 ;
        RECT 2042.535 1114.490 2042.865 1115.290 ;
      LAYER li1 ;
        RECT 2043.035 1114.660 2043.205 1115.510 ;
      LAYER li1 ;
        RECT 2043.375 1114.490 2043.705 1115.290 ;
      LAYER li1 ;
        RECT 2043.875 1114.660 2044.045 1115.510 ;
      LAYER li1 ;
        RECT 2044.215 1114.490 2044.545 1115.290 ;
      LAYER li1 ;
        RECT 2044.715 1114.660 2044.885 1115.510 ;
      LAYER li1 ;
        RECT 2045.135 1114.490 2045.305 1115.290 ;
        RECT 2045.475 1114.660 2045.805 1115.510 ;
        RECT 2045.975 1114.490 2046.145 1115.290 ;
        RECT 2046.315 1114.660 2046.645 1115.510 ;
        RECT 2046.825 1114.490 2047.115 1115.655 ;
        RECT 2047.675 1114.490 2048.005 1115.640 ;
      LAYER li1 ;
        RECT 2048.175 1115.510 2050.865 1115.680 ;
      LAYER li1 ;
        RECT 2051.125 1115.510 2052.625 1115.680 ;
      LAYER li1 ;
        RECT 2048.175 1114.660 2048.345 1115.510 ;
      LAYER li1 ;
        RECT 2048.515 1114.490 2048.845 1115.290 ;
      LAYER li1 ;
        RECT 2049.015 1114.660 2049.185 1115.510 ;
      LAYER li1 ;
        RECT 2049.355 1114.490 2049.685 1115.290 ;
      LAYER li1 ;
        RECT 2049.855 1114.660 2050.025 1115.510 ;
      LAYER li1 ;
        RECT 2050.195 1114.490 2050.525 1115.290 ;
      LAYER li1 ;
        RECT 2050.695 1114.660 2050.865 1115.510 ;
      LAYER li1 ;
        RECT 2051.115 1114.490 2051.285 1115.290 ;
        RECT 2051.455 1114.660 2051.785 1115.510 ;
        RECT 2051.955 1114.490 2052.125 1115.290 ;
        RECT 2052.295 1114.660 2052.625 1115.510 ;
        RECT 2052.805 1114.490 2053.095 1115.655 ;
        RECT 2053.655 1114.490 2053.985 1115.640 ;
      LAYER li1 ;
        RECT 2054.155 1115.510 2056.845 1115.680 ;
      LAYER li1 ;
        RECT 2057.105 1115.510 2058.605 1115.680 ;
      LAYER li1 ;
        RECT 2054.155 1114.660 2054.325 1115.510 ;
      LAYER li1 ;
        RECT 2054.495 1114.490 2054.825 1115.290 ;
      LAYER li1 ;
        RECT 2054.995 1114.660 2055.165 1115.510 ;
      LAYER li1 ;
        RECT 2055.335 1114.490 2055.665 1115.290 ;
      LAYER li1 ;
        RECT 2055.835 1114.660 2056.005 1115.510 ;
      LAYER li1 ;
        RECT 2056.175 1114.490 2056.505 1115.290 ;
      LAYER li1 ;
        RECT 2056.675 1114.660 2056.845 1115.510 ;
      LAYER li1 ;
        RECT 2057.095 1114.490 2057.265 1115.290 ;
        RECT 2057.435 1114.660 2057.765 1115.510 ;
        RECT 2057.935 1114.490 2058.105 1115.290 ;
        RECT 2058.275 1114.660 2058.605 1115.510 ;
        RECT 2058.785 1114.490 2059.075 1115.655 ;
        RECT 2059.635 1114.490 2059.965 1115.640 ;
      LAYER li1 ;
        RECT 2060.135 1115.510 2062.825 1115.680 ;
      LAYER li1 ;
        RECT 2063.085 1115.510 2064.585 1115.680 ;
      LAYER li1 ;
        RECT 2060.135 1114.660 2060.305 1115.510 ;
      LAYER li1 ;
        RECT 2060.475 1114.490 2060.805 1115.290 ;
      LAYER li1 ;
        RECT 2060.975 1114.660 2061.145 1115.510 ;
      LAYER li1 ;
        RECT 2061.315 1114.490 2061.645 1115.290 ;
      LAYER li1 ;
        RECT 2061.815 1114.660 2061.985 1115.510 ;
      LAYER li1 ;
        RECT 2062.155 1114.490 2062.485 1115.290 ;
      LAYER li1 ;
        RECT 2062.655 1114.660 2062.825 1115.510 ;
      LAYER li1 ;
        RECT 2063.075 1114.490 2063.245 1115.290 ;
        RECT 2063.415 1114.660 2063.745 1115.510 ;
        RECT 2063.915 1114.490 2064.085 1115.290 ;
        RECT 2064.255 1114.660 2064.585 1115.510 ;
        RECT 2064.765 1114.490 2065.055 1115.655 ;
        RECT 2065.615 1114.490 2065.945 1115.640 ;
      LAYER li1 ;
        RECT 2066.115 1115.510 2068.805 1115.680 ;
      LAYER li1 ;
        RECT 2069.065 1115.510 2070.565 1115.680 ;
      LAYER li1 ;
        RECT 2066.115 1114.660 2066.285 1115.510 ;
      LAYER li1 ;
        RECT 2066.455 1114.490 2066.785 1115.290 ;
      LAYER li1 ;
        RECT 2066.955 1114.660 2067.125 1115.510 ;
      LAYER li1 ;
        RECT 2067.295 1114.490 2067.625 1115.290 ;
      LAYER li1 ;
        RECT 2067.795 1114.660 2067.965 1115.510 ;
      LAYER li1 ;
        RECT 2068.135 1114.490 2068.465 1115.290 ;
      LAYER li1 ;
        RECT 2068.635 1114.660 2068.805 1115.510 ;
      LAYER li1 ;
        RECT 2069.055 1114.490 2069.225 1115.290 ;
        RECT 2069.395 1114.660 2069.725 1115.510 ;
        RECT 2069.895 1114.490 2070.065 1115.290 ;
        RECT 2070.235 1114.660 2070.565 1115.510 ;
        RECT 2070.745 1114.490 2071.035 1115.655 ;
        RECT 669.000 1114.320 669.145 1114.490 ;
        RECT 669.315 1114.320 669.605 1114.490 ;
        RECT 669.775 1114.320 670.065 1114.490 ;
        RECT 670.235 1114.320 670.525 1114.490 ;
        RECT 670.695 1114.320 670.985 1114.490 ;
        RECT 671.155 1114.320 671.445 1114.490 ;
        RECT 671.615 1114.320 671.905 1114.490 ;
        RECT 672.075 1114.320 672.365 1114.490 ;
        RECT 672.535 1114.320 672.825 1114.490 ;
        RECT 672.995 1114.320 673.285 1114.490 ;
        RECT 673.455 1114.320 673.745 1114.490 ;
        RECT 673.915 1114.320 674.205 1114.490 ;
        RECT 674.375 1114.320 674.665 1114.490 ;
        RECT 674.835 1114.320 675.125 1114.490 ;
        RECT 675.295 1114.320 675.585 1114.490 ;
        RECT 675.755 1114.320 676.045 1114.490 ;
        RECT 676.215 1114.320 676.505 1114.490 ;
        RECT 676.675 1114.320 676.965 1114.490 ;
        RECT 677.135 1114.320 677.425 1114.490 ;
        RECT 677.595 1114.320 677.885 1114.490 ;
        RECT 678.055 1114.320 678.345 1114.490 ;
        RECT 678.515 1114.320 678.805 1114.490 ;
        RECT 678.975 1114.320 679.265 1114.490 ;
        RECT 679.435 1114.320 679.725 1114.490 ;
        RECT 679.895 1114.320 680.185 1114.490 ;
        RECT 680.355 1114.320 680.645 1114.490 ;
        RECT 680.815 1114.320 681.105 1114.490 ;
        RECT 681.275 1114.320 681.565 1114.490 ;
        RECT 681.735 1114.320 682.025 1114.490 ;
        RECT 682.195 1114.320 682.485 1114.490 ;
        RECT 682.655 1114.320 682.945 1114.490 ;
        RECT 683.115 1114.320 683.405 1114.490 ;
        RECT 683.575 1114.320 683.865 1114.490 ;
        RECT 684.035 1114.320 684.325 1114.490 ;
        RECT 684.495 1114.320 684.785 1114.490 ;
        RECT 684.955 1114.320 685.245 1114.490 ;
        RECT 685.415 1114.320 685.705 1114.490 ;
        RECT 685.875 1114.320 686.165 1114.490 ;
        RECT 686.335 1114.320 686.625 1114.490 ;
        RECT 686.795 1114.320 687.085 1114.490 ;
        RECT 687.255 1114.320 687.545 1114.490 ;
        RECT 687.715 1114.320 688.005 1114.490 ;
        RECT 688.175 1114.320 688.465 1114.490 ;
        RECT 688.635 1114.320 688.925 1114.490 ;
        RECT 689.095 1114.320 689.385 1114.490 ;
        RECT 689.555 1114.320 689.845 1114.490 ;
        RECT 690.015 1114.320 690.305 1114.490 ;
        RECT 690.475 1114.320 690.765 1114.490 ;
        RECT 690.935 1114.320 691.225 1114.490 ;
        RECT 691.395 1114.320 691.685 1114.490 ;
        RECT 691.855 1114.320 692.145 1114.490 ;
        RECT 692.315 1114.320 692.605 1114.490 ;
        RECT 692.775 1114.320 693.065 1114.490 ;
        RECT 693.235 1114.320 693.525 1114.490 ;
        RECT 693.695 1114.320 693.985 1114.490 ;
        RECT 694.155 1114.320 694.445 1114.490 ;
        RECT 694.615 1114.320 694.905 1114.490 ;
        RECT 695.075 1114.320 695.365 1114.490 ;
        RECT 695.535 1114.320 695.825 1114.490 ;
        RECT 695.995 1114.320 696.285 1114.490 ;
        RECT 696.455 1114.320 696.745 1114.490 ;
        RECT 696.915 1114.320 697.205 1114.490 ;
        RECT 697.375 1114.320 697.665 1114.490 ;
        RECT 697.835 1114.320 698.125 1114.490 ;
        RECT 698.295 1114.320 698.585 1114.490 ;
        RECT 698.755 1114.320 699.045 1114.490 ;
        RECT 699.215 1114.320 699.505 1114.490 ;
        RECT 699.675 1114.320 699.965 1114.490 ;
        RECT 700.135 1114.320 700.425 1114.490 ;
        RECT 700.595 1114.320 700.885 1114.490 ;
        RECT 701.055 1114.320 701.345 1114.490 ;
        RECT 701.515 1114.320 701.805 1114.490 ;
        RECT 701.975 1114.320 702.265 1114.490 ;
        RECT 702.435 1114.320 702.725 1114.490 ;
        RECT 702.895 1114.320 703.185 1114.490 ;
        RECT 703.355 1114.320 703.645 1114.490 ;
        RECT 703.815 1114.320 704.105 1114.490 ;
        RECT 704.275 1114.320 704.565 1114.490 ;
        RECT 704.735 1114.320 705.025 1114.490 ;
        RECT 705.195 1114.320 705.485 1114.490 ;
        RECT 705.655 1114.320 705.945 1114.490 ;
        RECT 706.115 1114.320 706.405 1114.490 ;
        RECT 706.575 1114.320 706.865 1114.490 ;
        RECT 707.035 1114.320 707.325 1114.490 ;
        RECT 707.495 1114.320 707.785 1114.490 ;
        RECT 707.955 1114.320 708.245 1114.490 ;
        RECT 708.415 1114.320 708.705 1114.490 ;
        RECT 708.875 1114.320 709.165 1114.490 ;
        RECT 709.335 1114.320 709.625 1114.490 ;
        RECT 709.795 1114.320 710.085 1114.490 ;
        RECT 710.255 1114.320 710.545 1114.490 ;
        RECT 710.715 1114.320 711.005 1114.490 ;
        RECT 711.175 1114.320 711.465 1114.490 ;
        RECT 711.635 1114.320 711.925 1114.490 ;
        RECT 712.095 1114.320 712.385 1114.490 ;
        RECT 712.555 1114.320 712.845 1114.490 ;
        RECT 713.015 1114.320 713.305 1114.490 ;
        RECT 713.475 1114.320 713.765 1114.490 ;
        RECT 713.935 1114.320 714.225 1114.490 ;
        RECT 714.395 1114.320 714.685 1114.490 ;
        RECT 714.855 1114.320 715.145 1114.490 ;
        RECT 715.315 1114.320 715.605 1114.490 ;
        RECT 715.775 1114.320 716.065 1114.490 ;
        RECT 716.235 1114.320 716.525 1114.490 ;
        RECT 716.695 1114.320 716.985 1114.490 ;
        RECT 717.155 1114.320 717.445 1114.490 ;
        RECT 717.615 1114.320 717.905 1114.490 ;
        RECT 718.075 1114.320 718.365 1114.490 ;
        RECT 718.535 1114.320 718.825 1114.490 ;
        RECT 718.995 1114.320 719.285 1114.490 ;
        RECT 719.455 1114.320 719.745 1114.490 ;
        RECT 719.915 1114.320 720.205 1114.490 ;
        RECT 720.375 1114.320 720.665 1114.490 ;
        RECT 720.835 1114.320 721.125 1114.490 ;
        RECT 721.295 1114.320 721.585 1114.490 ;
        RECT 721.755 1114.320 722.045 1114.490 ;
        RECT 722.215 1114.320 722.505 1114.490 ;
        RECT 722.675 1114.320 722.965 1114.490 ;
        RECT 723.135 1114.320 723.425 1114.490 ;
        RECT 723.595 1114.320 723.885 1114.490 ;
        RECT 724.055 1114.320 724.345 1114.490 ;
        RECT 724.515 1114.320 724.805 1114.490 ;
        RECT 724.975 1114.320 725.265 1114.490 ;
        RECT 725.435 1114.320 725.725 1114.490 ;
        RECT 725.895 1114.320 726.185 1114.490 ;
        RECT 726.355 1114.320 726.645 1114.490 ;
        RECT 726.815 1114.320 727.105 1114.490 ;
        RECT 727.275 1114.320 727.565 1114.490 ;
        RECT 727.735 1114.320 728.025 1114.490 ;
        RECT 728.195 1114.320 728.485 1114.490 ;
        RECT 728.655 1114.320 728.945 1114.490 ;
        RECT 729.115 1114.320 729.405 1114.490 ;
        RECT 729.575 1114.320 729.865 1114.490 ;
        RECT 730.035 1114.320 730.325 1114.490 ;
        RECT 730.495 1114.320 730.785 1114.490 ;
        RECT 730.955 1114.320 731.245 1114.490 ;
        RECT 731.415 1114.320 731.705 1114.490 ;
        RECT 731.875 1114.320 732.165 1114.490 ;
        RECT 732.335 1114.320 732.625 1114.490 ;
        RECT 732.795 1114.320 733.085 1114.490 ;
        RECT 733.255 1114.320 733.545 1114.490 ;
        RECT 733.715 1114.320 734.005 1114.490 ;
        RECT 734.175 1114.320 734.465 1114.490 ;
        RECT 734.635 1114.320 734.925 1114.490 ;
        RECT 735.095 1114.320 735.385 1114.490 ;
        RECT 735.555 1114.320 735.845 1114.490 ;
        RECT 736.015 1114.320 736.305 1114.490 ;
        RECT 736.475 1114.320 736.765 1114.490 ;
        RECT 736.935 1114.320 737.225 1114.490 ;
        RECT 737.395 1114.320 737.685 1114.490 ;
        RECT 737.855 1114.320 738.145 1114.490 ;
        RECT 738.315 1114.320 738.605 1114.490 ;
        RECT 738.775 1114.320 739.065 1114.490 ;
        RECT 739.235 1114.320 739.525 1114.490 ;
        RECT 739.695 1114.320 739.985 1114.490 ;
        RECT 740.155 1114.320 740.445 1114.490 ;
        RECT 740.615 1114.320 740.905 1114.490 ;
        RECT 741.075 1114.320 741.365 1114.490 ;
        RECT 741.535 1114.320 741.825 1114.490 ;
        RECT 741.995 1114.320 742.285 1114.490 ;
        RECT 742.455 1114.320 742.745 1114.490 ;
        RECT 742.915 1114.320 743.205 1114.490 ;
        RECT 743.375 1114.320 743.665 1114.490 ;
        RECT 743.835 1114.320 744.125 1114.490 ;
        RECT 744.295 1114.320 744.585 1114.490 ;
        RECT 744.755 1114.320 745.045 1114.490 ;
        RECT 745.215 1114.320 745.505 1114.490 ;
        RECT 745.675 1114.320 745.965 1114.490 ;
        RECT 746.135 1114.320 746.425 1114.490 ;
        RECT 746.595 1114.320 746.885 1114.490 ;
        RECT 747.055 1114.320 747.345 1114.490 ;
        RECT 747.515 1114.320 747.805 1114.490 ;
        RECT 747.975 1114.320 748.265 1114.490 ;
        RECT 748.435 1114.320 748.725 1114.490 ;
        RECT 748.895 1114.320 749.185 1114.490 ;
        RECT 749.355 1114.320 749.645 1114.490 ;
        RECT 749.815 1114.320 750.105 1114.490 ;
        RECT 750.275 1114.320 750.565 1114.490 ;
        RECT 750.735 1114.320 751.025 1114.490 ;
        RECT 751.195 1114.320 751.485 1114.490 ;
        RECT 751.655 1114.320 751.945 1114.490 ;
        RECT 752.115 1114.320 752.405 1114.490 ;
        RECT 752.575 1114.320 752.865 1114.490 ;
        RECT 753.035 1114.320 753.325 1114.490 ;
        RECT 753.495 1114.320 753.785 1114.490 ;
        RECT 753.955 1114.320 754.245 1114.490 ;
        RECT 754.415 1114.320 754.705 1114.490 ;
        RECT 754.875 1114.320 755.165 1114.490 ;
        RECT 755.335 1114.320 755.625 1114.490 ;
        RECT 755.795 1114.320 756.085 1114.490 ;
        RECT 756.255 1114.320 756.545 1114.490 ;
        RECT 756.715 1114.320 757.005 1114.490 ;
        RECT 757.175 1114.320 757.465 1114.490 ;
        RECT 757.635 1114.320 757.925 1114.490 ;
        RECT 758.095 1114.320 758.385 1114.490 ;
        RECT 758.555 1114.320 758.845 1114.490 ;
        RECT 759.015 1114.320 759.305 1114.490 ;
        RECT 759.475 1114.320 759.765 1114.490 ;
        RECT 759.935 1114.320 760.225 1114.490 ;
        RECT 760.395 1114.320 760.685 1114.490 ;
        RECT 760.855 1114.320 761.145 1114.490 ;
        RECT 761.315 1114.320 761.605 1114.490 ;
        RECT 761.775 1114.320 762.065 1114.490 ;
        RECT 762.235 1114.320 762.525 1114.490 ;
        RECT 762.695 1114.320 762.985 1114.490 ;
        RECT 763.155 1114.320 763.445 1114.490 ;
        RECT 763.615 1114.320 763.905 1114.490 ;
        RECT 764.075 1114.320 764.365 1114.490 ;
        RECT 764.535 1114.320 764.825 1114.490 ;
        RECT 764.995 1114.320 765.285 1114.490 ;
        RECT 765.455 1114.320 765.745 1114.490 ;
        RECT 765.915 1114.320 766.205 1114.490 ;
        RECT 766.375 1114.320 766.665 1114.490 ;
        RECT 766.835 1114.320 767.125 1114.490 ;
        RECT 767.295 1114.320 767.585 1114.490 ;
        RECT 767.755 1114.320 768.045 1114.490 ;
        RECT 768.215 1114.320 768.505 1114.490 ;
        RECT 768.675 1114.320 768.965 1114.490 ;
        RECT 769.135 1114.320 769.425 1114.490 ;
        RECT 769.595 1114.320 769.885 1114.490 ;
        RECT 770.055 1114.320 770.345 1114.490 ;
        RECT 770.515 1114.320 770.805 1114.490 ;
        RECT 770.975 1114.320 771.120 1114.490 ;
        RECT 1969.000 1114.320 1969.145 1114.490 ;
        RECT 1969.315 1114.320 1969.605 1114.490 ;
        RECT 1969.775 1114.320 1970.065 1114.490 ;
        RECT 1970.235 1114.320 1970.525 1114.490 ;
        RECT 1970.695 1114.320 1970.985 1114.490 ;
        RECT 1971.155 1114.320 1971.445 1114.490 ;
        RECT 1971.615 1114.320 1971.905 1114.490 ;
        RECT 1972.075 1114.320 1972.365 1114.490 ;
        RECT 1972.535 1114.320 1972.825 1114.490 ;
        RECT 1972.995 1114.320 1973.285 1114.490 ;
        RECT 1973.455 1114.320 1973.745 1114.490 ;
        RECT 1973.915 1114.320 1974.205 1114.490 ;
        RECT 1974.375 1114.320 1974.665 1114.490 ;
        RECT 1974.835 1114.320 1975.125 1114.490 ;
        RECT 1975.295 1114.320 1975.585 1114.490 ;
        RECT 1975.755 1114.320 1976.045 1114.490 ;
        RECT 1976.215 1114.320 1976.505 1114.490 ;
        RECT 1976.675 1114.320 1976.965 1114.490 ;
        RECT 1977.135 1114.320 1977.425 1114.490 ;
        RECT 1977.595 1114.320 1977.885 1114.490 ;
        RECT 1978.055 1114.320 1978.345 1114.490 ;
        RECT 1978.515 1114.320 1978.805 1114.490 ;
        RECT 1978.975 1114.320 1979.265 1114.490 ;
        RECT 1979.435 1114.320 1979.725 1114.490 ;
        RECT 1979.895 1114.320 1980.185 1114.490 ;
        RECT 1980.355 1114.320 1980.645 1114.490 ;
        RECT 1980.815 1114.320 1981.105 1114.490 ;
        RECT 1981.275 1114.320 1981.565 1114.490 ;
        RECT 1981.735 1114.320 1982.025 1114.490 ;
        RECT 1982.195 1114.320 1982.485 1114.490 ;
        RECT 1982.655 1114.320 1982.945 1114.490 ;
        RECT 1983.115 1114.320 1983.405 1114.490 ;
        RECT 1983.575 1114.320 1983.865 1114.490 ;
        RECT 1984.035 1114.320 1984.325 1114.490 ;
        RECT 1984.495 1114.320 1984.785 1114.490 ;
        RECT 1984.955 1114.320 1985.245 1114.490 ;
        RECT 1985.415 1114.320 1985.705 1114.490 ;
        RECT 1985.875 1114.320 1986.165 1114.490 ;
        RECT 1986.335 1114.320 1986.625 1114.490 ;
        RECT 1986.795 1114.320 1987.085 1114.490 ;
        RECT 1987.255 1114.320 1987.545 1114.490 ;
        RECT 1987.715 1114.320 1988.005 1114.490 ;
        RECT 1988.175 1114.320 1988.465 1114.490 ;
        RECT 1988.635 1114.320 1988.925 1114.490 ;
        RECT 1989.095 1114.320 1989.385 1114.490 ;
        RECT 1989.555 1114.320 1989.845 1114.490 ;
        RECT 1990.015 1114.320 1990.305 1114.490 ;
        RECT 1990.475 1114.320 1990.765 1114.490 ;
        RECT 1990.935 1114.320 1991.225 1114.490 ;
        RECT 1991.395 1114.320 1991.685 1114.490 ;
        RECT 1991.855 1114.320 1992.145 1114.490 ;
        RECT 1992.315 1114.320 1992.605 1114.490 ;
        RECT 1992.775 1114.320 1993.065 1114.490 ;
        RECT 1993.235 1114.320 1993.525 1114.490 ;
        RECT 1993.695 1114.320 1993.985 1114.490 ;
        RECT 1994.155 1114.320 1994.445 1114.490 ;
        RECT 1994.615 1114.320 1994.905 1114.490 ;
        RECT 1995.075 1114.320 1995.365 1114.490 ;
        RECT 1995.535 1114.320 1995.825 1114.490 ;
        RECT 1995.995 1114.320 1996.285 1114.490 ;
        RECT 1996.455 1114.320 1996.745 1114.490 ;
        RECT 1996.915 1114.320 1997.205 1114.490 ;
        RECT 1997.375 1114.320 1997.665 1114.490 ;
        RECT 1997.835 1114.320 1998.125 1114.490 ;
        RECT 1998.295 1114.320 1998.585 1114.490 ;
        RECT 1998.755 1114.320 1999.045 1114.490 ;
        RECT 1999.215 1114.320 1999.505 1114.490 ;
        RECT 1999.675 1114.320 1999.965 1114.490 ;
        RECT 2000.135 1114.320 2000.425 1114.490 ;
        RECT 2000.595 1114.320 2000.885 1114.490 ;
        RECT 2001.055 1114.320 2001.345 1114.490 ;
        RECT 2001.515 1114.320 2001.805 1114.490 ;
        RECT 2001.975 1114.320 2002.265 1114.490 ;
        RECT 2002.435 1114.320 2002.725 1114.490 ;
        RECT 2002.895 1114.320 2003.185 1114.490 ;
        RECT 2003.355 1114.320 2003.645 1114.490 ;
        RECT 2003.815 1114.320 2004.105 1114.490 ;
        RECT 2004.275 1114.320 2004.565 1114.490 ;
        RECT 2004.735 1114.320 2005.025 1114.490 ;
        RECT 2005.195 1114.320 2005.485 1114.490 ;
        RECT 2005.655 1114.320 2005.945 1114.490 ;
        RECT 2006.115 1114.320 2006.405 1114.490 ;
        RECT 2006.575 1114.320 2006.865 1114.490 ;
        RECT 2007.035 1114.320 2007.325 1114.490 ;
        RECT 2007.495 1114.320 2007.785 1114.490 ;
        RECT 2007.955 1114.320 2008.245 1114.490 ;
        RECT 2008.415 1114.320 2008.705 1114.490 ;
        RECT 2008.875 1114.320 2009.165 1114.490 ;
        RECT 2009.335 1114.320 2009.625 1114.490 ;
        RECT 2009.795 1114.320 2010.085 1114.490 ;
        RECT 2010.255 1114.320 2010.545 1114.490 ;
        RECT 2010.715 1114.320 2011.005 1114.490 ;
        RECT 2011.175 1114.320 2011.465 1114.490 ;
        RECT 2011.635 1114.320 2011.925 1114.490 ;
        RECT 2012.095 1114.320 2012.385 1114.490 ;
        RECT 2012.555 1114.320 2012.845 1114.490 ;
        RECT 2013.015 1114.320 2013.305 1114.490 ;
        RECT 2013.475 1114.320 2013.765 1114.490 ;
        RECT 2013.935 1114.320 2014.225 1114.490 ;
        RECT 2014.395 1114.320 2014.685 1114.490 ;
        RECT 2014.855 1114.320 2015.145 1114.490 ;
        RECT 2015.315 1114.320 2015.605 1114.490 ;
        RECT 2015.775 1114.320 2016.065 1114.490 ;
        RECT 2016.235 1114.320 2016.525 1114.490 ;
        RECT 2016.695 1114.320 2016.985 1114.490 ;
        RECT 2017.155 1114.320 2017.445 1114.490 ;
        RECT 2017.615 1114.320 2017.905 1114.490 ;
        RECT 2018.075 1114.320 2018.365 1114.490 ;
        RECT 2018.535 1114.320 2018.825 1114.490 ;
        RECT 2018.995 1114.320 2019.285 1114.490 ;
        RECT 2019.455 1114.320 2019.745 1114.490 ;
        RECT 2019.915 1114.320 2020.205 1114.490 ;
        RECT 2020.375 1114.320 2020.665 1114.490 ;
        RECT 2020.835 1114.320 2021.125 1114.490 ;
        RECT 2021.295 1114.320 2021.585 1114.490 ;
        RECT 2021.755 1114.320 2022.045 1114.490 ;
        RECT 2022.215 1114.320 2022.505 1114.490 ;
        RECT 2022.675 1114.320 2022.965 1114.490 ;
        RECT 2023.135 1114.320 2023.425 1114.490 ;
        RECT 2023.595 1114.320 2023.885 1114.490 ;
        RECT 2024.055 1114.320 2024.345 1114.490 ;
        RECT 2024.515 1114.320 2024.805 1114.490 ;
        RECT 2024.975 1114.320 2025.265 1114.490 ;
        RECT 2025.435 1114.320 2025.725 1114.490 ;
        RECT 2025.895 1114.320 2026.185 1114.490 ;
        RECT 2026.355 1114.320 2026.645 1114.490 ;
        RECT 2026.815 1114.320 2027.105 1114.490 ;
        RECT 2027.275 1114.320 2027.565 1114.490 ;
        RECT 2027.735 1114.320 2028.025 1114.490 ;
        RECT 2028.195 1114.320 2028.485 1114.490 ;
        RECT 2028.655 1114.320 2028.945 1114.490 ;
        RECT 2029.115 1114.320 2029.405 1114.490 ;
        RECT 2029.575 1114.320 2029.865 1114.490 ;
        RECT 2030.035 1114.320 2030.325 1114.490 ;
        RECT 2030.495 1114.320 2030.785 1114.490 ;
        RECT 2030.955 1114.320 2031.245 1114.490 ;
        RECT 2031.415 1114.320 2031.705 1114.490 ;
        RECT 2031.875 1114.320 2032.165 1114.490 ;
        RECT 2032.335 1114.320 2032.625 1114.490 ;
        RECT 2032.795 1114.320 2033.085 1114.490 ;
        RECT 2033.255 1114.320 2033.545 1114.490 ;
        RECT 2033.715 1114.320 2034.005 1114.490 ;
        RECT 2034.175 1114.320 2034.465 1114.490 ;
        RECT 2034.635 1114.320 2034.925 1114.490 ;
        RECT 2035.095 1114.320 2035.385 1114.490 ;
        RECT 2035.555 1114.320 2035.845 1114.490 ;
        RECT 2036.015 1114.320 2036.305 1114.490 ;
        RECT 2036.475 1114.320 2036.765 1114.490 ;
        RECT 2036.935 1114.320 2037.225 1114.490 ;
        RECT 2037.395 1114.320 2037.685 1114.490 ;
        RECT 2037.855 1114.320 2038.145 1114.490 ;
        RECT 2038.315 1114.320 2038.605 1114.490 ;
        RECT 2038.775 1114.320 2039.065 1114.490 ;
        RECT 2039.235 1114.320 2039.525 1114.490 ;
        RECT 2039.695 1114.320 2039.985 1114.490 ;
        RECT 2040.155 1114.320 2040.445 1114.490 ;
        RECT 2040.615 1114.320 2040.905 1114.490 ;
        RECT 2041.075 1114.320 2041.365 1114.490 ;
        RECT 2041.535 1114.320 2041.825 1114.490 ;
        RECT 2041.995 1114.320 2042.285 1114.490 ;
        RECT 2042.455 1114.320 2042.745 1114.490 ;
        RECT 2042.915 1114.320 2043.205 1114.490 ;
        RECT 2043.375 1114.320 2043.665 1114.490 ;
        RECT 2043.835 1114.320 2044.125 1114.490 ;
        RECT 2044.295 1114.320 2044.585 1114.490 ;
        RECT 2044.755 1114.320 2045.045 1114.490 ;
        RECT 2045.215 1114.320 2045.505 1114.490 ;
        RECT 2045.675 1114.320 2045.965 1114.490 ;
        RECT 2046.135 1114.320 2046.425 1114.490 ;
        RECT 2046.595 1114.320 2046.885 1114.490 ;
        RECT 2047.055 1114.320 2047.345 1114.490 ;
        RECT 2047.515 1114.320 2047.805 1114.490 ;
        RECT 2047.975 1114.320 2048.265 1114.490 ;
        RECT 2048.435 1114.320 2048.725 1114.490 ;
        RECT 2048.895 1114.320 2049.185 1114.490 ;
        RECT 2049.355 1114.320 2049.645 1114.490 ;
        RECT 2049.815 1114.320 2050.105 1114.490 ;
        RECT 2050.275 1114.320 2050.565 1114.490 ;
        RECT 2050.735 1114.320 2051.025 1114.490 ;
        RECT 2051.195 1114.320 2051.485 1114.490 ;
        RECT 2051.655 1114.320 2051.945 1114.490 ;
        RECT 2052.115 1114.320 2052.405 1114.490 ;
        RECT 2052.575 1114.320 2052.865 1114.490 ;
        RECT 2053.035 1114.320 2053.325 1114.490 ;
        RECT 2053.495 1114.320 2053.785 1114.490 ;
        RECT 2053.955 1114.320 2054.245 1114.490 ;
        RECT 2054.415 1114.320 2054.705 1114.490 ;
        RECT 2054.875 1114.320 2055.165 1114.490 ;
        RECT 2055.335 1114.320 2055.625 1114.490 ;
        RECT 2055.795 1114.320 2056.085 1114.490 ;
        RECT 2056.255 1114.320 2056.545 1114.490 ;
        RECT 2056.715 1114.320 2057.005 1114.490 ;
        RECT 2057.175 1114.320 2057.465 1114.490 ;
        RECT 2057.635 1114.320 2057.925 1114.490 ;
        RECT 2058.095 1114.320 2058.385 1114.490 ;
        RECT 2058.555 1114.320 2058.845 1114.490 ;
        RECT 2059.015 1114.320 2059.305 1114.490 ;
        RECT 2059.475 1114.320 2059.765 1114.490 ;
        RECT 2059.935 1114.320 2060.225 1114.490 ;
        RECT 2060.395 1114.320 2060.685 1114.490 ;
        RECT 2060.855 1114.320 2061.145 1114.490 ;
        RECT 2061.315 1114.320 2061.605 1114.490 ;
        RECT 2061.775 1114.320 2062.065 1114.490 ;
        RECT 2062.235 1114.320 2062.525 1114.490 ;
        RECT 2062.695 1114.320 2062.985 1114.490 ;
        RECT 2063.155 1114.320 2063.445 1114.490 ;
        RECT 2063.615 1114.320 2063.905 1114.490 ;
        RECT 2064.075 1114.320 2064.365 1114.490 ;
        RECT 2064.535 1114.320 2064.825 1114.490 ;
        RECT 2064.995 1114.320 2065.285 1114.490 ;
        RECT 2065.455 1114.320 2065.745 1114.490 ;
        RECT 2065.915 1114.320 2066.205 1114.490 ;
        RECT 2066.375 1114.320 2066.665 1114.490 ;
        RECT 2066.835 1114.320 2067.125 1114.490 ;
        RECT 2067.295 1114.320 2067.585 1114.490 ;
        RECT 2067.755 1114.320 2068.045 1114.490 ;
        RECT 2068.215 1114.320 2068.505 1114.490 ;
        RECT 2068.675 1114.320 2068.965 1114.490 ;
        RECT 2069.135 1114.320 2069.425 1114.490 ;
        RECT 2069.595 1114.320 2069.885 1114.490 ;
        RECT 2070.055 1114.320 2070.345 1114.490 ;
        RECT 2070.515 1114.320 2070.805 1114.490 ;
        RECT 2070.975 1114.320 2071.120 1114.490 ;
        RECT 675.065 1113.155 675.355 1114.320 ;
        RECT 675.535 1113.300 675.865 1114.150 ;
        RECT 676.035 1113.520 676.205 1114.320 ;
        RECT 676.375 1113.300 676.705 1114.150 ;
        RECT 676.875 1113.520 677.045 1114.320 ;
      LAYER li1 ;
        RECT 677.295 1113.300 677.465 1114.150 ;
      LAYER li1 ;
        RECT 677.635 1113.520 677.965 1114.320 ;
      LAYER li1 ;
        RECT 678.135 1113.300 678.305 1114.150 ;
      LAYER li1 ;
        RECT 678.475 1113.520 678.805 1114.320 ;
      LAYER li1 ;
        RECT 678.975 1113.300 679.145 1114.150 ;
      LAYER li1 ;
        RECT 679.315 1113.520 679.645 1114.320 ;
      LAYER li1 ;
        RECT 679.815 1113.300 679.985 1114.150 ;
      LAYER li1 ;
        RECT 675.535 1113.130 677.035 1113.300 ;
      LAYER li1 ;
        RECT 677.295 1113.130 679.985 1113.300 ;
      LAYER li1 ;
        RECT 680.155 1113.170 680.485 1114.320 ;
        RECT 681.045 1113.155 681.335 1114.320 ;
        RECT 681.515 1113.300 681.845 1114.150 ;
        RECT 682.015 1113.520 682.185 1114.320 ;
        RECT 682.355 1113.300 682.685 1114.150 ;
        RECT 682.855 1113.520 683.025 1114.320 ;
      LAYER li1 ;
        RECT 683.275 1113.300 683.445 1114.150 ;
      LAYER li1 ;
        RECT 683.615 1113.520 683.945 1114.320 ;
      LAYER li1 ;
        RECT 684.115 1113.300 684.285 1114.150 ;
      LAYER li1 ;
        RECT 684.455 1113.520 684.785 1114.320 ;
      LAYER li1 ;
        RECT 684.955 1113.300 685.125 1114.150 ;
      LAYER li1 ;
        RECT 685.295 1113.520 685.625 1114.320 ;
      LAYER li1 ;
        RECT 685.795 1113.300 685.965 1114.150 ;
      LAYER li1 ;
        RECT 681.515 1113.130 683.015 1113.300 ;
      LAYER li1 ;
        RECT 683.275 1113.130 685.965 1113.300 ;
      LAYER li1 ;
        RECT 686.135 1113.170 686.465 1114.320 ;
        RECT 687.025 1113.155 687.315 1114.320 ;
        RECT 687.495 1113.300 687.825 1114.150 ;
        RECT 687.995 1113.520 688.165 1114.320 ;
        RECT 688.335 1113.300 688.665 1114.150 ;
        RECT 688.835 1113.520 689.005 1114.320 ;
      LAYER li1 ;
        RECT 689.255 1113.300 689.425 1114.150 ;
      LAYER li1 ;
        RECT 689.595 1113.520 689.925 1114.320 ;
      LAYER li1 ;
        RECT 690.095 1113.300 690.265 1114.150 ;
      LAYER li1 ;
        RECT 690.435 1113.520 690.765 1114.320 ;
      LAYER li1 ;
        RECT 690.935 1113.300 691.105 1114.150 ;
      LAYER li1 ;
        RECT 691.275 1113.520 691.605 1114.320 ;
      LAYER li1 ;
        RECT 691.775 1113.300 691.945 1114.150 ;
      LAYER li1 ;
        RECT 687.495 1113.130 688.995 1113.300 ;
      LAYER li1 ;
        RECT 689.255 1113.130 691.945 1113.300 ;
      LAYER li1 ;
        RECT 692.115 1113.170 692.445 1114.320 ;
        RECT 693.005 1113.155 693.295 1114.320 ;
        RECT 693.475 1113.300 693.805 1114.150 ;
        RECT 693.975 1113.520 694.145 1114.320 ;
        RECT 694.315 1113.300 694.645 1114.150 ;
        RECT 694.815 1113.520 694.985 1114.320 ;
      LAYER li1 ;
        RECT 695.235 1113.300 695.405 1114.150 ;
      LAYER li1 ;
        RECT 695.575 1113.520 695.905 1114.320 ;
      LAYER li1 ;
        RECT 696.075 1113.300 696.245 1114.150 ;
      LAYER li1 ;
        RECT 696.415 1113.520 696.745 1114.320 ;
      LAYER li1 ;
        RECT 696.915 1113.300 697.085 1114.150 ;
      LAYER li1 ;
        RECT 697.255 1113.520 697.585 1114.320 ;
      LAYER li1 ;
        RECT 697.755 1113.300 697.925 1114.150 ;
      LAYER li1 ;
        RECT 693.475 1113.130 694.975 1113.300 ;
      LAYER li1 ;
        RECT 695.235 1113.130 697.925 1113.300 ;
      LAYER li1 ;
        RECT 698.095 1113.170 698.425 1114.320 ;
        RECT 698.985 1113.155 699.275 1114.320 ;
        RECT 699.455 1113.300 699.785 1114.150 ;
        RECT 699.955 1113.520 700.125 1114.320 ;
        RECT 700.295 1113.300 700.625 1114.150 ;
        RECT 700.795 1113.520 700.965 1114.320 ;
      LAYER li1 ;
        RECT 701.215 1113.300 701.385 1114.150 ;
      LAYER li1 ;
        RECT 701.555 1113.520 701.885 1114.320 ;
      LAYER li1 ;
        RECT 702.055 1113.300 702.225 1114.150 ;
      LAYER li1 ;
        RECT 702.395 1113.520 702.725 1114.320 ;
      LAYER li1 ;
        RECT 702.895 1113.300 703.065 1114.150 ;
      LAYER li1 ;
        RECT 703.235 1113.520 703.565 1114.320 ;
      LAYER li1 ;
        RECT 703.735 1113.300 703.905 1114.150 ;
      LAYER li1 ;
        RECT 699.455 1113.130 700.955 1113.300 ;
      LAYER li1 ;
        RECT 701.215 1113.130 703.905 1113.300 ;
      LAYER li1 ;
        RECT 704.075 1113.170 704.405 1114.320 ;
        RECT 704.965 1113.155 705.255 1114.320 ;
        RECT 705.435 1113.300 705.765 1114.150 ;
        RECT 705.935 1113.520 706.105 1114.320 ;
        RECT 706.275 1113.300 706.605 1114.150 ;
        RECT 706.775 1113.520 706.945 1114.320 ;
      LAYER li1 ;
        RECT 707.195 1113.300 707.365 1114.150 ;
      LAYER li1 ;
        RECT 707.535 1113.520 707.865 1114.320 ;
      LAYER li1 ;
        RECT 708.035 1113.300 708.205 1114.150 ;
      LAYER li1 ;
        RECT 708.375 1113.520 708.705 1114.320 ;
      LAYER li1 ;
        RECT 708.875 1113.300 709.045 1114.150 ;
      LAYER li1 ;
        RECT 709.215 1113.520 709.545 1114.320 ;
      LAYER li1 ;
        RECT 709.715 1113.300 709.885 1114.150 ;
      LAYER li1 ;
        RECT 705.435 1113.130 706.935 1113.300 ;
      LAYER li1 ;
        RECT 707.195 1113.130 709.885 1113.300 ;
      LAYER li1 ;
        RECT 710.055 1113.170 710.385 1114.320 ;
        RECT 710.945 1113.155 711.235 1114.320 ;
        RECT 711.415 1113.300 711.745 1114.150 ;
        RECT 711.915 1113.520 712.085 1114.320 ;
        RECT 712.255 1113.300 712.585 1114.150 ;
        RECT 712.755 1113.520 712.925 1114.320 ;
      LAYER li1 ;
        RECT 713.175 1113.300 713.345 1114.150 ;
      LAYER li1 ;
        RECT 713.515 1113.520 713.845 1114.320 ;
      LAYER li1 ;
        RECT 714.015 1113.300 714.185 1114.150 ;
      LAYER li1 ;
        RECT 714.355 1113.520 714.685 1114.320 ;
      LAYER li1 ;
        RECT 714.855 1113.300 715.025 1114.150 ;
      LAYER li1 ;
        RECT 715.195 1113.520 715.525 1114.320 ;
      LAYER li1 ;
        RECT 715.695 1113.300 715.865 1114.150 ;
      LAYER li1 ;
        RECT 711.415 1113.130 712.915 1113.300 ;
      LAYER li1 ;
        RECT 713.175 1113.130 715.865 1113.300 ;
      LAYER li1 ;
        RECT 716.035 1113.170 716.365 1114.320 ;
        RECT 716.925 1113.155 717.215 1114.320 ;
        RECT 717.395 1113.300 717.725 1114.150 ;
        RECT 717.895 1113.520 718.065 1114.320 ;
        RECT 718.235 1113.300 718.565 1114.150 ;
        RECT 718.735 1113.520 718.905 1114.320 ;
      LAYER li1 ;
        RECT 719.155 1113.300 719.325 1114.150 ;
      LAYER li1 ;
        RECT 719.495 1113.520 719.825 1114.320 ;
      LAYER li1 ;
        RECT 719.995 1113.300 720.165 1114.150 ;
      LAYER li1 ;
        RECT 720.335 1113.520 720.665 1114.320 ;
      LAYER li1 ;
        RECT 720.835 1113.300 721.005 1114.150 ;
      LAYER li1 ;
        RECT 721.175 1113.520 721.505 1114.320 ;
      LAYER li1 ;
        RECT 721.675 1113.300 721.845 1114.150 ;
      LAYER li1 ;
        RECT 717.395 1113.130 718.895 1113.300 ;
      LAYER li1 ;
        RECT 719.155 1113.130 721.845 1113.300 ;
      LAYER li1 ;
        RECT 722.015 1113.170 722.345 1114.320 ;
        RECT 722.905 1113.155 723.195 1114.320 ;
        RECT 723.375 1113.300 723.705 1114.150 ;
        RECT 723.875 1113.520 724.045 1114.320 ;
        RECT 724.215 1113.300 724.545 1114.150 ;
        RECT 724.715 1113.520 724.885 1114.320 ;
      LAYER li1 ;
        RECT 725.135 1113.300 725.305 1114.150 ;
      LAYER li1 ;
        RECT 725.475 1113.520 725.805 1114.320 ;
      LAYER li1 ;
        RECT 725.975 1113.300 726.145 1114.150 ;
      LAYER li1 ;
        RECT 726.315 1113.520 726.645 1114.320 ;
      LAYER li1 ;
        RECT 726.815 1113.300 726.985 1114.150 ;
      LAYER li1 ;
        RECT 727.155 1113.520 727.485 1114.320 ;
      LAYER li1 ;
        RECT 727.655 1113.300 727.825 1114.150 ;
      LAYER li1 ;
        RECT 723.375 1113.130 724.875 1113.300 ;
      LAYER li1 ;
        RECT 725.135 1113.130 727.825 1113.300 ;
      LAYER li1 ;
        RECT 727.995 1113.170 728.325 1114.320 ;
        RECT 728.885 1113.155 729.175 1114.320 ;
        RECT 729.355 1113.300 729.685 1114.150 ;
        RECT 729.855 1113.520 730.025 1114.320 ;
        RECT 730.195 1113.300 730.525 1114.150 ;
        RECT 730.695 1113.520 730.865 1114.320 ;
      LAYER li1 ;
        RECT 731.115 1113.300 731.285 1114.150 ;
      LAYER li1 ;
        RECT 731.455 1113.520 731.785 1114.320 ;
      LAYER li1 ;
        RECT 731.955 1113.300 732.125 1114.150 ;
      LAYER li1 ;
        RECT 732.295 1113.520 732.625 1114.320 ;
      LAYER li1 ;
        RECT 732.795 1113.300 732.965 1114.150 ;
      LAYER li1 ;
        RECT 733.135 1113.520 733.465 1114.320 ;
      LAYER li1 ;
        RECT 733.635 1113.300 733.805 1114.150 ;
      LAYER li1 ;
        RECT 729.355 1113.130 730.855 1113.300 ;
      LAYER li1 ;
        RECT 731.115 1113.130 733.805 1113.300 ;
      LAYER li1 ;
        RECT 733.975 1113.170 734.305 1114.320 ;
        RECT 734.865 1113.155 735.155 1114.320 ;
        RECT 735.335 1113.300 735.665 1114.150 ;
        RECT 735.835 1113.520 736.005 1114.320 ;
        RECT 736.175 1113.300 736.505 1114.150 ;
        RECT 736.675 1113.520 736.845 1114.320 ;
      LAYER li1 ;
        RECT 737.095 1113.300 737.265 1114.150 ;
      LAYER li1 ;
        RECT 737.435 1113.520 737.765 1114.320 ;
      LAYER li1 ;
        RECT 737.935 1113.300 738.105 1114.150 ;
      LAYER li1 ;
        RECT 738.275 1113.520 738.605 1114.320 ;
      LAYER li1 ;
        RECT 738.775 1113.300 738.945 1114.150 ;
      LAYER li1 ;
        RECT 739.115 1113.520 739.445 1114.320 ;
      LAYER li1 ;
        RECT 739.615 1113.300 739.785 1114.150 ;
      LAYER li1 ;
        RECT 735.335 1113.130 736.835 1113.300 ;
      LAYER li1 ;
        RECT 737.095 1113.130 739.785 1113.300 ;
      LAYER li1 ;
        RECT 739.955 1113.170 740.285 1114.320 ;
        RECT 740.845 1113.155 741.135 1114.320 ;
        RECT 741.315 1113.300 741.645 1114.150 ;
        RECT 741.815 1113.520 741.985 1114.320 ;
        RECT 742.155 1113.300 742.485 1114.150 ;
        RECT 742.655 1113.520 742.825 1114.320 ;
      LAYER li1 ;
        RECT 743.075 1113.300 743.245 1114.150 ;
      LAYER li1 ;
        RECT 743.415 1113.520 743.745 1114.320 ;
      LAYER li1 ;
        RECT 743.915 1113.300 744.085 1114.150 ;
      LAYER li1 ;
        RECT 744.255 1113.520 744.585 1114.320 ;
      LAYER li1 ;
        RECT 744.755 1113.300 744.925 1114.150 ;
      LAYER li1 ;
        RECT 745.095 1113.520 745.425 1114.320 ;
      LAYER li1 ;
        RECT 745.595 1113.300 745.765 1114.150 ;
      LAYER li1 ;
        RECT 741.315 1113.130 742.815 1113.300 ;
      LAYER li1 ;
        RECT 743.075 1113.130 745.765 1113.300 ;
      LAYER li1 ;
        RECT 745.935 1113.170 746.265 1114.320 ;
        RECT 746.825 1113.155 747.115 1114.320 ;
        RECT 747.295 1113.300 747.625 1114.150 ;
        RECT 747.795 1113.520 747.965 1114.320 ;
        RECT 748.135 1113.300 748.465 1114.150 ;
        RECT 748.635 1113.520 748.805 1114.320 ;
      LAYER li1 ;
        RECT 749.055 1113.300 749.225 1114.150 ;
      LAYER li1 ;
        RECT 749.395 1113.520 749.725 1114.320 ;
      LAYER li1 ;
        RECT 749.895 1113.300 750.065 1114.150 ;
      LAYER li1 ;
        RECT 750.235 1113.520 750.565 1114.320 ;
      LAYER li1 ;
        RECT 750.735 1113.300 750.905 1114.150 ;
      LAYER li1 ;
        RECT 751.075 1113.520 751.405 1114.320 ;
      LAYER li1 ;
        RECT 751.575 1113.300 751.745 1114.150 ;
      LAYER li1 ;
        RECT 747.295 1113.130 748.795 1113.300 ;
      LAYER li1 ;
        RECT 749.055 1113.130 751.745 1113.300 ;
      LAYER li1 ;
        RECT 751.915 1113.170 752.245 1114.320 ;
        RECT 752.805 1113.155 753.095 1114.320 ;
        RECT 753.275 1113.300 753.605 1114.150 ;
        RECT 753.775 1113.520 753.945 1114.320 ;
        RECT 754.115 1113.300 754.445 1114.150 ;
        RECT 754.615 1113.520 754.785 1114.320 ;
      LAYER li1 ;
        RECT 755.035 1113.300 755.205 1114.150 ;
      LAYER li1 ;
        RECT 755.375 1113.520 755.705 1114.320 ;
      LAYER li1 ;
        RECT 755.875 1113.300 756.045 1114.150 ;
      LAYER li1 ;
        RECT 756.215 1113.520 756.545 1114.320 ;
      LAYER li1 ;
        RECT 756.715 1113.300 756.885 1114.150 ;
      LAYER li1 ;
        RECT 757.055 1113.520 757.385 1114.320 ;
      LAYER li1 ;
        RECT 757.555 1113.300 757.725 1114.150 ;
      LAYER li1 ;
        RECT 753.275 1113.130 754.775 1113.300 ;
      LAYER li1 ;
        RECT 755.035 1113.130 757.725 1113.300 ;
      LAYER li1 ;
        RECT 757.895 1113.170 758.225 1114.320 ;
        RECT 758.785 1113.155 759.075 1114.320 ;
        RECT 759.255 1113.300 759.585 1114.150 ;
        RECT 759.755 1113.520 759.925 1114.320 ;
        RECT 760.095 1113.300 760.425 1114.150 ;
        RECT 760.595 1113.520 760.765 1114.320 ;
      LAYER li1 ;
        RECT 761.015 1113.300 761.185 1114.150 ;
      LAYER li1 ;
        RECT 761.355 1113.520 761.685 1114.320 ;
      LAYER li1 ;
        RECT 761.855 1113.300 762.025 1114.150 ;
      LAYER li1 ;
        RECT 762.195 1113.520 762.525 1114.320 ;
      LAYER li1 ;
        RECT 762.695 1113.300 762.865 1114.150 ;
      LAYER li1 ;
        RECT 763.035 1113.520 763.365 1114.320 ;
      LAYER li1 ;
        RECT 763.535 1113.300 763.705 1114.150 ;
      LAYER li1 ;
        RECT 759.255 1113.130 760.755 1113.300 ;
      LAYER li1 ;
        RECT 761.015 1113.130 763.705 1113.300 ;
      LAYER li1 ;
        RECT 763.875 1113.170 764.205 1114.320 ;
        RECT 764.765 1113.155 765.055 1114.320 ;
        RECT 765.615 1113.170 765.945 1114.320 ;
        RECT 766.455 1113.520 766.785 1114.320 ;
        RECT 767.295 1113.520 767.625 1114.320 ;
        RECT 768.135 1113.520 768.465 1114.320 ;
        RECT 769.055 1113.520 769.225 1114.320 ;
        RECT 769.395 1113.300 769.725 1114.150 ;
        RECT 769.895 1113.520 770.065 1114.320 ;
        RECT 770.235 1113.300 770.565 1114.150 ;
      LAYER li1 ;
        RECT 675.580 1112.760 676.680 1112.960 ;
      LAYER li1 ;
        RECT 676.860 1112.930 677.035 1113.130 ;
        RECT 676.860 1112.760 679.485 1112.930 ;
        RECT 676.860 1112.590 677.035 1112.760 ;
      LAYER li1 ;
        RECT 679.730 1112.590 679.985 1113.130 ;
        RECT 681.560 1112.760 682.660 1112.960 ;
      LAYER li1 ;
        RECT 682.840 1112.930 683.015 1113.130 ;
        RECT 682.840 1112.760 685.465 1112.930 ;
        RECT 682.840 1112.590 683.015 1112.760 ;
      LAYER li1 ;
        RECT 685.710 1112.590 685.965 1113.130 ;
        RECT 687.540 1112.760 688.640 1112.960 ;
      LAYER li1 ;
        RECT 688.820 1112.930 688.995 1113.130 ;
        RECT 688.820 1112.760 691.445 1112.930 ;
        RECT 688.820 1112.590 688.995 1112.760 ;
      LAYER li1 ;
        RECT 691.690 1112.590 691.945 1113.130 ;
        RECT 693.520 1112.760 694.620 1112.960 ;
      LAYER li1 ;
        RECT 694.800 1112.930 694.975 1113.130 ;
        RECT 694.800 1112.760 697.425 1112.930 ;
        RECT 694.800 1112.590 694.975 1112.760 ;
      LAYER li1 ;
        RECT 697.670 1112.590 697.925 1113.130 ;
        RECT 699.500 1112.760 700.600 1112.960 ;
      LAYER li1 ;
        RECT 700.780 1112.930 700.955 1113.130 ;
        RECT 700.780 1112.760 703.405 1112.930 ;
        RECT 700.780 1112.590 700.955 1112.760 ;
      LAYER li1 ;
        RECT 703.650 1112.590 703.905 1113.130 ;
        RECT 705.480 1112.760 706.580 1112.960 ;
      LAYER li1 ;
        RECT 706.760 1112.930 706.935 1113.130 ;
        RECT 706.760 1112.760 709.385 1112.930 ;
        RECT 706.760 1112.590 706.935 1112.760 ;
      LAYER li1 ;
        RECT 709.630 1112.590 709.885 1113.130 ;
        RECT 711.460 1112.760 712.560 1112.960 ;
      LAYER li1 ;
        RECT 712.740 1112.930 712.915 1113.130 ;
        RECT 712.740 1112.760 715.365 1112.930 ;
        RECT 712.740 1112.590 712.915 1112.760 ;
      LAYER li1 ;
        RECT 715.610 1112.590 715.865 1113.130 ;
        RECT 717.440 1112.760 718.540 1112.960 ;
      LAYER li1 ;
        RECT 718.720 1112.930 718.895 1113.130 ;
        RECT 718.720 1112.760 721.345 1112.930 ;
        RECT 718.720 1112.590 718.895 1112.760 ;
      LAYER li1 ;
        RECT 721.590 1112.590 721.845 1113.130 ;
        RECT 723.420 1112.760 724.520 1112.960 ;
      LAYER li1 ;
        RECT 724.700 1112.930 724.875 1113.130 ;
        RECT 724.700 1112.760 727.325 1112.930 ;
        RECT 724.700 1112.590 724.875 1112.760 ;
      LAYER li1 ;
        RECT 727.570 1112.590 727.825 1113.130 ;
        RECT 729.400 1112.760 730.500 1112.960 ;
      LAYER li1 ;
        RECT 730.680 1112.930 730.855 1113.130 ;
        RECT 730.680 1112.760 733.305 1112.930 ;
        RECT 730.680 1112.590 730.855 1112.760 ;
      LAYER li1 ;
        RECT 733.550 1112.590 733.805 1113.130 ;
        RECT 735.380 1112.760 736.480 1112.960 ;
      LAYER li1 ;
        RECT 736.660 1112.930 736.835 1113.130 ;
        RECT 736.660 1112.760 739.285 1112.930 ;
        RECT 736.660 1112.590 736.835 1112.760 ;
      LAYER li1 ;
        RECT 739.530 1112.590 739.785 1113.130 ;
      LAYER li1 ;
        RECT 742.640 1112.930 742.815 1113.130 ;
        RECT 742.640 1112.760 745.265 1112.930 ;
        RECT 742.640 1112.590 742.815 1112.760 ;
      LAYER li1 ;
        RECT 745.510 1112.590 745.765 1113.130 ;
      LAYER li1 ;
        RECT 748.620 1112.930 748.795 1113.130 ;
        RECT 748.620 1112.760 751.245 1112.930 ;
        RECT 748.620 1112.590 748.795 1112.760 ;
      LAYER li1 ;
        RECT 751.490 1112.590 751.745 1113.130 ;
      LAYER li1 ;
        RECT 754.600 1112.930 754.775 1113.130 ;
        RECT 754.600 1112.760 757.225 1112.930 ;
        RECT 754.600 1112.590 754.775 1112.760 ;
      LAYER li1 ;
        RECT 757.470 1112.590 757.725 1113.130 ;
      LAYER li1 ;
        RECT 760.580 1112.930 760.755 1113.130 ;
        RECT 760.580 1112.760 763.205 1112.930 ;
        RECT 760.580 1112.590 760.755 1112.760 ;
      LAYER li1 ;
        RECT 763.450 1112.590 763.705 1113.130 ;
      LAYER li1 ;
        RECT 769.065 1113.130 770.565 1113.300 ;
        RECT 770.745 1113.155 771.035 1114.320 ;
        RECT 1975.065 1113.155 1975.355 1114.320 ;
        RECT 1975.535 1113.300 1975.865 1114.150 ;
        RECT 1976.035 1113.520 1976.205 1114.320 ;
        RECT 1976.375 1113.300 1976.705 1114.150 ;
        RECT 1976.875 1113.520 1977.045 1114.320 ;
        RECT 1977.635 1113.520 1977.965 1114.320 ;
        RECT 1978.475 1113.520 1978.805 1114.320 ;
        RECT 1979.315 1113.520 1979.645 1114.320 ;
        RECT 1975.535 1113.130 1977.035 1113.300 ;
        RECT 1980.155 1113.170 1980.485 1114.320 ;
        RECT 1981.045 1113.155 1981.335 1114.320 ;
        RECT 1981.515 1113.300 1981.845 1114.150 ;
        RECT 1982.015 1113.520 1982.185 1114.320 ;
        RECT 1982.355 1113.300 1982.685 1114.150 ;
        RECT 1982.855 1113.520 1983.025 1114.320 ;
        RECT 1983.615 1113.520 1983.945 1114.320 ;
        RECT 1984.455 1113.520 1984.785 1114.320 ;
        RECT 1985.295 1113.520 1985.625 1114.320 ;
        RECT 1981.515 1113.130 1983.015 1113.300 ;
        RECT 1986.135 1113.170 1986.465 1114.320 ;
        RECT 1987.025 1113.155 1987.315 1114.320 ;
        RECT 1987.495 1113.300 1987.825 1114.150 ;
        RECT 1987.995 1113.520 1988.165 1114.320 ;
        RECT 1988.335 1113.300 1988.665 1114.150 ;
        RECT 1988.835 1113.520 1989.005 1114.320 ;
        RECT 1989.595 1113.520 1989.925 1114.320 ;
        RECT 1990.435 1113.520 1990.765 1114.320 ;
        RECT 1991.275 1113.520 1991.605 1114.320 ;
        RECT 1987.495 1113.130 1988.995 1113.300 ;
        RECT 1992.115 1113.170 1992.445 1114.320 ;
        RECT 1993.005 1113.155 1993.295 1114.320 ;
        RECT 1993.475 1113.300 1993.805 1114.150 ;
        RECT 1993.975 1113.520 1994.145 1114.320 ;
        RECT 1994.315 1113.300 1994.645 1114.150 ;
        RECT 1994.815 1113.520 1994.985 1114.320 ;
        RECT 1995.575 1113.520 1995.905 1114.320 ;
        RECT 1996.415 1113.520 1996.745 1114.320 ;
        RECT 1997.255 1113.520 1997.585 1114.320 ;
        RECT 1993.475 1113.130 1994.975 1113.300 ;
        RECT 1998.095 1113.170 1998.425 1114.320 ;
        RECT 1998.985 1113.155 1999.275 1114.320 ;
        RECT 1999.455 1113.300 1999.785 1114.150 ;
        RECT 1999.955 1113.520 2000.125 1114.320 ;
        RECT 2000.295 1113.300 2000.625 1114.150 ;
        RECT 2000.795 1113.520 2000.965 1114.320 ;
        RECT 2001.555 1113.520 2001.885 1114.320 ;
        RECT 2002.395 1113.520 2002.725 1114.320 ;
        RECT 2003.235 1113.520 2003.565 1114.320 ;
        RECT 1999.455 1113.130 2000.955 1113.300 ;
        RECT 2004.075 1113.170 2004.405 1114.320 ;
        RECT 2004.965 1113.155 2005.255 1114.320 ;
        RECT 2005.435 1113.300 2005.765 1114.150 ;
        RECT 2005.935 1113.520 2006.105 1114.320 ;
        RECT 2006.275 1113.300 2006.605 1114.150 ;
        RECT 2006.775 1113.520 2006.945 1114.320 ;
        RECT 2007.535 1113.520 2007.865 1114.320 ;
        RECT 2008.375 1113.520 2008.705 1114.320 ;
        RECT 2009.215 1113.520 2009.545 1114.320 ;
        RECT 2005.435 1113.130 2006.935 1113.300 ;
        RECT 2010.055 1113.170 2010.385 1114.320 ;
        RECT 2010.945 1113.155 2011.235 1114.320 ;
        RECT 2011.415 1113.300 2011.745 1114.150 ;
        RECT 2011.915 1113.520 2012.085 1114.320 ;
        RECT 2012.255 1113.300 2012.585 1114.150 ;
        RECT 2012.755 1113.520 2012.925 1114.320 ;
        RECT 2013.515 1113.520 2013.845 1114.320 ;
        RECT 2014.355 1113.520 2014.685 1114.320 ;
        RECT 2015.195 1113.520 2015.525 1114.320 ;
        RECT 2011.415 1113.130 2012.915 1113.300 ;
        RECT 2016.035 1113.170 2016.365 1114.320 ;
        RECT 2016.925 1113.155 2017.215 1114.320 ;
        RECT 2017.395 1113.300 2017.725 1114.150 ;
        RECT 2017.895 1113.520 2018.065 1114.320 ;
        RECT 2018.235 1113.300 2018.565 1114.150 ;
        RECT 2018.735 1113.520 2018.905 1114.320 ;
        RECT 2019.495 1113.520 2019.825 1114.320 ;
        RECT 2020.335 1113.520 2020.665 1114.320 ;
        RECT 2021.175 1113.520 2021.505 1114.320 ;
        RECT 2017.395 1113.130 2018.895 1113.300 ;
        RECT 2022.015 1113.170 2022.345 1114.320 ;
        RECT 2022.905 1113.155 2023.195 1114.320 ;
        RECT 2023.375 1113.300 2023.705 1114.150 ;
        RECT 2023.875 1113.520 2024.045 1114.320 ;
        RECT 2024.215 1113.300 2024.545 1114.150 ;
        RECT 2024.715 1113.520 2024.885 1114.320 ;
        RECT 2025.475 1113.520 2025.805 1114.320 ;
        RECT 2026.315 1113.520 2026.645 1114.320 ;
        RECT 2027.155 1113.520 2027.485 1114.320 ;
        RECT 2023.375 1113.130 2024.875 1113.300 ;
        RECT 2027.995 1113.170 2028.325 1114.320 ;
        RECT 2028.885 1113.155 2029.175 1114.320 ;
        RECT 2029.355 1113.300 2029.685 1114.150 ;
        RECT 2029.855 1113.520 2030.025 1114.320 ;
        RECT 2030.195 1113.300 2030.525 1114.150 ;
        RECT 2030.695 1113.520 2030.865 1114.320 ;
        RECT 2031.455 1113.520 2031.785 1114.320 ;
        RECT 2032.295 1113.520 2032.625 1114.320 ;
        RECT 2033.135 1113.520 2033.465 1114.320 ;
        RECT 2029.355 1113.130 2030.855 1113.300 ;
        RECT 2033.975 1113.170 2034.305 1114.320 ;
        RECT 2034.865 1113.155 2035.155 1114.320 ;
        RECT 2035.335 1113.300 2035.665 1114.150 ;
        RECT 2035.835 1113.520 2036.005 1114.320 ;
        RECT 2036.175 1113.300 2036.505 1114.150 ;
        RECT 2036.675 1113.520 2036.845 1114.320 ;
      LAYER li1 ;
        RECT 2037.095 1113.300 2037.265 1114.150 ;
      LAYER li1 ;
        RECT 2037.435 1113.520 2037.765 1114.320 ;
      LAYER li1 ;
        RECT 2037.935 1113.300 2038.105 1114.150 ;
      LAYER li1 ;
        RECT 2038.275 1113.520 2038.605 1114.320 ;
      LAYER li1 ;
        RECT 2038.775 1113.300 2038.945 1114.150 ;
      LAYER li1 ;
        RECT 2039.115 1113.520 2039.445 1114.320 ;
      LAYER li1 ;
        RECT 2039.615 1113.300 2039.785 1114.150 ;
      LAYER li1 ;
        RECT 2035.335 1113.130 2036.835 1113.300 ;
      LAYER li1 ;
        RECT 2037.095 1113.130 2039.785 1113.300 ;
      LAYER li1 ;
        RECT 2039.955 1113.170 2040.285 1114.320 ;
        RECT 2040.845 1113.155 2041.135 1114.320 ;
        RECT 2041.315 1113.300 2041.645 1114.150 ;
        RECT 2041.815 1113.520 2041.985 1114.320 ;
        RECT 2042.155 1113.300 2042.485 1114.150 ;
        RECT 2042.655 1113.520 2042.825 1114.320 ;
        RECT 2043.415 1113.520 2043.745 1114.320 ;
        RECT 2044.255 1113.520 2044.585 1114.320 ;
        RECT 2045.095 1113.520 2045.425 1114.320 ;
        RECT 2041.315 1113.130 2042.815 1113.300 ;
        RECT 2045.935 1113.170 2046.265 1114.320 ;
        RECT 2046.825 1113.155 2047.115 1114.320 ;
        RECT 2047.295 1113.300 2047.625 1114.150 ;
        RECT 2047.795 1113.520 2047.965 1114.320 ;
        RECT 2048.135 1113.300 2048.465 1114.150 ;
        RECT 2048.635 1113.520 2048.805 1114.320 ;
        RECT 2049.395 1113.520 2049.725 1114.320 ;
        RECT 2050.235 1113.520 2050.565 1114.320 ;
        RECT 2051.075 1113.520 2051.405 1114.320 ;
        RECT 2047.295 1113.130 2048.795 1113.300 ;
        RECT 2051.915 1113.170 2052.245 1114.320 ;
        RECT 2052.805 1113.155 2053.095 1114.320 ;
        RECT 2053.275 1113.300 2053.605 1114.150 ;
        RECT 2053.775 1113.520 2053.945 1114.320 ;
        RECT 2054.115 1113.300 2054.445 1114.150 ;
        RECT 2054.615 1113.520 2054.785 1114.320 ;
        RECT 2055.375 1113.520 2055.705 1114.320 ;
        RECT 2056.215 1113.520 2056.545 1114.320 ;
        RECT 2057.055 1113.520 2057.385 1114.320 ;
        RECT 2053.275 1113.130 2054.775 1113.300 ;
        RECT 2057.895 1113.170 2058.225 1114.320 ;
        RECT 2058.785 1113.155 2059.075 1114.320 ;
        RECT 2059.255 1113.300 2059.585 1114.150 ;
        RECT 2059.755 1113.520 2059.925 1114.320 ;
        RECT 2060.095 1113.300 2060.425 1114.150 ;
        RECT 2060.595 1113.520 2060.765 1114.320 ;
        RECT 2061.355 1113.520 2061.685 1114.320 ;
        RECT 2062.195 1113.520 2062.525 1114.320 ;
        RECT 2063.035 1113.520 2063.365 1114.320 ;
        RECT 2059.255 1113.130 2060.755 1113.300 ;
        RECT 2063.875 1113.170 2064.205 1114.320 ;
        RECT 2064.765 1113.155 2065.055 1114.320 ;
        RECT 2065.615 1113.170 2065.945 1114.320 ;
      LAYER li1 ;
        RECT 2066.115 1113.300 2066.285 1114.150 ;
      LAYER li1 ;
        RECT 2066.455 1113.520 2066.785 1114.320 ;
      LAYER li1 ;
        RECT 2066.955 1113.300 2067.125 1114.150 ;
      LAYER li1 ;
        RECT 2067.295 1113.520 2067.625 1114.320 ;
      LAYER li1 ;
        RECT 2067.795 1113.300 2067.965 1114.150 ;
      LAYER li1 ;
        RECT 2068.135 1113.520 2068.465 1114.320 ;
      LAYER li1 ;
        RECT 2068.635 1113.300 2068.805 1114.150 ;
      LAYER li1 ;
        RECT 2069.055 1113.520 2069.225 1114.320 ;
        RECT 2069.395 1113.300 2069.725 1114.150 ;
        RECT 2069.895 1113.520 2070.065 1114.320 ;
        RECT 2070.235 1113.300 2070.565 1114.150 ;
        RECT 769.065 1112.930 769.240 1113.130 ;
        RECT 766.615 1112.760 769.240 1112.930 ;
      LAYER li1 ;
        RECT 769.420 1112.760 770.520 1112.960 ;
        RECT 1975.580 1112.760 1976.680 1112.960 ;
      LAYER li1 ;
        RECT 1976.860 1112.930 1977.035 1113.130 ;
        RECT 1976.860 1112.760 1979.485 1112.930 ;
      LAYER li1 ;
        RECT 1981.560 1112.760 1982.660 1112.960 ;
      LAYER li1 ;
        RECT 1982.840 1112.930 1983.015 1113.130 ;
        RECT 1982.840 1112.760 1985.465 1112.930 ;
      LAYER li1 ;
        RECT 1987.540 1112.760 1988.640 1112.960 ;
      LAYER li1 ;
        RECT 1988.820 1112.930 1988.995 1113.130 ;
        RECT 1988.820 1112.760 1991.445 1112.930 ;
      LAYER li1 ;
        RECT 1993.520 1112.760 1994.620 1112.960 ;
      LAYER li1 ;
        RECT 1994.800 1112.930 1994.975 1113.130 ;
        RECT 1994.800 1112.760 1997.425 1112.930 ;
      LAYER li1 ;
        RECT 1999.500 1112.760 2000.600 1112.960 ;
      LAYER li1 ;
        RECT 2000.780 1112.930 2000.955 1113.130 ;
        RECT 2000.780 1112.760 2003.405 1112.930 ;
      LAYER li1 ;
        RECT 2005.480 1112.760 2006.580 1112.960 ;
      LAYER li1 ;
        RECT 2006.760 1112.930 2006.935 1113.130 ;
        RECT 2006.760 1112.760 2009.385 1112.930 ;
      LAYER li1 ;
        RECT 2011.460 1112.760 2012.560 1112.960 ;
      LAYER li1 ;
        RECT 2012.740 1112.930 2012.915 1113.130 ;
        RECT 2012.740 1112.760 2015.365 1112.930 ;
      LAYER li1 ;
        RECT 2017.440 1112.760 2018.540 1112.960 ;
      LAYER li1 ;
        RECT 2018.720 1112.930 2018.895 1113.130 ;
        RECT 2018.720 1112.760 2021.345 1112.930 ;
      LAYER li1 ;
        RECT 2023.420 1112.760 2024.520 1112.960 ;
      LAYER li1 ;
        RECT 2024.700 1112.930 2024.875 1113.130 ;
        RECT 2024.700 1112.760 2027.325 1112.930 ;
      LAYER li1 ;
        RECT 2029.400 1112.760 2030.500 1112.960 ;
      LAYER li1 ;
        RECT 2030.680 1112.930 2030.855 1113.130 ;
        RECT 2030.680 1112.760 2033.305 1112.930 ;
      LAYER li1 ;
        RECT 2035.380 1112.760 2036.480 1112.960 ;
      LAYER li1 ;
        RECT 2036.660 1112.930 2036.835 1113.130 ;
        RECT 2036.660 1112.760 2039.285 1112.930 ;
        RECT 675.065 1111.770 675.355 1112.495 ;
        RECT 675.615 1112.420 677.035 1112.590 ;
      LAYER li1 ;
        RECT 677.295 1112.420 679.985 1112.590 ;
      LAYER li1 ;
        RECT 675.615 1111.940 675.785 1112.420 ;
        RECT 675.955 1111.770 676.285 1112.250 ;
        RECT 676.455 1111.945 676.625 1112.420 ;
        RECT 676.795 1111.770 677.125 1112.250 ;
      LAYER li1 ;
        RECT 677.295 1111.940 677.465 1112.420 ;
      LAYER li1 ;
        RECT 677.635 1111.770 677.965 1112.250 ;
      LAYER li1 ;
        RECT 678.135 1111.940 678.305 1112.420 ;
      LAYER li1 ;
        RECT 678.475 1111.770 678.805 1112.250 ;
      LAYER li1 ;
        RECT 678.975 1111.940 679.145 1112.420 ;
      LAYER li1 ;
        RECT 679.315 1111.770 679.645 1112.250 ;
      LAYER li1 ;
        RECT 679.815 1111.940 679.985 1112.420 ;
      LAYER li1 ;
        RECT 680.155 1111.770 680.485 1112.570 ;
        RECT 681.045 1111.770 681.335 1112.495 ;
        RECT 681.595 1112.420 683.015 1112.590 ;
      LAYER li1 ;
        RECT 683.275 1112.420 685.965 1112.590 ;
      LAYER li1 ;
        RECT 681.595 1111.940 681.765 1112.420 ;
        RECT 681.935 1111.770 682.265 1112.250 ;
        RECT 682.435 1111.945 682.605 1112.420 ;
        RECT 682.775 1111.770 683.105 1112.250 ;
      LAYER li1 ;
        RECT 683.275 1111.940 683.445 1112.420 ;
      LAYER li1 ;
        RECT 683.615 1111.770 683.945 1112.250 ;
      LAYER li1 ;
        RECT 684.115 1111.940 684.285 1112.420 ;
      LAYER li1 ;
        RECT 684.455 1111.770 684.785 1112.250 ;
      LAYER li1 ;
        RECT 684.955 1111.940 685.125 1112.420 ;
      LAYER li1 ;
        RECT 685.295 1111.770 685.625 1112.250 ;
      LAYER li1 ;
        RECT 685.795 1111.940 685.965 1112.420 ;
      LAYER li1 ;
        RECT 686.135 1111.770 686.465 1112.570 ;
        RECT 687.025 1111.770 687.315 1112.495 ;
        RECT 687.575 1112.420 688.995 1112.590 ;
      LAYER li1 ;
        RECT 689.255 1112.420 691.945 1112.590 ;
      LAYER li1 ;
        RECT 687.575 1111.940 687.745 1112.420 ;
        RECT 687.915 1111.770 688.245 1112.250 ;
        RECT 688.415 1111.945 688.585 1112.420 ;
        RECT 688.755 1111.770 689.085 1112.250 ;
      LAYER li1 ;
        RECT 689.255 1111.940 689.425 1112.420 ;
      LAYER li1 ;
        RECT 689.595 1111.770 689.925 1112.250 ;
      LAYER li1 ;
        RECT 690.095 1111.940 690.265 1112.420 ;
      LAYER li1 ;
        RECT 690.435 1111.770 690.765 1112.250 ;
      LAYER li1 ;
        RECT 690.935 1111.940 691.105 1112.420 ;
      LAYER li1 ;
        RECT 691.275 1111.770 691.605 1112.250 ;
      LAYER li1 ;
        RECT 691.775 1111.940 691.945 1112.420 ;
      LAYER li1 ;
        RECT 692.115 1111.770 692.445 1112.570 ;
        RECT 693.005 1111.770 693.295 1112.495 ;
        RECT 693.555 1112.420 694.975 1112.590 ;
      LAYER li1 ;
        RECT 695.235 1112.420 697.925 1112.590 ;
      LAYER li1 ;
        RECT 693.555 1111.940 693.725 1112.420 ;
        RECT 693.895 1111.770 694.225 1112.250 ;
        RECT 694.395 1111.945 694.565 1112.420 ;
        RECT 694.735 1111.770 695.065 1112.250 ;
      LAYER li1 ;
        RECT 695.235 1111.940 695.405 1112.420 ;
      LAYER li1 ;
        RECT 695.575 1111.770 695.905 1112.250 ;
      LAYER li1 ;
        RECT 696.075 1111.940 696.245 1112.420 ;
      LAYER li1 ;
        RECT 696.415 1111.770 696.745 1112.250 ;
      LAYER li1 ;
        RECT 696.915 1111.940 697.085 1112.420 ;
      LAYER li1 ;
        RECT 697.255 1111.770 697.585 1112.250 ;
      LAYER li1 ;
        RECT 697.755 1111.940 697.925 1112.420 ;
      LAYER li1 ;
        RECT 698.095 1111.770 698.425 1112.570 ;
        RECT 698.985 1111.770 699.275 1112.495 ;
        RECT 699.535 1112.420 700.955 1112.590 ;
      LAYER li1 ;
        RECT 701.215 1112.420 703.905 1112.590 ;
      LAYER li1 ;
        RECT 699.535 1111.940 699.705 1112.420 ;
        RECT 699.875 1111.770 700.205 1112.250 ;
        RECT 700.375 1111.945 700.545 1112.420 ;
        RECT 700.715 1111.770 701.045 1112.250 ;
      LAYER li1 ;
        RECT 701.215 1111.940 701.385 1112.420 ;
      LAYER li1 ;
        RECT 701.555 1111.770 701.885 1112.250 ;
      LAYER li1 ;
        RECT 702.055 1111.940 702.225 1112.420 ;
      LAYER li1 ;
        RECT 702.395 1111.770 702.725 1112.250 ;
      LAYER li1 ;
        RECT 702.895 1111.940 703.065 1112.420 ;
      LAYER li1 ;
        RECT 703.235 1111.770 703.565 1112.250 ;
      LAYER li1 ;
        RECT 703.735 1111.940 703.905 1112.420 ;
      LAYER li1 ;
        RECT 704.075 1111.770 704.405 1112.570 ;
        RECT 704.965 1111.770 705.255 1112.495 ;
        RECT 705.515 1112.420 706.935 1112.590 ;
      LAYER li1 ;
        RECT 707.195 1112.420 709.885 1112.590 ;
      LAYER li1 ;
        RECT 705.515 1111.940 705.685 1112.420 ;
        RECT 705.855 1111.770 706.185 1112.250 ;
        RECT 706.355 1111.945 706.525 1112.420 ;
        RECT 706.695 1111.770 707.025 1112.250 ;
      LAYER li1 ;
        RECT 707.195 1111.940 707.365 1112.420 ;
      LAYER li1 ;
        RECT 707.535 1111.770 707.865 1112.250 ;
      LAYER li1 ;
        RECT 708.035 1111.940 708.205 1112.420 ;
      LAYER li1 ;
        RECT 708.375 1111.770 708.705 1112.250 ;
      LAYER li1 ;
        RECT 708.875 1111.940 709.045 1112.420 ;
      LAYER li1 ;
        RECT 709.215 1111.770 709.545 1112.250 ;
      LAYER li1 ;
        RECT 709.715 1111.940 709.885 1112.420 ;
      LAYER li1 ;
        RECT 710.055 1111.770 710.385 1112.570 ;
        RECT 710.945 1111.770 711.235 1112.495 ;
        RECT 711.495 1112.420 712.915 1112.590 ;
      LAYER li1 ;
        RECT 713.175 1112.420 715.865 1112.590 ;
      LAYER li1 ;
        RECT 711.495 1111.940 711.665 1112.420 ;
        RECT 711.835 1111.770 712.165 1112.250 ;
        RECT 712.335 1111.945 712.505 1112.420 ;
        RECT 712.675 1111.770 713.005 1112.250 ;
      LAYER li1 ;
        RECT 713.175 1111.940 713.345 1112.420 ;
      LAYER li1 ;
        RECT 713.515 1111.770 713.845 1112.250 ;
      LAYER li1 ;
        RECT 714.015 1111.940 714.185 1112.420 ;
      LAYER li1 ;
        RECT 714.355 1111.770 714.685 1112.250 ;
      LAYER li1 ;
        RECT 714.855 1111.940 715.025 1112.420 ;
      LAYER li1 ;
        RECT 715.195 1111.770 715.525 1112.250 ;
      LAYER li1 ;
        RECT 715.695 1111.940 715.865 1112.420 ;
      LAYER li1 ;
        RECT 716.035 1111.770 716.365 1112.570 ;
        RECT 716.925 1111.770 717.215 1112.495 ;
        RECT 717.475 1112.420 718.895 1112.590 ;
      LAYER li1 ;
        RECT 719.155 1112.420 721.845 1112.590 ;
      LAYER li1 ;
        RECT 717.475 1111.940 717.645 1112.420 ;
        RECT 717.815 1111.770 718.145 1112.250 ;
        RECT 718.315 1111.945 718.485 1112.420 ;
        RECT 718.655 1111.770 718.985 1112.250 ;
      LAYER li1 ;
        RECT 719.155 1111.940 719.325 1112.420 ;
      LAYER li1 ;
        RECT 719.495 1111.770 719.825 1112.250 ;
      LAYER li1 ;
        RECT 719.995 1111.940 720.165 1112.420 ;
      LAYER li1 ;
        RECT 720.335 1111.770 720.665 1112.250 ;
      LAYER li1 ;
        RECT 720.835 1111.940 721.005 1112.420 ;
      LAYER li1 ;
        RECT 721.175 1111.770 721.505 1112.250 ;
      LAYER li1 ;
        RECT 721.675 1111.940 721.845 1112.420 ;
      LAYER li1 ;
        RECT 722.015 1111.770 722.345 1112.570 ;
        RECT 722.905 1111.770 723.195 1112.495 ;
        RECT 723.455 1112.420 724.875 1112.590 ;
      LAYER li1 ;
        RECT 725.135 1112.420 727.825 1112.590 ;
      LAYER li1 ;
        RECT 723.455 1111.940 723.625 1112.420 ;
        RECT 723.795 1111.770 724.125 1112.250 ;
        RECT 724.295 1111.945 724.465 1112.420 ;
        RECT 724.635 1111.770 724.965 1112.250 ;
      LAYER li1 ;
        RECT 725.135 1111.940 725.305 1112.420 ;
      LAYER li1 ;
        RECT 725.475 1111.770 725.805 1112.250 ;
      LAYER li1 ;
        RECT 725.975 1111.940 726.145 1112.420 ;
      LAYER li1 ;
        RECT 726.315 1111.770 726.645 1112.250 ;
      LAYER li1 ;
        RECT 726.815 1111.940 726.985 1112.420 ;
      LAYER li1 ;
        RECT 727.155 1111.770 727.485 1112.250 ;
      LAYER li1 ;
        RECT 727.655 1111.940 727.825 1112.420 ;
      LAYER li1 ;
        RECT 727.995 1111.770 728.325 1112.570 ;
        RECT 728.885 1111.770 729.175 1112.495 ;
        RECT 729.435 1112.420 730.855 1112.590 ;
      LAYER li1 ;
        RECT 731.115 1112.420 733.805 1112.590 ;
      LAYER li1 ;
        RECT 729.435 1111.940 729.605 1112.420 ;
        RECT 729.775 1111.770 730.105 1112.250 ;
        RECT 730.275 1111.945 730.445 1112.420 ;
        RECT 730.615 1111.770 730.945 1112.250 ;
      LAYER li1 ;
        RECT 731.115 1111.940 731.285 1112.420 ;
      LAYER li1 ;
        RECT 731.455 1111.770 731.785 1112.250 ;
      LAYER li1 ;
        RECT 731.955 1111.940 732.125 1112.420 ;
      LAYER li1 ;
        RECT 732.295 1111.770 732.625 1112.250 ;
      LAYER li1 ;
        RECT 732.795 1111.940 732.965 1112.420 ;
      LAYER li1 ;
        RECT 733.135 1111.770 733.465 1112.250 ;
      LAYER li1 ;
        RECT 733.635 1111.940 733.805 1112.420 ;
      LAYER li1 ;
        RECT 733.975 1111.770 734.305 1112.570 ;
        RECT 734.865 1111.770 735.155 1112.495 ;
        RECT 735.415 1112.420 736.835 1112.590 ;
      LAYER li1 ;
        RECT 737.095 1112.420 739.785 1112.590 ;
      LAYER li1 ;
        RECT 735.415 1111.940 735.585 1112.420 ;
        RECT 735.755 1111.770 736.085 1112.250 ;
        RECT 736.255 1111.945 736.425 1112.420 ;
        RECT 736.595 1111.770 736.925 1112.250 ;
      LAYER li1 ;
        RECT 737.095 1111.940 737.265 1112.420 ;
      LAYER li1 ;
        RECT 737.435 1111.770 737.765 1112.250 ;
      LAYER li1 ;
        RECT 737.935 1111.940 738.105 1112.420 ;
      LAYER li1 ;
        RECT 738.275 1111.770 738.605 1112.250 ;
      LAYER li1 ;
        RECT 738.775 1111.940 738.945 1112.420 ;
      LAYER li1 ;
        RECT 739.115 1111.770 739.445 1112.250 ;
      LAYER li1 ;
        RECT 739.615 1111.940 739.785 1112.420 ;
      LAYER li1 ;
        RECT 739.955 1111.770 740.285 1112.570 ;
        RECT 740.845 1111.770 741.135 1112.495 ;
        RECT 741.395 1112.420 742.815 1112.590 ;
      LAYER li1 ;
        RECT 743.075 1112.420 745.765 1112.590 ;
      LAYER li1 ;
        RECT 741.395 1111.940 741.565 1112.420 ;
        RECT 741.735 1111.770 742.065 1112.250 ;
        RECT 742.235 1111.945 742.405 1112.420 ;
        RECT 742.575 1111.770 742.905 1112.250 ;
      LAYER li1 ;
        RECT 743.075 1111.940 743.245 1112.420 ;
      LAYER li1 ;
        RECT 743.415 1111.770 743.745 1112.250 ;
      LAYER li1 ;
        RECT 743.915 1111.940 744.085 1112.420 ;
      LAYER li1 ;
        RECT 744.255 1111.770 744.585 1112.250 ;
      LAYER li1 ;
        RECT 744.755 1111.940 744.925 1112.420 ;
      LAYER li1 ;
        RECT 745.095 1111.770 745.425 1112.250 ;
      LAYER li1 ;
        RECT 745.595 1111.940 745.765 1112.420 ;
      LAYER li1 ;
        RECT 745.935 1111.770 746.265 1112.570 ;
        RECT 746.825 1111.770 747.115 1112.495 ;
        RECT 747.375 1112.420 748.795 1112.590 ;
      LAYER li1 ;
        RECT 749.055 1112.420 751.745 1112.590 ;
      LAYER li1 ;
        RECT 747.375 1111.940 747.545 1112.420 ;
        RECT 747.715 1111.770 748.045 1112.250 ;
        RECT 748.215 1111.945 748.385 1112.420 ;
        RECT 748.555 1111.770 748.885 1112.250 ;
      LAYER li1 ;
        RECT 749.055 1111.940 749.225 1112.420 ;
      LAYER li1 ;
        RECT 749.395 1111.770 749.725 1112.250 ;
      LAYER li1 ;
        RECT 749.895 1111.940 750.065 1112.420 ;
      LAYER li1 ;
        RECT 750.235 1111.770 750.565 1112.250 ;
      LAYER li1 ;
        RECT 750.735 1111.940 750.905 1112.420 ;
      LAYER li1 ;
        RECT 751.075 1111.770 751.405 1112.250 ;
      LAYER li1 ;
        RECT 751.575 1111.940 751.745 1112.420 ;
      LAYER li1 ;
        RECT 751.915 1111.770 752.245 1112.570 ;
        RECT 752.805 1111.770 753.095 1112.495 ;
        RECT 753.355 1112.420 754.775 1112.590 ;
      LAYER li1 ;
        RECT 755.035 1112.420 757.725 1112.590 ;
      LAYER li1 ;
        RECT 753.355 1111.940 753.525 1112.420 ;
        RECT 753.695 1111.770 754.025 1112.250 ;
        RECT 754.195 1111.945 754.365 1112.420 ;
        RECT 754.535 1111.770 754.865 1112.250 ;
      LAYER li1 ;
        RECT 755.035 1111.940 755.205 1112.420 ;
      LAYER li1 ;
        RECT 755.375 1111.770 755.705 1112.250 ;
      LAYER li1 ;
        RECT 755.875 1111.940 756.045 1112.420 ;
      LAYER li1 ;
        RECT 756.215 1111.770 756.545 1112.250 ;
      LAYER li1 ;
        RECT 756.715 1111.940 756.885 1112.420 ;
      LAYER li1 ;
        RECT 757.055 1111.770 757.385 1112.250 ;
      LAYER li1 ;
        RECT 757.555 1111.940 757.725 1112.420 ;
      LAYER li1 ;
        RECT 757.895 1111.770 758.225 1112.570 ;
        RECT 758.785 1111.770 759.075 1112.495 ;
        RECT 759.335 1112.420 760.755 1112.590 ;
      LAYER li1 ;
        RECT 761.015 1112.420 763.705 1112.590 ;
      LAYER li1 ;
        RECT 769.065 1112.590 769.240 1112.760 ;
        RECT 1976.860 1112.590 1977.035 1112.760 ;
        RECT 1982.840 1112.590 1983.015 1112.760 ;
        RECT 1988.820 1112.590 1988.995 1112.760 ;
        RECT 1994.800 1112.590 1994.975 1112.760 ;
        RECT 2000.780 1112.590 2000.955 1112.760 ;
        RECT 2006.760 1112.590 2006.935 1112.760 ;
        RECT 2012.740 1112.590 2012.915 1112.760 ;
        RECT 2018.720 1112.590 2018.895 1112.760 ;
        RECT 2024.700 1112.590 2024.875 1112.760 ;
        RECT 2030.680 1112.590 2030.855 1112.760 ;
        RECT 2036.660 1112.590 2036.835 1112.760 ;
      LAYER li1 ;
        RECT 2039.530 1112.590 2039.785 1113.130 ;
        RECT 2041.360 1112.760 2042.460 1112.960 ;
      LAYER li1 ;
        RECT 2042.640 1112.930 2042.815 1113.130 ;
        RECT 2042.640 1112.760 2045.265 1112.930 ;
      LAYER li1 ;
        RECT 2047.340 1112.760 2048.440 1112.960 ;
      LAYER li1 ;
        RECT 2048.620 1112.930 2048.795 1113.130 ;
        RECT 2048.620 1112.760 2051.245 1112.930 ;
      LAYER li1 ;
        RECT 2053.320 1112.760 2054.420 1112.960 ;
      LAYER li1 ;
        RECT 2054.600 1112.930 2054.775 1113.130 ;
        RECT 2054.600 1112.760 2057.225 1112.930 ;
      LAYER li1 ;
        RECT 2059.300 1112.760 2060.400 1112.960 ;
      LAYER li1 ;
        RECT 2060.580 1112.930 2060.755 1113.130 ;
      LAYER li1 ;
        RECT 2066.115 1113.130 2068.805 1113.300 ;
      LAYER li1 ;
        RECT 2069.065 1113.130 2070.565 1113.300 ;
        RECT 2070.745 1113.155 2071.035 1114.320 ;
        RECT 2060.580 1112.760 2063.205 1112.930 ;
        RECT 2042.640 1112.590 2042.815 1112.760 ;
        RECT 2048.620 1112.590 2048.795 1112.760 ;
        RECT 2054.600 1112.590 2054.775 1112.760 ;
        RECT 2060.580 1112.590 2060.755 1112.760 ;
        RECT 759.335 1111.940 759.505 1112.420 ;
        RECT 759.675 1111.770 760.005 1112.250 ;
        RECT 760.175 1111.945 760.345 1112.420 ;
        RECT 760.515 1111.770 760.845 1112.250 ;
      LAYER li1 ;
        RECT 761.015 1111.940 761.185 1112.420 ;
      LAYER li1 ;
        RECT 761.355 1111.770 761.685 1112.250 ;
      LAYER li1 ;
        RECT 761.855 1111.940 762.025 1112.420 ;
      LAYER li1 ;
        RECT 762.195 1111.770 762.525 1112.250 ;
      LAYER li1 ;
        RECT 762.695 1111.940 762.865 1112.420 ;
      LAYER li1 ;
        RECT 763.035 1111.770 763.365 1112.250 ;
      LAYER li1 ;
        RECT 763.535 1111.940 763.705 1112.420 ;
      LAYER li1 ;
        RECT 763.875 1111.770 764.205 1112.570 ;
        RECT 764.765 1111.770 765.055 1112.495 ;
        RECT 765.615 1111.770 765.945 1112.570 ;
        RECT 769.065 1112.420 770.485 1112.590 ;
        RECT 766.455 1111.770 766.785 1112.250 ;
        RECT 767.295 1111.770 767.625 1112.250 ;
        RECT 768.135 1111.770 768.465 1112.250 ;
        RECT 768.975 1111.770 769.305 1112.250 ;
        RECT 769.475 1111.945 769.645 1112.420 ;
        RECT 769.815 1111.770 770.145 1112.250 ;
        RECT 770.315 1111.940 770.485 1112.420 ;
        RECT 770.745 1111.770 771.035 1112.495 ;
        RECT 1975.065 1111.770 1975.355 1112.495 ;
        RECT 1975.615 1112.420 1977.035 1112.590 ;
        RECT 1975.615 1111.940 1975.785 1112.420 ;
        RECT 1975.955 1111.770 1976.285 1112.250 ;
        RECT 1976.455 1111.945 1976.625 1112.420 ;
        RECT 1976.795 1111.770 1977.125 1112.250 ;
        RECT 1977.635 1111.770 1977.965 1112.250 ;
        RECT 1978.475 1111.770 1978.805 1112.250 ;
        RECT 1979.315 1111.770 1979.645 1112.250 ;
        RECT 1980.155 1111.770 1980.485 1112.570 ;
        RECT 1981.045 1111.770 1981.335 1112.495 ;
        RECT 1981.595 1112.420 1983.015 1112.590 ;
        RECT 1981.595 1111.940 1981.765 1112.420 ;
        RECT 1981.935 1111.770 1982.265 1112.250 ;
        RECT 1982.435 1111.945 1982.605 1112.420 ;
        RECT 1982.775 1111.770 1983.105 1112.250 ;
        RECT 1983.615 1111.770 1983.945 1112.250 ;
        RECT 1984.455 1111.770 1984.785 1112.250 ;
        RECT 1985.295 1111.770 1985.625 1112.250 ;
        RECT 1986.135 1111.770 1986.465 1112.570 ;
        RECT 1987.025 1111.770 1987.315 1112.495 ;
        RECT 1987.575 1112.420 1988.995 1112.590 ;
        RECT 1987.575 1111.940 1987.745 1112.420 ;
        RECT 1987.915 1111.770 1988.245 1112.250 ;
        RECT 1988.415 1111.945 1988.585 1112.420 ;
        RECT 1988.755 1111.770 1989.085 1112.250 ;
        RECT 1989.595 1111.770 1989.925 1112.250 ;
        RECT 1990.435 1111.770 1990.765 1112.250 ;
        RECT 1991.275 1111.770 1991.605 1112.250 ;
        RECT 1992.115 1111.770 1992.445 1112.570 ;
        RECT 1993.005 1111.770 1993.295 1112.495 ;
        RECT 1993.555 1112.420 1994.975 1112.590 ;
        RECT 1993.555 1111.940 1993.725 1112.420 ;
        RECT 1993.895 1111.770 1994.225 1112.250 ;
        RECT 1994.395 1111.945 1994.565 1112.420 ;
        RECT 1994.735 1111.770 1995.065 1112.250 ;
        RECT 1995.575 1111.770 1995.905 1112.250 ;
        RECT 1996.415 1111.770 1996.745 1112.250 ;
        RECT 1997.255 1111.770 1997.585 1112.250 ;
        RECT 1998.095 1111.770 1998.425 1112.570 ;
        RECT 1998.985 1111.770 1999.275 1112.495 ;
        RECT 1999.535 1112.420 2000.955 1112.590 ;
        RECT 1999.535 1111.940 1999.705 1112.420 ;
        RECT 1999.875 1111.770 2000.205 1112.250 ;
        RECT 2000.375 1111.945 2000.545 1112.420 ;
        RECT 2000.715 1111.770 2001.045 1112.250 ;
        RECT 2001.555 1111.770 2001.885 1112.250 ;
        RECT 2002.395 1111.770 2002.725 1112.250 ;
        RECT 2003.235 1111.770 2003.565 1112.250 ;
        RECT 2004.075 1111.770 2004.405 1112.570 ;
        RECT 2004.965 1111.770 2005.255 1112.495 ;
        RECT 2005.515 1112.420 2006.935 1112.590 ;
        RECT 2005.515 1111.940 2005.685 1112.420 ;
        RECT 2005.855 1111.770 2006.185 1112.250 ;
        RECT 2006.355 1111.945 2006.525 1112.420 ;
        RECT 2006.695 1111.770 2007.025 1112.250 ;
        RECT 2007.535 1111.770 2007.865 1112.250 ;
        RECT 2008.375 1111.770 2008.705 1112.250 ;
        RECT 2009.215 1111.770 2009.545 1112.250 ;
        RECT 2010.055 1111.770 2010.385 1112.570 ;
        RECT 2010.945 1111.770 2011.235 1112.495 ;
        RECT 2011.495 1112.420 2012.915 1112.590 ;
        RECT 2011.495 1111.940 2011.665 1112.420 ;
        RECT 2011.835 1111.770 2012.165 1112.250 ;
        RECT 2012.335 1111.945 2012.505 1112.420 ;
        RECT 2012.675 1111.770 2013.005 1112.250 ;
        RECT 2013.515 1111.770 2013.845 1112.250 ;
        RECT 2014.355 1111.770 2014.685 1112.250 ;
        RECT 2015.195 1111.770 2015.525 1112.250 ;
        RECT 2016.035 1111.770 2016.365 1112.570 ;
        RECT 2016.925 1111.770 2017.215 1112.495 ;
        RECT 2017.475 1112.420 2018.895 1112.590 ;
        RECT 2017.475 1111.940 2017.645 1112.420 ;
        RECT 2017.815 1111.770 2018.145 1112.250 ;
        RECT 2018.315 1111.945 2018.485 1112.420 ;
        RECT 2018.655 1111.770 2018.985 1112.250 ;
        RECT 2019.495 1111.770 2019.825 1112.250 ;
        RECT 2020.335 1111.770 2020.665 1112.250 ;
        RECT 2021.175 1111.770 2021.505 1112.250 ;
        RECT 2022.015 1111.770 2022.345 1112.570 ;
        RECT 2022.905 1111.770 2023.195 1112.495 ;
        RECT 2023.455 1112.420 2024.875 1112.590 ;
        RECT 2023.455 1111.940 2023.625 1112.420 ;
        RECT 2023.795 1111.770 2024.125 1112.250 ;
        RECT 2024.295 1111.945 2024.465 1112.420 ;
        RECT 2024.635 1111.770 2024.965 1112.250 ;
        RECT 2025.475 1111.770 2025.805 1112.250 ;
        RECT 2026.315 1111.770 2026.645 1112.250 ;
        RECT 2027.155 1111.770 2027.485 1112.250 ;
        RECT 2027.995 1111.770 2028.325 1112.570 ;
        RECT 2028.885 1111.770 2029.175 1112.495 ;
        RECT 2029.435 1112.420 2030.855 1112.590 ;
        RECT 2029.435 1111.940 2029.605 1112.420 ;
        RECT 2029.775 1111.770 2030.105 1112.250 ;
        RECT 2030.275 1111.945 2030.445 1112.420 ;
        RECT 2030.615 1111.770 2030.945 1112.250 ;
        RECT 2031.455 1111.770 2031.785 1112.250 ;
        RECT 2032.295 1111.770 2032.625 1112.250 ;
        RECT 2033.135 1111.770 2033.465 1112.250 ;
        RECT 2033.975 1111.770 2034.305 1112.570 ;
        RECT 2034.865 1111.770 2035.155 1112.495 ;
        RECT 2035.415 1112.420 2036.835 1112.590 ;
      LAYER li1 ;
        RECT 2037.095 1112.420 2039.785 1112.590 ;
      LAYER li1 ;
        RECT 2035.415 1111.940 2035.585 1112.420 ;
        RECT 2035.755 1111.770 2036.085 1112.250 ;
        RECT 2036.255 1111.945 2036.425 1112.420 ;
        RECT 2036.595 1111.770 2036.925 1112.250 ;
      LAYER li1 ;
        RECT 2037.095 1111.940 2037.265 1112.420 ;
      LAYER li1 ;
        RECT 2037.435 1111.770 2037.765 1112.250 ;
      LAYER li1 ;
        RECT 2037.935 1111.940 2038.105 1112.420 ;
      LAYER li1 ;
        RECT 2038.275 1111.770 2038.605 1112.250 ;
      LAYER li1 ;
        RECT 2038.775 1111.940 2038.945 1112.420 ;
      LAYER li1 ;
        RECT 2039.115 1111.770 2039.445 1112.250 ;
      LAYER li1 ;
        RECT 2039.615 1111.940 2039.785 1112.420 ;
      LAYER li1 ;
        RECT 2039.955 1111.770 2040.285 1112.570 ;
        RECT 2040.845 1111.770 2041.135 1112.495 ;
        RECT 2041.395 1112.420 2042.815 1112.590 ;
        RECT 2041.395 1111.940 2041.565 1112.420 ;
        RECT 2041.735 1111.770 2042.065 1112.250 ;
        RECT 2042.235 1111.945 2042.405 1112.420 ;
        RECT 2042.575 1111.770 2042.905 1112.250 ;
        RECT 2043.415 1111.770 2043.745 1112.250 ;
        RECT 2044.255 1111.770 2044.585 1112.250 ;
        RECT 2045.095 1111.770 2045.425 1112.250 ;
        RECT 2045.935 1111.770 2046.265 1112.570 ;
        RECT 2046.825 1111.770 2047.115 1112.495 ;
        RECT 2047.375 1112.420 2048.795 1112.590 ;
        RECT 2047.375 1111.940 2047.545 1112.420 ;
        RECT 2047.715 1111.770 2048.045 1112.250 ;
        RECT 2048.215 1111.945 2048.385 1112.420 ;
        RECT 2048.555 1111.770 2048.885 1112.250 ;
        RECT 2049.395 1111.770 2049.725 1112.250 ;
        RECT 2050.235 1111.770 2050.565 1112.250 ;
        RECT 2051.075 1111.770 2051.405 1112.250 ;
        RECT 2051.915 1111.770 2052.245 1112.570 ;
        RECT 2052.805 1111.770 2053.095 1112.495 ;
        RECT 2053.355 1112.420 2054.775 1112.590 ;
        RECT 2053.355 1111.940 2053.525 1112.420 ;
        RECT 2053.695 1111.770 2054.025 1112.250 ;
        RECT 2054.195 1111.945 2054.365 1112.420 ;
        RECT 2054.535 1111.770 2054.865 1112.250 ;
        RECT 2055.375 1111.770 2055.705 1112.250 ;
        RECT 2056.215 1111.770 2056.545 1112.250 ;
        RECT 2057.055 1111.770 2057.385 1112.250 ;
        RECT 2057.895 1111.770 2058.225 1112.570 ;
        RECT 2058.785 1111.770 2059.075 1112.495 ;
        RECT 2059.335 1112.420 2060.755 1112.590 ;
      LAYER li1 ;
        RECT 2066.115 1112.590 2066.370 1113.130 ;
      LAYER li1 ;
        RECT 2069.065 1112.930 2069.240 1113.130 ;
        RECT 2066.615 1112.760 2069.240 1112.930 ;
        RECT 2069.065 1112.590 2069.240 1112.760 ;
        RECT 2059.335 1111.940 2059.505 1112.420 ;
        RECT 2059.675 1111.770 2060.005 1112.250 ;
        RECT 2060.175 1111.945 2060.345 1112.420 ;
        RECT 2060.515 1111.770 2060.845 1112.250 ;
        RECT 2061.355 1111.770 2061.685 1112.250 ;
        RECT 2062.195 1111.770 2062.525 1112.250 ;
        RECT 2063.035 1111.770 2063.365 1112.250 ;
        RECT 2063.875 1111.770 2064.205 1112.570 ;
        RECT 2064.765 1111.770 2065.055 1112.495 ;
        RECT 2065.615 1111.770 2065.945 1112.570 ;
      LAYER li1 ;
        RECT 2066.115 1112.420 2068.805 1112.590 ;
      LAYER li1 ;
        RECT 2069.065 1112.420 2070.485 1112.590 ;
      LAYER li1 ;
        RECT 2066.115 1111.940 2066.285 1112.420 ;
      LAYER li1 ;
        RECT 2066.455 1111.770 2066.785 1112.250 ;
      LAYER li1 ;
        RECT 2066.955 1111.940 2067.125 1112.420 ;
      LAYER li1 ;
        RECT 2067.295 1111.770 2067.625 1112.250 ;
      LAYER li1 ;
        RECT 2067.795 1111.940 2067.965 1112.420 ;
      LAYER li1 ;
        RECT 2068.135 1111.770 2068.465 1112.250 ;
      LAYER li1 ;
        RECT 2068.635 1111.940 2068.805 1112.420 ;
      LAYER li1 ;
        RECT 2068.975 1111.770 2069.305 1112.250 ;
        RECT 2069.475 1111.945 2069.645 1112.420 ;
        RECT 2069.815 1111.770 2070.145 1112.250 ;
        RECT 2070.315 1111.940 2070.485 1112.420 ;
        RECT 2070.745 1111.770 2071.035 1112.495 ;
        RECT 674.980 1111.600 675.125 1111.770 ;
        RECT 675.295 1111.600 675.585 1111.770 ;
        RECT 675.755 1111.600 676.045 1111.770 ;
        RECT 676.215 1111.600 676.505 1111.770 ;
        RECT 676.675 1111.600 676.965 1111.770 ;
        RECT 677.135 1111.600 677.425 1111.770 ;
        RECT 677.595 1111.600 677.885 1111.770 ;
        RECT 678.055 1111.600 678.345 1111.770 ;
        RECT 678.515 1111.600 678.805 1111.770 ;
        RECT 678.975 1111.600 679.265 1111.770 ;
        RECT 679.435 1111.600 679.725 1111.770 ;
        RECT 679.895 1111.600 680.185 1111.770 ;
        RECT 680.355 1111.600 680.645 1111.770 ;
        RECT 680.815 1111.600 681.105 1111.770 ;
        RECT 681.275 1111.600 681.565 1111.770 ;
        RECT 681.735 1111.600 682.025 1111.770 ;
        RECT 682.195 1111.600 682.485 1111.770 ;
        RECT 682.655 1111.600 682.945 1111.770 ;
        RECT 683.115 1111.600 683.405 1111.770 ;
        RECT 683.575 1111.600 683.865 1111.770 ;
        RECT 684.035 1111.600 684.325 1111.770 ;
        RECT 684.495 1111.600 684.785 1111.770 ;
        RECT 684.955 1111.600 685.245 1111.770 ;
        RECT 685.415 1111.600 685.705 1111.770 ;
        RECT 685.875 1111.600 686.165 1111.770 ;
        RECT 686.335 1111.600 686.625 1111.770 ;
        RECT 686.795 1111.600 687.085 1111.770 ;
        RECT 687.255 1111.600 687.545 1111.770 ;
        RECT 687.715 1111.600 688.005 1111.770 ;
        RECT 688.175 1111.600 688.465 1111.770 ;
        RECT 688.635 1111.600 688.925 1111.770 ;
        RECT 689.095 1111.600 689.385 1111.770 ;
        RECT 689.555 1111.600 689.845 1111.770 ;
        RECT 690.015 1111.600 690.305 1111.770 ;
        RECT 690.475 1111.600 690.765 1111.770 ;
        RECT 690.935 1111.600 691.225 1111.770 ;
        RECT 691.395 1111.600 691.685 1111.770 ;
        RECT 691.855 1111.600 692.145 1111.770 ;
        RECT 692.315 1111.600 692.605 1111.770 ;
        RECT 692.775 1111.600 693.065 1111.770 ;
        RECT 693.235 1111.600 693.525 1111.770 ;
        RECT 693.695 1111.600 693.985 1111.770 ;
        RECT 694.155 1111.600 694.445 1111.770 ;
        RECT 694.615 1111.600 694.905 1111.770 ;
        RECT 695.075 1111.600 695.365 1111.770 ;
        RECT 695.535 1111.600 695.825 1111.770 ;
        RECT 695.995 1111.600 696.285 1111.770 ;
        RECT 696.455 1111.600 696.745 1111.770 ;
        RECT 696.915 1111.600 697.205 1111.770 ;
        RECT 697.375 1111.600 697.665 1111.770 ;
        RECT 697.835 1111.600 698.125 1111.770 ;
        RECT 698.295 1111.600 698.585 1111.770 ;
        RECT 698.755 1111.600 699.045 1111.770 ;
        RECT 699.215 1111.600 699.505 1111.770 ;
        RECT 699.675 1111.600 699.965 1111.770 ;
        RECT 700.135 1111.600 700.425 1111.770 ;
        RECT 700.595 1111.600 700.885 1111.770 ;
        RECT 701.055 1111.600 701.345 1111.770 ;
        RECT 701.515 1111.600 701.805 1111.770 ;
        RECT 701.975 1111.600 702.265 1111.770 ;
        RECT 702.435 1111.600 702.725 1111.770 ;
        RECT 702.895 1111.600 703.185 1111.770 ;
        RECT 703.355 1111.600 703.645 1111.770 ;
        RECT 703.815 1111.600 704.105 1111.770 ;
        RECT 704.275 1111.600 704.565 1111.770 ;
        RECT 704.735 1111.600 705.025 1111.770 ;
        RECT 705.195 1111.600 705.485 1111.770 ;
        RECT 705.655 1111.600 705.945 1111.770 ;
        RECT 706.115 1111.600 706.405 1111.770 ;
        RECT 706.575 1111.600 706.865 1111.770 ;
        RECT 707.035 1111.600 707.325 1111.770 ;
        RECT 707.495 1111.600 707.785 1111.770 ;
        RECT 707.955 1111.600 708.245 1111.770 ;
        RECT 708.415 1111.600 708.705 1111.770 ;
        RECT 708.875 1111.600 709.165 1111.770 ;
        RECT 709.335 1111.600 709.625 1111.770 ;
        RECT 709.795 1111.600 710.085 1111.770 ;
        RECT 710.255 1111.600 710.545 1111.770 ;
        RECT 710.715 1111.600 711.005 1111.770 ;
        RECT 711.175 1111.600 711.465 1111.770 ;
        RECT 711.635 1111.600 711.925 1111.770 ;
        RECT 712.095 1111.600 712.385 1111.770 ;
        RECT 712.555 1111.600 712.845 1111.770 ;
        RECT 713.015 1111.600 713.305 1111.770 ;
        RECT 713.475 1111.600 713.765 1111.770 ;
        RECT 713.935 1111.600 714.225 1111.770 ;
        RECT 714.395 1111.600 714.685 1111.770 ;
        RECT 714.855 1111.600 715.145 1111.770 ;
        RECT 715.315 1111.600 715.605 1111.770 ;
        RECT 715.775 1111.600 716.065 1111.770 ;
        RECT 716.235 1111.600 716.525 1111.770 ;
        RECT 716.695 1111.600 716.985 1111.770 ;
        RECT 717.155 1111.600 717.445 1111.770 ;
        RECT 717.615 1111.600 717.905 1111.770 ;
        RECT 718.075 1111.600 718.365 1111.770 ;
        RECT 718.535 1111.600 718.825 1111.770 ;
        RECT 718.995 1111.600 719.285 1111.770 ;
        RECT 719.455 1111.600 719.745 1111.770 ;
        RECT 719.915 1111.600 720.205 1111.770 ;
        RECT 720.375 1111.600 720.665 1111.770 ;
        RECT 720.835 1111.600 721.125 1111.770 ;
        RECT 721.295 1111.600 721.585 1111.770 ;
        RECT 721.755 1111.600 722.045 1111.770 ;
        RECT 722.215 1111.600 722.505 1111.770 ;
        RECT 722.675 1111.600 722.965 1111.770 ;
        RECT 723.135 1111.600 723.425 1111.770 ;
        RECT 723.595 1111.600 723.885 1111.770 ;
        RECT 724.055 1111.600 724.345 1111.770 ;
        RECT 724.515 1111.600 724.805 1111.770 ;
        RECT 724.975 1111.600 725.265 1111.770 ;
        RECT 725.435 1111.600 725.725 1111.770 ;
        RECT 725.895 1111.600 726.185 1111.770 ;
        RECT 726.355 1111.600 726.645 1111.770 ;
        RECT 726.815 1111.600 727.105 1111.770 ;
        RECT 727.275 1111.600 727.565 1111.770 ;
        RECT 727.735 1111.600 728.025 1111.770 ;
        RECT 728.195 1111.600 728.485 1111.770 ;
        RECT 728.655 1111.600 728.945 1111.770 ;
        RECT 729.115 1111.600 729.405 1111.770 ;
        RECT 729.575 1111.600 729.865 1111.770 ;
        RECT 730.035 1111.600 730.325 1111.770 ;
        RECT 730.495 1111.600 730.785 1111.770 ;
        RECT 730.955 1111.600 731.245 1111.770 ;
        RECT 731.415 1111.600 731.705 1111.770 ;
        RECT 731.875 1111.600 732.165 1111.770 ;
        RECT 732.335 1111.600 732.625 1111.770 ;
        RECT 732.795 1111.600 733.085 1111.770 ;
        RECT 733.255 1111.600 733.545 1111.770 ;
        RECT 733.715 1111.600 734.005 1111.770 ;
        RECT 734.175 1111.600 734.465 1111.770 ;
        RECT 734.635 1111.600 734.925 1111.770 ;
        RECT 735.095 1111.600 735.385 1111.770 ;
        RECT 735.555 1111.600 735.845 1111.770 ;
        RECT 736.015 1111.600 736.305 1111.770 ;
        RECT 736.475 1111.600 736.765 1111.770 ;
        RECT 736.935 1111.600 737.225 1111.770 ;
        RECT 737.395 1111.600 737.685 1111.770 ;
        RECT 737.855 1111.600 738.145 1111.770 ;
        RECT 738.315 1111.600 738.605 1111.770 ;
        RECT 738.775 1111.600 739.065 1111.770 ;
        RECT 739.235 1111.600 739.525 1111.770 ;
        RECT 739.695 1111.600 739.985 1111.770 ;
        RECT 740.155 1111.600 740.445 1111.770 ;
        RECT 740.615 1111.600 740.905 1111.770 ;
        RECT 741.075 1111.600 741.365 1111.770 ;
        RECT 741.535 1111.600 741.825 1111.770 ;
        RECT 741.995 1111.600 742.285 1111.770 ;
        RECT 742.455 1111.600 742.745 1111.770 ;
        RECT 742.915 1111.600 743.205 1111.770 ;
        RECT 743.375 1111.600 743.665 1111.770 ;
        RECT 743.835 1111.600 744.125 1111.770 ;
        RECT 744.295 1111.600 744.585 1111.770 ;
        RECT 744.755 1111.600 745.045 1111.770 ;
        RECT 745.215 1111.600 745.505 1111.770 ;
        RECT 745.675 1111.600 745.965 1111.770 ;
        RECT 746.135 1111.600 746.425 1111.770 ;
        RECT 746.595 1111.600 746.885 1111.770 ;
        RECT 747.055 1111.600 747.345 1111.770 ;
        RECT 747.515 1111.600 747.805 1111.770 ;
        RECT 747.975 1111.600 748.265 1111.770 ;
        RECT 748.435 1111.600 748.725 1111.770 ;
        RECT 748.895 1111.600 749.185 1111.770 ;
        RECT 749.355 1111.600 749.645 1111.770 ;
        RECT 749.815 1111.600 750.105 1111.770 ;
        RECT 750.275 1111.600 750.565 1111.770 ;
        RECT 750.735 1111.600 751.025 1111.770 ;
        RECT 751.195 1111.600 751.485 1111.770 ;
        RECT 751.655 1111.600 751.945 1111.770 ;
        RECT 752.115 1111.600 752.405 1111.770 ;
        RECT 752.575 1111.600 752.865 1111.770 ;
        RECT 753.035 1111.600 753.325 1111.770 ;
        RECT 753.495 1111.600 753.785 1111.770 ;
        RECT 753.955 1111.600 754.245 1111.770 ;
        RECT 754.415 1111.600 754.705 1111.770 ;
        RECT 754.875 1111.600 755.165 1111.770 ;
        RECT 755.335 1111.600 755.625 1111.770 ;
        RECT 755.795 1111.600 756.085 1111.770 ;
        RECT 756.255 1111.600 756.545 1111.770 ;
        RECT 756.715 1111.600 757.005 1111.770 ;
        RECT 757.175 1111.600 757.465 1111.770 ;
        RECT 757.635 1111.600 757.925 1111.770 ;
        RECT 758.095 1111.600 758.385 1111.770 ;
        RECT 758.555 1111.600 758.845 1111.770 ;
        RECT 759.015 1111.600 759.305 1111.770 ;
        RECT 759.475 1111.600 759.765 1111.770 ;
        RECT 759.935 1111.600 760.225 1111.770 ;
        RECT 760.395 1111.600 760.685 1111.770 ;
        RECT 760.855 1111.600 761.145 1111.770 ;
        RECT 761.315 1111.600 761.605 1111.770 ;
        RECT 761.775 1111.600 762.065 1111.770 ;
        RECT 762.235 1111.600 762.525 1111.770 ;
        RECT 762.695 1111.600 762.985 1111.770 ;
        RECT 763.155 1111.600 763.445 1111.770 ;
        RECT 763.615 1111.600 763.905 1111.770 ;
        RECT 764.075 1111.600 764.365 1111.770 ;
        RECT 764.535 1111.600 764.825 1111.770 ;
        RECT 764.995 1111.600 765.285 1111.770 ;
        RECT 765.455 1111.600 765.745 1111.770 ;
        RECT 765.915 1111.600 766.205 1111.770 ;
        RECT 766.375 1111.600 766.665 1111.770 ;
        RECT 766.835 1111.600 767.125 1111.770 ;
        RECT 767.295 1111.600 767.585 1111.770 ;
        RECT 767.755 1111.600 768.045 1111.770 ;
        RECT 768.215 1111.600 768.505 1111.770 ;
        RECT 768.675 1111.600 768.965 1111.770 ;
        RECT 769.135 1111.600 769.425 1111.770 ;
        RECT 769.595 1111.600 769.885 1111.770 ;
        RECT 770.055 1111.600 770.345 1111.770 ;
        RECT 770.515 1111.600 770.805 1111.770 ;
        RECT 770.975 1111.600 771.120 1111.770 ;
        RECT 1974.980 1111.600 1975.125 1111.770 ;
        RECT 1975.295 1111.600 1975.585 1111.770 ;
        RECT 1975.755 1111.600 1976.045 1111.770 ;
        RECT 1976.215 1111.600 1976.505 1111.770 ;
        RECT 1976.675 1111.600 1976.965 1111.770 ;
        RECT 1977.135 1111.600 1977.425 1111.770 ;
        RECT 1977.595 1111.600 1977.885 1111.770 ;
        RECT 1978.055 1111.600 1978.345 1111.770 ;
        RECT 1978.515 1111.600 1978.805 1111.770 ;
        RECT 1978.975 1111.600 1979.265 1111.770 ;
        RECT 1979.435 1111.600 1979.725 1111.770 ;
        RECT 1979.895 1111.600 1980.185 1111.770 ;
        RECT 1980.355 1111.600 1980.645 1111.770 ;
        RECT 1980.815 1111.600 1981.105 1111.770 ;
        RECT 1981.275 1111.600 1981.565 1111.770 ;
        RECT 1981.735 1111.600 1982.025 1111.770 ;
        RECT 1982.195 1111.600 1982.485 1111.770 ;
        RECT 1982.655 1111.600 1982.945 1111.770 ;
        RECT 1983.115 1111.600 1983.405 1111.770 ;
        RECT 1983.575 1111.600 1983.865 1111.770 ;
        RECT 1984.035 1111.600 1984.325 1111.770 ;
        RECT 1984.495 1111.600 1984.785 1111.770 ;
        RECT 1984.955 1111.600 1985.245 1111.770 ;
        RECT 1985.415 1111.600 1985.705 1111.770 ;
        RECT 1985.875 1111.600 1986.165 1111.770 ;
        RECT 1986.335 1111.600 1986.625 1111.770 ;
        RECT 1986.795 1111.600 1987.085 1111.770 ;
        RECT 1987.255 1111.600 1987.545 1111.770 ;
        RECT 1987.715 1111.600 1988.005 1111.770 ;
        RECT 1988.175 1111.600 1988.465 1111.770 ;
        RECT 1988.635 1111.600 1988.925 1111.770 ;
        RECT 1989.095 1111.600 1989.385 1111.770 ;
        RECT 1989.555 1111.600 1989.845 1111.770 ;
        RECT 1990.015 1111.600 1990.305 1111.770 ;
        RECT 1990.475 1111.600 1990.765 1111.770 ;
        RECT 1990.935 1111.600 1991.225 1111.770 ;
        RECT 1991.395 1111.600 1991.685 1111.770 ;
        RECT 1991.855 1111.600 1992.145 1111.770 ;
        RECT 1992.315 1111.600 1992.605 1111.770 ;
        RECT 1992.775 1111.600 1993.065 1111.770 ;
        RECT 1993.235 1111.600 1993.525 1111.770 ;
        RECT 1993.695 1111.600 1993.985 1111.770 ;
        RECT 1994.155 1111.600 1994.445 1111.770 ;
        RECT 1994.615 1111.600 1994.905 1111.770 ;
        RECT 1995.075 1111.600 1995.365 1111.770 ;
        RECT 1995.535 1111.600 1995.825 1111.770 ;
        RECT 1995.995 1111.600 1996.285 1111.770 ;
        RECT 1996.455 1111.600 1996.745 1111.770 ;
        RECT 1996.915 1111.600 1997.205 1111.770 ;
        RECT 1997.375 1111.600 1997.665 1111.770 ;
        RECT 1997.835 1111.600 1998.125 1111.770 ;
        RECT 1998.295 1111.600 1998.585 1111.770 ;
        RECT 1998.755 1111.600 1999.045 1111.770 ;
        RECT 1999.215 1111.600 1999.505 1111.770 ;
        RECT 1999.675 1111.600 1999.965 1111.770 ;
        RECT 2000.135 1111.600 2000.425 1111.770 ;
        RECT 2000.595 1111.600 2000.885 1111.770 ;
        RECT 2001.055 1111.600 2001.345 1111.770 ;
        RECT 2001.515 1111.600 2001.805 1111.770 ;
        RECT 2001.975 1111.600 2002.265 1111.770 ;
        RECT 2002.435 1111.600 2002.725 1111.770 ;
        RECT 2002.895 1111.600 2003.185 1111.770 ;
        RECT 2003.355 1111.600 2003.645 1111.770 ;
        RECT 2003.815 1111.600 2004.105 1111.770 ;
        RECT 2004.275 1111.600 2004.565 1111.770 ;
        RECT 2004.735 1111.600 2005.025 1111.770 ;
        RECT 2005.195 1111.600 2005.485 1111.770 ;
        RECT 2005.655 1111.600 2005.945 1111.770 ;
        RECT 2006.115 1111.600 2006.405 1111.770 ;
        RECT 2006.575 1111.600 2006.865 1111.770 ;
        RECT 2007.035 1111.600 2007.325 1111.770 ;
        RECT 2007.495 1111.600 2007.785 1111.770 ;
        RECT 2007.955 1111.600 2008.245 1111.770 ;
        RECT 2008.415 1111.600 2008.705 1111.770 ;
        RECT 2008.875 1111.600 2009.165 1111.770 ;
        RECT 2009.335 1111.600 2009.625 1111.770 ;
        RECT 2009.795 1111.600 2010.085 1111.770 ;
        RECT 2010.255 1111.600 2010.545 1111.770 ;
        RECT 2010.715 1111.600 2011.005 1111.770 ;
        RECT 2011.175 1111.600 2011.465 1111.770 ;
        RECT 2011.635 1111.600 2011.925 1111.770 ;
        RECT 2012.095 1111.600 2012.385 1111.770 ;
        RECT 2012.555 1111.600 2012.845 1111.770 ;
        RECT 2013.015 1111.600 2013.305 1111.770 ;
        RECT 2013.475 1111.600 2013.765 1111.770 ;
        RECT 2013.935 1111.600 2014.225 1111.770 ;
        RECT 2014.395 1111.600 2014.685 1111.770 ;
        RECT 2014.855 1111.600 2015.145 1111.770 ;
        RECT 2015.315 1111.600 2015.605 1111.770 ;
        RECT 2015.775 1111.600 2016.065 1111.770 ;
        RECT 2016.235 1111.600 2016.525 1111.770 ;
        RECT 2016.695 1111.600 2016.985 1111.770 ;
        RECT 2017.155 1111.600 2017.445 1111.770 ;
        RECT 2017.615 1111.600 2017.905 1111.770 ;
        RECT 2018.075 1111.600 2018.365 1111.770 ;
        RECT 2018.535 1111.600 2018.825 1111.770 ;
        RECT 2018.995 1111.600 2019.285 1111.770 ;
        RECT 2019.455 1111.600 2019.745 1111.770 ;
        RECT 2019.915 1111.600 2020.205 1111.770 ;
        RECT 2020.375 1111.600 2020.665 1111.770 ;
        RECT 2020.835 1111.600 2021.125 1111.770 ;
        RECT 2021.295 1111.600 2021.585 1111.770 ;
        RECT 2021.755 1111.600 2022.045 1111.770 ;
        RECT 2022.215 1111.600 2022.505 1111.770 ;
        RECT 2022.675 1111.600 2022.965 1111.770 ;
        RECT 2023.135 1111.600 2023.425 1111.770 ;
        RECT 2023.595 1111.600 2023.885 1111.770 ;
        RECT 2024.055 1111.600 2024.345 1111.770 ;
        RECT 2024.515 1111.600 2024.805 1111.770 ;
        RECT 2024.975 1111.600 2025.265 1111.770 ;
        RECT 2025.435 1111.600 2025.725 1111.770 ;
        RECT 2025.895 1111.600 2026.185 1111.770 ;
        RECT 2026.355 1111.600 2026.645 1111.770 ;
        RECT 2026.815 1111.600 2027.105 1111.770 ;
        RECT 2027.275 1111.600 2027.565 1111.770 ;
        RECT 2027.735 1111.600 2028.025 1111.770 ;
        RECT 2028.195 1111.600 2028.485 1111.770 ;
        RECT 2028.655 1111.600 2028.945 1111.770 ;
        RECT 2029.115 1111.600 2029.405 1111.770 ;
        RECT 2029.575 1111.600 2029.865 1111.770 ;
        RECT 2030.035 1111.600 2030.325 1111.770 ;
        RECT 2030.495 1111.600 2030.785 1111.770 ;
        RECT 2030.955 1111.600 2031.245 1111.770 ;
        RECT 2031.415 1111.600 2031.705 1111.770 ;
        RECT 2031.875 1111.600 2032.165 1111.770 ;
        RECT 2032.335 1111.600 2032.625 1111.770 ;
        RECT 2032.795 1111.600 2033.085 1111.770 ;
        RECT 2033.255 1111.600 2033.545 1111.770 ;
        RECT 2033.715 1111.600 2034.005 1111.770 ;
        RECT 2034.175 1111.600 2034.465 1111.770 ;
        RECT 2034.635 1111.600 2034.925 1111.770 ;
        RECT 2035.095 1111.600 2035.385 1111.770 ;
        RECT 2035.555 1111.600 2035.845 1111.770 ;
        RECT 2036.015 1111.600 2036.305 1111.770 ;
        RECT 2036.475 1111.600 2036.765 1111.770 ;
        RECT 2036.935 1111.600 2037.225 1111.770 ;
        RECT 2037.395 1111.600 2037.685 1111.770 ;
        RECT 2037.855 1111.600 2038.145 1111.770 ;
        RECT 2038.315 1111.600 2038.605 1111.770 ;
        RECT 2038.775 1111.600 2039.065 1111.770 ;
        RECT 2039.235 1111.600 2039.525 1111.770 ;
        RECT 2039.695 1111.600 2039.985 1111.770 ;
        RECT 2040.155 1111.600 2040.445 1111.770 ;
        RECT 2040.615 1111.600 2040.905 1111.770 ;
        RECT 2041.075 1111.600 2041.365 1111.770 ;
        RECT 2041.535 1111.600 2041.825 1111.770 ;
        RECT 2041.995 1111.600 2042.285 1111.770 ;
        RECT 2042.455 1111.600 2042.745 1111.770 ;
        RECT 2042.915 1111.600 2043.205 1111.770 ;
        RECT 2043.375 1111.600 2043.665 1111.770 ;
        RECT 2043.835 1111.600 2044.125 1111.770 ;
        RECT 2044.295 1111.600 2044.585 1111.770 ;
        RECT 2044.755 1111.600 2045.045 1111.770 ;
        RECT 2045.215 1111.600 2045.505 1111.770 ;
        RECT 2045.675 1111.600 2045.965 1111.770 ;
        RECT 2046.135 1111.600 2046.425 1111.770 ;
        RECT 2046.595 1111.600 2046.885 1111.770 ;
        RECT 2047.055 1111.600 2047.345 1111.770 ;
        RECT 2047.515 1111.600 2047.805 1111.770 ;
        RECT 2047.975 1111.600 2048.265 1111.770 ;
        RECT 2048.435 1111.600 2048.725 1111.770 ;
        RECT 2048.895 1111.600 2049.185 1111.770 ;
        RECT 2049.355 1111.600 2049.645 1111.770 ;
        RECT 2049.815 1111.600 2050.105 1111.770 ;
        RECT 2050.275 1111.600 2050.565 1111.770 ;
        RECT 2050.735 1111.600 2051.025 1111.770 ;
        RECT 2051.195 1111.600 2051.485 1111.770 ;
        RECT 2051.655 1111.600 2051.945 1111.770 ;
        RECT 2052.115 1111.600 2052.405 1111.770 ;
        RECT 2052.575 1111.600 2052.865 1111.770 ;
        RECT 2053.035 1111.600 2053.325 1111.770 ;
        RECT 2053.495 1111.600 2053.785 1111.770 ;
        RECT 2053.955 1111.600 2054.245 1111.770 ;
        RECT 2054.415 1111.600 2054.705 1111.770 ;
        RECT 2054.875 1111.600 2055.165 1111.770 ;
        RECT 2055.335 1111.600 2055.625 1111.770 ;
        RECT 2055.795 1111.600 2056.085 1111.770 ;
        RECT 2056.255 1111.600 2056.545 1111.770 ;
        RECT 2056.715 1111.600 2057.005 1111.770 ;
        RECT 2057.175 1111.600 2057.465 1111.770 ;
        RECT 2057.635 1111.600 2057.925 1111.770 ;
        RECT 2058.095 1111.600 2058.385 1111.770 ;
        RECT 2058.555 1111.600 2058.845 1111.770 ;
        RECT 2059.015 1111.600 2059.305 1111.770 ;
        RECT 2059.475 1111.600 2059.765 1111.770 ;
        RECT 2059.935 1111.600 2060.225 1111.770 ;
        RECT 2060.395 1111.600 2060.685 1111.770 ;
        RECT 2060.855 1111.600 2061.145 1111.770 ;
        RECT 2061.315 1111.600 2061.605 1111.770 ;
        RECT 2061.775 1111.600 2062.065 1111.770 ;
        RECT 2062.235 1111.600 2062.525 1111.770 ;
        RECT 2062.695 1111.600 2062.985 1111.770 ;
        RECT 2063.155 1111.600 2063.445 1111.770 ;
        RECT 2063.615 1111.600 2063.905 1111.770 ;
        RECT 2064.075 1111.600 2064.365 1111.770 ;
        RECT 2064.535 1111.600 2064.825 1111.770 ;
        RECT 2064.995 1111.600 2065.285 1111.770 ;
        RECT 2065.455 1111.600 2065.745 1111.770 ;
        RECT 2065.915 1111.600 2066.205 1111.770 ;
        RECT 2066.375 1111.600 2066.665 1111.770 ;
        RECT 2066.835 1111.600 2067.125 1111.770 ;
        RECT 2067.295 1111.600 2067.585 1111.770 ;
        RECT 2067.755 1111.600 2068.045 1111.770 ;
        RECT 2068.215 1111.600 2068.505 1111.770 ;
        RECT 2068.675 1111.600 2068.965 1111.770 ;
        RECT 2069.135 1111.600 2069.425 1111.770 ;
        RECT 2069.595 1111.600 2069.885 1111.770 ;
        RECT 2070.055 1111.600 2070.345 1111.770 ;
        RECT 2070.515 1111.600 2070.805 1111.770 ;
        RECT 2070.975 1111.600 2071.120 1111.770 ;
      LAYER mcon ;
        RECT 3384.350 3537.580 3385.200 3537.750 ;
        RECT 3387.750 3536.670 3387.920 3537.760 ;
        RECT 199.875 3018.240 200.045 3019.330 ;
        RECT 202.595 3019.150 203.445 3019.320 ;
        RECT 199.875 3012.260 200.045 3013.350 ;
        RECT 202.595 3013.170 203.445 3013.340 ;
        RECT 199.875 3006.280 200.045 3007.370 ;
        RECT 202.595 3007.190 203.445 3007.360 ;
        RECT 199.875 3000.300 200.045 3001.390 ;
        RECT 202.595 3001.210 203.445 3001.380 ;
        RECT 199.875 2994.320 200.045 2995.410 ;
        RECT 202.595 2995.230 203.445 2995.400 ;
        RECT 199.875 2988.340 200.045 2989.430 ;
        RECT 202.595 2989.250 203.445 2989.420 ;
        RECT 3384.690 2237.180 3384.860 2238.270 ;
        RECT 199.645 1731.475 200.495 1731.645 ;
        RECT 203.045 1731.965 203.215 1733.055 ;
        RECT 199.985 1727.335 200.155 1728.425 ;
        RECT 202.705 1728.245 203.555 1728.415 ;
        RECT 199.645 1725.495 200.495 1725.665 ;
        RECT 203.045 1725.985 203.215 1727.075 ;
        RECT 199.985 1721.355 200.155 1722.445 ;
        RECT 202.705 1722.265 203.555 1722.435 ;
        RECT 199.645 1719.515 200.495 1719.685 ;
        RECT 203.045 1720.005 203.215 1721.095 ;
        RECT 199.985 1715.375 200.155 1716.465 ;
        RECT 202.705 1716.285 203.555 1716.455 ;
        RECT 199.645 1713.535 200.495 1713.705 ;
        RECT 203.045 1714.025 203.215 1715.115 ;
        RECT 199.985 1709.395 200.155 1710.485 ;
        RECT 202.705 1710.305 203.555 1710.475 ;
        RECT 199.645 1707.555 200.495 1707.725 ;
        RECT 203.045 1708.045 203.215 1709.135 ;
        RECT 199.985 1703.415 200.155 1704.505 ;
        RECT 202.705 1704.325 203.555 1704.495 ;
        RECT 199.645 1701.575 200.495 1701.745 ;
        RECT 203.045 1702.065 203.215 1703.155 ;
        RECT 199.985 1697.435 200.155 1698.525 ;
        RECT 202.705 1698.345 203.555 1698.515 ;
        RECT 199.985 1691.455 200.155 1692.545 ;
        RECT 202.705 1692.365 203.555 1692.535 ;
        RECT 199.985 1685.475 200.155 1686.565 ;
        RECT 202.705 1686.385 203.555 1686.555 ;
        RECT 199.985 1679.495 200.155 1680.585 ;
        RECT 202.705 1680.405 203.555 1680.575 ;
        RECT 199.985 1673.515 200.155 1674.605 ;
        RECT 202.705 1674.425 203.555 1674.595 ;
        RECT 670.520 1115.510 670.690 1116.360 ;
        RECT 674.240 1115.850 675.330 1116.020 ;
        RECT 676.500 1115.510 676.670 1116.360 ;
        RECT 680.220 1115.850 681.310 1116.020 ;
        RECT 682.480 1115.510 682.650 1116.360 ;
        RECT 686.200 1115.850 687.290 1116.020 ;
        RECT 688.460 1115.510 688.630 1116.360 ;
        RECT 692.180 1115.850 693.270 1116.020 ;
        RECT 694.440 1115.510 694.610 1116.360 ;
        RECT 698.160 1115.850 699.250 1116.020 ;
        RECT 700.420 1115.510 700.590 1116.360 ;
        RECT 704.140 1115.850 705.230 1116.020 ;
        RECT 706.400 1115.510 706.570 1116.360 ;
        RECT 710.120 1115.850 711.210 1116.020 ;
        RECT 712.380 1115.510 712.550 1116.360 ;
        RECT 716.100 1115.850 717.190 1116.020 ;
        RECT 718.360 1115.510 718.530 1116.360 ;
        RECT 722.080 1115.850 723.170 1116.020 ;
        RECT 724.340 1115.510 724.510 1116.360 ;
        RECT 728.060 1115.850 729.150 1116.020 ;
        RECT 740.020 1115.850 741.110 1116.020 ;
        RECT 746.000 1115.850 747.090 1116.020 ;
        RECT 751.980 1115.850 753.070 1116.020 ;
        RECT 757.960 1115.850 759.050 1116.020 ;
        RECT 763.940 1115.850 765.030 1116.020 ;
        RECT 769.920 1115.850 771.010 1116.020 ;
        RECT 1970.520 1115.510 1970.690 1116.360 ;
        RECT 1976.500 1115.510 1976.670 1116.360 ;
        RECT 1982.480 1115.510 1982.650 1116.360 ;
        RECT 1988.460 1115.510 1988.630 1116.360 ;
        RECT 1994.440 1115.510 1994.610 1116.360 ;
        RECT 2000.420 1115.510 2000.590 1116.360 ;
        RECT 2006.400 1115.510 2006.570 1116.360 ;
        RECT 2012.380 1115.510 2012.550 1116.360 ;
        RECT 2018.360 1115.510 2018.530 1116.360 ;
        RECT 2024.340 1115.510 2024.510 1116.360 ;
        RECT 2036.300 1115.510 2036.470 1116.360 ;
        RECT 2042.280 1115.510 2042.450 1116.360 ;
        RECT 2048.260 1115.510 2048.430 1116.360 ;
        RECT 2054.240 1115.510 2054.410 1116.360 ;
        RECT 2060.220 1115.510 2060.390 1116.360 ;
        RECT 2066.200 1115.510 2066.370 1116.360 ;
        RECT 675.590 1112.790 676.680 1112.960 ;
        RECT 679.730 1112.450 679.900 1113.300 ;
        RECT 681.570 1112.790 682.660 1112.960 ;
        RECT 685.710 1112.450 685.880 1113.300 ;
        RECT 687.550 1112.790 688.640 1112.960 ;
        RECT 691.690 1112.450 691.860 1113.300 ;
        RECT 693.530 1112.790 694.620 1112.960 ;
        RECT 697.670 1112.450 697.840 1113.300 ;
        RECT 699.510 1112.790 700.600 1112.960 ;
        RECT 703.650 1112.450 703.820 1113.300 ;
        RECT 705.490 1112.790 706.580 1112.960 ;
        RECT 709.630 1112.450 709.800 1113.300 ;
        RECT 711.470 1112.790 712.560 1112.960 ;
        RECT 715.610 1112.450 715.780 1113.300 ;
        RECT 717.450 1112.790 718.540 1112.960 ;
        RECT 721.590 1112.450 721.760 1113.300 ;
        RECT 723.430 1112.790 724.520 1112.960 ;
        RECT 727.570 1112.450 727.740 1113.300 ;
        RECT 729.410 1112.790 730.500 1112.960 ;
        RECT 733.550 1112.450 733.720 1113.300 ;
        RECT 745.510 1112.450 745.680 1113.300 ;
        RECT 751.490 1112.450 751.660 1113.300 ;
        RECT 757.470 1112.450 757.640 1113.300 ;
        RECT 763.450 1112.450 763.620 1113.300 ;
        RECT 769.420 1112.790 770.510 1112.960 ;
        RECT 1975.590 1112.790 1976.680 1112.960 ;
        RECT 1981.570 1112.790 1982.660 1112.960 ;
        RECT 1987.550 1112.790 1988.640 1112.960 ;
        RECT 1993.530 1112.790 1994.620 1112.960 ;
        RECT 1999.510 1112.790 2000.600 1112.960 ;
        RECT 2005.490 1112.790 2006.580 1112.960 ;
        RECT 2011.470 1112.790 2012.560 1112.960 ;
        RECT 2017.450 1112.790 2018.540 1112.960 ;
        RECT 2023.430 1112.790 2024.520 1112.960 ;
        RECT 2029.410 1112.790 2030.500 1112.960 ;
        RECT 2041.370 1112.790 2042.460 1112.960 ;
        RECT 2047.350 1112.790 2048.440 1112.960 ;
        RECT 2053.330 1112.790 2054.420 1112.960 ;
        RECT 2059.310 1112.790 2060.400 1112.960 ;
        RECT 2066.200 1112.450 2066.370 1113.300 ;
      LAYER met1 ;
        RECT 3381.780 3537.550 3382.040 3537.870 ;
        RECT 3381.620 3537.250 3381.760 3537.275 ;
        RECT 3381.500 3536.930 3381.760 3537.250 ;
        RECT 199.835 3018.180 200.095 3019.390 ;
        RECT 202.535 3019.100 203.505 3019.360 ;
        RECT 205.875 3019.120 206.135 3019.440 ;
        RECT 199.835 3012.200 200.095 3013.410 ;
        RECT 202.535 3013.120 203.505 3013.380 ;
        RECT 199.835 3006.220 200.095 3007.430 ;
        RECT 202.535 3007.140 203.505 3007.400 ;
        RECT 199.835 3000.240 200.095 3001.450 ;
        RECT 202.535 3001.160 203.505 3001.420 ;
        RECT 199.835 2994.260 200.095 2995.470 ;
        RECT 202.535 2995.180 203.505 2995.440 ;
        RECT 199.835 2988.280 200.095 2989.490 ;
        RECT 202.535 2989.200 203.505 2989.460 ;
        RECT 203.005 1731.905 203.265 1733.115 ;
        RECT 205.875 1732.750 206.015 3019.120 ;
        RECT 205.755 1732.430 206.015 1732.750 ;
        RECT 206.155 3018.500 206.415 3018.820 ;
        RECT 206.155 1731.780 206.295 3018.500 ;
        RECT 199.585 1731.425 200.555 1731.685 ;
        RECT 206.035 1731.460 206.295 1731.780 ;
        RECT 206.435 3013.140 206.695 3013.460 ;
        RECT 199.945 1727.275 200.205 1728.485 ;
        RECT 202.645 1728.195 203.615 1728.455 ;
        RECT 205.735 1728.215 205.995 1728.535 ;
        RECT 203.005 1725.925 203.265 1727.135 ;
        RECT 199.585 1725.445 200.555 1725.705 ;
        RECT 199.945 1721.295 200.205 1722.505 ;
        RECT 202.645 1722.215 203.615 1722.475 ;
        RECT 203.005 1719.945 203.265 1721.155 ;
        RECT 199.585 1719.465 200.555 1719.725 ;
        RECT 199.945 1715.315 200.205 1716.525 ;
        RECT 202.645 1716.235 203.615 1716.495 ;
        RECT 203.005 1713.965 203.265 1715.175 ;
        RECT 199.585 1713.485 200.555 1713.745 ;
        RECT 199.945 1709.335 200.205 1710.545 ;
        RECT 202.645 1710.255 203.615 1710.515 ;
        RECT 203.005 1707.985 203.265 1709.195 ;
        RECT 199.585 1707.505 200.555 1707.765 ;
        RECT 199.945 1703.355 200.205 1704.565 ;
        RECT 202.645 1704.275 203.615 1704.535 ;
        RECT 203.005 1702.005 203.265 1703.215 ;
        RECT 199.585 1701.525 200.555 1701.785 ;
        RECT 199.945 1697.375 200.205 1698.585 ;
        RECT 202.645 1698.295 203.615 1698.555 ;
        RECT 199.945 1691.395 200.205 1692.605 ;
        RECT 202.645 1692.315 203.615 1692.575 ;
        RECT 199.945 1685.415 200.205 1686.625 ;
        RECT 202.645 1686.335 203.615 1686.595 ;
        RECT 199.945 1679.435 200.205 1680.645 ;
        RECT 202.645 1680.355 203.615 1680.615 ;
        RECT 199.945 1673.455 200.205 1674.665 ;
        RECT 202.645 1674.375 203.615 1674.635 ;
        RECT 205.735 1121.260 205.875 1728.215 ;
        RECT 206.015 1727.595 206.275 1727.915 ;
        RECT 206.015 1121.540 206.155 1727.595 ;
        RECT 206.435 1726.770 206.575 3013.140 ;
        RECT 206.315 1726.450 206.575 1726.770 ;
        RECT 206.715 3012.520 206.975 3012.840 ;
        RECT 206.715 1725.800 206.855 3012.520 ;
        RECT 206.595 1725.480 206.855 1725.800 ;
        RECT 206.995 3007.160 207.255 3007.480 ;
        RECT 206.295 1722.235 206.555 1722.555 ;
        RECT 206.295 1121.820 206.435 1722.235 ;
        RECT 206.575 1721.615 206.835 1721.935 ;
        RECT 206.575 1122.100 206.715 1721.615 ;
        RECT 206.995 1720.790 207.135 3007.160 ;
        RECT 206.875 1720.470 207.135 1720.790 ;
        RECT 207.275 3006.540 207.535 3006.860 ;
        RECT 207.275 1719.820 207.415 3006.540 ;
        RECT 207.155 1719.500 207.415 1719.820 ;
        RECT 207.555 3001.180 207.815 3001.500 ;
        RECT 206.855 1716.255 207.115 1716.575 ;
        RECT 206.855 1122.380 206.995 1716.255 ;
        RECT 207.135 1715.635 207.395 1715.955 ;
        RECT 207.135 1122.660 207.275 1715.635 ;
        RECT 207.555 1714.810 207.695 3001.180 ;
        RECT 207.435 1714.490 207.695 1714.810 ;
        RECT 207.835 3000.560 208.095 3000.880 ;
        RECT 207.835 1713.840 207.975 3000.560 ;
        RECT 207.715 1713.520 207.975 1713.840 ;
        RECT 208.115 2995.200 208.375 2995.520 ;
        RECT 207.415 1710.275 207.675 1710.595 ;
        RECT 207.415 1122.940 207.555 1710.275 ;
        RECT 207.695 1709.655 207.955 1709.975 ;
        RECT 207.695 1123.220 207.835 1709.655 ;
        RECT 208.115 1708.830 208.255 2995.200 ;
        RECT 207.995 1708.510 208.255 1708.830 ;
        RECT 208.395 2994.580 208.655 2994.900 ;
        RECT 208.395 1707.860 208.535 2994.580 ;
        RECT 208.275 1707.540 208.535 1707.860 ;
        RECT 208.675 2989.220 208.935 2989.540 ;
        RECT 207.975 1704.295 208.235 1704.615 ;
        RECT 207.975 1123.500 208.115 1704.295 ;
        RECT 208.255 1703.675 208.515 1703.995 ;
        RECT 208.255 1123.780 208.395 1703.675 ;
        RECT 208.675 1702.850 208.815 2989.220 ;
        RECT 208.555 1702.530 208.815 1702.850 ;
        RECT 208.955 2988.600 209.215 2988.920 ;
        RECT 208.955 1701.880 209.095 2988.600 ;
        RECT 3381.620 2275.540 3381.760 3536.930 ;
        RECT 3381.480 2275.395 3381.760 2275.540 ;
        RECT 3381.480 2236.995 3381.620 2275.395 ;
        RECT 3381.900 2275.250 3382.040 3537.550 ;
        RECT 3384.290 3537.530 3385.260 3537.790 ;
        RECT 3387.700 3536.610 3387.960 3537.820 ;
        RECT 3381.760 2275.100 3382.040 2275.250 ;
        RECT 3381.760 2237.965 3381.900 2275.100 ;
        RECT 3381.760 2237.645 3382.020 2237.965 ;
        RECT 3384.640 2237.120 3384.900 2238.330 ;
        RECT 3381.480 2236.675 3381.740 2236.995 ;
        RECT 3387.350 2236.640 3388.320 2236.900 ;
        RECT 208.835 1701.560 209.095 1701.880 ;
        RECT 208.535 1698.315 208.795 1698.635 ;
        RECT 208.535 1124.060 208.675 1698.315 ;
        RECT 208.815 1697.695 209.075 1698.015 ;
        RECT 208.815 1124.340 208.955 1697.695 ;
        RECT 209.095 1692.335 209.355 1692.655 ;
        RECT 209.095 1124.620 209.235 1692.335 ;
        RECT 209.375 1691.715 209.635 1692.035 ;
        RECT 209.375 1124.900 209.515 1691.715 ;
        RECT 209.655 1686.355 209.915 1686.675 ;
        RECT 209.655 1125.180 209.795 1686.355 ;
        RECT 209.935 1685.735 210.195 1686.055 ;
        RECT 209.935 1125.460 210.075 1685.735 ;
        RECT 210.215 1680.375 210.475 1680.695 ;
        RECT 210.215 1125.740 210.355 1680.375 ;
        RECT 210.495 1679.755 210.755 1680.075 ;
        RECT 210.495 1126.020 210.635 1679.755 ;
        RECT 210.775 1674.395 211.035 1674.715 ;
        RECT 210.775 1126.300 210.915 1674.395 ;
        RECT 211.055 1673.775 211.315 1674.095 ;
        RECT 211.055 1126.580 211.195 1673.775 ;
        RECT 1970.490 1126.720 1970.810 1126.840 ;
        RECT 670.490 1126.580 670.810 1126.700 ;
        RECT 211.055 1126.440 670.810 1126.580 ;
        RECT 674.705 1126.580 1970.810 1126.720 ;
        RECT 674.705 1126.460 675.025 1126.580 ;
        RECT 1975.850 1126.440 1976.170 1126.560 ;
        RECT 675.850 1126.300 676.170 1126.420 ;
        RECT 210.775 1126.160 676.170 1126.300 ;
        RECT 679.715 1126.300 1976.170 1126.440 ;
        RECT 679.715 1126.180 680.035 1126.300 ;
        RECT 1976.470 1126.160 1976.790 1126.280 ;
        RECT 676.470 1126.020 676.790 1126.140 ;
        RECT 210.495 1125.880 676.790 1126.020 ;
        RECT 680.685 1126.020 1976.790 1126.160 ;
        RECT 680.685 1125.900 681.005 1126.020 ;
        RECT 1981.830 1125.880 1982.150 1126.000 ;
        RECT 681.830 1125.740 682.150 1125.860 ;
        RECT 210.215 1125.600 682.150 1125.740 ;
        RECT 685.695 1125.740 1982.150 1125.880 ;
        RECT 685.695 1125.620 686.015 1125.740 ;
        RECT 1982.450 1125.600 1982.770 1125.720 ;
        RECT 682.450 1125.460 682.770 1125.580 ;
        RECT 209.935 1125.320 682.770 1125.460 ;
        RECT 686.665 1125.460 1982.770 1125.600 ;
        RECT 686.665 1125.340 686.985 1125.460 ;
        RECT 1987.810 1125.320 1988.130 1125.440 ;
        RECT 687.810 1125.180 688.130 1125.300 ;
        RECT 209.655 1125.040 688.130 1125.180 ;
        RECT 691.675 1125.180 1988.130 1125.320 ;
        RECT 691.675 1125.060 691.995 1125.180 ;
        RECT 1988.430 1125.040 1988.750 1125.160 ;
        RECT 688.430 1124.900 688.750 1125.020 ;
        RECT 209.375 1124.760 688.750 1124.900 ;
        RECT 692.645 1124.900 1988.750 1125.040 ;
        RECT 692.645 1124.780 692.965 1124.900 ;
        RECT 1993.790 1124.760 1994.110 1124.880 ;
        RECT 693.790 1124.620 694.110 1124.740 ;
        RECT 209.095 1124.480 694.110 1124.620 ;
        RECT 697.655 1124.620 1994.110 1124.760 ;
        RECT 697.655 1124.500 697.975 1124.620 ;
        RECT 1994.410 1124.480 1994.730 1124.600 ;
        RECT 694.410 1124.340 694.730 1124.460 ;
        RECT 208.815 1124.200 694.730 1124.340 ;
        RECT 698.625 1124.340 1994.730 1124.480 ;
        RECT 698.625 1124.220 698.945 1124.340 ;
        RECT 1999.770 1124.200 2000.090 1124.320 ;
        RECT 699.770 1124.060 700.090 1124.180 ;
        RECT 208.535 1123.920 700.090 1124.060 ;
        RECT 703.635 1124.060 2000.090 1124.200 ;
        RECT 703.635 1123.940 703.955 1124.060 ;
        RECT 2000.390 1123.920 2000.710 1124.040 ;
        RECT 700.390 1123.780 700.710 1123.900 ;
        RECT 208.255 1123.640 700.710 1123.780 ;
        RECT 704.485 1123.780 2000.710 1123.920 ;
        RECT 704.485 1123.660 704.805 1123.780 ;
        RECT 2005.750 1123.640 2006.070 1123.760 ;
        RECT 705.750 1123.500 706.070 1123.620 ;
        RECT 207.975 1123.360 706.070 1123.500 ;
        RECT 709.615 1123.500 2006.070 1123.640 ;
        RECT 709.615 1123.380 709.935 1123.500 ;
        RECT 2006.370 1123.360 2006.690 1123.480 ;
        RECT 706.370 1123.220 706.690 1123.340 ;
        RECT 207.695 1123.080 706.690 1123.220 ;
        RECT 710.585 1123.220 2006.690 1123.360 ;
        RECT 710.585 1123.100 710.905 1123.220 ;
        RECT 2011.730 1123.080 2012.050 1123.200 ;
        RECT 711.730 1122.940 712.050 1123.060 ;
        RECT 207.415 1122.800 712.050 1122.940 ;
        RECT 715.595 1122.940 2012.050 1123.080 ;
        RECT 715.595 1122.820 715.915 1122.940 ;
        RECT 2012.350 1122.800 2012.670 1122.920 ;
        RECT 712.350 1122.660 712.670 1122.780 ;
        RECT 207.135 1122.520 712.670 1122.660 ;
        RECT 716.445 1122.660 2012.670 1122.800 ;
        RECT 716.445 1122.540 716.765 1122.660 ;
        RECT 2017.710 1122.520 2018.030 1122.640 ;
        RECT 717.710 1122.380 718.030 1122.500 ;
        RECT 206.855 1122.240 718.030 1122.380 ;
        RECT 721.575 1122.380 2018.030 1122.520 ;
        RECT 721.575 1122.260 721.895 1122.380 ;
        RECT 2018.330 1122.240 2018.650 1122.360 ;
        RECT 718.330 1122.100 718.650 1122.220 ;
        RECT 206.575 1121.960 718.650 1122.100 ;
        RECT 722.545 1122.100 2018.650 1122.240 ;
        RECT 722.545 1121.980 722.865 1122.100 ;
        RECT 2023.690 1121.960 2024.010 1122.080 ;
        RECT 723.690 1121.820 724.010 1121.940 ;
        RECT 206.295 1121.680 724.010 1121.820 ;
        RECT 727.555 1121.820 2024.010 1121.960 ;
        RECT 727.555 1121.700 727.875 1121.820 ;
        RECT 2024.310 1121.680 2024.630 1121.800 ;
        RECT 724.310 1121.540 724.630 1121.660 ;
        RECT 206.015 1121.400 724.630 1121.540 ;
        RECT 728.525 1121.540 2024.630 1121.680 ;
        RECT 728.525 1121.420 728.845 1121.540 ;
        RECT 2029.670 1121.400 2029.990 1121.520 ;
        RECT 729.670 1121.260 729.990 1121.380 ;
        RECT 733.000 1121.260 2029.990 1121.400 ;
        RECT 205.735 1121.120 729.990 1121.260 ;
        RECT 733.535 1121.140 733.855 1121.260 ;
        RECT 2036.270 1121.120 2036.590 1121.240 ;
        RECT 740.485 1120.980 2036.590 1121.120 ;
        RECT 740.485 1120.860 740.805 1120.980 ;
        RECT 2041.630 1120.840 2041.950 1120.960 ;
        RECT 745.495 1120.700 2041.950 1120.840 ;
        RECT 745.495 1120.580 745.815 1120.700 ;
        RECT 2042.250 1120.560 2042.570 1120.680 ;
        RECT 746.465 1120.420 2042.570 1120.560 ;
        RECT 746.465 1120.300 746.785 1120.420 ;
        RECT 2047.610 1120.280 2047.930 1120.400 ;
        RECT 751.475 1120.140 2047.930 1120.280 ;
        RECT 751.475 1120.020 751.795 1120.140 ;
        RECT 2048.230 1120.000 2048.550 1120.120 ;
        RECT 752.325 1119.860 2048.550 1120.000 ;
        RECT 752.325 1119.740 752.645 1119.860 ;
        RECT 2053.590 1119.720 2053.910 1119.840 ;
        RECT 757.455 1119.580 2053.910 1119.720 ;
        RECT 757.455 1119.460 757.775 1119.580 ;
        RECT 2054.210 1119.440 2054.530 1119.560 ;
        RECT 758.425 1119.300 2054.530 1119.440 ;
        RECT 758.425 1119.180 758.745 1119.300 ;
        RECT 2059.570 1119.160 2059.890 1119.280 ;
        RECT 763.435 1119.020 2059.890 1119.160 ;
        RECT 763.435 1118.900 763.755 1119.020 ;
        RECT 2060.190 1118.880 2060.510 1119.000 ;
        RECT 764.285 1118.740 2060.510 1118.880 ;
        RECT 764.285 1118.620 764.605 1118.740 ;
        RECT 2065.550 1118.600 2065.870 1118.720 ;
        RECT 769.415 1118.460 2065.870 1118.600 ;
        RECT 769.415 1118.340 769.735 1118.460 ;
        RECT 2066.170 1118.320 2066.490 1118.440 ;
        RECT 770.385 1118.180 2066.490 1118.320 ;
        RECT 770.385 1118.060 770.705 1118.180 ;
        RECT 670.470 1115.450 670.730 1116.420 ;
        RECT 674.180 1115.810 675.390 1116.070 ;
        RECT 676.450 1115.450 676.710 1116.420 ;
        RECT 680.160 1115.810 681.370 1116.070 ;
        RECT 682.430 1115.450 682.690 1116.420 ;
        RECT 686.140 1115.810 687.350 1116.070 ;
        RECT 688.410 1115.450 688.670 1116.420 ;
        RECT 692.120 1115.810 693.330 1116.070 ;
        RECT 694.390 1115.450 694.650 1116.420 ;
        RECT 698.100 1115.810 699.310 1116.070 ;
        RECT 700.370 1115.450 700.630 1116.420 ;
        RECT 704.080 1115.810 705.290 1116.070 ;
        RECT 706.350 1115.450 706.610 1116.420 ;
        RECT 710.060 1115.810 711.270 1116.070 ;
        RECT 712.330 1115.450 712.590 1116.420 ;
        RECT 716.040 1115.810 717.250 1116.070 ;
        RECT 718.310 1115.450 718.570 1116.420 ;
        RECT 722.020 1115.810 723.230 1116.070 ;
        RECT 724.290 1115.450 724.550 1116.420 ;
        RECT 728.000 1115.810 729.210 1116.070 ;
        RECT 739.960 1115.810 741.170 1116.070 ;
        RECT 745.940 1115.810 747.150 1116.070 ;
        RECT 751.920 1115.810 753.130 1116.070 ;
        RECT 757.900 1115.810 759.110 1116.070 ;
        RECT 763.880 1115.810 765.090 1116.070 ;
        RECT 769.860 1115.810 771.070 1116.070 ;
        RECT 1970.470 1115.450 1970.730 1116.420 ;
        RECT 1976.450 1115.450 1976.710 1116.420 ;
        RECT 1982.430 1115.450 1982.690 1116.420 ;
        RECT 1988.410 1115.450 1988.670 1116.420 ;
        RECT 1994.390 1115.450 1994.650 1116.420 ;
        RECT 2000.370 1115.450 2000.630 1116.420 ;
        RECT 2006.350 1115.450 2006.610 1116.420 ;
        RECT 2012.330 1115.450 2012.590 1116.420 ;
        RECT 2018.310 1115.450 2018.570 1116.420 ;
        RECT 2024.290 1115.450 2024.550 1116.420 ;
        RECT 2036.250 1115.450 2036.510 1116.420 ;
        RECT 2042.230 1115.450 2042.490 1116.420 ;
        RECT 2048.210 1115.450 2048.470 1116.420 ;
        RECT 2054.190 1115.450 2054.450 1116.420 ;
        RECT 2060.170 1115.450 2060.430 1116.420 ;
        RECT 2066.150 1115.450 2066.410 1116.420 ;
        RECT 675.530 1112.750 676.740 1113.010 ;
        RECT 679.680 1112.390 679.940 1113.360 ;
        RECT 681.510 1112.750 682.720 1113.010 ;
        RECT 685.660 1112.390 685.920 1113.360 ;
        RECT 687.490 1112.750 688.700 1113.010 ;
        RECT 691.640 1112.390 691.900 1113.360 ;
        RECT 693.470 1112.750 694.680 1113.010 ;
        RECT 697.620 1112.390 697.880 1113.360 ;
        RECT 699.450 1112.750 700.660 1113.010 ;
        RECT 703.600 1112.390 703.860 1113.360 ;
        RECT 705.430 1112.750 706.640 1113.010 ;
        RECT 709.580 1112.390 709.840 1113.360 ;
        RECT 711.410 1112.750 712.620 1113.010 ;
        RECT 715.560 1112.390 715.820 1113.360 ;
        RECT 717.390 1112.750 718.600 1113.010 ;
        RECT 721.540 1112.390 721.800 1113.360 ;
        RECT 723.370 1112.750 724.580 1113.010 ;
        RECT 727.520 1112.390 727.780 1113.360 ;
        RECT 729.350 1112.750 730.560 1113.010 ;
        RECT 733.500 1112.390 733.760 1113.360 ;
        RECT 745.460 1112.390 745.720 1113.360 ;
        RECT 751.440 1112.390 751.700 1113.360 ;
        RECT 757.420 1112.390 757.680 1113.360 ;
        RECT 763.400 1112.390 763.660 1113.360 ;
        RECT 769.360 1112.750 770.570 1113.010 ;
        RECT 1975.530 1112.750 1976.740 1113.010 ;
        RECT 1981.510 1112.750 1982.720 1113.010 ;
        RECT 1987.490 1112.750 1988.700 1113.010 ;
        RECT 1993.470 1112.750 1994.680 1113.010 ;
        RECT 1999.450 1112.750 2000.660 1113.010 ;
        RECT 2005.430 1112.750 2006.640 1113.010 ;
        RECT 2011.410 1112.750 2012.620 1113.010 ;
        RECT 2017.390 1112.750 2018.600 1113.010 ;
        RECT 2023.370 1112.750 2024.580 1113.010 ;
        RECT 2029.350 1112.750 2030.560 1113.010 ;
        RECT 2041.310 1112.750 2042.520 1113.010 ;
        RECT 2047.290 1112.750 2048.500 1113.010 ;
        RECT 2053.270 1112.750 2054.480 1113.010 ;
        RECT 2059.250 1112.750 2060.460 1113.010 ;
        RECT 2066.160 1112.390 2066.420 1113.360 ;
      LAYER via ;
        RECT 3381.780 3537.580 3382.040 3537.840 ;
        RECT 3381.500 3536.960 3381.760 3537.220 ;
        RECT 199.835 3018.240 200.095 3019.330 ;
        RECT 202.595 3019.100 203.445 3019.360 ;
        RECT 205.875 3019.150 206.135 3019.410 ;
        RECT 199.835 3012.260 200.095 3013.350 ;
        RECT 202.595 3013.120 203.445 3013.380 ;
        RECT 199.835 3006.280 200.095 3007.370 ;
        RECT 202.595 3007.140 203.445 3007.400 ;
        RECT 199.835 3000.300 200.095 3001.390 ;
        RECT 202.595 3001.160 203.445 3001.420 ;
        RECT 199.835 2994.320 200.095 2995.410 ;
        RECT 202.595 2995.180 203.445 2995.440 ;
        RECT 199.835 2988.340 200.095 2989.430 ;
        RECT 202.595 2989.200 203.445 2989.460 ;
        RECT 203.005 1731.965 203.265 1733.055 ;
        RECT 205.755 1732.460 206.015 1732.720 ;
        RECT 206.155 3018.530 206.415 3018.790 ;
        RECT 199.645 1731.425 200.495 1731.685 ;
        RECT 206.035 1731.490 206.295 1731.750 ;
        RECT 206.435 3013.170 206.695 3013.430 ;
        RECT 199.945 1727.335 200.205 1728.425 ;
        RECT 202.705 1728.195 203.555 1728.455 ;
        RECT 205.735 1728.245 205.995 1728.505 ;
        RECT 203.005 1725.985 203.265 1727.075 ;
        RECT 199.645 1725.445 200.495 1725.705 ;
        RECT 199.945 1721.355 200.205 1722.445 ;
        RECT 202.705 1722.215 203.555 1722.475 ;
        RECT 203.005 1720.005 203.265 1721.095 ;
        RECT 199.645 1719.465 200.495 1719.725 ;
        RECT 199.945 1715.375 200.205 1716.465 ;
        RECT 202.705 1716.235 203.555 1716.495 ;
        RECT 203.005 1714.025 203.265 1715.115 ;
        RECT 199.645 1713.485 200.495 1713.745 ;
        RECT 199.945 1709.395 200.205 1710.485 ;
        RECT 202.705 1710.255 203.555 1710.515 ;
        RECT 203.005 1708.045 203.265 1709.135 ;
        RECT 199.645 1707.505 200.495 1707.765 ;
        RECT 199.945 1703.415 200.205 1704.505 ;
        RECT 202.705 1704.275 203.555 1704.535 ;
        RECT 203.005 1702.065 203.265 1703.155 ;
        RECT 199.645 1701.525 200.495 1701.785 ;
        RECT 199.945 1697.435 200.205 1698.525 ;
        RECT 202.705 1698.295 203.555 1698.555 ;
        RECT 199.945 1691.455 200.205 1692.545 ;
        RECT 202.705 1692.315 203.555 1692.575 ;
        RECT 199.945 1685.475 200.205 1686.565 ;
        RECT 202.705 1686.335 203.555 1686.595 ;
        RECT 199.945 1679.495 200.205 1680.585 ;
        RECT 202.705 1680.355 203.555 1680.615 ;
        RECT 199.945 1673.515 200.205 1674.605 ;
        RECT 202.705 1674.375 203.555 1674.635 ;
        RECT 206.015 1727.625 206.275 1727.885 ;
        RECT 206.315 1726.480 206.575 1726.740 ;
        RECT 206.715 3012.550 206.975 3012.810 ;
        RECT 206.595 1725.510 206.855 1725.770 ;
        RECT 206.995 3007.190 207.255 3007.450 ;
        RECT 206.295 1722.265 206.555 1722.525 ;
        RECT 206.575 1721.645 206.835 1721.905 ;
        RECT 206.875 1720.500 207.135 1720.760 ;
        RECT 207.275 3006.570 207.535 3006.830 ;
        RECT 207.155 1719.530 207.415 1719.790 ;
        RECT 207.555 3001.210 207.815 3001.470 ;
        RECT 206.855 1716.285 207.115 1716.545 ;
        RECT 207.135 1715.665 207.395 1715.925 ;
        RECT 207.435 1714.520 207.695 1714.780 ;
        RECT 207.835 3000.590 208.095 3000.850 ;
        RECT 207.715 1713.550 207.975 1713.810 ;
        RECT 208.115 2995.230 208.375 2995.490 ;
        RECT 207.415 1710.305 207.675 1710.565 ;
        RECT 207.695 1709.685 207.955 1709.945 ;
        RECT 207.995 1708.540 208.255 1708.800 ;
        RECT 208.395 2994.610 208.655 2994.870 ;
        RECT 208.275 1707.570 208.535 1707.830 ;
        RECT 208.675 2989.250 208.935 2989.510 ;
        RECT 207.975 1704.325 208.235 1704.585 ;
        RECT 208.255 1703.705 208.515 1703.965 ;
        RECT 208.555 1702.560 208.815 1702.820 ;
        RECT 208.955 2988.630 209.215 2988.890 ;
        RECT 3384.350 3537.530 3385.200 3537.790 ;
        RECT 3387.700 3536.670 3387.960 3537.760 ;
        RECT 3381.760 2237.675 3382.020 2237.935 ;
        RECT 3384.640 2237.180 3384.900 2238.270 ;
        RECT 3381.480 2236.705 3381.740 2236.965 ;
        RECT 3387.410 2236.640 3388.260 2236.900 ;
        RECT 208.835 1701.590 209.095 1701.850 ;
        RECT 208.535 1698.345 208.795 1698.605 ;
        RECT 208.815 1697.725 209.075 1697.985 ;
        RECT 209.095 1692.365 209.355 1692.625 ;
        RECT 209.375 1691.745 209.635 1692.005 ;
        RECT 209.655 1686.385 209.915 1686.645 ;
        RECT 209.935 1685.765 210.195 1686.025 ;
        RECT 210.215 1680.405 210.475 1680.665 ;
        RECT 210.495 1679.785 210.755 1680.045 ;
        RECT 210.775 1674.425 211.035 1674.685 ;
        RECT 211.055 1673.805 211.315 1674.065 ;
        RECT 670.520 1126.440 670.780 1126.700 ;
        RECT 674.735 1126.460 674.995 1126.720 ;
        RECT 1970.520 1126.580 1970.780 1126.840 ;
        RECT 675.880 1126.160 676.140 1126.420 ;
        RECT 679.745 1126.180 680.005 1126.440 ;
        RECT 1975.880 1126.300 1976.140 1126.560 ;
        RECT 676.500 1125.880 676.760 1126.140 ;
        RECT 680.715 1125.900 680.975 1126.160 ;
        RECT 1976.500 1126.020 1976.760 1126.280 ;
        RECT 681.860 1125.600 682.120 1125.860 ;
        RECT 685.725 1125.620 685.985 1125.880 ;
        RECT 1981.860 1125.740 1982.120 1126.000 ;
        RECT 682.480 1125.320 682.740 1125.580 ;
        RECT 686.695 1125.340 686.955 1125.600 ;
        RECT 1982.480 1125.460 1982.740 1125.720 ;
        RECT 687.840 1125.040 688.100 1125.300 ;
        RECT 691.705 1125.060 691.965 1125.320 ;
        RECT 1987.840 1125.180 1988.100 1125.440 ;
        RECT 688.460 1124.760 688.720 1125.020 ;
        RECT 692.675 1124.780 692.935 1125.040 ;
        RECT 1988.460 1124.900 1988.720 1125.160 ;
        RECT 693.820 1124.480 694.080 1124.740 ;
        RECT 697.685 1124.500 697.945 1124.760 ;
        RECT 1993.820 1124.620 1994.080 1124.880 ;
        RECT 694.440 1124.200 694.700 1124.460 ;
        RECT 698.655 1124.220 698.915 1124.480 ;
        RECT 1994.440 1124.340 1994.700 1124.600 ;
        RECT 699.800 1123.920 700.060 1124.180 ;
        RECT 703.665 1123.940 703.925 1124.200 ;
        RECT 1999.800 1124.060 2000.060 1124.320 ;
        RECT 700.420 1123.640 700.680 1123.900 ;
        RECT 704.515 1123.660 704.775 1123.920 ;
        RECT 2000.420 1123.780 2000.680 1124.040 ;
        RECT 705.780 1123.360 706.040 1123.620 ;
        RECT 709.645 1123.380 709.905 1123.640 ;
        RECT 2005.780 1123.500 2006.040 1123.760 ;
        RECT 706.400 1123.080 706.660 1123.340 ;
        RECT 710.615 1123.100 710.875 1123.360 ;
        RECT 2006.400 1123.220 2006.660 1123.480 ;
        RECT 711.760 1122.800 712.020 1123.060 ;
        RECT 715.625 1122.820 715.885 1123.080 ;
        RECT 2011.760 1122.940 2012.020 1123.200 ;
        RECT 712.380 1122.520 712.640 1122.780 ;
        RECT 716.475 1122.540 716.735 1122.800 ;
        RECT 2012.380 1122.660 2012.640 1122.920 ;
        RECT 717.740 1122.240 718.000 1122.500 ;
        RECT 721.605 1122.260 721.865 1122.520 ;
        RECT 2017.740 1122.380 2018.000 1122.640 ;
        RECT 718.360 1121.960 718.620 1122.220 ;
        RECT 722.575 1121.980 722.835 1122.240 ;
        RECT 2018.360 1122.100 2018.620 1122.360 ;
        RECT 723.720 1121.680 723.980 1121.940 ;
        RECT 727.585 1121.700 727.845 1121.960 ;
        RECT 2023.720 1121.820 2023.980 1122.080 ;
        RECT 724.340 1121.400 724.600 1121.660 ;
        RECT 728.555 1121.420 728.815 1121.680 ;
        RECT 2024.340 1121.540 2024.600 1121.800 ;
        RECT 729.700 1121.120 729.960 1121.380 ;
        RECT 733.565 1121.140 733.825 1121.400 ;
        RECT 2029.700 1121.260 2029.960 1121.520 ;
        RECT 740.515 1120.860 740.775 1121.120 ;
        RECT 2036.300 1120.980 2036.560 1121.240 ;
        RECT 745.525 1120.580 745.785 1120.840 ;
        RECT 2041.660 1120.700 2041.920 1120.960 ;
        RECT 746.495 1120.300 746.755 1120.560 ;
        RECT 2042.280 1120.420 2042.540 1120.680 ;
        RECT 751.505 1120.020 751.765 1120.280 ;
        RECT 2047.640 1120.140 2047.900 1120.400 ;
        RECT 752.355 1119.740 752.615 1120.000 ;
        RECT 2048.260 1119.860 2048.520 1120.120 ;
        RECT 757.485 1119.460 757.745 1119.720 ;
        RECT 2053.620 1119.580 2053.880 1119.840 ;
        RECT 758.455 1119.180 758.715 1119.440 ;
        RECT 2054.240 1119.300 2054.500 1119.560 ;
        RECT 763.465 1118.900 763.725 1119.160 ;
        RECT 2059.600 1119.020 2059.860 1119.280 ;
        RECT 764.315 1118.620 764.575 1118.880 ;
        RECT 2060.220 1118.740 2060.480 1119.000 ;
        RECT 769.445 1118.340 769.705 1118.600 ;
        RECT 2065.580 1118.460 2065.840 1118.720 ;
        RECT 770.415 1118.060 770.675 1118.320 ;
        RECT 2066.200 1118.180 2066.460 1118.440 ;
        RECT 670.470 1115.510 670.730 1116.360 ;
        RECT 674.240 1115.810 675.330 1116.070 ;
        RECT 676.450 1115.510 676.710 1116.360 ;
        RECT 680.220 1115.810 681.310 1116.070 ;
        RECT 682.430 1115.510 682.690 1116.360 ;
        RECT 686.200 1115.810 687.290 1116.070 ;
        RECT 688.410 1115.510 688.670 1116.360 ;
        RECT 692.180 1115.810 693.270 1116.070 ;
        RECT 694.390 1115.510 694.650 1116.360 ;
        RECT 698.160 1115.810 699.250 1116.070 ;
        RECT 700.370 1115.510 700.630 1116.360 ;
        RECT 704.140 1115.810 705.230 1116.070 ;
        RECT 706.350 1115.510 706.610 1116.360 ;
        RECT 710.120 1115.810 711.210 1116.070 ;
        RECT 712.330 1115.510 712.590 1116.360 ;
        RECT 716.100 1115.810 717.190 1116.070 ;
        RECT 718.310 1115.510 718.570 1116.360 ;
        RECT 722.080 1115.810 723.170 1116.070 ;
        RECT 724.290 1115.510 724.550 1116.360 ;
        RECT 728.060 1115.810 729.150 1116.070 ;
        RECT 740.020 1115.810 741.110 1116.070 ;
        RECT 746.000 1115.810 747.090 1116.070 ;
        RECT 751.980 1115.810 753.070 1116.070 ;
        RECT 757.960 1115.810 759.050 1116.070 ;
        RECT 763.940 1115.810 765.030 1116.070 ;
        RECT 769.920 1115.810 771.010 1116.070 ;
        RECT 1970.470 1115.510 1970.730 1116.360 ;
        RECT 1976.450 1115.510 1976.710 1116.360 ;
        RECT 1982.430 1115.510 1982.690 1116.360 ;
        RECT 1988.410 1115.510 1988.670 1116.360 ;
        RECT 1994.390 1115.510 1994.650 1116.360 ;
        RECT 2000.370 1115.510 2000.630 1116.360 ;
        RECT 2006.350 1115.510 2006.610 1116.360 ;
        RECT 2012.330 1115.510 2012.590 1116.360 ;
        RECT 2018.310 1115.510 2018.570 1116.360 ;
        RECT 2024.290 1115.510 2024.550 1116.360 ;
        RECT 2036.250 1115.510 2036.510 1116.360 ;
        RECT 2042.230 1115.510 2042.490 1116.360 ;
        RECT 2048.210 1115.510 2048.470 1116.360 ;
        RECT 2054.190 1115.510 2054.450 1116.360 ;
        RECT 2060.170 1115.510 2060.430 1116.360 ;
        RECT 2066.150 1115.510 2066.410 1116.360 ;
        RECT 675.590 1112.750 676.680 1113.010 ;
        RECT 679.680 1112.450 679.940 1113.300 ;
        RECT 681.570 1112.750 682.660 1113.010 ;
        RECT 685.660 1112.450 685.920 1113.300 ;
        RECT 687.550 1112.750 688.640 1113.010 ;
        RECT 691.640 1112.450 691.900 1113.300 ;
        RECT 693.530 1112.750 694.620 1113.010 ;
        RECT 697.620 1112.450 697.880 1113.300 ;
        RECT 699.510 1112.750 700.600 1113.010 ;
        RECT 703.600 1112.450 703.860 1113.300 ;
        RECT 705.490 1112.750 706.580 1113.010 ;
        RECT 709.580 1112.450 709.840 1113.300 ;
        RECT 711.470 1112.750 712.560 1113.010 ;
        RECT 715.560 1112.450 715.820 1113.300 ;
        RECT 717.450 1112.750 718.540 1113.010 ;
        RECT 721.540 1112.450 721.800 1113.300 ;
        RECT 723.430 1112.750 724.520 1113.010 ;
        RECT 727.520 1112.450 727.780 1113.300 ;
        RECT 729.410 1112.750 730.500 1113.010 ;
        RECT 733.500 1112.450 733.760 1113.300 ;
        RECT 745.460 1112.450 745.720 1113.300 ;
        RECT 751.440 1112.450 751.700 1113.300 ;
        RECT 757.420 1112.450 757.680 1113.300 ;
        RECT 763.400 1112.450 763.660 1113.300 ;
        RECT 769.420 1112.750 770.510 1113.010 ;
        RECT 1975.590 1112.750 1976.680 1113.010 ;
        RECT 1981.570 1112.750 1982.660 1113.010 ;
        RECT 1987.550 1112.750 1988.640 1113.010 ;
        RECT 1993.530 1112.750 1994.620 1113.010 ;
        RECT 1999.510 1112.750 2000.600 1113.010 ;
        RECT 2005.490 1112.750 2006.580 1113.010 ;
        RECT 2011.470 1112.750 2012.560 1113.010 ;
        RECT 2017.450 1112.750 2018.540 1113.010 ;
        RECT 2023.430 1112.750 2024.520 1113.010 ;
        RECT 2029.410 1112.750 2030.500 1113.010 ;
        RECT 2041.370 1112.750 2042.460 1113.010 ;
        RECT 2047.350 1112.750 2048.440 1113.010 ;
        RECT 2053.330 1112.750 2054.420 1113.010 ;
        RECT 2059.310 1112.750 2060.400 1113.010 ;
        RECT 2066.160 1112.450 2066.420 1113.300 ;
      LAYER met2 ;
        RECT 3381.750 3537.720 3382.070 3537.840 ;
        RECT 3384.350 3537.720 3385.200 3537.820 ;
        RECT 3381.310 3537.580 3385.200 3537.720 ;
        RECT 3384.350 3537.500 3385.200 3537.580 ;
        RECT 3381.470 3537.100 3381.790 3537.220 ;
        RECT 3387.670 3537.100 3387.990 3537.760 ;
        RECT 3381.310 3536.960 3387.990 3537.100 ;
        RECT 3387.670 3536.670 3387.990 3536.960 ;
        RECT 199.805 3018.670 200.125 3019.330 ;
        RECT 202.595 3019.290 203.445 3019.390 ;
        RECT 205.845 3019.290 206.165 3019.410 ;
        RECT 202.595 3019.150 209.300 3019.290 ;
        RECT 202.595 3019.070 203.445 3019.150 ;
        RECT 206.125 3018.670 206.445 3018.790 ;
        RECT 199.805 3018.530 209.300 3018.670 ;
        RECT 199.805 3018.240 200.125 3018.530 ;
        RECT 199.805 3012.690 200.125 3013.350 ;
        RECT 202.595 3013.310 203.445 3013.410 ;
        RECT 206.405 3013.310 206.725 3013.430 ;
        RECT 202.595 3013.170 209.300 3013.310 ;
        RECT 202.595 3013.090 203.445 3013.170 ;
        RECT 206.685 3012.690 207.005 3012.810 ;
        RECT 199.805 3012.550 209.300 3012.690 ;
        RECT 199.805 3012.260 200.125 3012.550 ;
        RECT 199.805 3006.710 200.125 3007.370 ;
        RECT 202.595 3007.330 203.445 3007.430 ;
        RECT 206.965 3007.330 207.285 3007.450 ;
        RECT 202.595 3007.190 209.300 3007.330 ;
        RECT 202.595 3007.110 203.445 3007.190 ;
        RECT 207.245 3006.710 207.565 3006.830 ;
        RECT 199.805 3006.570 209.300 3006.710 ;
        RECT 199.805 3006.280 200.125 3006.570 ;
        RECT 199.805 3000.730 200.125 3001.390 ;
        RECT 202.595 3001.350 203.445 3001.450 ;
        RECT 207.525 3001.350 207.845 3001.470 ;
        RECT 202.595 3001.210 209.300 3001.350 ;
        RECT 202.595 3001.130 203.445 3001.210 ;
        RECT 207.805 3000.730 208.125 3000.850 ;
        RECT 199.805 3000.590 209.300 3000.730 ;
        RECT 199.805 3000.300 200.125 3000.590 ;
        RECT 199.805 2994.750 200.125 2995.410 ;
        RECT 202.595 2995.370 203.445 2995.470 ;
        RECT 208.085 2995.370 208.405 2995.490 ;
        RECT 202.595 2995.230 209.300 2995.370 ;
        RECT 202.595 2995.150 203.445 2995.230 ;
        RECT 208.365 2994.750 208.685 2994.870 ;
        RECT 199.805 2994.610 209.300 2994.750 ;
        RECT 199.805 2994.320 200.125 2994.610 ;
        RECT 199.805 2988.770 200.125 2989.430 ;
        RECT 202.595 2989.390 203.445 2989.490 ;
        RECT 208.645 2989.390 208.965 2989.510 ;
        RECT 202.595 2989.250 209.300 2989.390 ;
        RECT 202.595 2989.170 203.445 2989.250 ;
        RECT 208.925 2988.770 209.245 2988.890 ;
        RECT 199.805 2988.630 209.300 2988.770 ;
        RECT 199.805 2988.340 200.125 2988.630 ;
        RECT 3381.730 2237.815 3382.050 2237.935 ;
        RECT 3384.610 2237.815 3384.930 2238.270 ;
        RECT 3377.950 2237.675 3384.930 2237.815 ;
        RECT 3384.610 2237.180 3384.930 2237.675 ;
        RECT 3381.450 2236.845 3381.770 2236.965 ;
        RECT 3387.410 2236.845 3388.260 2236.930 ;
        RECT 3377.950 2236.705 3388.260 2236.845 ;
        RECT 3387.410 2236.610 3388.260 2236.705 ;
        RECT 202.975 1732.600 203.295 1733.055 ;
        RECT 205.725 1732.600 206.045 1732.720 ;
        RECT 202.975 1732.460 211.440 1732.600 ;
        RECT 202.975 1731.965 203.295 1732.460 ;
        RECT 199.645 1731.630 200.495 1731.715 ;
        RECT 206.005 1731.630 206.325 1731.750 ;
        RECT 199.645 1731.490 211.440 1731.630 ;
        RECT 199.645 1731.395 200.495 1731.490 ;
        RECT 199.915 1727.765 200.235 1728.425 ;
        RECT 202.705 1728.385 203.555 1728.485 ;
        RECT 205.705 1728.385 206.025 1728.505 ;
        RECT 202.705 1728.245 211.440 1728.385 ;
        RECT 202.705 1728.165 203.555 1728.245 ;
        RECT 205.985 1727.765 206.305 1727.885 ;
        RECT 199.915 1727.625 211.440 1727.765 ;
        RECT 199.915 1727.335 200.235 1727.625 ;
        RECT 202.975 1726.620 203.295 1727.075 ;
        RECT 206.285 1726.620 206.605 1726.740 ;
        RECT 202.975 1726.480 211.440 1726.620 ;
        RECT 202.975 1725.985 203.295 1726.480 ;
        RECT 199.645 1725.650 200.495 1725.735 ;
        RECT 206.565 1725.650 206.885 1725.770 ;
        RECT 199.645 1725.510 211.440 1725.650 ;
        RECT 199.645 1725.415 200.495 1725.510 ;
        RECT 199.915 1721.785 200.235 1722.445 ;
        RECT 202.705 1722.405 203.555 1722.505 ;
        RECT 206.265 1722.405 206.585 1722.525 ;
        RECT 202.705 1722.265 211.440 1722.405 ;
        RECT 202.705 1722.185 203.555 1722.265 ;
        RECT 206.545 1721.785 206.865 1721.905 ;
        RECT 199.915 1721.645 211.440 1721.785 ;
        RECT 199.915 1721.355 200.235 1721.645 ;
        RECT 202.975 1720.640 203.295 1721.095 ;
        RECT 206.845 1720.640 207.165 1720.760 ;
        RECT 202.975 1720.500 211.440 1720.640 ;
        RECT 202.975 1720.005 203.295 1720.500 ;
        RECT 199.645 1719.670 200.495 1719.755 ;
        RECT 207.125 1719.670 207.445 1719.790 ;
        RECT 199.645 1719.530 211.440 1719.670 ;
        RECT 199.645 1719.435 200.495 1719.530 ;
        RECT 199.915 1715.805 200.235 1716.465 ;
        RECT 202.705 1716.425 203.555 1716.525 ;
        RECT 206.825 1716.425 207.145 1716.545 ;
        RECT 202.705 1716.285 211.440 1716.425 ;
        RECT 202.705 1716.205 203.555 1716.285 ;
        RECT 207.105 1715.805 207.425 1715.925 ;
        RECT 199.915 1715.665 211.440 1715.805 ;
        RECT 199.915 1715.375 200.235 1715.665 ;
        RECT 202.975 1714.660 203.295 1715.115 ;
        RECT 207.405 1714.660 207.725 1714.780 ;
        RECT 202.975 1714.520 211.440 1714.660 ;
        RECT 202.975 1714.025 203.295 1714.520 ;
        RECT 199.645 1713.690 200.495 1713.775 ;
        RECT 207.685 1713.690 208.005 1713.810 ;
        RECT 199.645 1713.550 211.440 1713.690 ;
        RECT 199.645 1713.455 200.495 1713.550 ;
        RECT 199.915 1709.825 200.235 1710.485 ;
        RECT 202.705 1710.445 203.555 1710.545 ;
        RECT 207.385 1710.445 207.705 1710.565 ;
        RECT 202.705 1710.305 211.440 1710.445 ;
        RECT 202.705 1710.225 203.555 1710.305 ;
        RECT 207.665 1709.825 207.985 1709.945 ;
        RECT 199.915 1709.685 211.440 1709.825 ;
        RECT 199.915 1709.395 200.235 1709.685 ;
        RECT 202.975 1708.680 203.295 1709.135 ;
        RECT 207.965 1708.680 208.285 1708.800 ;
        RECT 202.975 1708.540 211.440 1708.680 ;
        RECT 202.975 1708.045 203.295 1708.540 ;
        RECT 199.645 1707.710 200.495 1707.795 ;
        RECT 208.245 1707.710 208.565 1707.830 ;
        RECT 199.645 1707.570 211.440 1707.710 ;
        RECT 199.645 1707.475 200.495 1707.570 ;
        RECT 199.915 1703.845 200.235 1704.505 ;
        RECT 202.705 1704.465 203.555 1704.565 ;
        RECT 207.945 1704.465 208.265 1704.585 ;
        RECT 202.705 1704.325 211.440 1704.465 ;
        RECT 202.705 1704.245 203.555 1704.325 ;
        RECT 208.225 1703.845 208.545 1703.965 ;
        RECT 199.915 1703.705 211.440 1703.845 ;
        RECT 199.915 1703.415 200.235 1703.705 ;
        RECT 202.975 1702.700 203.295 1703.155 ;
        RECT 208.525 1702.700 208.845 1702.820 ;
        RECT 202.975 1702.560 211.440 1702.700 ;
        RECT 202.975 1702.065 203.295 1702.560 ;
        RECT 199.645 1701.730 200.495 1701.815 ;
        RECT 208.805 1701.730 209.125 1701.850 ;
        RECT 199.645 1701.590 211.440 1701.730 ;
        RECT 199.645 1701.495 200.495 1701.590 ;
        RECT 199.915 1697.865 200.235 1698.525 ;
        RECT 202.705 1698.485 203.555 1698.585 ;
        RECT 208.505 1698.485 208.825 1698.605 ;
        RECT 202.705 1698.345 211.440 1698.485 ;
        RECT 202.705 1698.265 203.555 1698.345 ;
        RECT 208.785 1697.865 209.105 1697.985 ;
        RECT 199.915 1697.725 211.440 1697.865 ;
        RECT 199.915 1697.435 200.235 1697.725 ;
        RECT 199.915 1691.885 200.235 1692.545 ;
        RECT 202.705 1692.505 203.555 1692.605 ;
        RECT 209.065 1692.505 209.385 1692.625 ;
        RECT 202.705 1692.365 211.440 1692.505 ;
        RECT 202.705 1692.285 203.555 1692.365 ;
        RECT 209.345 1691.885 209.665 1692.005 ;
        RECT 199.915 1691.745 211.440 1691.885 ;
        RECT 199.915 1691.455 200.235 1691.745 ;
        RECT 199.915 1685.905 200.235 1686.565 ;
        RECT 202.705 1686.525 203.555 1686.625 ;
        RECT 209.625 1686.525 209.945 1686.645 ;
        RECT 202.705 1686.385 211.440 1686.525 ;
        RECT 202.705 1686.305 203.555 1686.385 ;
        RECT 209.905 1685.905 210.225 1686.025 ;
        RECT 199.915 1685.765 211.440 1685.905 ;
        RECT 199.915 1685.475 200.235 1685.765 ;
        RECT 199.915 1679.925 200.235 1680.585 ;
        RECT 202.705 1680.545 203.555 1680.645 ;
        RECT 210.185 1680.545 210.505 1680.665 ;
        RECT 202.705 1680.405 211.440 1680.545 ;
        RECT 202.705 1680.325 203.555 1680.405 ;
        RECT 210.465 1679.925 210.785 1680.045 ;
        RECT 199.915 1679.785 211.440 1679.925 ;
        RECT 199.915 1679.495 200.235 1679.785 ;
        RECT 199.915 1673.945 200.235 1674.605 ;
        RECT 202.705 1674.565 203.555 1674.665 ;
        RECT 210.745 1674.565 211.065 1674.685 ;
        RECT 202.705 1674.425 211.440 1674.565 ;
        RECT 202.705 1674.345 203.555 1674.425 ;
        RECT 211.025 1673.945 211.345 1674.065 ;
        RECT 199.915 1673.805 211.440 1673.945 ;
        RECT 199.915 1673.515 200.235 1673.805 ;
        RECT 1970.520 1126.870 1970.660 1126.965 ;
        RECT 670.520 1126.730 670.660 1126.825 ;
        RECT 674.735 1126.750 674.875 1126.825 ;
        RECT 670.520 1126.410 670.780 1126.730 ;
        RECT 674.735 1126.430 674.995 1126.750 ;
        RECT 675.880 1126.450 676.020 1126.825 ;
        RECT 670.520 1116.360 670.660 1126.410 ;
        RECT 670.440 1115.510 670.760 1116.360 ;
        RECT 674.735 1116.100 674.875 1126.430 ;
        RECT 675.880 1126.130 676.140 1126.450 ;
        RECT 676.500 1126.170 676.640 1126.825 ;
        RECT 679.745 1126.470 679.885 1126.825 ;
        RECT 674.240 1115.780 675.330 1116.100 ;
        RECT 675.880 1113.040 676.020 1126.130 ;
        RECT 676.500 1125.850 676.760 1126.170 ;
        RECT 679.745 1126.150 680.005 1126.470 ;
        RECT 680.715 1126.190 680.855 1126.825 ;
        RECT 676.500 1116.360 676.640 1125.850 ;
        RECT 676.420 1115.510 676.740 1116.360 ;
        RECT 679.745 1113.300 679.885 1126.150 ;
        RECT 680.715 1125.870 680.975 1126.190 ;
        RECT 681.860 1125.890 682.000 1126.825 ;
        RECT 680.715 1116.100 680.855 1125.870 ;
        RECT 681.860 1125.570 682.120 1125.890 ;
        RECT 682.480 1125.610 682.620 1126.825 ;
        RECT 685.725 1125.910 685.865 1126.825 ;
        RECT 680.220 1115.780 681.310 1116.100 ;
        RECT 675.590 1112.720 676.680 1113.040 ;
        RECT 679.650 1112.450 679.970 1113.300 ;
        RECT 681.860 1113.040 682.000 1125.570 ;
        RECT 682.480 1125.290 682.740 1125.610 ;
        RECT 685.725 1125.590 685.985 1125.910 ;
        RECT 686.695 1125.630 686.835 1126.825 ;
        RECT 682.480 1116.360 682.620 1125.290 ;
        RECT 682.400 1115.510 682.720 1116.360 ;
        RECT 685.725 1113.300 685.865 1125.590 ;
        RECT 686.695 1125.310 686.955 1125.630 ;
        RECT 687.840 1125.330 687.980 1126.825 ;
        RECT 686.695 1116.100 686.835 1125.310 ;
        RECT 687.840 1125.010 688.100 1125.330 ;
        RECT 688.460 1125.050 688.600 1126.825 ;
        RECT 691.705 1125.350 691.845 1126.825 ;
        RECT 686.200 1115.780 687.290 1116.100 ;
        RECT 681.570 1112.720 682.660 1113.040 ;
        RECT 685.630 1112.450 685.950 1113.300 ;
        RECT 687.840 1113.040 687.980 1125.010 ;
        RECT 688.460 1124.730 688.720 1125.050 ;
        RECT 691.705 1125.030 691.965 1125.350 ;
        RECT 692.675 1125.070 692.815 1126.825 ;
        RECT 688.460 1116.360 688.600 1124.730 ;
        RECT 688.380 1115.510 688.700 1116.360 ;
        RECT 691.705 1113.300 691.845 1125.030 ;
        RECT 692.675 1124.750 692.935 1125.070 ;
        RECT 693.820 1124.770 693.960 1126.825 ;
        RECT 692.675 1116.100 692.815 1124.750 ;
        RECT 693.820 1124.450 694.080 1124.770 ;
        RECT 694.440 1124.490 694.580 1126.825 ;
        RECT 697.685 1124.790 697.825 1126.825 ;
        RECT 692.180 1115.780 693.270 1116.100 ;
        RECT 687.550 1112.720 688.640 1113.040 ;
        RECT 691.610 1112.450 691.930 1113.300 ;
        RECT 693.820 1113.040 693.960 1124.450 ;
        RECT 694.440 1124.170 694.700 1124.490 ;
        RECT 697.685 1124.470 697.945 1124.790 ;
        RECT 698.655 1124.510 698.795 1126.825 ;
        RECT 694.440 1116.360 694.580 1124.170 ;
        RECT 694.360 1115.510 694.680 1116.360 ;
        RECT 697.685 1113.300 697.825 1124.470 ;
        RECT 698.655 1124.190 698.915 1124.510 ;
        RECT 699.800 1124.210 699.940 1126.825 ;
        RECT 698.655 1116.100 698.795 1124.190 ;
        RECT 699.800 1123.890 700.060 1124.210 ;
        RECT 700.420 1123.930 700.560 1126.825 ;
        RECT 703.665 1124.230 703.805 1126.825 ;
        RECT 698.160 1115.780 699.250 1116.100 ;
        RECT 693.530 1112.720 694.620 1113.040 ;
        RECT 697.590 1112.450 697.910 1113.300 ;
        RECT 699.800 1113.040 699.940 1123.890 ;
        RECT 700.420 1123.610 700.680 1123.930 ;
        RECT 703.665 1123.910 703.925 1124.230 ;
        RECT 704.635 1123.950 704.775 1126.825 ;
        RECT 700.420 1116.360 700.560 1123.610 ;
        RECT 700.340 1115.510 700.660 1116.360 ;
        RECT 703.665 1113.300 703.805 1123.910 ;
        RECT 704.515 1123.630 704.775 1123.950 ;
        RECT 704.635 1116.100 704.775 1123.630 ;
        RECT 705.780 1123.650 705.920 1126.825 ;
        RECT 705.780 1123.330 706.040 1123.650 ;
        RECT 706.400 1123.370 706.540 1126.825 ;
        RECT 709.645 1123.670 709.785 1126.825 ;
        RECT 704.140 1115.780 705.230 1116.100 ;
        RECT 699.510 1112.720 700.600 1113.040 ;
        RECT 703.570 1112.450 703.890 1113.300 ;
        RECT 705.780 1113.040 705.920 1123.330 ;
        RECT 706.400 1123.050 706.660 1123.370 ;
        RECT 709.645 1123.350 709.905 1123.670 ;
        RECT 710.615 1123.390 710.755 1126.825 ;
        RECT 706.400 1116.360 706.540 1123.050 ;
        RECT 706.320 1115.510 706.640 1116.360 ;
        RECT 709.645 1113.300 709.785 1123.350 ;
        RECT 710.615 1123.070 710.875 1123.390 ;
        RECT 711.760 1123.090 711.900 1126.825 ;
        RECT 710.615 1116.100 710.755 1123.070 ;
        RECT 711.760 1122.770 712.020 1123.090 ;
        RECT 712.380 1122.810 712.520 1126.825 ;
        RECT 715.625 1123.110 715.765 1126.825 ;
        RECT 710.120 1115.780 711.210 1116.100 ;
        RECT 705.490 1112.720 706.580 1113.040 ;
        RECT 709.550 1112.450 709.870 1113.300 ;
        RECT 711.760 1113.040 711.900 1122.770 ;
        RECT 712.380 1122.490 712.640 1122.810 ;
        RECT 715.625 1122.790 715.885 1123.110 ;
        RECT 716.595 1122.830 716.735 1126.825 ;
        RECT 712.380 1116.360 712.520 1122.490 ;
        RECT 712.300 1115.510 712.620 1116.360 ;
        RECT 715.625 1113.300 715.765 1122.790 ;
        RECT 716.475 1122.510 716.735 1122.830 ;
        RECT 716.595 1116.100 716.735 1122.510 ;
        RECT 717.740 1122.530 717.880 1126.825 ;
        RECT 717.740 1122.210 718.000 1122.530 ;
        RECT 718.360 1122.250 718.500 1126.825 ;
        RECT 721.605 1122.550 721.745 1126.825 ;
        RECT 716.100 1115.780 717.190 1116.100 ;
        RECT 711.470 1112.720 712.560 1113.040 ;
        RECT 715.530 1112.450 715.850 1113.300 ;
        RECT 717.740 1113.040 717.880 1122.210 ;
        RECT 718.360 1121.930 718.620 1122.250 ;
        RECT 721.605 1122.230 721.865 1122.550 ;
        RECT 722.575 1122.270 722.715 1126.825 ;
        RECT 718.360 1116.360 718.500 1121.930 ;
        RECT 718.280 1115.510 718.600 1116.360 ;
        RECT 721.605 1113.300 721.745 1122.230 ;
        RECT 722.575 1121.950 722.835 1122.270 ;
        RECT 723.720 1121.970 723.860 1126.825 ;
        RECT 722.575 1116.100 722.715 1121.950 ;
        RECT 723.720 1121.650 723.980 1121.970 ;
        RECT 724.340 1121.690 724.480 1126.825 ;
        RECT 727.585 1121.990 727.725 1126.825 ;
        RECT 722.080 1115.780 723.170 1116.100 ;
        RECT 717.450 1112.720 718.540 1113.040 ;
        RECT 721.510 1112.450 721.830 1113.300 ;
        RECT 723.720 1113.040 723.860 1121.650 ;
        RECT 724.340 1121.370 724.600 1121.690 ;
        RECT 727.585 1121.670 727.845 1121.990 ;
        RECT 728.555 1121.710 728.695 1126.825 ;
        RECT 724.340 1116.360 724.480 1121.370 ;
        RECT 724.260 1115.510 724.580 1116.360 ;
        RECT 727.585 1113.300 727.725 1121.670 ;
        RECT 728.555 1121.390 728.815 1121.710 ;
        RECT 729.700 1121.410 729.840 1126.825 ;
        RECT 733.565 1121.430 733.705 1126.825 ;
        RECT 728.555 1116.100 728.695 1121.390 ;
        RECT 729.700 1121.090 729.960 1121.410 ;
        RECT 733.565 1121.110 733.825 1121.430 ;
        RECT 740.515 1121.150 740.655 1126.825 ;
        RECT 728.060 1115.780 729.150 1116.100 ;
        RECT 723.430 1112.720 724.520 1113.040 ;
        RECT 727.490 1112.450 727.810 1113.300 ;
        RECT 729.700 1113.040 729.840 1121.090 ;
        RECT 733.565 1113.300 733.705 1121.110 ;
        RECT 740.515 1120.830 740.775 1121.150 ;
        RECT 745.525 1120.870 745.665 1126.825 ;
        RECT 740.515 1116.100 740.655 1120.830 ;
        RECT 745.525 1120.550 745.785 1120.870 ;
        RECT 746.495 1120.590 746.635 1126.825 ;
        RECT 740.020 1115.780 741.110 1116.100 ;
        RECT 745.525 1113.300 745.665 1120.550 ;
        RECT 746.495 1120.270 746.755 1120.590 ;
        RECT 751.505 1120.310 751.645 1126.825 ;
        RECT 746.495 1116.100 746.635 1120.270 ;
        RECT 751.505 1119.990 751.765 1120.310 ;
        RECT 752.475 1120.030 752.615 1126.825 ;
        RECT 746.000 1115.780 747.090 1116.100 ;
        RECT 751.505 1113.300 751.645 1119.990 ;
        RECT 752.355 1119.710 752.615 1120.030 ;
        RECT 752.475 1116.100 752.615 1119.710 ;
        RECT 757.485 1119.750 757.625 1126.825 ;
        RECT 757.485 1119.430 757.745 1119.750 ;
        RECT 758.455 1119.470 758.595 1126.825 ;
        RECT 751.980 1115.780 753.070 1116.100 ;
        RECT 757.485 1113.300 757.625 1119.430 ;
        RECT 758.455 1119.150 758.715 1119.470 ;
        RECT 763.465 1119.190 763.605 1126.825 ;
        RECT 758.455 1116.100 758.595 1119.150 ;
        RECT 763.465 1118.870 763.725 1119.190 ;
        RECT 764.435 1118.910 764.575 1126.825 ;
        RECT 757.960 1115.780 759.050 1116.100 ;
        RECT 763.465 1113.300 763.605 1118.870 ;
        RECT 764.315 1118.590 764.575 1118.910 ;
        RECT 764.435 1116.100 764.575 1118.590 ;
        RECT 769.445 1118.630 769.585 1126.825 ;
        RECT 769.445 1118.310 769.705 1118.630 ;
        RECT 770.415 1118.350 770.555 1126.825 ;
        RECT 1970.520 1126.550 1970.780 1126.870 ;
        RECT 1975.880 1126.590 1976.020 1126.965 ;
        RECT 763.940 1115.780 765.030 1116.100 ;
        RECT 769.445 1114.240 769.585 1118.310 ;
        RECT 770.415 1118.030 770.675 1118.350 ;
        RECT 770.415 1116.100 770.555 1118.030 ;
        RECT 1970.520 1116.360 1970.660 1126.550 ;
        RECT 1975.880 1126.270 1976.140 1126.590 ;
        RECT 1976.500 1126.310 1976.640 1126.965 ;
        RECT 769.920 1115.780 771.010 1116.100 ;
        RECT 1970.440 1115.510 1970.760 1116.360 ;
        RECT 769.445 1114.100 770.220 1114.240 ;
        RECT 729.410 1112.720 730.500 1113.040 ;
        RECT 733.470 1112.450 733.790 1113.300 ;
        RECT 745.430 1112.450 745.750 1113.300 ;
        RECT 751.410 1112.450 751.730 1113.300 ;
        RECT 757.390 1112.450 757.710 1113.300 ;
        RECT 763.370 1112.450 763.690 1113.300 ;
        RECT 770.080 1113.040 770.220 1114.100 ;
        RECT 1975.880 1113.040 1976.020 1126.270 ;
        RECT 1976.500 1125.990 1976.760 1126.310 ;
        RECT 1981.860 1126.030 1982.000 1126.965 ;
        RECT 1976.500 1116.360 1976.640 1125.990 ;
        RECT 1981.860 1125.710 1982.120 1126.030 ;
        RECT 1982.480 1125.750 1982.620 1126.965 ;
        RECT 1976.420 1115.510 1976.740 1116.360 ;
        RECT 1981.860 1113.040 1982.000 1125.710 ;
        RECT 1982.480 1125.430 1982.740 1125.750 ;
        RECT 1987.840 1125.470 1987.980 1126.965 ;
        RECT 1982.480 1116.360 1982.620 1125.430 ;
        RECT 1987.840 1125.150 1988.100 1125.470 ;
        RECT 1988.460 1125.190 1988.600 1126.965 ;
        RECT 1982.400 1115.510 1982.720 1116.360 ;
        RECT 1987.840 1113.040 1987.980 1125.150 ;
        RECT 1988.460 1124.870 1988.720 1125.190 ;
        RECT 1993.820 1124.910 1993.960 1126.965 ;
        RECT 1988.460 1116.360 1988.600 1124.870 ;
        RECT 1993.820 1124.590 1994.080 1124.910 ;
        RECT 1994.440 1124.630 1994.580 1126.965 ;
        RECT 1988.380 1115.510 1988.700 1116.360 ;
        RECT 1993.820 1113.040 1993.960 1124.590 ;
        RECT 1994.440 1124.310 1994.700 1124.630 ;
        RECT 1999.800 1124.350 1999.940 1126.965 ;
        RECT 1994.440 1116.360 1994.580 1124.310 ;
        RECT 1999.800 1124.030 2000.060 1124.350 ;
        RECT 2000.420 1124.070 2000.560 1126.965 ;
        RECT 1994.360 1115.510 1994.680 1116.360 ;
        RECT 1999.800 1113.040 1999.940 1124.030 ;
        RECT 2000.420 1123.750 2000.680 1124.070 ;
        RECT 2005.780 1123.790 2005.920 1126.965 ;
        RECT 2000.420 1116.360 2000.560 1123.750 ;
        RECT 2005.780 1123.470 2006.040 1123.790 ;
        RECT 2006.400 1123.510 2006.540 1126.965 ;
        RECT 2000.340 1115.510 2000.660 1116.360 ;
        RECT 2005.780 1113.040 2005.920 1123.470 ;
        RECT 2006.400 1123.190 2006.660 1123.510 ;
        RECT 2011.760 1123.230 2011.900 1126.965 ;
        RECT 2006.400 1116.360 2006.540 1123.190 ;
        RECT 2011.760 1122.910 2012.020 1123.230 ;
        RECT 2012.380 1122.950 2012.520 1126.965 ;
        RECT 2006.320 1115.510 2006.640 1116.360 ;
        RECT 2011.760 1113.040 2011.900 1122.910 ;
        RECT 2012.380 1122.630 2012.640 1122.950 ;
        RECT 2017.740 1122.670 2017.880 1126.965 ;
        RECT 2012.380 1116.360 2012.520 1122.630 ;
        RECT 2017.740 1122.350 2018.000 1122.670 ;
        RECT 2018.360 1122.390 2018.500 1126.965 ;
        RECT 2012.300 1115.510 2012.620 1116.360 ;
        RECT 2017.740 1113.040 2017.880 1122.350 ;
        RECT 2018.360 1122.070 2018.620 1122.390 ;
        RECT 2023.720 1122.110 2023.860 1126.965 ;
        RECT 2018.360 1116.360 2018.500 1122.070 ;
        RECT 2023.720 1121.790 2023.980 1122.110 ;
        RECT 2024.340 1121.830 2024.480 1126.965 ;
        RECT 2018.280 1115.510 2018.600 1116.360 ;
        RECT 2023.720 1113.040 2023.860 1121.790 ;
        RECT 2024.340 1121.510 2024.600 1121.830 ;
        RECT 2029.700 1121.550 2029.840 1126.965 ;
        RECT 2024.340 1116.360 2024.480 1121.510 ;
        RECT 2029.700 1121.230 2029.960 1121.550 ;
        RECT 2036.300 1121.270 2036.440 1126.965 ;
        RECT 2024.260 1115.510 2024.580 1116.360 ;
        RECT 2029.700 1113.040 2029.840 1121.230 ;
        RECT 2036.300 1120.950 2036.560 1121.270 ;
        RECT 2041.660 1120.990 2041.800 1126.965 ;
        RECT 2036.300 1116.360 2036.440 1120.950 ;
        RECT 2041.660 1120.670 2041.920 1120.990 ;
        RECT 2042.280 1120.710 2042.420 1126.965 ;
        RECT 2036.220 1115.510 2036.540 1116.360 ;
        RECT 2041.660 1113.040 2041.800 1120.670 ;
        RECT 2042.280 1120.390 2042.540 1120.710 ;
        RECT 2047.640 1120.430 2047.780 1126.965 ;
        RECT 2042.280 1116.360 2042.420 1120.390 ;
        RECT 2047.640 1120.110 2047.900 1120.430 ;
        RECT 2048.260 1120.150 2048.400 1126.965 ;
        RECT 2042.200 1115.510 2042.520 1116.360 ;
        RECT 2047.640 1113.040 2047.780 1120.110 ;
        RECT 2048.260 1119.830 2048.520 1120.150 ;
        RECT 2053.620 1119.870 2053.760 1126.965 ;
        RECT 2048.260 1116.360 2048.400 1119.830 ;
        RECT 2053.620 1119.550 2053.880 1119.870 ;
        RECT 2054.240 1119.590 2054.380 1126.965 ;
        RECT 2048.180 1115.510 2048.500 1116.360 ;
        RECT 2053.620 1113.040 2053.760 1119.550 ;
        RECT 2054.240 1119.270 2054.500 1119.590 ;
        RECT 2059.600 1119.310 2059.740 1126.965 ;
        RECT 2054.240 1116.360 2054.380 1119.270 ;
        RECT 2059.600 1118.990 2059.860 1119.310 ;
        RECT 2060.220 1119.030 2060.360 1126.965 ;
        RECT 2054.160 1115.510 2054.480 1116.360 ;
        RECT 2059.600 1113.040 2059.740 1118.990 ;
        RECT 2060.220 1118.710 2060.480 1119.030 ;
        RECT 2065.580 1118.750 2065.720 1126.965 ;
        RECT 2060.220 1116.360 2060.360 1118.710 ;
        RECT 2065.580 1118.430 2065.840 1118.750 ;
        RECT 2066.200 1118.470 2066.340 1126.965 ;
        RECT 2060.140 1115.510 2060.460 1116.360 ;
        RECT 2065.580 1114.170 2065.720 1118.430 ;
        RECT 2066.200 1118.150 2066.460 1118.470 ;
        RECT 2066.200 1116.360 2066.340 1118.150 ;
        RECT 2066.120 1115.510 2066.440 1116.360 ;
        RECT 2065.580 1114.030 2066.355 1114.170 ;
        RECT 2066.215 1113.300 2066.355 1114.030 ;
        RECT 769.420 1112.720 770.510 1113.040 ;
        RECT 1975.590 1112.720 1976.680 1113.040 ;
        RECT 1981.570 1112.720 1982.660 1113.040 ;
        RECT 1987.550 1112.720 1988.640 1113.040 ;
        RECT 1993.530 1112.720 1994.620 1113.040 ;
        RECT 1999.510 1112.720 2000.600 1113.040 ;
        RECT 2005.490 1112.720 2006.580 1113.040 ;
        RECT 2011.470 1112.720 2012.560 1113.040 ;
        RECT 2017.450 1112.720 2018.540 1113.040 ;
        RECT 2023.430 1112.720 2024.520 1113.040 ;
        RECT 2029.410 1112.720 2030.500 1113.040 ;
        RECT 2041.370 1112.720 2042.460 1113.040 ;
        RECT 2047.350 1112.720 2048.440 1113.040 ;
        RECT 2053.330 1112.720 2054.420 1113.040 ;
        RECT 2059.310 1112.720 2060.400 1113.040 ;
        RECT 2066.130 1112.450 2066.450 1113.300 ;
  END
END gpio_signal_buffering_alt
END LIBRARY

