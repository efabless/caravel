magic
tech sky130A
magscale 1 2
timestamp 1665680517
<< nwell >>
rect 1066 29637 422870 30203
rect 1066 28549 422870 29115
rect 1066 27461 422870 28027
rect 1066 26373 422870 26939
rect 1066 25285 422870 25851
rect 1066 24197 422870 24763
rect 1066 23109 422870 23675
rect 1066 22021 422870 22587
rect 1066 20933 422870 21499
rect 1066 19845 422870 20411
rect 1066 18757 422870 19323
rect 1066 17669 422870 18235
rect 1066 16581 422870 17147
rect 1066 15493 133714 16059
rect 1066 14405 133714 14971
rect 1066 13317 133714 13883
rect 1066 12229 133714 12795
rect 1066 11386 133714 11707
rect 1066 11141 64070 11386
rect 1066 10053 64070 10619
rect 1066 8965 64070 9531
rect 1066 7877 64070 8443
rect 1066 6789 64070 7355
rect 1066 5701 64070 6267
rect 1066 4613 422870 5179
rect 1066 3525 422870 4091
rect 1066 2437 422870 3003
rect 1066 1349 422870 1915
<< obsli1 >>
rect 1104 1071 422832 30481
<< obsm1 >>
rect 1104 8 422832 30728
<< metal2 >>
rect 9126 31200 9182 32400
rect 9954 31200 10010 32400
rect 10782 31200 10838 32400
rect 11610 31200 11666 32400
rect 12438 31200 12494 32400
rect 13266 31200 13322 32400
rect 14094 31200 14150 32400
rect 14922 31200 14978 32400
rect 15750 31200 15806 32400
rect 16578 31200 16634 32400
rect 17406 31200 17462 32400
rect 18234 31200 18290 32400
rect 19062 31200 19118 32400
rect 19890 31200 19946 32400
rect 20718 31200 20774 32400
rect 21546 31200 21602 32400
rect 22374 31200 22430 32400
rect 23202 31200 23258 32400
rect 24030 31200 24086 32400
rect 24858 31200 24914 32400
rect 25686 31200 25742 32400
rect 26514 31200 26570 32400
rect 27342 31200 27398 32400
rect 28170 31200 28226 32400
rect 28998 31200 29054 32400
rect 29826 31200 29882 32400
rect 30654 31200 30710 32400
rect 31482 31200 31538 32400
rect 32310 31200 32366 32400
rect 33138 31200 33194 32400
rect 33966 31200 34022 32400
rect 34794 31200 34850 32400
rect 35622 31200 35678 32400
rect 36450 31200 36506 32400
rect 37278 31200 37334 32400
rect 38106 31200 38162 32400
rect 38934 31200 38990 32400
rect 39762 31200 39818 32400
rect 40590 31200 40646 32400
rect 41418 31200 41474 32400
rect 42246 31200 42302 32400
rect 43074 31200 43130 32400
rect 43902 31200 43958 32400
rect 44730 31200 44786 32400
rect 45558 31200 45614 32400
rect 46386 31200 46442 32400
rect 47214 31200 47270 32400
rect 48042 31200 48098 32400
rect 48870 31200 48926 32400
rect 49698 31200 49754 32400
rect 50526 31200 50582 32400
rect 51354 31200 51410 32400
rect 52182 31200 52238 32400
rect 53010 31200 53066 32400
rect 53838 31200 53894 32400
rect 54666 31200 54722 32400
rect 55494 31200 55550 32400
rect 56322 31200 56378 32400
rect 57150 31200 57206 32400
rect 57978 31200 58034 32400
rect 58806 31200 58862 32400
rect 59634 31200 59690 32400
rect 60462 31200 60518 32400
rect 61290 31200 61346 32400
rect 62118 31200 62174 32400
rect 62946 31200 63002 32400
rect 63774 31200 63830 32400
rect 64602 31200 64658 32400
rect 65430 31200 65486 32400
rect 66258 31200 66314 32400
rect 67086 31200 67142 32400
rect 67914 31200 67970 32400
rect 68742 31200 68798 32400
rect 69570 31200 69626 32400
rect 70398 31200 70454 32400
rect 71226 31200 71282 32400
rect 72054 31200 72110 32400
rect 72882 31200 72938 32400
rect 73710 31200 73766 32400
rect 74538 31200 74594 32400
rect 75366 31200 75422 32400
rect 76194 31200 76250 32400
rect 77022 31200 77078 32400
rect 77850 31200 77906 32400
rect 78678 31200 78734 32400
rect 79506 31200 79562 32400
rect 80334 31200 80390 32400
rect 81162 31200 81218 32400
rect 81990 31200 82046 32400
rect 82818 31200 82874 32400
rect 83646 31200 83702 32400
rect 84474 31200 84530 32400
rect 85302 31200 85358 32400
rect 86130 31200 86186 32400
rect 86958 31200 87014 32400
rect 87786 31200 87842 32400
rect 88614 31200 88670 32400
rect 89442 31200 89498 32400
rect 90270 31200 90326 32400
rect 91098 31200 91154 32400
rect 91926 31200 91982 32400
rect 92754 31200 92810 32400
rect 93582 31200 93638 32400
rect 94410 31200 94466 32400
rect 95238 31200 95294 32400
rect 96066 31200 96122 32400
rect 96894 31200 96950 32400
rect 97722 31200 97778 32400
rect 98550 31200 98606 32400
rect 99378 31200 99434 32400
rect 100206 31200 100262 32400
rect 101034 31200 101090 32400
rect 101862 31200 101918 32400
rect 102690 31200 102746 32400
rect 103518 31200 103574 32400
rect 104346 31200 104402 32400
rect 105174 31200 105230 32400
rect 106002 31200 106058 32400
rect 106830 31200 106886 32400
rect 107658 31200 107714 32400
rect 108486 31200 108542 32400
rect 109314 31200 109370 32400
rect 110142 31200 110198 32400
rect 110970 31200 111026 32400
rect 111798 31200 111854 32400
rect 112626 31200 112682 32400
rect 113454 31200 113510 32400
rect 114282 31200 114338 32400
rect 115110 31200 115166 32400
rect 115938 31200 115994 32400
rect 116766 31200 116822 32400
rect 117594 31200 117650 32400
rect 118422 31200 118478 32400
rect 119250 31200 119306 32400
rect 120078 31200 120134 32400
rect 120906 31200 120962 32400
rect 121734 31200 121790 32400
rect 122562 31200 122618 32400
rect 123390 31200 123446 32400
rect 124218 31200 124274 32400
rect 125046 31200 125102 32400
rect 125874 31200 125930 32400
rect 126702 31200 126758 32400
rect 127530 31200 127586 32400
rect 128358 31200 128414 32400
rect 129186 31200 129242 32400
rect 130014 31200 130070 32400
rect 130842 31200 130898 32400
rect 131670 31200 131726 32400
rect 132498 31200 132554 32400
rect 133326 31200 133382 32400
rect 134154 31200 134210 32400
rect 134982 31200 135038 32400
rect 135810 31200 135866 32400
rect 136638 31200 136694 32400
rect 137466 31200 137522 32400
rect 138294 31200 138350 32400
rect 139122 31200 139178 32400
rect 139950 31200 140006 32400
rect 140778 31200 140834 32400
rect 141606 31200 141662 32400
rect 142434 31200 142490 32400
rect 143262 31200 143318 32400
rect 144090 31200 144146 32400
rect 144918 31200 144974 32400
rect 145746 31200 145802 32400
rect 146574 31200 146630 32400
rect 147402 31200 147458 32400
rect 148230 31200 148286 32400
rect 149058 31200 149114 32400
rect 149886 31200 149942 32400
rect 150714 31200 150770 32400
rect 151542 31200 151598 32400
rect 152370 31200 152426 32400
rect 153198 31200 153254 32400
rect 154026 31200 154082 32400
rect 154854 31200 154910 32400
rect 155682 31200 155738 32400
rect 156510 31200 156566 32400
rect 157338 31200 157394 32400
rect 158166 31200 158222 32400
rect 158994 31200 159050 32400
rect 159822 31200 159878 32400
rect 160650 31200 160706 32400
rect 161478 31200 161534 32400
rect 162306 31200 162362 32400
rect 163134 31200 163190 32400
rect 163962 31200 164018 32400
rect 164790 31200 164846 32400
rect 165618 31200 165674 32400
rect 166446 31200 166502 32400
rect 167274 31200 167330 32400
rect 168102 31200 168158 32400
rect 168930 31200 168986 32400
rect 169758 31200 169814 32400
rect 170586 31200 170642 32400
rect 171414 31200 171470 32400
rect 172242 31200 172298 32400
rect 173070 31200 173126 32400
rect 173898 31200 173954 32400
rect 174726 31200 174782 32400
rect 175554 31200 175610 32400
rect 176382 31200 176438 32400
rect 177210 31200 177266 32400
rect 178038 31200 178094 32400
rect 178866 31200 178922 32400
rect 179694 31200 179750 32400
rect 180522 31200 180578 32400
rect 181350 31200 181406 32400
rect 182178 31200 182234 32400
rect 183006 31200 183062 32400
rect 183834 31200 183890 32400
rect 184662 31200 184718 32400
rect 185490 31200 185546 32400
rect 186318 31200 186374 32400
rect 187146 31200 187202 32400
rect 187974 31200 188030 32400
rect 188802 31200 188858 32400
rect 189630 31200 189686 32400
rect 190458 31200 190514 32400
rect 191286 31200 191342 32400
rect 192114 31200 192170 32400
rect 192942 31200 192998 32400
rect 193770 31200 193826 32400
rect 194598 31200 194654 32400
rect 195426 31200 195482 32400
rect 196254 31200 196310 32400
rect 197082 31200 197138 32400
rect 197910 31200 197966 32400
rect 198738 31200 198794 32400
rect 199566 31200 199622 32400
rect 200394 31200 200450 32400
rect 201222 31200 201278 32400
rect 202050 31200 202106 32400
rect 202878 31200 202934 32400
rect 203706 31200 203762 32400
rect 204534 31200 204590 32400
rect 205362 31200 205418 32400
rect 206190 31200 206246 32400
rect 207018 31200 207074 32400
rect 207846 31200 207902 32400
rect 208674 31200 208730 32400
rect 209502 31200 209558 32400
rect 210330 31200 210386 32400
rect 211158 31200 211214 32400
rect 211986 31200 212042 32400
rect 212814 31200 212870 32400
rect 213642 31200 213698 32400
rect 214470 31200 214526 32400
rect 215298 31200 215354 32400
rect 216126 31200 216182 32400
rect 216954 31200 217010 32400
rect 217782 31200 217838 32400
rect 218610 31200 218666 32400
rect 219438 31200 219494 32400
rect 220266 31200 220322 32400
rect 221094 31200 221150 32400
rect 221922 31200 221978 32400
rect 222750 31200 222806 32400
rect 223578 31200 223634 32400
rect 224406 31200 224462 32400
rect 225234 31200 225290 32400
rect 226062 31200 226118 32400
rect 226890 31200 226946 32400
rect 227718 31200 227774 32400
rect 228546 31200 228602 32400
rect 229374 31200 229430 32400
rect 230202 31200 230258 32400
rect 231030 31200 231086 32400
rect 231858 31200 231914 32400
rect 232686 31200 232742 32400
rect 233514 31200 233570 32400
rect 234342 31200 234398 32400
rect 235170 31200 235226 32400
rect 235998 31200 236054 32400
rect 236826 31200 236882 32400
rect 237654 31200 237710 32400
rect 238482 31200 238538 32400
rect 239310 31200 239366 32400
rect 240138 31200 240194 32400
rect 240966 31200 241022 32400
rect 241794 31200 241850 32400
rect 242622 31200 242678 32400
rect 243450 31200 243506 32400
rect 244278 31200 244334 32400
rect 245106 31200 245162 32400
rect 245934 31200 245990 32400
rect 246762 31200 246818 32400
rect 247590 31200 247646 32400
rect 248418 31200 248474 32400
rect 249246 31200 249302 32400
rect 250074 31200 250130 32400
rect 250902 31200 250958 32400
rect 251730 31200 251786 32400
rect 252558 31200 252614 32400
rect 253386 31200 253442 32400
rect 254214 31200 254270 32400
rect 255042 31200 255098 32400
rect 255870 31200 255926 32400
rect 256698 31200 256754 32400
rect 257526 31200 257582 32400
rect 258354 31200 258410 32400
rect 259182 31200 259238 32400
rect 260010 31200 260066 32400
rect 260838 31200 260894 32400
rect 261666 31200 261722 32400
rect 262494 31200 262550 32400
rect 263322 31200 263378 32400
rect 264150 31200 264206 32400
rect 264978 31200 265034 32400
rect 265806 31200 265862 32400
rect 266634 31200 266690 32400
rect 267462 31200 267518 32400
rect 268290 31200 268346 32400
rect 269118 31200 269174 32400
rect 269946 31200 270002 32400
rect 270774 31200 270830 32400
rect 271602 31200 271658 32400
rect 272430 31200 272486 32400
rect 273258 31200 273314 32400
rect 274086 31200 274142 32400
rect 274914 31200 274970 32400
rect 275742 31200 275798 32400
rect 276570 31200 276626 32400
rect 277398 31200 277454 32400
rect 278226 31200 278282 32400
rect 279054 31200 279110 32400
rect 279882 31200 279938 32400
rect 280710 31200 280766 32400
rect 281538 31200 281594 32400
rect 282366 31200 282422 32400
rect 283194 31200 283250 32400
rect 284022 31200 284078 32400
rect 284850 31200 284906 32400
rect 285678 31200 285734 32400
rect 286506 31200 286562 32400
rect 287334 31200 287390 32400
rect 288162 31200 288218 32400
rect 288990 31200 289046 32400
rect 289818 31200 289874 32400
rect 290646 31200 290702 32400
rect 291474 31200 291530 32400
rect 292302 31200 292358 32400
rect 293130 31200 293186 32400
rect 293958 31200 294014 32400
rect 294786 31200 294842 32400
rect 295614 31200 295670 32400
rect 296442 31200 296498 32400
rect 297270 31200 297326 32400
rect 298098 31200 298154 32400
rect 298926 31200 298982 32400
rect 299754 31200 299810 32400
rect 300582 31200 300638 32400
rect 301410 31200 301466 32400
rect 302238 31200 302294 32400
rect 303066 31200 303122 32400
rect 303894 31200 303950 32400
rect 304722 31200 304778 32400
rect 305550 31200 305606 32400
rect 306378 31200 306434 32400
rect 307206 31200 307262 32400
rect 308034 31200 308090 32400
rect 308862 31200 308918 32400
rect 309690 31200 309746 32400
rect 310518 31200 310574 32400
rect 311346 31200 311402 32400
rect 312174 31200 312230 32400
rect 313002 31200 313058 32400
rect 313830 31200 313886 32400
rect 314658 31200 314714 32400
rect 315486 31200 315542 32400
rect 316314 31200 316370 32400
rect 317142 31200 317198 32400
rect 317970 31200 318026 32400
rect 318798 31200 318854 32400
rect 319626 31200 319682 32400
rect 320454 31200 320510 32400
rect 321282 31200 321338 32400
rect 322110 31200 322166 32400
rect 322938 31200 322994 32400
rect 323766 31200 323822 32400
rect 324594 31200 324650 32400
rect 325422 31200 325478 32400
rect 326250 31200 326306 32400
rect 327078 31200 327134 32400
rect 327906 31200 327962 32400
rect 328734 31200 328790 32400
rect 329562 31200 329618 32400
rect 330390 31200 330446 32400
rect 331218 31200 331274 32400
rect 332046 31200 332102 32400
rect 332874 31200 332930 32400
rect 333702 31200 333758 32400
rect 334530 31200 334586 32400
rect 335358 31200 335414 32400
rect 336186 31200 336242 32400
rect 337014 31200 337070 32400
rect 337842 31200 337898 32400
rect 338670 31200 338726 32400
rect 339498 31200 339554 32400
rect 340326 31200 340382 32400
rect 341154 31200 341210 32400
rect 341982 31200 342038 32400
rect 342810 31200 342866 32400
rect 343638 31200 343694 32400
rect 344466 31200 344522 32400
rect 345294 31200 345350 32400
rect 346122 31200 346178 32400
rect 346950 31200 347006 32400
rect 347778 31200 347834 32400
rect 348606 31200 348662 32400
rect 349434 31200 349490 32400
rect 350262 31200 350318 32400
rect 351090 31200 351146 32400
rect 351918 31200 351974 32400
rect 352746 31200 352802 32400
rect 353574 31200 353630 32400
rect 354402 31200 354458 32400
rect 355230 31200 355286 32400
rect 356058 31200 356114 32400
rect 356886 31200 356942 32400
rect 357714 31200 357770 32400
rect 358542 31200 358598 32400
rect 359370 31200 359426 32400
rect 360198 31200 360254 32400
rect 361026 31200 361082 32400
rect 361854 31200 361910 32400
rect 362682 31200 362738 32400
rect 363510 31200 363566 32400
rect 364338 31200 364394 32400
rect 365166 31200 365222 32400
rect 365994 31200 366050 32400
rect 366822 31200 366878 32400
rect 367650 31200 367706 32400
rect 368478 31200 368534 32400
rect 369306 31200 369362 32400
rect 370134 31200 370190 32400
rect 370962 31200 371018 32400
rect 371790 31200 371846 32400
rect 372618 31200 372674 32400
rect 373446 31200 373502 32400
rect 374274 31200 374330 32400
rect 375102 31200 375158 32400
rect 375930 31200 375986 32400
rect 376758 31200 376814 32400
rect 377586 31200 377642 32400
rect 378414 31200 378470 32400
rect 379242 31200 379298 32400
rect 380070 31200 380126 32400
rect 380898 31200 380954 32400
rect 381726 31200 381782 32400
rect 382554 31200 382610 32400
rect 383382 31200 383438 32400
rect 384210 31200 384266 32400
rect 385038 31200 385094 32400
rect 385866 31200 385922 32400
rect 386694 31200 386750 32400
rect 387522 31200 387578 32400
rect 388350 31200 388406 32400
rect 389178 31200 389234 32400
rect 390006 31200 390062 32400
rect 390834 31200 390890 32400
rect 391662 31200 391718 32400
rect 392490 31200 392546 32400
rect 393318 31200 393374 32400
rect 394146 31200 394202 32400
rect 394974 31200 395030 32400
rect 395802 31200 395858 32400
rect 396630 31200 396686 32400
rect 397458 31200 397514 32400
rect 398286 31200 398342 32400
rect 399114 31200 399170 32400
rect 399942 31200 399998 32400
rect 400770 31200 400826 32400
rect 401598 31200 401654 32400
rect 402426 31200 402482 32400
rect 403254 31200 403310 32400
rect 404082 31200 404138 32400
rect 404910 31200 404966 32400
rect 405738 31200 405794 32400
rect 406566 31200 406622 32400
rect 407394 31200 407450 32400
rect 408222 31200 408278 32400
rect 409050 31200 409106 32400
rect 409878 31200 409934 32400
rect 410706 31200 410762 32400
rect 411534 31200 411590 32400
rect 412362 31200 412418 32400
rect 413190 31200 413246 32400
rect 414018 31200 414074 32400
rect 414846 31200 414902 32400
rect 16210 -400 16266 800
rect 16854 -400 16910 800
rect 17498 -400 17554 800
rect 18142 -400 18198 800
rect 18786 -400 18842 800
rect 19430 -400 19486 800
rect 20074 -400 20130 800
rect 20718 -400 20774 800
rect 21362 -400 21418 800
rect 22006 -400 22062 800
rect 22650 -400 22706 800
rect 23294 -400 23350 800
rect 23938 -400 23994 800
rect 24582 -400 24638 800
rect 25226 -400 25282 800
rect 25870 -400 25926 800
rect 26514 -400 26570 800
rect 27158 -400 27214 800
rect 27802 -400 27858 800
rect 28446 -400 28502 800
rect 29090 -400 29146 800
rect 29734 -400 29790 800
rect 30378 -400 30434 800
rect 31022 -400 31078 800
rect 31666 -400 31722 800
rect 32310 -400 32366 800
rect 32954 -400 33010 800
rect 33598 -400 33654 800
rect 34242 -400 34298 800
rect 34886 -400 34942 800
rect 35530 -400 35586 800
rect 36174 -400 36230 800
rect 36818 -400 36874 800
rect 37462 -400 37518 800
rect 38106 -400 38162 800
rect 38750 -400 38806 800
rect 39394 -400 39450 800
rect 40038 -400 40094 800
rect 40682 -400 40738 800
rect 41326 -400 41382 800
rect 41970 -400 42026 800
rect 42614 -400 42670 800
rect 43258 -400 43314 800
rect 43902 -400 43958 800
rect 44546 -400 44602 800
rect 45190 -400 45246 800
rect 45834 -400 45890 800
rect 46478 -400 46534 800
rect 47122 -400 47178 800
rect 47766 -400 47822 800
rect 48410 -400 48466 800
rect 49054 -400 49110 800
rect 49698 -400 49754 800
rect 50342 -400 50398 800
rect 50986 -400 51042 800
rect 51630 -400 51686 800
rect 52274 -400 52330 800
rect 52918 -400 52974 800
rect 53562 -400 53618 800
rect 54206 -400 54262 800
rect 54850 -400 54906 800
rect 55494 -400 55550 800
rect 56138 -400 56194 800
rect 56782 -400 56838 800
rect 57426 -400 57482 800
rect 58070 -400 58126 800
rect 58714 -400 58770 800
rect 59358 -400 59414 800
rect 60002 -400 60058 800
rect 60646 -400 60702 800
rect 61290 -400 61346 800
rect 61934 -400 61990 800
rect 62578 -400 62634 800
rect 63222 -400 63278 800
rect 63866 -400 63922 800
rect 64510 -400 64566 800
rect 65154 -400 65210 800
rect 65798 -400 65854 800
rect 66442 -400 66498 800
rect 67086 -400 67142 800
rect 67730 -400 67786 800
rect 68374 -400 68430 800
rect 69018 -400 69074 800
rect 69662 -400 69718 800
rect 70306 -400 70362 800
rect 70950 -400 71006 800
rect 71594 -400 71650 800
rect 72238 -400 72294 800
rect 72882 -400 72938 800
rect 73526 -400 73582 800
rect 74170 -400 74226 800
rect 74814 -400 74870 800
rect 75458 -400 75514 800
rect 76102 -400 76158 800
rect 76746 -400 76802 800
rect 77390 -400 77446 800
rect 78034 -400 78090 800
rect 78678 -400 78734 800
rect 79322 -400 79378 800
rect 79966 -400 80022 800
rect 80610 -400 80666 800
rect 81254 -400 81310 800
rect 81898 -400 81954 800
rect 82542 -400 82598 800
rect 83186 -400 83242 800
rect 83830 -400 83886 800
rect 84474 -400 84530 800
rect 85118 -400 85174 800
rect 85762 -400 85818 800
rect 86406 -400 86462 800
rect 87050 -400 87106 800
rect 87694 -400 87750 800
rect 88338 -400 88394 800
rect 88982 -400 89038 800
rect 89626 -400 89682 800
rect 90270 -400 90326 800
rect 90914 -400 90970 800
rect 91558 -400 91614 800
rect 92202 -400 92258 800
rect 92846 -400 92902 800
rect 93490 -400 93546 800
rect 94134 -400 94190 800
rect 94778 -400 94834 800
rect 95422 -400 95478 800
rect 96066 -400 96122 800
rect 96710 -400 96766 800
rect 97354 -400 97410 800
rect 97998 -400 98054 800
rect 98642 -400 98698 800
rect 99286 -400 99342 800
rect 99930 -400 99986 800
rect 100574 -400 100630 800
rect 101218 -400 101274 800
rect 101862 -400 101918 800
rect 102506 -400 102562 800
rect 103150 -400 103206 800
rect 103794 -400 103850 800
rect 104438 -400 104494 800
rect 105082 -400 105138 800
rect 105726 -400 105782 800
rect 106370 -400 106426 800
rect 107014 -400 107070 800
rect 107658 -400 107714 800
rect 108302 -400 108358 800
rect 108946 -400 109002 800
rect 109590 -400 109646 800
rect 110234 -400 110290 800
rect 110878 -400 110934 800
rect 111522 -400 111578 800
rect 112166 -400 112222 800
rect 112810 -400 112866 800
rect 113454 -400 113510 800
rect 114098 -400 114154 800
rect 114742 -400 114798 800
rect 115386 -400 115442 800
rect 116030 -400 116086 800
rect 116674 -400 116730 800
rect 117318 -400 117374 800
rect 117962 -400 118018 800
rect 118606 -400 118662 800
rect 119250 -400 119306 800
rect 119894 -400 119950 800
rect 120538 -400 120594 800
rect 121182 -400 121238 800
rect 121826 -400 121882 800
rect 122470 -400 122526 800
rect 123114 -400 123170 800
rect 123758 -400 123814 800
rect 124402 -400 124458 800
rect 125046 -400 125102 800
rect 125690 -400 125746 800
rect 126334 -400 126390 800
rect 126978 -400 127034 800
rect 127622 -400 127678 800
rect 128266 -400 128322 800
rect 128910 -400 128966 800
rect 129554 -400 129610 800
rect 130198 -400 130254 800
rect 130842 -400 130898 800
rect 131486 -400 131542 800
rect 132130 -400 132186 800
rect 132774 -400 132830 800
rect 133418 -400 133474 800
rect 134062 -400 134118 800
rect 134706 -400 134762 800
rect 135350 -400 135406 800
rect 135994 -400 136050 800
rect 136638 -400 136694 800
rect 137282 -400 137338 800
rect 137926 -400 137982 800
rect 138570 -400 138626 800
rect 139214 -400 139270 800
rect 139858 -400 139914 800
rect 140502 -400 140558 800
rect 141146 -400 141202 800
rect 141790 -400 141846 800
rect 142434 -400 142490 800
rect 143078 -400 143134 800
rect 143722 -400 143778 800
rect 144366 -400 144422 800
rect 145010 -400 145066 800
rect 145654 -400 145710 800
rect 146298 -400 146354 800
rect 146942 -400 146998 800
rect 147586 -400 147642 800
rect 148230 -400 148286 800
rect 148874 -400 148930 800
rect 149518 -400 149574 800
rect 150162 -400 150218 800
rect 150806 -400 150862 800
rect 151450 -400 151506 800
rect 152094 -400 152150 800
rect 152738 -400 152794 800
rect 153382 -400 153438 800
rect 154026 -400 154082 800
rect 154670 -400 154726 800
rect 155314 -400 155370 800
rect 155958 -400 156014 800
rect 156602 -400 156658 800
rect 157246 -400 157302 800
rect 157890 -400 157946 800
rect 158534 -400 158590 800
rect 159178 -400 159234 800
rect 159822 -400 159878 800
rect 160466 -400 160522 800
rect 161110 -400 161166 800
rect 161754 -400 161810 800
rect 162398 -400 162454 800
rect 163042 -400 163098 800
rect 163686 -400 163742 800
rect 164330 -400 164386 800
rect 164974 -400 165030 800
rect 165618 -400 165674 800
rect 166262 -400 166318 800
rect 166906 -400 166962 800
rect 167550 -400 167606 800
rect 168194 -400 168250 800
rect 168838 -400 168894 800
rect 169482 -400 169538 800
rect 170126 -400 170182 800
rect 170770 -400 170826 800
rect 171414 -400 171470 800
rect 172058 -400 172114 800
rect 172702 -400 172758 800
rect 173346 -400 173402 800
rect 173990 -400 174046 800
rect 174634 -400 174690 800
rect 175278 -400 175334 800
rect 175922 -400 175978 800
rect 176566 -400 176622 800
rect 177210 -400 177266 800
rect 177854 -400 177910 800
rect 178498 -400 178554 800
rect 179142 -400 179198 800
rect 179786 -400 179842 800
rect 180430 -400 180486 800
rect 181074 -400 181130 800
rect 181718 -400 181774 800
rect 182362 -400 182418 800
rect 183006 -400 183062 800
rect 183650 -400 183706 800
rect 184294 -400 184350 800
rect 184938 -400 184994 800
rect 185582 -400 185638 800
rect 186226 -400 186282 800
rect 186870 -400 186926 800
rect 187514 -400 187570 800
rect 188158 -400 188214 800
rect 188802 -400 188858 800
rect 189446 -400 189502 800
rect 190090 -400 190146 800
rect 190734 -400 190790 800
rect 191378 -400 191434 800
rect 192022 -400 192078 800
rect 192666 -400 192722 800
rect 193310 -400 193366 800
rect 193954 -400 194010 800
rect 194598 -400 194654 800
rect 195242 -400 195298 800
rect 195886 -400 195942 800
rect 196530 -400 196586 800
rect 197174 -400 197230 800
rect 197818 -400 197874 800
rect 198462 -400 198518 800
rect 199106 -400 199162 800
rect 199750 -400 199806 800
rect 200394 -400 200450 800
rect 201038 -400 201094 800
rect 201682 -400 201738 800
rect 202326 -400 202382 800
rect 202970 -400 203026 800
rect 203614 -400 203670 800
rect 204258 -400 204314 800
rect 204902 -400 204958 800
rect 205546 -400 205602 800
rect 206190 -400 206246 800
rect 206834 -400 206890 800
rect 207478 -400 207534 800
rect 208122 -400 208178 800
rect 208766 -400 208822 800
rect 209410 -400 209466 800
rect 210054 -400 210110 800
rect 210698 -400 210754 800
rect 211342 -400 211398 800
rect 211986 -400 212042 800
rect 212630 -400 212686 800
rect 213274 -400 213330 800
rect 213918 -400 213974 800
rect 214562 -400 214618 800
rect 215206 -400 215262 800
rect 215850 -400 215906 800
rect 216494 -400 216550 800
rect 217138 -400 217194 800
rect 217782 -400 217838 800
rect 218426 -400 218482 800
rect 219070 -400 219126 800
rect 219714 -400 219770 800
rect 220358 -400 220414 800
rect 221002 -400 221058 800
rect 221646 -400 221702 800
rect 222290 -400 222346 800
rect 222934 -400 222990 800
rect 223578 -400 223634 800
rect 224222 -400 224278 800
rect 224866 -400 224922 800
rect 225510 -400 225566 800
rect 226154 -400 226210 800
rect 226798 -400 226854 800
rect 227442 -400 227498 800
rect 228086 -400 228142 800
rect 228730 -400 228786 800
rect 229374 -400 229430 800
rect 230018 -400 230074 800
rect 230662 -400 230718 800
rect 231306 -400 231362 800
rect 231950 -400 232006 800
rect 232594 -400 232650 800
rect 233238 -400 233294 800
rect 233882 -400 233938 800
rect 234526 -400 234582 800
rect 235170 -400 235226 800
rect 235814 -400 235870 800
rect 236458 -400 236514 800
rect 237102 -400 237158 800
rect 237746 -400 237802 800
rect 238390 -400 238446 800
rect 239034 -400 239090 800
rect 239678 -400 239734 800
rect 240322 -400 240378 800
rect 240966 -400 241022 800
rect 241610 -400 241666 800
rect 242254 -400 242310 800
rect 242898 -400 242954 800
rect 243542 -400 243598 800
rect 244186 -400 244242 800
rect 244830 -400 244886 800
rect 245474 -400 245530 800
rect 246118 -400 246174 800
rect 246762 -400 246818 800
rect 247406 -400 247462 800
rect 248050 -400 248106 800
rect 248694 -400 248750 800
rect 249338 -400 249394 800
rect 249982 -400 250038 800
rect 250626 -400 250682 800
rect 251270 -400 251326 800
rect 251914 -400 251970 800
rect 252558 -400 252614 800
rect 253202 -400 253258 800
rect 253846 -400 253902 800
rect 254490 -400 254546 800
rect 255134 -400 255190 800
rect 255778 -400 255834 800
rect 256422 -400 256478 800
rect 257066 -400 257122 800
rect 257710 -400 257766 800
rect 258354 -400 258410 800
rect 258998 -400 259054 800
rect 259642 -400 259698 800
rect 260286 -400 260342 800
rect 260930 -400 260986 800
rect 261574 -400 261630 800
rect 262218 -400 262274 800
rect 262862 -400 262918 800
rect 263506 -400 263562 800
rect 264150 -400 264206 800
rect 264794 -400 264850 800
rect 265438 -400 265494 800
rect 266082 -400 266138 800
rect 266726 -400 266782 800
rect 267370 -400 267426 800
rect 268014 -400 268070 800
rect 268658 -400 268714 800
rect 269302 -400 269358 800
rect 269946 -400 270002 800
rect 270590 -400 270646 800
rect 271234 -400 271290 800
rect 271878 -400 271934 800
rect 272522 -400 272578 800
rect 273166 -400 273222 800
rect 273810 -400 273866 800
rect 274454 -400 274510 800
rect 275098 -400 275154 800
rect 275742 -400 275798 800
rect 276386 -400 276442 800
rect 277030 -400 277086 800
rect 277674 -400 277730 800
rect 278318 -400 278374 800
rect 278962 -400 279018 800
rect 279606 -400 279662 800
rect 280250 -400 280306 800
rect 280894 -400 280950 800
rect 281538 -400 281594 800
rect 282182 -400 282238 800
rect 282826 -400 282882 800
rect 283470 -400 283526 800
rect 284114 -400 284170 800
rect 284758 -400 284814 800
rect 285402 -400 285458 800
rect 286046 -400 286102 800
rect 286690 -400 286746 800
rect 287334 -400 287390 800
rect 287978 -400 288034 800
rect 288622 -400 288678 800
rect 289266 -400 289322 800
rect 289910 -400 289966 800
rect 290554 -400 290610 800
rect 291198 -400 291254 800
rect 291842 -400 291898 800
rect 292486 -400 292542 800
rect 293130 -400 293186 800
rect 293774 -400 293830 800
rect 294418 -400 294474 800
rect 295062 -400 295118 800
rect 295706 -400 295762 800
rect 296350 -400 296406 800
rect 296994 -400 297050 800
rect 297638 -400 297694 800
rect 298282 -400 298338 800
rect 298926 -400 298982 800
rect 299570 -400 299626 800
rect 300214 -400 300270 800
rect 300858 -400 300914 800
rect 301502 -400 301558 800
rect 302146 -400 302202 800
rect 302790 -400 302846 800
rect 303434 -400 303490 800
rect 304078 -400 304134 800
rect 304722 -400 304778 800
rect 305366 -400 305422 800
rect 306010 -400 306066 800
rect 306654 -400 306710 800
rect 307298 -400 307354 800
rect 307942 -400 307998 800
rect 308586 -400 308642 800
rect 309230 -400 309286 800
rect 309874 -400 309930 800
rect 310518 -400 310574 800
rect 311162 -400 311218 800
rect 311806 -400 311862 800
rect 312450 -400 312506 800
rect 313094 -400 313150 800
rect 313738 -400 313794 800
rect 314382 -400 314438 800
rect 315026 -400 315082 800
rect 315670 -400 315726 800
rect 316314 -400 316370 800
rect 316958 -400 317014 800
rect 317602 -400 317658 800
rect 318246 -400 318302 800
rect 318890 -400 318946 800
rect 319534 -400 319590 800
rect 320178 -400 320234 800
rect 320822 -400 320878 800
rect 321466 -400 321522 800
rect 322110 -400 322166 800
rect 322754 -400 322810 800
rect 323398 -400 323454 800
rect 324042 -400 324098 800
rect 324686 -400 324742 800
rect 325330 -400 325386 800
rect 325974 -400 326030 800
rect 326618 -400 326674 800
rect 327262 -400 327318 800
rect 327906 -400 327962 800
rect 328550 -400 328606 800
rect 329194 -400 329250 800
rect 329838 -400 329894 800
rect 330482 -400 330538 800
rect 331126 -400 331182 800
rect 331770 -400 331826 800
rect 332414 -400 332470 800
rect 333058 -400 333114 800
rect 333702 -400 333758 800
rect 334346 -400 334402 800
rect 334990 -400 335046 800
rect 335634 -400 335690 800
rect 336278 -400 336334 800
rect 336922 -400 336978 800
rect 337566 -400 337622 800
rect 338210 -400 338266 800
rect 338854 -400 338910 800
rect 339498 -400 339554 800
rect 340142 -400 340198 800
rect 340786 -400 340842 800
rect 341430 -400 341486 800
rect 342074 -400 342130 800
rect 342718 -400 342774 800
rect 343362 -400 343418 800
rect 344006 -400 344062 800
rect 344650 -400 344706 800
rect 345294 -400 345350 800
rect 345938 -400 345994 800
rect 346582 -400 346638 800
rect 347226 -400 347282 800
rect 347870 -400 347926 800
rect 348514 -400 348570 800
rect 349158 -400 349214 800
rect 349802 -400 349858 800
rect 350446 -400 350502 800
rect 351090 -400 351146 800
rect 351734 -400 351790 800
rect 352378 -400 352434 800
rect 353022 -400 353078 800
rect 353666 -400 353722 800
rect 354310 -400 354366 800
rect 354954 -400 355010 800
rect 355598 -400 355654 800
rect 356242 -400 356298 800
rect 356886 -400 356942 800
rect 357530 -400 357586 800
rect 358174 -400 358230 800
rect 358818 -400 358874 800
rect 359462 -400 359518 800
rect 360106 -400 360162 800
rect 360750 -400 360806 800
rect 361394 -400 361450 800
rect 362038 -400 362094 800
rect 362682 -400 362738 800
rect 363326 -400 363382 800
rect 363970 -400 364026 800
rect 364614 -400 364670 800
rect 365258 -400 365314 800
rect 365902 -400 365958 800
rect 366546 -400 366602 800
rect 367190 -400 367246 800
rect 367834 -400 367890 800
rect 368478 -400 368534 800
rect 369122 -400 369178 800
rect 369766 -400 369822 800
rect 370410 -400 370466 800
rect 371054 -400 371110 800
rect 371698 -400 371754 800
rect 372342 -400 372398 800
rect 372986 -400 373042 800
rect 373630 -400 373686 800
rect 374274 -400 374330 800
rect 374918 -400 374974 800
rect 375562 -400 375618 800
rect 376206 -400 376262 800
rect 376850 -400 376906 800
rect 377494 -400 377550 800
rect 378138 -400 378194 800
rect 378782 -400 378838 800
rect 379426 -400 379482 800
rect 380070 -400 380126 800
rect 380714 -400 380770 800
rect 381358 -400 381414 800
rect 382002 -400 382058 800
rect 382646 -400 382702 800
rect 383290 -400 383346 800
rect 383934 -400 383990 800
rect 384578 -400 384634 800
rect 385222 -400 385278 800
rect 385866 -400 385922 800
rect 386510 -400 386566 800
rect 387154 -400 387210 800
rect 387798 -400 387854 800
rect 388442 -400 388498 800
rect 389086 -400 389142 800
rect 389730 -400 389786 800
rect 390374 -400 390430 800
rect 391018 -400 391074 800
rect 391662 -400 391718 800
rect 392306 -400 392362 800
rect 392950 -400 393006 800
rect 393594 -400 393650 800
rect 394238 -400 394294 800
rect 394882 -400 394938 800
rect 395526 -400 395582 800
rect 396170 -400 396226 800
rect 396814 -400 396870 800
rect 397458 -400 397514 800
rect 398102 -400 398158 800
rect 398746 -400 398802 800
rect 399390 -400 399446 800
rect 400034 -400 400090 800
rect 400678 -400 400734 800
rect 401322 -400 401378 800
rect 401966 -400 402022 800
rect 402610 -400 402666 800
rect 403254 -400 403310 800
rect 403898 -400 403954 800
rect 404542 -400 404598 800
rect 405186 -400 405242 800
rect 405830 -400 405886 800
rect 406474 -400 406530 800
rect 407118 -400 407174 800
rect 407762 -400 407818 800
<< obsm2 >>
rect 5036 31144 9070 31362
rect 9238 31144 9898 31362
rect 10066 31144 10726 31362
rect 10894 31144 11554 31362
rect 11722 31144 12382 31362
rect 12550 31144 13210 31362
rect 13378 31144 14038 31362
rect 14206 31144 14866 31362
rect 15034 31144 15694 31362
rect 15862 31144 16522 31362
rect 16690 31144 17350 31362
rect 17518 31144 18178 31362
rect 18346 31144 19006 31362
rect 19174 31144 19834 31362
rect 20002 31144 20662 31362
rect 20830 31144 21490 31362
rect 21658 31144 22318 31362
rect 22486 31144 23146 31362
rect 23314 31144 23974 31362
rect 24142 31144 24802 31362
rect 24970 31144 25630 31362
rect 25798 31144 26458 31362
rect 26626 31144 27286 31362
rect 27454 31144 28114 31362
rect 28282 31144 28942 31362
rect 29110 31144 29770 31362
rect 29938 31144 30598 31362
rect 30766 31144 31426 31362
rect 31594 31144 32254 31362
rect 32422 31144 33082 31362
rect 33250 31144 33910 31362
rect 34078 31144 34738 31362
rect 34906 31144 35566 31362
rect 35734 31144 36394 31362
rect 36562 31144 37222 31362
rect 37390 31144 38050 31362
rect 38218 31144 38878 31362
rect 39046 31144 39706 31362
rect 39874 31144 40534 31362
rect 40702 31144 41362 31362
rect 41530 31144 42190 31362
rect 42358 31144 43018 31362
rect 43186 31144 43846 31362
rect 44014 31144 44674 31362
rect 44842 31144 45502 31362
rect 45670 31144 46330 31362
rect 46498 31144 47158 31362
rect 47326 31144 47986 31362
rect 48154 31144 48814 31362
rect 48982 31144 49642 31362
rect 49810 31144 50470 31362
rect 50638 31144 51298 31362
rect 51466 31144 52126 31362
rect 52294 31144 52954 31362
rect 53122 31144 53782 31362
rect 53950 31144 54610 31362
rect 54778 31144 55438 31362
rect 55606 31144 56266 31362
rect 56434 31144 57094 31362
rect 57262 31144 57922 31362
rect 58090 31144 58750 31362
rect 58918 31144 59578 31362
rect 59746 31144 60406 31362
rect 60574 31144 61234 31362
rect 61402 31144 62062 31362
rect 62230 31144 62890 31362
rect 63058 31144 63718 31362
rect 63886 31144 64546 31362
rect 64714 31144 65374 31362
rect 65542 31144 66202 31362
rect 66370 31144 67030 31362
rect 67198 31144 67858 31362
rect 68026 31144 68686 31362
rect 68854 31144 69514 31362
rect 69682 31144 70342 31362
rect 70510 31144 71170 31362
rect 71338 31144 71998 31362
rect 72166 31144 72826 31362
rect 72994 31144 73654 31362
rect 73822 31144 74482 31362
rect 74650 31144 75310 31362
rect 75478 31144 76138 31362
rect 76306 31144 76966 31362
rect 77134 31144 77794 31362
rect 77962 31144 78622 31362
rect 78790 31144 79450 31362
rect 79618 31144 80278 31362
rect 80446 31144 81106 31362
rect 81274 31144 81934 31362
rect 82102 31144 82762 31362
rect 82930 31144 83590 31362
rect 83758 31144 84418 31362
rect 84586 31144 85246 31362
rect 85414 31144 86074 31362
rect 86242 31144 86902 31362
rect 87070 31144 87730 31362
rect 87898 31144 88558 31362
rect 88726 31144 89386 31362
rect 89554 31144 90214 31362
rect 90382 31144 91042 31362
rect 91210 31144 91870 31362
rect 92038 31144 92698 31362
rect 92866 31144 93526 31362
rect 93694 31144 94354 31362
rect 94522 31144 95182 31362
rect 95350 31144 96010 31362
rect 96178 31144 96838 31362
rect 97006 31144 97666 31362
rect 97834 31144 98494 31362
rect 98662 31144 99322 31362
rect 99490 31144 100150 31362
rect 100318 31144 100978 31362
rect 101146 31144 101806 31362
rect 101974 31144 102634 31362
rect 102802 31144 103462 31362
rect 103630 31144 104290 31362
rect 104458 31144 105118 31362
rect 105286 31144 105946 31362
rect 106114 31144 106774 31362
rect 106942 31144 107602 31362
rect 107770 31144 108430 31362
rect 108598 31144 109258 31362
rect 109426 31144 110086 31362
rect 110254 31144 110914 31362
rect 111082 31144 111742 31362
rect 111910 31144 112570 31362
rect 112738 31144 113398 31362
rect 113566 31144 114226 31362
rect 114394 31144 115054 31362
rect 115222 31144 115882 31362
rect 116050 31144 116710 31362
rect 116878 31144 117538 31362
rect 117706 31144 118366 31362
rect 118534 31144 119194 31362
rect 119362 31144 120022 31362
rect 120190 31144 120850 31362
rect 121018 31144 121678 31362
rect 121846 31144 122506 31362
rect 122674 31144 123334 31362
rect 123502 31144 124162 31362
rect 124330 31144 124990 31362
rect 125158 31144 125818 31362
rect 125986 31144 126646 31362
rect 126814 31144 127474 31362
rect 127642 31144 128302 31362
rect 128470 31144 129130 31362
rect 129298 31144 129958 31362
rect 130126 31144 130786 31362
rect 130954 31144 131614 31362
rect 131782 31144 132442 31362
rect 132610 31144 133270 31362
rect 133438 31144 134098 31362
rect 134266 31144 134926 31362
rect 135094 31144 135754 31362
rect 135922 31144 136582 31362
rect 136750 31144 137410 31362
rect 137578 31144 138238 31362
rect 138406 31144 139066 31362
rect 139234 31144 139894 31362
rect 140062 31144 140722 31362
rect 140890 31144 141550 31362
rect 141718 31144 142378 31362
rect 142546 31144 143206 31362
rect 143374 31144 144034 31362
rect 144202 31144 144862 31362
rect 145030 31144 145690 31362
rect 145858 31144 146518 31362
rect 146686 31144 147346 31362
rect 147514 31144 148174 31362
rect 148342 31144 149002 31362
rect 149170 31144 149830 31362
rect 149998 31144 150658 31362
rect 150826 31144 151486 31362
rect 151654 31144 152314 31362
rect 152482 31144 153142 31362
rect 153310 31144 153970 31362
rect 154138 31144 154798 31362
rect 154966 31144 155626 31362
rect 155794 31144 156454 31362
rect 156622 31144 157282 31362
rect 157450 31144 158110 31362
rect 158278 31144 158938 31362
rect 159106 31144 159766 31362
rect 159934 31144 160594 31362
rect 160762 31144 161422 31362
rect 161590 31144 162250 31362
rect 162418 31144 163078 31362
rect 163246 31144 163906 31362
rect 164074 31144 164734 31362
rect 164902 31144 165562 31362
rect 165730 31144 166390 31362
rect 166558 31144 167218 31362
rect 167386 31144 168046 31362
rect 168214 31144 168874 31362
rect 169042 31144 169702 31362
rect 169870 31144 170530 31362
rect 170698 31144 171358 31362
rect 171526 31144 172186 31362
rect 172354 31144 173014 31362
rect 173182 31144 173842 31362
rect 174010 31144 174670 31362
rect 174838 31144 175498 31362
rect 175666 31144 176326 31362
rect 176494 31144 177154 31362
rect 177322 31144 177982 31362
rect 178150 31144 178810 31362
rect 178978 31144 179638 31362
rect 179806 31144 180466 31362
rect 180634 31144 181294 31362
rect 181462 31144 182122 31362
rect 182290 31144 182950 31362
rect 183118 31144 183778 31362
rect 183946 31144 184606 31362
rect 184774 31144 185434 31362
rect 185602 31144 186262 31362
rect 186430 31144 187090 31362
rect 187258 31144 187918 31362
rect 188086 31144 188746 31362
rect 188914 31144 189574 31362
rect 189742 31144 190402 31362
rect 190570 31144 191230 31362
rect 191398 31144 192058 31362
rect 192226 31144 192886 31362
rect 193054 31144 193714 31362
rect 193882 31144 194542 31362
rect 194710 31144 195370 31362
rect 195538 31144 196198 31362
rect 196366 31144 197026 31362
rect 197194 31144 197854 31362
rect 198022 31144 198682 31362
rect 198850 31144 199510 31362
rect 199678 31144 200338 31362
rect 200506 31144 201166 31362
rect 201334 31144 201994 31362
rect 202162 31144 202822 31362
rect 202990 31144 203650 31362
rect 203818 31144 204478 31362
rect 204646 31144 205306 31362
rect 205474 31144 206134 31362
rect 206302 31144 206962 31362
rect 207130 31144 207790 31362
rect 207958 31144 208618 31362
rect 208786 31144 209446 31362
rect 209614 31144 210274 31362
rect 210442 31144 211102 31362
rect 211270 31144 211930 31362
rect 212098 31144 212758 31362
rect 212926 31144 213586 31362
rect 213754 31144 214414 31362
rect 214582 31144 215242 31362
rect 215410 31144 216070 31362
rect 216238 31144 216898 31362
rect 217066 31144 217726 31362
rect 217894 31144 218554 31362
rect 218722 31144 219382 31362
rect 219550 31144 220210 31362
rect 220378 31144 221038 31362
rect 221206 31144 221866 31362
rect 222034 31144 222694 31362
rect 222862 31144 223522 31362
rect 223690 31144 224350 31362
rect 224518 31144 225178 31362
rect 225346 31144 226006 31362
rect 226174 31144 226834 31362
rect 227002 31144 227662 31362
rect 227830 31144 228490 31362
rect 228658 31144 229318 31362
rect 229486 31144 230146 31362
rect 230314 31144 230974 31362
rect 231142 31144 231802 31362
rect 231970 31144 232630 31362
rect 232798 31144 233458 31362
rect 233626 31144 234286 31362
rect 234454 31144 235114 31362
rect 235282 31144 235942 31362
rect 236110 31144 236770 31362
rect 236938 31144 237598 31362
rect 237766 31144 238426 31362
rect 238594 31144 239254 31362
rect 239422 31144 240082 31362
rect 240250 31144 240910 31362
rect 241078 31144 241738 31362
rect 241906 31144 242566 31362
rect 242734 31144 243394 31362
rect 243562 31144 244222 31362
rect 244390 31144 245050 31362
rect 245218 31144 245878 31362
rect 246046 31144 246706 31362
rect 246874 31144 247534 31362
rect 247702 31144 248362 31362
rect 248530 31144 249190 31362
rect 249358 31144 250018 31362
rect 250186 31144 250846 31362
rect 251014 31144 251674 31362
rect 251842 31144 252502 31362
rect 252670 31144 253330 31362
rect 253498 31144 254158 31362
rect 254326 31144 254986 31362
rect 255154 31144 255814 31362
rect 255982 31144 256642 31362
rect 256810 31144 257470 31362
rect 257638 31144 258298 31362
rect 258466 31144 259126 31362
rect 259294 31144 259954 31362
rect 260122 31144 260782 31362
rect 260950 31144 261610 31362
rect 261778 31144 262438 31362
rect 262606 31144 263266 31362
rect 263434 31144 264094 31362
rect 264262 31144 264922 31362
rect 265090 31144 265750 31362
rect 265918 31144 266578 31362
rect 266746 31144 267406 31362
rect 267574 31144 268234 31362
rect 268402 31144 269062 31362
rect 269230 31144 269890 31362
rect 270058 31144 270718 31362
rect 270886 31144 271546 31362
rect 271714 31144 272374 31362
rect 272542 31144 273202 31362
rect 273370 31144 274030 31362
rect 274198 31144 274858 31362
rect 275026 31144 275686 31362
rect 275854 31144 276514 31362
rect 276682 31144 277342 31362
rect 277510 31144 278170 31362
rect 278338 31144 278998 31362
rect 279166 31144 279826 31362
rect 279994 31144 280654 31362
rect 280822 31144 281482 31362
rect 281650 31144 282310 31362
rect 282478 31144 283138 31362
rect 283306 31144 283966 31362
rect 284134 31144 284794 31362
rect 284962 31144 285622 31362
rect 285790 31144 286450 31362
rect 286618 31144 287278 31362
rect 287446 31144 288106 31362
rect 288274 31144 288934 31362
rect 289102 31144 289762 31362
rect 289930 31144 290590 31362
rect 290758 31144 291418 31362
rect 291586 31144 292246 31362
rect 292414 31144 293074 31362
rect 293242 31144 293902 31362
rect 294070 31144 294730 31362
rect 294898 31144 295558 31362
rect 295726 31144 296386 31362
rect 296554 31144 297214 31362
rect 297382 31144 298042 31362
rect 298210 31144 298870 31362
rect 299038 31144 299698 31362
rect 299866 31144 300526 31362
rect 300694 31144 301354 31362
rect 301522 31144 302182 31362
rect 302350 31144 303010 31362
rect 303178 31144 303838 31362
rect 304006 31144 304666 31362
rect 304834 31144 305494 31362
rect 305662 31144 306322 31362
rect 306490 31144 307150 31362
rect 307318 31144 307978 31362
rect 308146 31144 308806 31362
rect 308974 31144 309634 31362
rect 309802 31144 310462 31362
rect 310630 31144 311290 31362
rect 311458 31144 312118 31362
rect 312286 31144 312946 31362
rect 313114 31144 313774 31362
rect 313942 31144 314602 31362
rect 314770 31144 315430 31362
rect 315598 31144 316258 31362
rect 316426 31144 317086 31362
rect 317254 31144 317914 31362
rect 318082 31144 318742 31362
rect 318910 31144 319570 31362
rect 319738 31144 320398 31362
rect 320566 31144 321226 31362
rect 321394 31144 322054 31362
rect 322222 31144 322882 31362
rect 323050 31144 323710 31362
rect 323878 31144 324538 31362
rect 324706 31144 325366 31362
rect 325534 31144 326194 31362
rect 326362 31144 327022 31362
rect 327190 31144 327850 31362
rect 328018 31144 328678 31362
rect 328846 31144 329506 31362
rect 329674 31144 330334 31362
rect 330502 31144 331162 31362
rect 331330 31144 331990 31362
rect 332158 31144 332818 31362
rect 332986 31144 333646 31362
rect 333814 31144 334474 31362
rect 334642 31144 335302 31362
rect 335470 31144 336130 31362
rect 336298 31144 336958 31362
rect 337126 31144 337786 31362
rect 337954 31144 338614 31362
rect 338782 31144 339442 31362
rect 339610 31144 340270 31362
rect 340438 31144 341098 31362
rect 341266 31144 341926 31362
rect 342094 31144 342754 31362
rect 342922 31144 343582 31362
rect 343750 31144 344410 31362
rect 344578 31144 345238 31362
rect 345406 31144 346066 31362
rect 346234 31144 346894 31362
rect 347062 31144 347722 31362
rect 347890 31144 348550 31362
rect 348718 31144 349378 31362
rect 349546 31144 350206 31362
rect 350374 31144 351034 31362
rect 351202 31144 351862 31362
rect 352030 31144 352690 31362
rect 352858 31144 353518 31362
rect 353686 31144 354346 31362
rect 354514 31144 355174 31362
rect 355342 31144 356002 31362
rect 356170 31144 356830 31362
rect 356998 31144 357658 31362
rect 357826 31144 358486 31362
rect 358654 31144 359314 31362
rect 359482 31144 360142 31362
rect 360310 31144 360970 31362
rect 361138 31144 361798 31362
rect 361966 31144 362626 31362
rect 362794 31144 363454 31362
rect 363622 31144 364282 31362
rect 364450 31144 365110 31362
rect 365278 31144 365938 31362
rect 366106 31144 366766 31362
rect 366934 31144 367594 31362
rect 367762 31144 368422 31362
rect 368590 31144 369250 31362
rect 369418 31144 370078 31362
rect 370246 31144 370906 31362
rect 371074 31144 371734 31362
rect 371902 31144 372562 31362
rect 372730 31144 373390 31362
rect 373558 31144 374218 31362
rect 374386 31144 375046 31362
rect 375214 31144 375874 31362
rect 376042 31144 376702 31362
rect 376870 31144 377530 31362
rect 377698 31144 378358 31362
rect 378526 31144 379186 31362
rect 379354 31144 380014 31362
rect 380182 31144 380842 31362
rect 381010 31144 381670 31362
rect 381838 31144 382498 31362
rect 382666 31144 383326 31362
rect 383494 31144 384154 31362
rect 384322 31144 384982 31362
rect 385150 31144 385810 31362
rect 385978 31144 386638 31362
rect 386806 31144 387466 31362
rect 387634 31144 388294 31362
rect 388462 31144 389122 31362
rect 389290 31144 389950 31362
rect 390118 31144 390778 31362
rect 390946 31144 391606 31362
rect 391774 31144 392434 31362
rect 392602 31144 393262 31362
rect 393430 31144 394090 31362
rect 394258 31144 394918 31362
rect 395086 31144 395746 31362
rect 395914 31144 396574 31362
rect 396742 31144 397402 31362
rect 397570 31144 398230 31362
rect 398398 31144 399058 31362
rect 399226 31144 399886 31362
rect 400054 31144 400714 31362
rect 400882 31144 401542 31362
rect 401710 31144 402370 31362
rect 402538 31144 403198 31362
rect 403366 31144 404026 31362
rect 404194 31144 404854 31362
rect 405022 31144 405682 31362
rect 405850 31144 406510 31362
rect 406678 31144 407338 31362
rect 407506 31144 408166 31362
rect 408334 31144 408994 31362
rect 409162 31144 409822 31362
rect 409990 31144 410650 31362
rect 410818 31144 411478 31362
rect 411646 31144 412306 31362
rect 412474 31144 413134 31362
rect 413302 31144 413962 31362
rect 414130 31144 414790 31362
rect 414958 31144 422444 31362
rect 5036 856 422444 31144
rect 5036 2 16154 856
rect 16322 2 16798 856
rect 16966 2 17442 856
rect 17610 2 18086 856
rect 18254 2 18730 856
rect 18898 2 19374 856
rect 19542 2 20018 856
rect 20186 2 20662 856
rect 20830 2 21306 856
rect 21474 2 21950 856
rect 22118 2 22594 856
rect 22762 2 23238 856
rect 23406 2 23882 856
rect 24050 2 24526 856
rect 24694 2 25170 856
rect 25338 2 25814 856
rect 25982 2 26458 856
rect 26626 2 27102 856
rect 27270 2 27746 856
rect 27914 2 28390 856
rect 28558 2 29034 856
rect 29202 2 29678 856
rect 29846 2 30322 856
rect 30490 2 30966 856
rect 31134 2 31610 856
rect 31778 2 32254 856
rect 32422 2 32898 856
rect 33066 2 33542 856
rect 33710 2 34186 856
rect 34354 2 34830 856
rect 34998 2 35474 856
rect 35642 2 36118 856
rect 36286 2 36762 856
rect 36930 2 37406 856
rect 37574 2 38050 856
rect 38218 2 38694 856
rect 38862 2 39338 856
rect 39506 2 39982 856
rect 40150 2 40626 856
rect 40794 2 41270 856
rect 41438 2 41914 856
rect 42082 2 42558 856
rect 42726 2 43202 856
rect 43370 2 43846 856
rect 44014 2 44490 856
rect 44658 2 45134 856
rect 45302 2 45778 856
rect 45946 2 46422 856
rect 46590 2 47066 856
rect 47234 2 47710 856
rect 47878 2 48354 856
rect 48522 2 48998 856
rect 49166 2 49642 856
rect 49810 2 50286 856
rect 50454 2 50930 856
rect 51098 2 51574 856
rect 51742 2 52218 856
rect 52386 2 52862 856
rect 53030 2 53506 856
rect 53674 2 54150 856
rect 54318 2 54794 856
rect 54962 2 55438 856
rect 55606 2 56082 856
rect 56250 2 56726 856
rect 56894 2 57370 856
rect 57538 2 58014 856
rect 58182 2 58658 856
rect 58826 2 59302 856
rect 59470 2 59946 856
rect 60114 2 60590 856
rect 60758 2 61234 856
rect 61402 2 61878 856
rect 62046 2 62522 856
rect 62690 2 63166 856
rect 63334 2 63810 856
rect 63978 2 64454 856
rect 64622 2 65098 856
rect 65266 2 65742 856
rect 65910 2 66386 856
rect 66554 2 67030 856
rect 67198 2 67674 856
rect 67842 2 68318 856
rect 68486 2 68962 856
rect 69130 2 69606 856
rect 69774 2 70250 856
rect 70418 2 70894 856
rect 71062 2 71538 856
rect 71706 2 72182 856
rect 72350 2 72826 856
rect 72994 2 73470 856
rect 73638 2 74114 856
rect 74282 2 74758 856
rect 74926 2 75402 856
rect 75570 2 76046 856
rect 76214 2 76690 856
rect 76858 2 77334 856
rect 77502 2 77978 856
rect 78146 2 78622 856
rect 78790 2 79266 856
rect 79434 2 79910 856
rect 80078 2 80554 856
rect 80722 2 81198 856
rect 81366 2 81842 856
rect 82010 2 82486 856
rect 82654 2 83130 856
rect 83298 2 83774 856
rect 83942 2 84418 856
rect 84586 2 85062 856
rect 85230 2 85706 856
rect 85874 2 86350 856
rect 86518 2 86994 856
rect 87162 2 87638 856
rect 87806 2 88282 856
rect 88450 2 88926 856
rect 89094 2 89570 856
rect 89738 2 90214 856
rect 90382 2 90858 856
rect 91026 2 91502 856
rect 91670 2 92146 856
rect 92314 2 92790 856
rect 92958 2 93434 856
rect 93602 2 94078 856
rect 94246 2 94722 856
rect 94890 2 95366 856
rect 95534 2 96010 856
rect 96178 2 96654 856
rect 96822 2 97298 856
rect 97466 2 97942 856
rect 98110 2 98586 856
rect 98754 2 99230 856
rect 99398 2 99874 856
rect 100042 2 100518 856
rect 100686 2 101162 856
rect 101330 2 101806 856
rect 101974 2 102450 856
rect 102618 2 103094 856
rect 103262 2 103738 856
rect 103906 2 104382 856
rect 104550 2 105026 856
rect 105194 2 105670 856
rect 105838 2 106314 856
rect 106482 2 106958 856
rect 107126 2 107602 856
rect 107770 2 108246 856
rect 108414 2 108890 856
rect 109058 2 109534 856
rect 109702 2 110178 856
rect 110346 2 110822 856
rect 110990 2 111466 856
rect 111634 2 112110 856
rect 112278 2 112754 856
rect 112922 2 113398 856
rect 113566 2 114042 856
rect 114210 2 114686 856
rect 114854 2 115330 856
rect 115498 2 115974 856
rect 116142 2 116618 856
rect 116786 2 117262 856
rect 117430 2 117906 856
rect 118074 2 118550 856
rect 118718 2 119194 856
rect 119362 2 119838 856
rect 120006 2 120482 856
rect 120650 2 121126 856
rect 121294 2 121770 856
rect 121938 2 122414 856
rect 122582 2 123058 856
rect 123226 2 123702 856
rect 123870 2 124346 856
rect 124514 2 124990 856
rect 125158 2 125634 856
rect 125802 2 126278 856
rect 126446 2 126922 856
rect 127090 2 127566 856
rect 127734 2 128210 856
rect 128378 2 128854 856
rect 129022 2 129498 856
rect 129666 2 130142 856
rect 130310 2 130786 856
rect 130954 2 131430 856
rect 131598 2 132074 856
rect 132242 2 132718 856
rect 132886 2 133362 856
rect 133530 2 134006 856
rect 134174 2 134650 856
rect 134818 2 135294 856
rect 135462 2 135938 856
rect 136106 2 136582 856
rect 136750 2 137226 856
rect 137394 2 137870 856
rect 138038 2 138514 856
rect 138682 2 139158 856
rect 139326 2 139802 856
rect 139970 2 140446 856
rect 140614 2 141090 856
rect 141258 2 141734 856
rect 141902 2 142378 856
rect 142546 2 143022 856
rect 143190 2 143666 856
rect 143834 2 144310 856
rect 144478 2 144954 856
rect 145122 2 145598 856
rect 145766 2 146242 856
rect 146410 2 146886 856
rect 147054 2 147530 856
rect 147698 2 148174 856
rect 148342 2 148818 856
rect 148986 2 149462 856
rect 149630 2 150106 856
rect 150274 2 150750 856
rect 150918 2 151394 856
rect 151562 2 152038 856
rect 152206 2 152682 856
rect 152850 2 153326 856
rect 153494 2 153970 856
rect 154138 2 154614 856
rect 154782 2 155258 856
rect 155426 2 155902 856
rect 156070 2 156546 856
rect 156714 2 157190 856
rect 157358 2 157834 856
rect 158002 2 158478 856
rect 158646 2 159122 856
rect 159290 2 159766 856
rect 159934 2 160410 856
rect 160578 2 161054 856
rect 161222 2 161698 856
rect 161866 2 162342 856
rect 162510 2 162986 856
rect 163154 2 163630 856
rect 163798 2 164274 856
rect 164442 2 164918 856
rect 165086 2 165562 856
rect 165730 2 166206 856
rect 166374 2 166850 856
rect 167018 2 167494 856
rect 167662 2 168138 856
rect 168306 2 168782 856
rect 168950 2 169426 856
rect 169594 2 170070 856
rect 170238 2 170714 856
rect 170882 2 171358 856
rect 171526 2 172002 856
rect 172170 2 172646 856
rect 172814 2 173290 856
rect 173458 2 173934 856
rect 174102 2 174578 856
rect 174746 2 175222 856
rect 175390 2 175866 856
rect 176034 2 176510 856
rect 176678 2 177154 856
rect 177322 2 177798 856
rect 177966 2 178442 856
rect 178610 2 179086 856
rect 179254 2 179730 856
rect 179898 2 180374 856
rect 180542 2 181018 856
rect 181186 2 181662 856
rect 181830 2 182306 856
rect 182474 2 182950 856
rect 183118 2 183594 856
rect 183762 2 184238 856
rect 184406 2 184882 856
rect 185050 2 185526 856
rect 185694 2 186170 856
rect 186338 2 186814 856
rect 186982 2 187458 856
rect 187626 2 188102 856
rect 188270 2 188746 856
rect 188914 2 189390 856
rect 189558 2 190034 856
rect 190202 2 190678 856
rect 190846 2 191322 856
rect 191490 2 191966 856
rect 192134 2 192610 856
rect 192778 2 193254 856
rect 193422 2 193898 856
rect 194066 2 194542 856
rect 194710 2 195186 856
rect 195354 2 195830 856
rect 195998 2 196474 856
rect 196642 2 197118 856
rect 197286 2 197762 856
rect 197930 2 198406 856
rect 198574 2 199050 856
rect 199218 2 199694 856
rect 199862 2 200338 856
rect 200506 2 200982 856
rect 201150 2 201626 856
rect 201794 2 202270 856
rect 202438 2 202914 856
rect 203082 2 203558 856
rect 203726 2 204202 856
rect 204370 2 204846 856
rect 205014 2 205490 856
rect 205658 2 206134 856
rect 206302 2 206778 856
rect 206946 2 207422 856
rect 207590 2 208066 856
rect 208234 2 208710 856
rect 208878 2 209354 856
rect 209522 2 209998 856
rect 210166 2 210642 856
rect 210810 2 211286 856
rect 211454 2 211930 856
rect 212098 2 212574 856
rect 212742 2 213218 856
rect 213386 2 213862 856
rect 214030 2 214506 856
rect 214674 2 215150 856
rect 215318 2 215794 856
rect 215962 2 216438 856
rect 216606 2 217082 856
rect 217250 2 217726 856
rect 217894 2 218370 856
rect 218538 2 219014 856
rect 219182 2 219658 856
rect 219826 2 220302 856
rect 220470 2 220946 856
rect 221114 2 221590 856
rect 221758 2 222234 856
rect 222402 2 222878 856
rect 223046 2 223522 856
rect 223690 2 224166 856
rect 224334 2 224810 856
rect 224978 2 225454 856
rect 225622 2 226098 856
rect 226266 2 226742 856
rect 226910 2 227386 856
rect 227554 2 228030 856
rect 228198 2 228674 856
rect 228842 2 229318 856
rect 229486 2 229962 856
rect 230130 2 230606 856
rect 230774 2 231250 856
rect 231418 2 231894 856
rect 232062 2 232538 856
rect 232706 2 233182 856
rect 233350 2 233826 856
rect 233994 2 234470 856
rect 234638 2 235114 856
rect 235282 2 235758 856
rect 235926 2 236402 856
rect 236570 2 237046 856
rect 237214 2 237690 856
rect 237858 2 238334 856
rect 238502 2 238978 856
rect 239146 2 239622 856
rect 239790 2 240266 856
rect 240434 2 240910 856
rect 241078 2 241554 856
rect 241722 2 242198 856
rect 242366 2 242842 856
rect 243010 2 243486 856
rect 243654 2 244130 856
rect 244298 2 244774 856
rect 244942 2 245418 856
rect 245586 2 246062 856
rect 246230 2 246706 856
rect 246874 2 247350 856
rect 247518 2 247994 856
rect 248162 2 248638 856
rect 248806 2 249282 856
rect 249450 2 249926 856
rect 250094 2 250570 856
rect 250738 2 251214 856
rect 251382 2 251858 856
rect 252026 2 252502 856
rect 252670 2 253146 856
rect 253314 2 253790 856
rect 253958 2 254434 856
rect 254602 2 255078 856
rect 255246 2 255722 856
rect 255890 2 256366 856
rect 256534 2 257010 856
rect 257178 2 257654 856
rect 257822 2 258298 856
rect 258466 2 258942 856
rect 259110 2 259586 856
rect 259754 2 260230 856
rect 260398 2 260874 856
rect 261042 2 261518 856
rect 261686 2 262162 856
rect 262330 2 262806 856
rect 262974 2 263450 856
rect 263618 2 264094 856
rect 264262 2 264738 856
rect 264906 2 265382 856
rect 265550 2 266026 856
rect 266194 2 266670 856
rect 266838 2 267314 856
rect 267482 2 267958 856
rect 268126 2 268602 856
rect 268770 2 269246 856
rect 269414 2 269890 856
rect 270058 2 270534 856
rect 270702 2 271178 856
rect 271346 2 271822 856
rect 271990 2 272466 856
rect 272634 2 273110 856
rect 273278 2 273754 856
rect 273922 2 274398 856
rect 274566 2 275042 856
rect 275210 2 275686 856
rect 275854 2 276330 856
rect 276498 2 276974 856
rect 277142 2 277618 856
rect 277786 2 278262 856
rect 278430 2 278906 856
rect 279074 2 279550 856
rect 279718 2 280194 856
rect 280362 2 280838 856
rect 281006 2 281482 856
rect 281650 2 282126 856
rect 282294 2 282770 856
rect 282938 2 283414 856
rect 283582 2 284058 856
rect 284226 2 284702 856
rect 284870 2 285346 856
rect 285514 2 285990 856
rect 286158 2 286634 856
rect 286802 2 287278 856
rect 287446 2 287922 856
rect 288090 2 288566 856
rect 288734 2 289210 856
rect 289378 2 289854 856
rect 290022 2 290498 856
rect 290666 2 291142 856
rect 291310 2 291786 856
rect 291954 2 292430 856
rect 292598 2 293074 856
rect 293242 2 293718 856
rect 293886 2 294362 856
rect 294530 2 295006 856
rect 295174 2 295650 856
rect 295818 2 296294 856
rect 296462 2 296938 856
rect 297106 2 297582 856
rect 297750 2 298226 856
rect 298394 2 298870 856
rect 299038 2 299514 856
rect 299682 2 300158 856
rect 300326 2 300802 856
rect 300970 2 301446 856
rect 301614 2 302090 856
rect 302258 2 302734 856
rect 302902 2 303378 856
rect 303546 2 304022 856
rect 304190 2 304666 856
rect 304834 2 305310 856
rect 305478 2 305954 856
rect 306122 2 306598 856
rect 306766 2 307242 856
rect 307410 2 307886 856
rect 308054 2 308530 856
rect 308698 2 309174 856
rect 309342 2 309818 856
rect 309986 2 310462 856
rect 310630 2 311106 856
rect 311274 2 311750 856
rect 311918 2 312394 856
rect 312562 2 313038 856
rect 313206 2 313682 856
rect 313850 2 314326 856
rect 314494 2 314970 856
rect 315138 2 315614 856
rect 315782 2 316258 856
rect 316426 2 316902 856
rect 317070 2 317546 856
rect 317714 2 318190 856
rect 318358 2 318834 856
rect 319002 2 319478 856
rect 319646 2 320122 856
rect 320290 2 320766 856
rect 320934 2 321410 856
rect 321578 2 322054 856
rect 322222 2 322698 856
rect 322866 2 323342 856
rect 323510 2 323986 856
rect 324154 2 324630 856
rect 324798 2 325274 856
rect 325442 2 325918 856
rect 326086 2 326562 856
rect 326730 2 327206 856
rect 327374 2 327850 856
rect 328018 2 328494 856
rect 328662 2 329138 856
rect 329306 2 329782 856
rect 329950 2 330426 856
rect 330594 2 331070 856
rect 331238 2 331714 856
rect 331882 2 332358 856
rect 332526 2 333002 856
rect 333170 2 333646 856
rect 333814 2 334290 856
rect 334458 2 334934 856
rect 335102 2 335578 856
rect 335746 2 336222 856
rect 336390 2 336866 856
rect 337034 2 337510 856
rect 337678 2 338154 856
rect 338322 2 338798 856
rect 338966 2 339442 856
rect 339610 2 340086 856
rect 340254 2 340730 856
rect 340898 2 341374 856
rect 341542 2 342018 856
rect 342186 2 342662 856
rect 342830 2 343306 856
rect 343474 2 343950 856
rect 344118 2 344594 856
rect 344762 2 345238 856
rect 345406 2 345882 856
rect 346050 2 346526 856
rect 346694 2 347170 856
rect 347338 2 347814 856
rect 347982 2 348458 856
rect 348626 2 349102 856
rect 349270 2 349746 856
rect 349914 2 350390 856
rect 350558 2 351034 856
rect 351202 2 351678 856
rect 351846 2 352322 856
rect 352490 2 352966 856
rect 353134 2 353610 856
rect 353778 2 354254 856
rect 354422 2 354898 856
rect 355066 2 355542 856
rect 355710 2 356186 856
rect 356354 2 356830 856
rect 356998 2 357474 856
rect 357642 2 358118 856
rect 358286 2 358762 856
rect 358930 2 359406 856
rect 359574 2 360050 856
rect 360218 2 360694 856
rect 360862 2 361338 856
rect 361506 2 361982 856
rect 362150 2 362626 856
rect 362794 2 363270 856
rect 363438 2 363914 856
rect 364082 2 364558 856
rect 364726 2 365202 856
rect 365370 2 365846 856
rect 366014 2 366490 856
rect 366658 2 367134 856
rect 367302 2 367778 856
rect 367946 2 368422 856
rect 368590 2 369066 856
rect 369234 2 369710 856
rect 369878 2 370354 856
rect 370522 2 370998 856
rect 371166 2 371642 856
rect 371810 2 372286 856
rect 372454 2 372930 856
rect 373098 2 373574 856
rect 373742 2 374218 856
rect 374386 2 374862 856
rect 375030 2 375506 856
rect 375674 2 376150 856
rect 376318 2 376794 856
rect 376962 2 377438 856
rect 377606 2 378082 856
rect 378250 2 378726 856
rect 378894 2 379370 856
rect 379538 2 380014 856
rect 380182 2 380658 856
rect 380826 2 381302 856
rect 381470 2 381946 856
rect 382114 2 382590 856
rect 382758 2 383234 856
rect 383402 2 383878 856
rect 384046 2 384522 856
rect 384690 2 385166 856
rect 385334 2 385810 856
rect 385978 2 386454 856
rect 386622 2 387098 856
rect 387266 2 387742 856
rect 387910 2 388386 856
rect 388554 2 389030 856
rect 389198 2 389674 856
rect 389842 2 390318 856
rect 390486 2 390962 856
rect 391130 2 391606 856
rect 391774 2 392250 856
rect 392418 2 392894 856
rect 393062 2 393538 856
rect 393706 2 394182 856
rect 394350 2 394826 856
rect 394994 2 395470 856
rect 395638 2 396114 856
rect 396282 2 396758 856
rect 396926 2 397402 856
rect 397570 2 398046 856
rect 398214 2 398690 856
rect 398858 2 399334 856
rect 399502 2 399978 856
rect 400146 2 400622 856
rect 400790 2 401266 856
rect 401434 2 401910 856
rect 402078 2 402554 856
rect 402722 2 403198 856
rect 403366 2 403842 856
rect 404010 2 404486 856
rect 404654 2 405130 856
rect 405298 2 405774 856
rect 405942 2 406418 856
rect 406586 2 407062 856
rect 407230 2 407706 856
rect 407874 2 422444 856
<< metal3 >>
rect 423200 29928 424400 30048
rect 423200 28704 424400 28824
rect 423200 27480 424400 27600
rect 423200 26256 424400 26376
rect 423200 25032 424400 25152
rect 423200 23808 424400 23928
rect 423200 22584 424400 22704
rect 423200 21360 424400 21480
rect 423200 20136 424400 20256
rect 423200 18912 424400 19032
rect 423200 17688 424400 17808
rect 423200 16464 424400 16584
rect 423200 15240 424400 15360
rect 423200 14016 424400 14136
rect 423200 12792 424400 12912
rect 423200 11568 424400 11688
rect 423200 10344 424400 10464
rect 423200 9120 424400 9240
rect 423200 7896 424400 8016
rect 423200 6672 424400 6792
rect 423200 5448 424400 5568
rect 423200 4224 424400 4344
rect 423200 3000 424400 3120
rect 423200 1776 424400 1896
<< obsm3 >>
rect 5026 30128 423200 30497
rect 5026 29848 423120 30128
rect 5026 28904 423200 29848
rect 5026 28624 423120 28904
rect 5026 27680 423200 28624
rect 5026 27400 423120 27680
rect 5026 26456 423200 27400
rect 5026 26176 423120 26456
rect 5026 25232 423200 26176
rect 5026 24952 423120 25232
rect 5026 24008 423200 24952
rect 5026 23728 423120 24008
rect 5026 22784 423200 23728
rect 5026 22504 423120 22784
rect 5026 21560 423200 22504
rect 5026 21280 423120 21560
rect 5026 20336 423200 21280
rect 5026 20056 423120 20336
rect 5026 19112 423200 20056
rect 5026 18832 423120 19112
rect 5026 17888 423200 18832
rect 5026 17608 423120 17888
rect 5026 16664 423200 17608
rect 5026 16384 423120 16664
rect 5026 15440 423200 16384
rect 5026 15160 423120 15440
rect 5026 14216 423200 15160
rect 5026 13936 423120 14216
rect 5026 12992 423200 13936
rect 5026 12712 423120 12992
rect 5026 11768 423200 12712
rect 5026 11488 423120 11768
rect 5026 10544 423200 11488
rect 5026 10264 423120 10544
rect 5026 9320 423200 10264
rect 5026 9040 423120 9320
rect 5026 8096 423200 9040
rect 5026 7816 423120 8096
rect 5026 6872 423200 7816
rect 5026 6592 423120 6872
rect 5026 5648 423200 6592
rect 5026 5368 423120 5648
rect 5026 4424 423200 5368
rect 5026 4144 423120 4424
rect 5026 3200 423200 4144
rect 5026 2920 423120 3200
rect 5026 1976 423200 2920
rect 5026 1696 423120 1976
rect 5026 35 423200 1696
<< metal4 >>
rect 5014 1040 5194 30512
rect 12394 1040 12574 30512
rect 20064 1040 20244 30512
rect 27444 1040 27624 30512
rect 35114 1040 35294 30512
rect 42494 1040 42674 30512
rect 50164 1040 50344 30512
rect 57544 1040 57724 30512
rect 65214 1040 65394 30512
rect 66854 1040 67034 30512
rect 71034 1040 71214 30512
rect 72594 1040 72774 30512
rect 76854 1040 77034 30512
rect 80264 1040 80444 30512
rect 81034 1040 81214 30512
rect 87644 1040 87824 30512
rect 95314 1040 95494 30512
rect 102694 1040 102874 30512
rect 110364 1040 110544 30512
rect 117744 1040 117924 30512
rect 125414 1040 125594 30512
rect 132794 1040 132974 30512
rect 140464 1040 140644 30512
rect 141284 1040 141464 30512
rect 147844 1040 148024 30512
rect 148664 1040 148844 30512
rect 155514 1040 155694 30512
rect 156334 1040 156514 30512
rect 162894 1040 163074 30512
rect 163714 1040 163894 30512
rect 170564 1040 170744 30512
rect 171384 1040 171564 30512
rect 177944 1040 178124 30512
rect 178764 1040 178944 30512
rect 185614 1040 185794 30512
rect 186434 1040 186614 30512
rect 192994 1040 193174 30512
rect 193814 1040 193994 30512
rect 200664 1040 200844 30512
rect 208044 1040 208224 30512
rect 215714 1040 215894 30512
rect 223094 1040 223274 30512
rect 230764 1040 230944 30512
rect 238144 1040 238324 30512
rect 245814 1040 245994 30512
rect 253194 1040 253374 30512
rect 255814 1040 255994 30512
rect 256614 1040 256794 30512
rect 260864 1040 261044 30512
rect 263194 1040 263374 30512
rect 263994 1040 264174 30512
rect 268244 1040 268424 30512
rect 270864 1040 271044 30512
rect 271664 1040 271844 30512
rect 275914 1040 276094 30512
rect 278244 1040 278424 30512
rect 279044 1040 279224 30512
rect 283294 1040 283474 30512
rect 290964 1040 291144 30512
rect 298344 1040 298524 30512
rect 306014 1040 306194 30512
rect 313394 1040 313574 30512
rect 321064 1040 321244 30512
rect 328444 1040 328624 30512
rect 336114 1040 336294 30512
rect 343494 1040 343674 30512
rect 351164 1040 351344 30512
rect 358544 1040 358724 30512
rect 366214 1040 366394 30512
rect 373594 1040 373774 30512
rect 381264 1040 381444 30512
rect 388644 1040 388824 30512
rect 396314 1040 396494 30512
rect 403694 1040 403874 30512
rect 411364 1040 411544 30512
rect 418744 1040 418924 30512
<< obsm4 >>
rect 12194 960 12314 30512
rect 12654 960 19984 30512
rect 20324 960 27364 30512
rect 27704 960 35034 30512
rect 35374 960 42414 30512
rect 42754 960 50084 30512
rect 50424 960 57464 30512
rect 57804 960 65134 30512
rect 65474 960 66774 30512
rect 67114 960 70954 30512
rect 71294 960 72514 30512
rect 72854 960 76774 30512
rect 77114 960 80184 30512
rect 80524 960 80954 30512
rect 81294 960 87564 30512
rect 87904 960 95234 30512
rect 95574 960 102614 30512
rect 102954 960 110284 30512
rect 110624 960 117664 30512
rect 118004 960 125334 30512
rect 125674 960 132714 30512
rect 133054 960 140384 30512
rect 140724 960 141204 30512
rect 141544 960 147764 30512
rect 148104 960 148584 30512
rect 148924 960 155434 30512
rect 155774 960 156254 30512
rect 156594 960 162814 30512
rect 163154 960 163634 30512
rect 163974 960 170484 30512
rect 170824 960 171304 30512
rect 171644 960 177864 30512
rect 178204 960 178684 30512
rect 179024 960 185534 30512
rect 185874 960 186354 30512
rect 186694 960 192914 30512
rect 193254 960 193734 30512
rect 194074 960 200584 30512
rect 200924 960 207964 30512
rect 208304 960 215634 30512
rect 215974 960 223014 30512
rect 223354 960 230684 30512
rect 231024 960 238064 30512
rect 238404 960 245734 30512
rect 246074 960 253114 30512
rect 253454 960 255734 30512
rect 256074 960 256534 30512
rect 256874 960 260784 30512
rect 261124 960 263114 30512
rect 263454 960 263914 30512
rect 264254 960 268164 30512
rect 268504 960 270784 30512
rect 271124 960 271584 30512
rect 271924 960 275834 30512
rect 276174 960 278164 30512
rect 278504 960 278964 30512
rect 279304 960 283214 30512
rect 283554 960 290884 30512
rect 291224 960 298264 30512
rect 298604 960 305934 30512
rect 306274 960 313314 30512
rect 313654 960 320984 30512
rect 321324 960 328364 30512
rect 328704 960 336034 30512
rect 336374 960 343414 30512
rect 343754 960 351084 30512
rect 351424 960 358464 30512
rect 358804 960 366134 30512
rect 366474 960 373514 30512
rect 373854 960 373974 30512
rect 12194 35 373974 960
<< labels >>
rlabel metal3 s 423200 15240 424400 15360 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s 423200 16464 424400 16584 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s 423200 17688 424400 17808 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 96894 31200 96950 32400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 345294 31200 345350 32400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 347778 31200 347834 32400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 350262 31200 350318 32400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 352746 31200 352802 32400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 355230 31200 355286 32400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 357714 31200 357770 32400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 360198 31200 360254 32400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 362682 31200 362738 32400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 365166 31200 365222 32400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 367650 31200 367706 32400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 121734 31200 121790 32400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 370134 31200 370190 32400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 372618 31200 372674 32400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 375102 31200 375158 32400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 377586 31200 377642 32400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 380070 31200 380126 32400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 382554 31200 382610 32400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 385038 31200 385094 32400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 387522 31200 387578 32400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 390006 31200 390062 32400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 392490 31200 392546 32400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 124218 31200 124274 32400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 394974 31200 395030 32400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 397458 31200 397514 32400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 399942 31200 399998 32400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 402426 31200 402482 32400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 404910 31200 404966 32400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 407394 31200 407450 32400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 409878 31200 409934 32400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 412362 31200 412418 32400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 126702 31200 126758 32400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 129186 31200 129242 32400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 131670 31200 131726 32400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 134154 31200 134210 32400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 136638 31200 136694 32400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 139122 31200 139178 32400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 141606 31200 141662 32400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 144090 31200 144146 32400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 99378 31200 99434 32400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 146574 31200 146630 32400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 149058 31200 149114 32400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 151542 31200 151598 32400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 154026 31200 154082 32400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 156510 31200 156566 32400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 158994 31200 159050 32400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 161478 31200 161534 32400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 163962 31200 164018 32400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 166446 31200 166502 32400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 168930 31200 168986 32400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 101862 31200 101918 32400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 171414 31200 171470 32400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 173898 31200 173954 32400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 176382 31200 176438 32400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 178866 31200 178922 32400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 181350 31200 181406 32400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 183834 31200 183890 32400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 186318 31200 186374 32400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 188802 31200 188858 32400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 191286 31200 191342 32400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 193770 31200 193826 32400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 104346 31200 104402 32400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 196254 31200 196310 32400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 198738 31200 198794 32400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 201222 31200 201278 32400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 203706 31200 203762 32400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 206190 31200 206246 32400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 208674 31200 208730 32400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 211158 31200 211214 32400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 213642 31200 213698 32400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 216126 31200 216182 32400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 218610 31200 218666 32400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 106830 31200 106886 32400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 221094 31200 221150 32400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 223578 31200 223634 32400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 226062 31200 226118 32400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 228546 31200 228602 32400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 231030 31200 231086 32400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 233514 31200 233570 32400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 235998 31200 236054 32400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 238482 31200 238538 32400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 240966 31200 241022 32400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 243450 31200 243506 32400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 109314 31200 109370 32400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 245934 31200 245990 32400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 248418 31200 248474 32400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 250902 31200 250958 32400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 253386 31200 253442 32400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 255870 31200 255926 32400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 258354 31200 258410 32400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 260838 31200 260894 32400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 263322 31200 263378 32400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 265806 31200 265862 32400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 268290 31200 268346 32400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 111798 31200 111854 32400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 270774 31200 270830 32400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 273258 31200 273314 32400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 275742 31200 275798 32400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 278226 31200 278282 32400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 280710 31200 280766 32400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 283194 31200 283250 32400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 285678 31200 285734 32400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 288162 31200 288218 32400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 290646 31200 290702 32400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 293130 31200 293186 32400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 114282 31200 114338 32400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 295614 31200 295670 32400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 298098 31200 298154 32400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 300582 31200 300638 32400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 303066 31200 303122 32400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 305550 31200 305606 32400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 308034 31200 308090 32400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 310518 31200 310574 32400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 313002 31200 313058 32400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 315486 31200 315542 32400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 317970 31200 318026 32400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 116766 31200 116822 32400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 320454 31200 320510 32400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 322938 31200 322994 32400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 325422 31200 325478 32400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 327906 31200 327962 32400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 330390 31200 330446 32400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 332874 31200 332930 32400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 335358 31200 335414 32400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 337842 31200 337898 32400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 340326 31200 340382 32400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 342810 31200 342866 32400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 119250 31200 119306 32400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 16210 -400 16266 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 273810 -400 273866 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 276386 -400 276442 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 278962 -400 279018 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 281538 -400 281594 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 284114 -400 284170 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 286690 -400 286746 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 289266 -400 289322 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 291842 -400 291898 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 294418 -400 294474 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 296994 -400 297050 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 41970 -400 42026 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 299570 -400 299626 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 302146 -400 302202 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 304722 -400 304778 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 307298 -400 307354 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 309874 -400 309930 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 312450 -400 312506 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 315026 -400 315082 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 317602 -400 317658 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 320178 -400 320234 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 322754 -400 322810 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 44546 -400 44602 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 325330 -400 325386 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 327906 -400 327962 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 330482 -400 330538 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 333058 -400 333114 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 335634 -400 335690 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 338210 -400 338266 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 340786 -400 340842 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 343362 -400 343418 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 47122 -400 47178 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 49698 -400 49754 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 52274 -400 52330 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 54850 -400 54906 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 57426 -400 57482 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 60002 -400 60058 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 62578 -400 62634 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 65154 -400 65210 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 18786 -400 18842 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 67730 -400 67786 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 70306 -400 70362 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 72882 -400 72938 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 75458 -400 75514 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 78034 -400 78090 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 80610 -400 80666 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 83186 -400 83242 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 85762 -400 85818 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 88338 -400 88394 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 90914 -400 90970 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 21362 -400 21418 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 93490 -400 93546 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 96066 -400 96122 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 98642 -400 98698 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 101218 -400 101274 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 103794 -400 103850 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 106370 -400 106426 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 108946 -400 109002 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 111522 -400 111578 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 114098 -400 114154 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 116674 -400 116730 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 23938 -400 23994 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 119250 -400 119306 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 121826 -400 121882 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 124402 -400 124458 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 126978 -400 127034 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 129554 -400 129610 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 132130 -400 132186 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 134706 -400 134762 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 137282 -400 137338 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 139858 -400 139914 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 142434 -400 142490 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 26514 -400 26570 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 145010 -400 145066 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 147586 -400 147642 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 150162 -400 150218 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 152738 -400 152794 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 155314 -400 155370 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 157890 -400 157946 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 160466 -400 160522 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 163042 -400 163098 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 165618 -400 165674 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 168194 -400 168250 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 29090 -400 29146 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 170770 -400 170826 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 173346 -400 173402 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 175922 -400 175978 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 178498 -400 178554 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 181074 -400 181130 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 183650 -400 183706 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 186226 -400 186282 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 188802 -400 188858 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 191378 -400 191434 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 193954 -400 194010 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 31666 -400 31722 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 196530 -400 196586 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 199106 -400 199162 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 201682 -400 201738 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 204258 -400 204314 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 206834 -400 206890 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 209410 -400 209466 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 211986 -400 212042 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 214562 -400 214618 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 217138 -400 217194 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 219714 -400 219770 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 34242 -400 34298 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 222290 -400 222346 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 224866 -400 224922 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 227442 -400 227498 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 230018 -400 230074 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 232594 -400 232650 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 235170 -400 235226 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 237746 -400 237802 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 240322 -400 240378 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 242898 -400 242954 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 245474 -400 245530 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 36818 -400 36874 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 248050 -400 248106 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 250626 -400 250682 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 253202 -400 253258 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 255778 -400 255834 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 258354 -400 258410 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 260930 -400 260986 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 263506 -400 263562 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 266082 -400 266138 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 268658 -400 268714 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 271234 -400 271290 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 39394 -400 39450 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 97722 31200 97778 32400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 346122 31200 346178 32400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 348606 31200 348662 32400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 351090 31200 351146 32400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 353574 31200 353630 32400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 356058 31200 356114 32400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 358542 31200 358598 32400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 361026 31200 361082 32400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 363510 31200 363566 32400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 365994 31200 366050 32400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 368478 31200 368534 32400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 122562 31200 122618 32400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 370962 31200 371018 32400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 373446 31200 373502 32400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 375930 31200 375986 32400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 378414 31200 378470 32400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 380898 31200 380954 32400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 383382 31200 383438 32400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 385866 31200 385922 32400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 388350 31200 388406 32400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 390834 31200 390890 32400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 393318 31200 393374 32400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 125046 31200 125102 32400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 395802 31200 395858 32400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 398286 31200 398342 32400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 400770 31200 400826 32400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 403254 31200 403310 32400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 405738 31200 405794 32400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 408222 31200 408278 32400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 410706 31200 410762 32400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 413190 31200 413246 32400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 127530 31200 127586 32400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 130014 31200 130070 32400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 132498 31200 132554 32400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 134982 31200 135038 32400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 137466 31200 137522 32400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 139950 31200 140006 32400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 142434 31200 142490 32400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 144918 31200 144974 32400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 100206 31200 100262 32400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 147402 31200 147458 32400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 149886 31200 149942 32400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 152370 31200 152426 32400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 154854 31200 154910 32400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 157338 31200 157394 32400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 159822 31200 159878 32400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 162306 31200 162362 32400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 164790 31200 164846 32400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 167274 31200 167330 32400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 169758 31200 169814 32400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 102690 31200 102746 32400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 172242 31200 172298 32400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 174726 31200 174782 32400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 177210 31200 177266 32400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 179694 31200 179750 32400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 182178 31200 182234 32400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 184662 31200 184718 32400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 187146 31200 187202 32400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 189630 31200 189686 32400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 192114 31200 192170 32400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 194598 31200 194654 32400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 105174 31200 105230 32400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 197082 31200 197138 32400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 199566 31200 199622 32400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 202050 31200 202106 32400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 204534 31200 204590 32400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 207018 31200 207074 32400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 209502 31200 209558 32400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 211986 31200 212042 32400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 214470 31200 214526 32400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 216954 31200 217010 32400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 219438 31200 219494 32400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 107658 31200 107714 32400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 221922 31200 221978 32400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 224406 31200 224462 32400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 226890 31200 226946 32400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 229374 31200 229430 32400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 231858 31200 231914 32400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 234342 31200 234398 32400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 236826 31200 236882 32400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 239310 31200 239366 32400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 241794 31200 241850 32400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 244278 31200 244334 32400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 110142 31200 110198 32400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 246762 31200 246818 32400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 249246 31200 249302 32400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 251730 31200 251786 32400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 254214 31200 254270 32400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 256698 31200 256754 32400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 259182 31200 259238 32400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 261666 31200 261722 32400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 264150 31200 264206 32400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 266634 31200 266690 32400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 269118 31200 269174 32400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 112626 31200 112682 32400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 271602 31200 271658 32400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 274086 31200 274142 32400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 276570 31200 276626 32400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 279054 31200 279110 32400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 281538 31200 281594 32400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 284022 31200 284078 32400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 286506 31200 286562 32400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 288990 31200 289046 32400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 291474 31200 291530 32400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 293958 31200 294014 32400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 115110 31200 115166 32400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 296442 31200 296498 32400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 298926 31200 298982 32400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 301410 31200 301466 32400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 303894 31200 303950 32400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 306378 31200 306434 32400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 308862 31200 308918 32400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 311346 31200 311402 32400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 313830 31200 313886 32400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 316314 31200 316370 32400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 318798 31200 318854 32400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 117594 31200 117650 32400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 321282 31200 321338 32400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 323766 31200 323822 32400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 326250 31200 326306 32400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 328734 31200 328790 32400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 331218 31200 331274 32400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 333702 31200 333758 32400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 336186 31200 336242 32400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 338670 31200 338726 32400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 341154 31200 341210 32400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 343638 31200 343694 32400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 120078 31200 120134 32400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 16854 -400 16910 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 274454 -400 274510 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 277030 -400 277086 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 279606 -400 279662 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 282182 -400 282238 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 284758 -400 284814 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 287334 -400 287390 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 289910 -400 289966 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 292486 -400 292542 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 295062 -400 295118 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 297638 -400 297694 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 42614 -400 42670 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 300214 -400 300270 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 302790 -400 302846 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 305366 -400 305422 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 307942 -400 307998 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 310518 -400 310574 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 313094 -400 313150 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 315670 -400 315726 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 318246 -400 318302 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 320822 -400 320878 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 323398 -400 323454 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 45190 -400 45246 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 325974 -400 326030 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 328550 -400 328606 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 331126 -400 331182 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 333702 -400 333758 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 336278 -400 336334 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 338854 -400 338910 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 341430 -400 341486 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 344006 -400 344062 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 47766 -400 47822 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 50342 -400 50398 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 52918 -400 52974 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 55494 -400 55550 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 58070 -400 58126 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 60646 -400 60702 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 63222 -400 63278 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 65798 -400 65854 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 19430 -400 19486 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 68374 -400 68430 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 70950 -400 71006 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 73526 -400 73582 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 76102 -400 76158 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 78678 -400 78734 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 81254 -400 81310 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 83830 -400 83886 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 86406 -400 86462 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 88982 -400 89038 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 91558 -400 91614 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 22006 -400 22062 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 94134 -400 94190 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 96710 -400 96766 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 99286 -400 99342 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 101862 -400 101918 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 104438 -400 104494 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 107014 -400 107070 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 109590 -400 109646 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 112166 -400 112222 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 114742 -400 114798 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 117318 -400 117374 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 24582 -400 24638 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 119894 -400 119950 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 122470 -400 122526 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 125046 -400 125102 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 127622 -400 127678 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 130198 -400 130254 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 132774 -400 132830 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 135350 -400 135406 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 137926 -400 137982 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 140502 -400 140558 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 143078 -400 143134 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 27158 -400 27214 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 145654 -400 145710 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 148230 -400 148286 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 150806 -400 150862 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 153382 -400 153438 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 155958 -400 156014 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 158534 -400 158590 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 161110 -400 161166 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 163686 -400 163742 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 166262 -400 166318 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 168838 -400 168894 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 29734 -400 29790 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 171414 -400 171470 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 173990 -400 174046 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 176566 -400 176622 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 179142 -400 179198 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 181718 -400 181774 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 184294 -400 184350 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 186870 -400 186926 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 189446 -400 189502 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 192022 -400 192078 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 194598 -400 194654 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 32310 -400 32366 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 197174 -400 197230 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 199750 -400 199806 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 202326 -400 202382 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 204902 -400 204958 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 207478 -400 207534 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 210054 -400 210110 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 212630 -400 212686 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 215206 -400 215262 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 217782 -400 217838 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 220358 -400 220414 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 34886 -400 34942 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 222934 -400 222990 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 225510 -400 225566 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 228086 -400 228142 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 230662 -400 230718 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 233238 -400 233294 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 235814 -400 235870 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 238390 -400 238446 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 240966 -400 241022 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 243542 -400 243598 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 246118 -400 246174 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 37462 -400 37518 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 248694 -400 248750 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 251270 -400 251326 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 253846 -400 253902 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 256422 -400 256478 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 258998 -400 259054 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 261574 -400 261630 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 264150 -400 264206 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 266726 -400 266782 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 269302 -400 269358 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 271878 -400 271934 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 40038 -400 40094 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 17498 -400 17554 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 275098 -400 275154 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 277674 -400 277730 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 280250 -400 280306 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 282826 -400 282882 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 285402 -400 285458 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 287978 -400 288034 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 290554 -400 290610 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 293130 -400 293186 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 295706 -400 295762 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 298282 -400 298338 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 43258 -400 43314 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 300858 -400 300914 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 303434 -400 303490 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 306010 -400 306066 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 308586 -400 308642 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 311162 -400 311218 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 313738 -400 313794 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 316314 -400 316370 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 318890 -400 318946 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 321466 -400 321522 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 324042 -400 324098 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 45834 -400 45890 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 326618 -400 326674 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 329194 -400 329250 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 331770 -400 331826 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 334346 -400 334402 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 336922 -400 336978 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 339498 -400 339554 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 342074 -400 342130 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 344650 -400 344706 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 48410 -400 48466 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 50986 -400 51042 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 53562 -400 53618 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 56138 -400 56194 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 58714 -400 58770 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 61290 -400 61346 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 63866 -400 63922 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 66442 -400 66498 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 20074 -400 20130 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 69018 -400 69074 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 71594 -400 71650 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 74170 -400 74226 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 76746 -400 76802 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 79322 -400 79378 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 81898 -400 81954 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 84474 -400 84530 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 87050 -400 87106 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 89626 -400 89682 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 92202 -400 92258 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 22650 -400 22706 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 94778 -400 94834 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 97354 -400 97410 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 99930 -400 99986 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 102506 -400 102562 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 105082 -400 105138 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 107658 -400 107714 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 110234 -400 110290 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 112810 -400 112866 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 115386 -400 115442 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 117962 -400 118018 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 25226 -400 25282 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 120538 -400 120594 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 123114 -400 123170 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 125690 -400 125746 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 128266 -400 128322 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 130842 -400 130898 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 133418 -400 133474 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 135994 -400 136050 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 138570 -400 138626 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 141146 -400 141202 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 143722 -400 143778 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 27802 -400 27858 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 146298 -400 146354 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 148874 -400 148930 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 151450 -400 151506 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 154026 -400 154082 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 156602 -400 156658 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 159178 -400 159234 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 161754 -400 161810 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 164330 -400 164386 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 166906 -400 166962 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 169482 -400 169538 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 30378 -400 30434 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 172058 -400 172114 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 174634 -400 174690 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 177210 -400 177266 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 179786 -400 179842 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 182362 -400 182418 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 184938 -400 184994 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 187514 -400 187570 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 190090 -400 190146 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 192666 -400 192722 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 195242 -400 195298 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 32954 -400 33010 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 197818 -400 197874 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 200394 -400 200450 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 202970 -400 203026 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 205546 -400 205602 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 208122 -400 208178 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 210698 -400 210754 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 213274 -400 213330 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 215850 -400 215906 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 218426 -400 218482 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 221002 -400 221058 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 35530 -400 35586 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 223578 -400 223634 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 226154 -400 226210 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 228730 -400 228786 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 231306 -400 231362 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 233882 -400 233938 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 236458 -400 236514 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 239034 -400 239090 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 241610 -400 241666 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 244186 -400 244242 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 246762 -400 246818 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 38106 -400 38162 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 249338 -400 249394 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 251914 -400 251970 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 254490 -400 254546 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 257066 -400 257122 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 259642 -400 259698 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 262218 -400 262274 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 264794 -400 264850 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 267370 -400 267426 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 269946 -400 270002 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 272522 -400 272578 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 40682 -400 40738 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 98550 31200 98606 32400 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 346950 31200 347006 32400 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 349434 31200 349490 32400 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 351918 31200 351974 32400 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 354402 31200 354458 32400 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 356886 31200 356942 32400 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 359370 31200 359426 32400 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 361854 31200 361910 32400 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 364338 31200 364394 32400 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 366822 31200 366878 32400 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 369306 31200 369362 32400 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 123390 31200 123446 32400 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 371790 31200 371846 32400 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 374274 31200 374330 32400 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 376758 31200 376814 32400 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 379242 31200 379298 32400 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 381726 31200 381782 32400 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 384210 31200 384266 32400 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 386694 31200 386750 32400 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 389178 31200 389234 32400 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 391662 31200 391718 32400 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 394146 31200 394202 32400 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 125874 31200 125930 32400 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 396630 31200 396686 32400 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 399114 31200 399170 32400 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 401598 31200 401654 32400 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 404082 31200 404138 32400 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 406566 31200 406622 32400 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 409050 31200 409106 32400 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 411534 31200 411590 32400 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 414018 31200 414074 32400 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 128358 31200 128414 32400 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 130842 31200 130898 32400 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 133326 31200 133382 32400 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 135810 31200 135866 32400 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 138294 31200 138350 32400 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 140778 31200 140834 32400 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 143262 31200 143318 32400 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 145746 31200 145802 32400 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 101034 31200 101090 32400 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 148230 31200 148286 32400 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 150714 31200 150770 32400 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 153198 31200 153254 32400 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 155682 31200 155738 32400 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 158166 31200 158222 32400 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 160650 31200 160706 32400 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 163134 31200 163190 32400 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 165618 31200 165674 32400 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 168102 31200 168158 32400 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 170586 31200 170642 32400 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 103518 31200 103574 32400 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 173070 31200 173126 32400 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 175554 31200 175610 32400 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 178038 31200 178094 32400 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 180522 31200 180578 32400 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 183006 31200 183062 32400 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 185490 31200 185546 32400 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 187974 31200 188030 32400 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 190458 31200 190514 32400 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 192942 31200 192998 32400 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 195426 31200 195482 32400 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 106002 31200 106058 32400 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 197910 31200 197966 32400 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 200394 31200 200450 32400 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 202878 31200 202934 32400 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 205362 31200 205418 32400 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 207846 31200 207902 32400 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 210330 31200 210386 32400 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 212814 31200 212870 32400 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 215298 31200 215354 32400 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 217782 31200 217838 32400 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 220266 31200 220322 32400 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 108486 31200 108542 32400 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 222750 31200 222806 32400 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 225234 31200 225290 32400 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 227718 31200 227774 32400 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 230202 31200 230258 32400 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 232686 31200 232742 32400 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 235170 31200 235226 32400 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 237654 31200 237710 32400 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 240138 31200 240194 32400 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 242622 31200 242678 32400 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 245106 31200 245162 32400 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 110970 31200 111026 32400 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 247590 31200 247646 32400 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 250074 31200 250130 32400 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 252558 31200 252614 32400 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 255042 31200 255098 32400 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 257526 31200 257582 32400 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 260010 31200 260066 32400 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 262494 31200 262550 32400 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 264978 31200 265034 32400 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 267462 31200 267518 32400 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 269946 31200 270002 32400 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 113454 31200 113510 32400 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 272430 31200 272486 32400 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 274914 31200 274970 32400 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 277398 31200 277454 32400 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 279882 31200 279938 32400 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 282366 31200 282422 32400 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 284850 31200 284906 32400 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 287334 31200 287390 32400 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 289818 31200 289874 32400 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 292302 31200 292358 32400 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 294786 31200 294842 32400 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 115938 31200 115994 32400 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 297270 31200 297326 32400 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 299754 31200 299810 32400 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 302238 31200 302294 32400 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 304722 31200 304778 32400 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 307206 31200 307262 32400 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 309690 31200 309746 32400 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 312174 31200 312230 32400 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 314658 31200 314714 32400 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 317142 31200 317198 32400 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 319626 31200 319682 32400 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 118422 31200 118478 32400 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 322110 31200 322166 32400 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 324594 31200 324650 32400 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 327078 31200 327134 32400 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 329562 31200 329618 32400 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 332046 31200 332102 32400 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 334530 31200 334586 32400 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 337014 31200 337070 32400 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 339498 31200 339554 32400 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 341982 31200 342038 32400 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 344466 31200 344522 32400 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 120906 31200 120962 32400 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 18142 -400 18198 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 275742 -400 275798 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 278318 -400 278374 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 280894 -400 280950 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 283470 -400 283526 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 286046 -400 286102 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 288622 -400 288678 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 291198 -400 291254 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 293774 -400 293830 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 296350 -400 296406 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 298926 -400 298982 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 43902 -400 43958 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 301502 -400 301558 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 304078 -400 304134 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 306654 -400 306710 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 309230 -400 309286 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 311806 -400 311862 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 314382 -400 314438 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 316958 -400 317014 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 319534 -400 319590 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 322110 -400 322166 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 324686 -400 324742 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 46478 -400 46534 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 327262 -400 327318 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 329838 -400 329894 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 332414 -400 332470 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 334990 -400 335046 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 337566 -400 337622 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 340142 -400 340198 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 342718 -400 342774 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 345294 -400 345350 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 49054 -400 49110 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 51630 -400 51686 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 54206 -400 54262 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 56782 -400 56838 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 59358 -400 59414 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 61934 -400 61990 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 64510 -400 64566 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 67086 -400 67142 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 20718 -400 20774 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 69662 -400 69718 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 72238 -400 72294 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 74814 -400 74870 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 77390 -400 77446 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 79966 -400 80022 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 82542 -400 82598 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 85118 -400 85174 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 87694 -400 87750 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 90270 -400 90326 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 92846 -400 92902 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 23294 -400 23350 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 95422 -400 95478 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 97998 -400 98054 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 100574 -400 100630 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 103150 -400 103206 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 105726 -400 105782 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 108302 -400 108358 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 110878 -400 110934 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 113454 -400 113510 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 116030 -400 116086 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 118606 -400 118662 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 25870 -400 25926 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 121182 -400 121238 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 123758 -400 123814 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 126334 -400 126390 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 128910 -400 128966 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 131486 -400 131542 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 134062 -400 134118 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 136638 -400 136694 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 139214 -400 139270 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 141790 -400 141846 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 144366 -400 144422 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 28446 -400 28502 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 146942 -400 146998 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 149518 -400 149574 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 152094 -400 152150 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 154670 -400 154726 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 157246 -400 157302 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 159822 -400 159878 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 162398 -400 162454 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 164974 -400 165030 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 167550 -400 167606 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 170126 -400 170182 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 31022 -400 31078 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 172702 -400 172758 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 175278 -400 175334 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 177854 -400 177910 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 180430 -400 180486 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 183006 -400 183062 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 185582 -400 185638 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 188158 -400 188214 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 190734 -400 190790 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 193310 -400 193366 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 195886 -400 195942 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 33598 -400 33654 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 198462 -400 198518 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 201038 -400 201094 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 203614 -400 203670 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 206190 -400 206246 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 208766 -400 208822 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 211342 -400 211398 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 213918 -400 213974 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 216494 -400 216550 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 219070 -400 219126 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 221646 -400 221702 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 36174 -400 36230 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 224222 -400 224278 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 226798 -400 226854 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 229374 -400 229430 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 231950 -400 232006 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 234526 -400 234582 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 237102 -400 237158 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 239678 -400 239734 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 242254 -400 242310 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 244830 -400 244886 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 247406 -400 247462 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 38750 -400 38806 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 249982 -400 250038 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 252558 -400 252614 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 255134 -400 255190 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 257710 -400 257766 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 260286 -400 260342 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 262862 -400 262918 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 265438 -400 265494 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 268014 -400 268070 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 270590 -400 270646 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 273166 -400 273222 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 41326 -400 41382 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal3 s 423200 5448 424400 5568 6 mprj_ack_i_core
port 900 nsew signal output
rlabel metal2 s 10782 31200 10838 32400 6 mprj_ack_i_user
port 901 nsew signal input
rlabel metal2 s 345938 -400 345994 800 6 mprj_adr_o_core[0]
port 902 nsew signal input
rlabel metal2 s 352378 -400 352434 800 6 mprj_adr_o_core[10]
port 903 nsew signal input
rlabel metal2 s 353022 -400 353078 800 6 mprj_adr_o_core[11]
port 904 nsew signal input
rlabel metal2 s 353666 -400 353722 800 6 mprj_adr_o_core[12]
port 905 nsew signal input
rlabel metal2 s 354310 -400 354366 800 6 mprj_adr_o_core[13]
port 906 nsew signal input
rlabel metal2 s 354954 -400 355010 800 6 mprj_adr_o_core[14]
port 907 nsew signal input
rlabel metal2 s 355598 -400 355654 800 6 mprj_adr_o_core[15]
port 908 nsew signal input
rlabel metal2 s 356242 -400 356298 800 6 mprj_adr_o_core[16]
port 909 nsew signal input
rlabel metal2 s 356886 -400 356942 800 6 mprj_adr_o_core[17]
port 910 nsew signal input
rlabel metal2 s 357530 -400 357586 800 6 mprj_adr_o_core[18]
port 911 nsew signal input
rlabel metal2 s 358174 -400 358230 800 6 mprj_adr_o_core[19]
port 912 nsew signal input
rlabel metal2 s 346582 -400 346638 800 6 mprj_adr_o_core[1]
port 913 nsew signal input
rlabel metal2 s 358818 -400 358874 800 6 mprj_adr_o_core[20]
port 914 nsew signal input
rlabel metal2 s 359462 -400 359518 800 6 mprj_adr_o_core[21]
port 915 nsew signal input
rlabel metal2 s 360106 -400 360162 800 6 mprj_adr_o_core[22]
port 916 nsew signal input
rlabel metal2 s 360750 -400 360806 800 6 mprj_adr_o_core[23]
port 917 nsew signal input
rlabel metal2 s 361394 -400 361450 800 6 mprj_adr_o_core[24]
port 918 nsew signal input
rlabel metal2 s 362038 -400 362094 800 6 mprj_adr_o_core[25]
port 919 nsew signal input
rlabel metal2 s 362682 -400 362738 800 6 mprj_adr_o_core[26]
port 920 nsew signal input
rlabel metal2 s 363326 -400 363382 800 6 mprj_adr_o_core[27]
port 921 nsew signal input
rlabel metal2 s 363970 -400 364026 800 6 mprj_adr_o_core[28]
port 922 nsew signal input
rlabel metal2 s 364614 -400 364670 800 6 mprj_adr_o_core[29]
port 923 nsew signal input
rlabel metal2 s 347226 -400 347282 800 6 mprj_adr_o_core[2]
port 924 nsew signal input
rlabel metal2 s 365258 -400 365314 800 6 mprj_adr_o_core[30]
port 925 nsew signal input
rlabel metal2 s 365902 -400 365958 800 6 mprj_adr_o_core[31]
port 926 nsew signal input
rlabel metal2 s 347870 -400 347926 800 6 mprj_adr_o_core[3]
port 927 nsew signal input
rlabel metal2 s 348514 -400 348570 800 6 mprj_adr_o_core[4]
port 928 nsew signal input
rlabel metal2 s 349158 -400 349214 800 6 mprj_adr_o_core[5]
port 929 nsew signal input
rlabel metal2 s 349802 -400 349858 800 6 mprj_adr_o_core[6]
port 930 nsew signal input
rlabel metal2 s 350446 -400 350502 800 6 mprj_adr_o_core[7]
port 931 nsew signal input
rlabel metal2 s 351090 -400 351146 800 6 mprj_adr_o_core[8]
port 932 nsew signal input
rlabel metal2 s 351734 -400 351790 800 6 mprj_adr_o_core[9]
port 933 nsew signal input
rlabel metal2 s 14094 31200 14150 32400 6 mprj_adr_o_user[0]
port 934 nsew signal output
rlabel metal2 s 42246 31200 42302 32400 6 mprj_adr_o_user[10]
port 935 nsew signal output
rlabel metal2 s 44730 31200 44786 32400 6 mprj_adr_o_user[11]
port 936 nsew signal output
rlabel metal2 s 47214 31200 47270 32400 6 mprj_adr_o_user[12]
port 937 nsew signal output
rlabel metal2 s 49698 31200 49754 32400 6 mprj_adr_o_user[13]
port 938 nsew signal output
rlabel metal2 s 52182 31200 52238 32400 6 mprj_adr_o_user[14]
port 939 nsew signal output
rlabel metal2 s 54666 31200 54722 32400 6 mprj_adr_o_user[15]
port 940 nsew signal output
rlabel metal2 s 57150 31200 57206 32400 6 mprj_adr_o_user[16]
port 941 nsew signal output
rlabel metal2 s 59634 31200 59690 32400 6 mprj_adr_o_user[17]
port 942 nsew signal output
rlabel metal2 s 62118 31200 62174 32400 6 mprj_adr_o_user[18]
port 943 nsew signal output
rlabel metal2 s 64602 31200 64658 32400 6 mprj_adr_o_user[19]
port 944 nsew signal output
rlabel metal2 s 17406 31200 17462 32400 6 mprj_adr_o_user[1]
port 945 nsew signal output
rlabel metal2 s 67086 31200 67142 32400 6 mprj_adr_o_user[20]
port 946 nsew signal output
rlabel metal2 s 69570 31200 69626 32400 6 mprj_adr_o_user[21]
port 947 nsew signal output
rlabel metal2 s 72054 31200 72110 32400 6 mprj_adr_o_user[22]
port 948 nsew signal output
rlabel metal2 s 74538 31200 74594 32400 6 mprj_adr_o_user[23]
port 949 nsew signal output
rlabel metal2 s 77022 31200 77078 32400 6 mprj_adr_o_user[24]
port 950 nsew signal output
rlabel metal2 s 79506 31200 79562 32400 6 mprj_adr_o_user[25]
port 951 nsew signal output
rlabel metal2 s 81990 31200 82046 32400 6 mprj_adr_o_user[26]
port 952 nsew signal output
rlabel metal2 s 84474 31200 84530 32400 6 mprj_adr_o_user[27]
port 953 nsew signal output
rlabel metal2 s 86958 31200 87014 32400 6 mprj_adr_o_user[28]
port 954 nsew signal output
rlabel metal2 s 89442 31200 89498 32400 6 mprj_adr_o_user[29]
port 955 nsew signal output
rlabel metal2 s 20718 31200 20774 32400 6 mprj_adr_o_user[2]
port 956 nsew signal output
rlabel metal2 s 91926 31200 91982 32400 6 mprj_adr_o_user[30]
port 957 nsew signal output
rlabel metal2 s 94410 31200 94466 32400 6 mprj_adr_o_user[31]
port 958 nsew signal output
rlabel metal2 s 24030 31200 24086 32400 6 mprj_adr_o_user[3]
port 959 nsew signal output
rlabel metal2 s 27342 31200 27398 32400 6 mprj_adr_o_user[4]
port 960 nsew signal output
rlabel metal2 s 29826 31200 29882 32400 6 mprj_adr_o_user[5]
port 961 nsew signal output
rlabel metal2 s 32310 31200 32366 32400 6 mprj_adr_o_user[6]
port 962 nsew signal output
rlabel metal2 s 34794 31200 34850 32400 6 mprj_adr_o_user[7]
port 963 nsew signal output
rlabel metal2 s 37278 31200 37334 32400 6 mprj_adr_o_user[8]
port 964 nsew signal output
rlabel metal2 s 39762 31200 39818 32400 6 mprj_adr_o_user[9]
port 965 nsew signal output
rlabel metal3 s 423200 1776 424400 1896 6 mprj_cyc_o_core
port 966 nsew signal input
rlabel metal2 s 11610 31200 11666 32400 6 mprj_cyc_o_user
port 967 nsew signal output
rlabel metal2 s 366546 -400 366602 800 6 mprj_dat_i_core[0]
port 968 nsew signal output
rlabel metal2 s 372986 -400 373042 800 6 mprj_dat_i_core[10]
port 969 nsew signal output
rlabel metal2 s 373630 -400 373686 800 6 mprj_dat_i_core[11]
port 970 nsew signal output
rlabel metal2 s 374274 -400 374330 800 6 mprj_dat_i_core[12]
port 971 nsew signal output
rlabel metal2 s 374918 -400 374974 800 6 mprj_dat_i_core[13]
port 972 nsew signal output
rlabel metal2 s 375562 -400 375618 800 6 mprj_dat_i_core[14]
port 973 nsew signal output
rlabel metal2 s 376206 -400 376262 800 6 mprj_dat_i_core[15]
port 974 nsew signal output
rlabel metal2 s 376850 -400 376906 800 6 mprj_dat_i_core[16]
port 975 nsew signal output
rlabel metal2 s 377494 -400 377550 800 6 mprj_dat_i_core[17]
port 976 nsew signal output
rlabel metal2 s 378138 -400 378194 800 6 mprj_dat_i_core[18]
port 977 nsew signal output
rlabel metal2 s 378782 -400 378838 800 6 mprj_dat_i_core[19]
port 978 nsew signal output
rlabel metal2 s 367190 -400 367246 800 6 mprj_dat_i_core[1]
port 979 nsew signal output
rlabel metal2 s 379426 -400 379482 800 6 mprj_dat_i_core[20]
port 980 nsew signal output
rlabel metal2 s 380070 -400 380126 800 6 mprj_dat_i_core[21]
port 981 nsew signal output
rlabel metal2 s 380714 -400 380770 800 6 mprj_dat_i_core[22]
port 982 nsew signal output
rlabel metal2 s 381358 -400 381414 800 6 mprj_dat_i_core[23]
port 983 nsew signal output
rlabel metal2 s 382002 -400 382058 800 6 mprj_dat_i_core[24]
port 984 nsew signal output
rlabel metal2 s 382646 -400 382702 800 6 mprj_dat_i_core[25]
port 985 nsew signal output
rlabel metal2 s 383290 -400 383346 800 6 mprj_dat_i_core[26]
port 986 nsew signal output
rlabel metal2 s 383934 -400 383990 800 6 mprj_dat_i_core[27]
port 987 nsew signal output
rlabel metal2 s 384578 -400 384634 800 6 mprj_dat_i_core[28]
port 988 nsew signal output
rlabel metal2 s 385222 -400 385278 800 6 mprj_dat_i_core[29]
port 989 nsew signal output
rlabel metal2 s 367834 -400 367890 800 6 mprj_dat_i_core[2]
port 990 nsew signal output
rlabel metal2 s 385866 -400 385922 800 6 mprj_dat_i_core[30]
port 991 nsew signal output
rlabel metal2 s 386510 -400 386566 800 6 mprj_dat_i_core[31]
port 992 nsew signal output
rlabel metal2 s 368478 -400 368534 800 6 mprj_dat_i_core[3]
port 993 nsew signal output
rlabel metal2 s 369122 -400 369178 800 6 mprj_dat_i_core[4]
port 994 nsew signal output
rlabel metal2 s 369766 -400 369822 800 6 mprj_dat_i_core[5]
port 995 nsew signal output
rlabel metal2 s 370410 -400 370466 800 6 mprj_dat_i_core[6]
port 996 nsew signal output
rlabel metal2 s 371054 -400 371110 800 6 mprj_dat_i_core[7]
port 997 nsew signal output
rlabel metal2 s 371698 -400 371754 800 6 mprj_dat_i_core[8]
port 998 nsew signal output
rlabel metal2 s 372342 -400 372398 800 6 mprj_dat_i_core[9]
port 999 nsew signal output
rlabel metal2 s 14922 31200 14978 32400 6 mprj_dat_i_user[0]
port 1000 nsew signal input
rlabel metal2 s 43074 31200 43130 32400 6 mprj_dat_i_user[10]
port 1001 nsew signal input
rlabel metal2 s 45558 31200 45614 32400 6 mprj_dat_i_user[11]
port 1002 nsew signal input
rlabel metal2 s 48042 31200 48098 32400 6 mprj_dat_i_user[12]
port 1003 nsew signal input
rlabel metal2 s 50526 31200 50582 32400 6 mprj_dat_i_user[13]
port 1004 nsew signal input
rlabel metal2 s 53010 31200 53066 32400 6 mprj_dat_i_user[14]
port 1005 nsew signal input
rlabel metal2 s 55494 31200 55550 32400 6 mprj_dat_i_user[15]
port 1006 nsew signal input
rlabel metal2 s 57978 31200 58034 32400 6 mprj_dat_i_user[16]
port 1007 nsew signal input
rlabel metal2 s 60462 31200 60518 32400 6 mprj_dat_i_user[17]
port 1008 nsew signal input
rlabel metal2 s 62946 31200 63002 32400 6 mprj_dat_i_user[18]
port 1009 nsew signal input
rlabel metal2 s 65430 31200 65486 32400 6 mprj_dat_i_user[19]
port 1010 nsew signal input
rlabel metal2 s 18234 31200 18290 32400 6 mprj_dat_i_user[1]
port 1011 nsew signal input
rlabel metal2 s 67914 31200 67970 32400 6 mprj_dat_i_user[20]
port 1012 nsew signal input
rlabel metal2 s 70398 31200 70454 32400 6 mprj_dat_i_user[21]
port 1013 nsew signal input
rlabel metal2 s 72882 31200 72938 32400 6 mprj_dat_i_user[22]
port 1014 nsew signal input
rlabel metal2 s 75366 31200 75422 32400 6 mprj_dat_i_user[23]
port 1015 nsew signal input
rlabel metal2 s 77850 31200 77906 32400 6 mprj_dat_i_user[24]
port 1016 nsew signal input
rlabel metal2 s 80334 31200 80390 32400 6 mprj_dat_i_user[25]
port 1017 nsew signal input
rlabel metal2 s 82818 31200 82874 32400 6 mprj_dat_i_user[26]
port 1018 nsew signal input
rlabel metal2 s 85302 31200 85358 32400 6 mprj_dat_i_user[27]
port 1019 nsew signal input
rlabel metal2 s 87786 31200 87842 32400 6 mprj_dat_i_user[28]
port 1020 nsew signal input
rlabel metal2 s 90270 31200 90326 32400 6 mprj_dat_i_user[29]
port 1021 nsew signal input
rlabel metal2 s 21546 31200 21602 32400 6 mprj_dat_i_user[2]
port 1022 nsew signal input
rlabel metal2 s 92754 31200 92810 32400 6 mprj_dat_i_user[30]
port 1023 nsew signal input
rlabel metal2 s 95238 31200 95294 32400 6 mprj_dat_i_user[31]
port 1024 nsew signal input
rlabel metal2 s 24858 31200 24914 32400 6 mprj_dat_i_user[3]
port 1025 nsew signal input
rlabel metal2 s 28170 31200 28226 32400 6 mprj_dat_i_user[4]
port 1026 nsew signal input
rlabel metal2 s 30654 31200 30710 32400 6 mprj_dat_i_user[5]
port 1027 nsew signal input
rlabel metal2 s 33138 31200 33194 32400 6 mprj_dat_i_user[6]
port 1028 nsew signal input
rlabel metal2 s 35622 31200 35678 32400 6 mprj_dat_i_user[7]
port 1029 nsew signal input
rlabel metal2 s 38106 31200 38162 32400 6 mprj_dat_i_user[8]
port 1030 nsew signal input
rlabel metal2 s 40590 31200 40646 32400 6 mprj_dat_i_user[9]
port 1031 nsew signal input
rlabel metal2 s 387154 -400 387210 800 6 mprj_dat_o_core[0]
port 1032 nsew signal input
rlabel metal2 s 393594 -400 393650 800 6 mprj_dat_o_core[10]
port 1033 nsew signal input
rlabel metal2 s 394238 -400 394294 800 6 mprj_dat_o_core[11]
port 1034 nsew signal input
rlabel metal2 s 394882 -400 394938 800 6 mprj_dat_o_core[12]
port 1035 nsew signal input
rlabel metal2 s 395526 -400 395582 800 6 mprj_dat_o_core[13]
port 1036 nsew signal input
rlabel metal2 s 396170 -400 396226 800 6 mprj_dat_o_core[14]
port 1037 nsew signal input
rlabel metal2 s 396814 -400 396870 800 6 mprj_dat_o_core[15]
port 1038 nsew signal input
rlabel metal2 s 397458 -400 397514 800 6 mprj_dat_o_core[16]
port 1039 nsew signal input
rlabel metal2 s 398102 -400 398158 800 6 mprj_dat_o_core[17]
port 1040 nsew signal input
rlabel metal2 s 398746 -400 398802 800 6 mprj_dat_o_core[18]
port 1041 nsew signal input
rlabel metal2 s 399390 -400 399446 800 6 mprj_dat_o_core[19]
port 1042 nsew signal input
rlabel metal2 s 387798 -400 387854 800 6 mprj_dat_o_core[1]
port 1043 nsew signal input
rlabel metal2 s 400034 -400 400090 800 6 mprj_dat_o_core[20]
port 1044 nsew signal input
rlabel metal2 s 400678 -400 400734 800 6 mprj_dat_o_core[21]
port 1045 nsew signal input
rlabel metal2 s 401322 -400 401378 800 6 mprj_dat_o_core[22]
port 1046 nsew signal input
rlabel metal2 s 401966 -400 402022 800 6 mprj_dat_o_core[23]
port 1047 nsew signal input
rlabel metal2 s 402610 -400 402666 800 6 mprj_dat_o_core[24]
port 1048 nsew signal input
rlabel metal2 s 403254 -400 403310 800 6 mprj_dat_o_core[25]
port 1049 nsew signal input
rlabel metal2 s 403898 -400 403954 800 6 mprj_dat_o_core[26]
port 1050 nsew signal input
rlabel metal2 s 404542 -400 404598 800 6 mprj_dat_o_core[27]
port 1051 nsew signal input
rlabel metal2 s 405186 -400 405242 800 6 mprj_dat_o_core[28]
port 1052 nsew signal input
rlabel metal2 s 405830 -400 405886 800 6 mprj_dat_o_core[29]
port 1053 nsew signal input
rlabel metal2 s 388442 -400 388498 800 6 mprj_dat_o_core[2]
port 1054 nsew signal input
rlabel metal2 s 406474 -400 406530 800 6 mprj_dat_o_core[30]
port 1055 nsew signal input
rlabel metal2 s 407118 -400 407174 800 6 mprj_dat_o_core[31]
port 1056 nsew signal input
rlabel metal2 s 389086 -400 389142 800 6 mprj_dat_o_core[3]
port 1057 nsew signal input
rlabel metal2 s 389730 -400 389786 800 6 mprj_dat_o_core[4]
port 1058 nsew signal input
rlabel metal2 s 390374 -400 390430 800 6 mprj_dat_o_core[5]
port 1059 nsew signal input
rlabel metal2 s 391018 -400 391074 800 6 mprj_dat_o_core[6]
port 1060 nsew signal input
rlabel metal2 s 391662 -400 391718 800 6 mprj_dat_o_core[7]
port 1061 nsew signal input
rlabel metal2 s 392306 -400 392362 800 6 mprj_dat_o_core[8]
port 1062 nsew signal input
rlabel metal2 s 392950 -400 393006 800 6 mprj_dat_o_core[9]
port 1063 nsew signal input
rlabel metal2 s 15750 31200 15806 32400 6 mprj_dat_o_user[0]
port 1064 nsew signal output
rlabel metal2 s 43902 31200 43958 32400 6 mprj_dat_o_user[10]
port 1065 nsew signal output
rlabel metal2 s 46386 31200 46442 32400 6 mprj_dat_o_user[11]
port 1066 nsew signal output
rlabel metal2 s 48870 31200 48926 32400 6 mprj_dat_o_user[12]
port 1067 nsew signal output
rlabel metal2 s 51354 31200 51410 32400 6 mprj_dat_o_user[13]
port 1068 nsew signal output
rlabel metal2 s 53838 31200 53894 32400 6 mprj_dat_o_user[14]
port 1069 nsew signal output
rlabel metal2 s 56322 31200 56378 32400 6 mprj_dat_o_user[15]
port 1070 nsew signal output
rlabel metal2 s 58806 31200 58862 32400 6 mprj_dat_o_user[16]
port 1071 nsew signal output
rlabel metal2 s 61290 31200 61346 32400 6 mprj_dat_o_user[17]
port 1072 nsew signal output
rlabel metal2 s 63774 31200 63830 32400 6 mprj_dat_o_user[18]
port 1073 nsew signal output
rlabel metal2 s 66258 31200 66314 32400 6 mprj_dat_o_user[19]
port 1074 nsew signal output
rlabel metal2 s 19062 31200 19118 32400 6 mprj_dat_o_user[1]
port 1075 nsew signal output
rlabel metal2 s 68742 31200 68798 32400 6 mprj_dat_o_user[20]
port 1076 nsew signal output
rlabel metal2 s 71226 31200 71282 32400 6 mprj_dat_o_user[21]
port 1077 nsew signal output
rlabel metal2 s 73710 31200 73766 32400 6 mprj_dat_o_user[22]
port 1078 nsew signal output
rlabel metal2 s 76194 31200 76250 32400 6 mprj_dat_o_user[23]
port 1079 nsew signal output
rlabel metal2 s 78678 31200 78734 32400 6 mprj_dat_o_user[24]
port 1080 nsew signal output
rlabel metal2 s 81162 31200 81218 32400 6 mprj_dat_o_user[25]
port 1081 nsew signal output
rlabel metal2 s 83646 31200 83702 32400 6 mprj_dat_o_user[26]
port 1082 nsew signal output
rlabel metal2 s 86130 31200 86186 32400 6 mprj_dat_o_user[27]
port 1083 nsew signal output
rlabel metal2 s 88614 31200 88670 32400 6 mprj_dat_o_user[28]
port 1084 nsew signal output
rlabel metal2 s 91098 31200 91154 32400 6 mprj_dat_o_user[29]
port 1085 nsew signal output
rlabel metal2 s 22374 31200 22430 32400 6 mprj_dat_o_user[2]
port 1086 nsew signal output
rlabel metal2 s 93582 31200 93638 32400 6 mprj_dat_o_user[30]
port 1087 nsew signal output
rlabel metal2 s 96066 31200 96122 32400 6 mprj_dat_o_user[31]
port 1088 nsew signal output
rlabel metal2 s 25686 31200 25742 32400 6 mprj_dat_o_user[3]
port 1089 nsew signal output
rlabel metal2 s 28998 31200 29054 32400 6 mprj_dat_o_user[4]
port 1090 nsew signal output
rlabel metal2 s 31482 31200 31538 32400 6 mprj_dat_o_user[5]
port 1091 nsew signal output
rlabel metal2 s 33966 31200 34022 32400 6 mprj_dat_o_user[6]
port 1092 nsew signal output
rlabel metal2 s 36450 31200 36506 32400 6 mprj_dat_o_user[7]
port 1093 nsew signal output
rlabel metal2 s 38934 31200 38990 32400 6 mprj_dat_o_user[8]
port 1094 nsew signal output
rlabel metal2 s 41418 31200 41474 32400 6 mprj_dat_o_user[9]
port 1095 nsew signal output
rlabel metal2 s 407762 -400 407818 800 6 mprj_iena_wb
port 1096 nsew signal input
rlabel metal3 s 423200 6672 424400 6792 6 mprj_sel_o_core[0]
port 1097 nsew signal input
rlabel metal3 s 423200 7896 424400 8016 6 mprj_sel_o_core[1]
port 1098 nsew signal input
rlabel metal3 s 423200 9120 424400 9240 6 mprj_sel_o_core[2]
port 1099 nsew signal input
rlabel metal3 s 423200 10344 424400 10464 6 mprj_sel_o_core[3]
port 1100 nsew signal input
rlabel metal2 s 16578 31200 16634 32400 6 mprj_sel_o_user[0]
port 1101 nsew signal output
rlabel metal2 s 19890 31200 19946 32400 6 mprj_sel_o_user[1]
port 1102 nsew signal output
rlabel metal2 s 23202 31200 23258 32400 6 mprj_sel_o_user[2]
port 1103 nsew signal output
rlabel metal2 s 26514 31200 26570 32400 6 mprj_sel_o_user[3]
port 1104 nsew signal output
rlabel metal3 s 423200 3000 424400 3120 6 mprj_stb_o_core
port 1105 nsew signal input
rlabel metal2 s 12438 31200 12494 32400 6 mprj_stb_o_user
port 1106 nsew signal output
rlabel metal3 s 423200 4224 424400 4344 6 mprj_we_o_core
port 1107 nsew signal input
rlabel metal2 s 13266 31200 13322 32400 6 mprj_we_o_user
port 1108 nsew signal output
rlabel metal3 s 423200 18912 424400 19032 6 user1_vcc_powergood
port 1109 nsew signal output
rlabel metal3 s 423200 20136 424400 20256 6 user1_vdd_powergood
port 1110 nsew signal output
rlabel metal3 s 423200 21360 424400 21480 6 user2_vcc_powergood
port 1111 nsew signal output
rlabel metal3 s 423200 22584 424400 22704 6 user2_vdd_powergood
port 1112 nsew signal output
rlabel metal2 s 9126 31200 9182 32400 6 user_clock
port 1113 nsew signal output
rlabel metal2 s 414846 31200 414902 32400 6 user_clock2
port 1114 nsew signal output
rlabel metal3 s 423200 23808 424400 23928 6 user_irq[0]
port 1115 nsew signal output
rlabel metal3 s 423200 25032 424400 25152 6 user_irq[1]
port 1116 nsew signal output
rlabel metal3 s 423200 26256 424400 26376 6 user_irq[2]
port 1117 nsew signal output
rlabel metal3 s 423200 11568 424400 11688 6 user_irq_core[0]
port 1118 nsew signal input
rlabel metal3 s 423200 12792 424400 12912 6 user_irq_core[1]
port 1119 nsew signal input
rlabel metal3 s 423200 14016 424400 14136 6 user_irq_core[2]
port 1120 nsew signal input
rlabel metal3 s 423200 27480 424400 27600 6 user_irq_ena[0]
port 1121 nsew signal input
rlabel metal3 s 423200 28704 424400 28824 6 user_irq_ena[1]
port 1122 nsew signal input
rlabel metal3 s 423200 29928 424400 30048 6 user_irq_ena[2]
port 1123 nsew signal input
rlabel metal2 s 9954 31200 10010 32400 6 user_reset
port 1124 nsew signal output
rlabel metal4 s 5014 1040 5194 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 20064 1040 20244 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 35114 1040 35294 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 50164 1040 50344 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 65214 1040 65394 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 80264 1040 80444 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 95314 1040 95494 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 110364 1040 110544 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 125414 1040 125594 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 140464 1040 140644 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 155514 1040 155694 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 170564 1040 170744 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 185614 1040 185794 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 200664 1040 200844 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 215714 1040 215894 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 230764 1040 230944 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 245814 1040 245994 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 260864 1040 261044 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 275914 1040 276094 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 290964 1040 291144 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 306014 1040 306194 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 321064 1040 321244 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 336114 1040 336294 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 351164 1040 351344 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 366214 1040 366394 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 381264 1040 381444 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 396314 1040 396494 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 411364 1040 411544 30512 6 vccd
port 1125 nsew power bidirectional
rlabel metal4 s 141284 1040 141464 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 156334 1040 156514 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 171384 1040 171564 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 186434 1040 186614 30512 6 vccd1
port 1126 nsew power bidirectional
rlabel metal4 s 66854 1040 67034 30512 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 76854 1040 77034 30512 6 vccd2
port 1127 nsew power bidirectional
rlabel metal4 s 255814 1040 255994 30512 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 270864 1040 271044 30512 6 vdda1
port 1128 nsew power bidirectional
rlabel metal4 s 256614 1040 256794 30512 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 271664 1040 271844 30512 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 263194 1040 263374 30512 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 278244 1040 278424 30512 6 vssa1
port 1130 nsew ground bidirectional
rlabel metal4 s 263994 1040 264174 30512 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 279044 1040 279224 30512 6 vssa2
port 1131 nsew ground bidirectional
rlabel metal4 s 12394 1040 12574 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 27444 1040 27624 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 42494 1040 42674 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 57544 1040 57724 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 72594 1040 72774 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 87644 1040 87824 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 102694 1040 102874 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 117744 1040 117924 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 132794 1040 132974 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 147844 1040 148024 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 162894 1040 163074 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 177944 1040 178124 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 192994 1040 193174 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 208044 1040 208224 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 223094 1040 223274 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 238144 1040 238324 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 253194 1040 253374 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 268244 1040 268424 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 283294 1040 283474 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 298344 1040 298524 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 313394 1040 313574 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 328444 1040 328624 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 343494 1040 343674 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 358544 1040 358724 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 373594 1040 373774 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 388644 1040 388824 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 403694 1040 403874 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 418744 1040 418924 30512 6 vssd
port 1132 nsew ground bidirectional
rlabel metal4 s 148664 1040 148844 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 163714 1040 163894 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 178764 1040 178944 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 193814 1040 193994 30512 6 vssd1
port 1133 nsew ground bidirectional
rlabel metal4 s 71034 1040 71214 30512 6 vssd2
port 1134 nsew ground bidirectional
rlabel metal4 s 81034 1040 81214 30512 6 vssd2
port 1134 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 424000 32000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16423370
string GDS_FILE /home/hosni/My_forks/FINAL/caravel/openlane/mgmt_protect/runs/22_10_13_09_37/results/signoff/mgmt_protect.magic.gds
string GDS_START 687500
<< end >>

