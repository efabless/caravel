magic
tech sky130A
magscale 1 2
timestamp 1665958328
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 510338 1007156 510344 1007208
rect 510396 1007196 510402 1007208
rect 518158 1007196 518164 1007208
rect 510396 1007168 518164 1007196
rect 510396 1007156 510402 1007168
rect 518158 1007156 518164 1007168
rect 518216 1007156 518222 1007208
rect 431678 1007088 431684 1007140
rect 431736 1007128 431742 1007140
rect 434622 1007128 434628 1007140
rect 431736 1007100 434628 1007128
rect 431736 1007088 431742 1007100
rect 434622 1007088 434628 1007100
rect 434680 1007088 434686 1007140
rect 505002 1007020 505008 1007072
rect 505060 1007060 505066 1007072
rect 515582 1007060 515588 1007072
rect 505060 1007032 515588 1007060
rect 505060 1007020 505066 1007032
rect 515582 1007020 515588 1007032
rect 515640 1007020 515646 1007072
rect 427998 1006952 428004 1007004
rect 428056 1006992 428062 1007004
rect 428056 1006964 441614 1006992
rect 428056 1006952 428062 1006964
rect 359734 1006884 359740 1006936
rect 359792 1006924 359798 1006936
rect 374638 1006924 374644 1006936
rect 359792 1006896 374644 1006924
rect 359792 1006884 359798 1006896
rect 374638 1006884 374644 1006896
rect 374696 1006884 374702 1006936
rect 428366 1006816 428372 1006868
rect 428424 1006856 428430 1006868
rect 436738 1006856 436744 1006868
rect 428424 1006828 436744 1006856
rect 428424 1006816 428430 1006828
rect 436738 1006816 436744 1006828
rect 436796 1006816 436802 1006868
rect 145558 1006748 145564 1006800
rect 145616 1006788 145622 1006800
rect 151722 1006788 151728 1006800
rect 145616 1006760 151728 1006788
rect 145616 1006748 145622 1006760
rect 151722 1006748 151728 1006760
rect 151780 1006748 151786 1006800
rect 359366 1006748 359372 1006800
rect 359424 1006788 359430 1006800
rect 369118 1006788 369124 1006800
rect 359424 1006760 369124 1006788
rect 359424 1006748 359430 1006760
rect 369118 1006748 369124 1006760
rect 369176 1006748 369182 1006800
rect 429194 1006680 429200 1006732
rect 429252 1006720 429258 1006732
rect 441586 1006720 441614 1006964
rect 552290 1006952 552296 1007004
rect 552348 1006992 552354 1007004
rect 568022 1006992 568028 1007004
rect 552348 1006964 568028 1006992
rect 552348 1006952 552354 1006964
rect 568022 1006952 568028 1006964
rect 568080 1006952 568086 1007004
rect 505370 1006884 505376 1006936
rect 505428 1006924 505434 1006936
rect 510338 1006924 510344 1006936
rect 505428 1006896 510344 1006924
rect 505428 1006884 505434 1006896
rect 510338 1006884 510344 1006896
rect 510396 1006884 510402 1006936
rect 510522 1006816 510528 1006868
rect 510580 1006856 510586 1006868
rect 520918 1006856 520924 1006868
rect 510580 1006828 520924 1006856
rect 510580 1006816 510586 1006828
rect 520918 1006816 520924 1006828
rect 520976 1006816 520982 1006868
rect 557166 1006748 557172 1006800
rect 557224 1006788 557230 1006800
rect 565262 1006788 565268 1006800
rect 557224 1006760 565268 1006788
rect 557224 1006748 557230 1006760
rect 565262 1006748 565268 1006760
rect 565320 1006748 565326 1006800
rect 451826 1006720 451832 1006732
rect 429252 1006692 431954 1006720
rect 441586 1006692 451832 1006720
rect 429252 1006680 429258 1006692
rect 145742 1006612 145748 1006664
rect 145800 1006652 145806 1006664
rect 145800 1006624 151814 1006652
rect 145800 1006612 145806 1006624
rect 151786 1006584 151814 1006624
rect 360562 1006612 360568 1006664
rect 360620 1006652 360626 1006664
rect 371878 1006652 371884 1006664
rect 360620 1006624 371884 1006652
rect 360620 1006612 360626 1006624
rect 371878 1006612 371884 1006624
rect 371936 1006612 371942 1006664
rect 152090 1006584 152096 1006596
rect 151786 1006556 152096 1006584
rect 152090 1006544 152096 1006556
rect 152148 1006544 152154 1006596
rect 157426 1006544 157432 1006596
rect 157484 1006584 157490 1006596
rect 166258 1006584 166264 1006596
rect 157484 1006556 166264 1006584
rect 157484 1006544 157490 1006556
rect 166258 1006544 166264 1006556
rect 166316 1006544 166322 1006596
rect 431926 1006584 431954 1006692
rect 451826 1006680 451832 1006692
rect 451884 1006680 451890 1006732
rect 505370 1006612 505376 1006664
rect 505428 1006652 505434 1006664
rect 514202 1006652 514208 1006664
rect 505428 1006624 514208 1006652
rect 505428 1006612 505434 1006624
rect 514202 1006612 514208 1006624
rect 514260 1006612 514266 1006664
rect 553118 1006612 553124 1006664
rect 553176 1006652 553182 1006664
rect 562502 1006652 562508 1006664
rect 553176 1006624 562508 1006652
rect 553176 1006612 553182 1006624
rect 562502 1006612 562508 1006624
rect 562560 1006612 562566 1006664
rect 469858 1006584 469864 1006596
rect 431926 1006556 469864 1006584
rect 469858 1006544 469864 1006556
rect 469916 1006544 469922 1006596
rect 144178 1006476 144184 1006528
rect 144236 1006516 144242 1006528
rect 151262 1006516 151268 1006528
rect 144236 1006488 151268 1006516
rect 144236 1006476 144242 1006488
rect 151262 1006476 151268 1006488
rect 151320 1006476 151326 1006528
rect 551094 1006476 551100 1006528
rect 551152 1006516 551158 1006528
rect 556614 1006516 556620 1006528
rect 551152 1006488 556620 1006516
rect 551152 1006476 551158 1006488
rect 556614 1006476 556620 1006488
rect 556672 1006476 556678 1006528
rect 556798 1006476 556804 1006528
rect 556856 1006516 556862 1006528
rect 564434 1006516 564440 1006528
rect 556856 1006488 564440 1006516
rect 556856 1006476 556862 1006488
rect 564434 1006476 564440 1006488
rect 564492 1006476 564498 1006528
rect 94682 1006408 94688 1006460
rect 94740 1006448 94746 1006460
rect 101122 1006448 101128 1006460
rect 94740 1006420 101128 1006448
rect 94740 1006408 94746 1006420
rect 101122 1006408 101128 1006420
rect 101180 1006408 101186 1006460
rect 158622 1006408 158628 1006460
rect 158680 1006448 158686 1006460
rect 173158 1006448 173164 1006460
rect 158680 1006420 173164 1006448
rect 158680 1006408 158686 1006420
rect 173158 1006408 173164 1006420
rect 173216 1006408 173222 1006460
rect 249242 1006408 249248 1006460
rect 249300 1006448 249306 1006460
rect 255314 1006448 255320 1006460
rect 249300 1006420 255320 1006448
rect 249300 1006408 249306 1006420
rect 255314 1006408 255320 1006420
rect 255372 1006408 255378 1006460
rect 361390 1006408 361396 1006460
rect 361448 1006448 361454 1006460
rect 376754 1006448 376760 1006460
rect 361448 1006420 376760 1006448
rect 361448 1006408 361454 1006420
rect 376754 1006408 376760 1006420
rect 376812 1006408 376818 1006460
rect 422662 1006408 422668 1006460
rect 422720 1006448 422726 1006460
rect 422720 1006420 431954 1006448
rect 422720 1006408 422726 1006420
rect 148502 1006340 148508 1006392
rect 148560 1006380 148566 1006392
rect 148560 1006352 151814 1006380
rect 148560 1006340 148566 1006352
rect 96062 1006272 96068 1006324
rect 96120 1006312 96126 1006324
rect 101950 1006312 101956 1006324
rect 96120 1006284 101956 1006312
rect 96120 1006272 96126 1006284
rect 101950 1006272 101956 1006284
rect 102008 1006272 102014 1006324
rect 108482 1006272 108488 1006324
rect 108540 1006312 108546 1006324
rect 126238 1006312 126244 1006324
rect 108540 1006284 126244 1006312
rect 108540 1006272 108546 1006284
rect 126238 1006272 126244 1006284
rect 126296 1006272 126302 1006324
rect 144362 1006204 144368 1006256
rect 144420 1006244 144426 1006256
rect 150894 1006244 150900 1006256
rect 144420 1006216 150900 1006244
rect 144420 1006204 144426 1006216
rect 150894 1006204 150900 1006216
rect 150952 1006204 150958 1006256
rect 93302 1006136 93308 1006188
rect 93360 1006176 93366 1006188
rect 99466 1006176 99472 1006188
rect 93360 1006148 99472 1006176
rect 93360 1006136 93366 1006148
rect 99466 1006136 99472 1006148
rect 99524 1006136 99530 1006188
rect 102962 1006136 102968 1006188
rect 103020 1006176 103026 1006188
rect 104802 1006176 104808 1006188
rect 103020 1006148 104808 1006176
rect 103020 1006136 103026 1006148
rect 104802 1006136 104808 1006148
rect 104860 1006136 104866 1006188
rect 106826 1006136 106832 1006188
rect 106884 1006176 106890 1006188
rect 113818 1006176 113824 1006188
rect 106884 1006148 113824 1006176
rect 106884 1006136 106890 1006148
rect 113818 1006136 113824 1006148
rect 113876 1006136 113882 1006188
rect 151786 1006176 151814 1006352
rect 153930 1006272 153936 1006324
rect 153988 1006312 153994 1006324
rect 158254 1006312 158260 1006324
rect 153988 1006284 158260 1006312
rect 153988 1006272 153994 1006284
rect 158254 1006272 158260 1006284
rect 158312 1006272 158318 1006324
rect 159450 1006272 159456 1006324
rect 159508 1006312 159514 1006324
rect 177298 1006312 177304 1006324
rect 159508 1006284 177304 1006312
rect 159508 1006272 159514 1006284
rect 177298 1006272 177304 1006284
rect 177356 1006272 177362 1006324
rect 249058 1006272 249064 1006324
rect 249116 1006312 249122 1006324
rect 254118 1006312 254124 1006324
rect 249116 1006284 254124 1006312
rect 249116 1006272 249122 1006284
rect 254118 1006272 254124 1006284
rect 254176 1006272 254182 1006324
rect 301498 1006272 301504 1006324
rect 301556 1006312 301562 1006324
rect 306926 1006312 306932 1006324
rect 301556 1006284 306932 1006312
rect 301556 1006272 301562 1006284
rect 306926 1006272 306932 1006284
rect 306984 1006272 306990 1006324
rect 314654 1006272 314660 1006324
rect 314712 1006312 314718 1006324
rect 319438 1006312 319444 1006324
rect 314712 1006284 319444 1006312
rect 314712 1006272 314718 1006284
rect 319438 1006272 319444 1006284
rect 319496 1006272 319502 1006324
rect 354858 1006272 354864 1006324
rect 354916 1006312 354922 1006324
rect 354916 1006284 367968 1006312
rect 354916 1006272 354922 1006284
rect 153746 1006176 153752 1006188
rect 151786 1006148 153752 1006176
rect 153746 1006136 153752 1006148
rect 153804 1006136 153810 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 164878 1006176 164884 1006188
rect 160336 1006148 164884 1006176
rect 160336 1006136 160342 1006148
rect 164878 1006136 164884 1006148
rect 164936 1006136 164942 1006188
rect 166258 1006136 166264 1006188
rect 166316 1006176 166322 1006188
rect 175918 1006176 175924 1006188
rect 166316 1006148 175924 1006176
rect 166316 1006136 166322 1006148
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 210418 1006136 210424 1006188
rect 210476 1006176 210482 1006188
rect 228358 1006176 228364 1006188
rect 210476 1006148 228364 1006176
rect 210476 1006136 210482 1006148
rect 228358 1006136 228364 1006148
rect 228416 1006136 228422 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 279418 1006176 279424 1006188
rect 262732 1006148 279424 1006176
rect 262732 1006136 262738 1006148
rect 279418 1006136 279424 1006148
rect 279476 1006136 279482 1006188
rect 298738 1006136 298744 1006188
rect 298796 1006176 298802 1006188
rect 304902 1006176 304908 1006188
rect 298796 1006148 304908 1006176
rect 298796 1006136 298802 1006148
rect 304902 1006136 304908 1006148
rect 304960 1006136 304966 1006188
rect 355686 1006136 355692 1006188
rect 355744 1006176 355750 1006188
rect 363598 1006176 363604 1006188
rect 355744 1006148 363604 1006176
rect 355744 1006136 355750 1006148
rect 363598 1006136 363604 1006148
rect 363656 1006136 363662 1006188
rect 365070 1006136 365076 1006188
rect 365128 1006176 365134 1006188
rect 367738 1006176 367744 1006188
rect 365128 1006148 367744 1006176
rect 365128 1006136 365134 1006148
rect 367738 1006136 367744 1006148
rect 367796 1006136 367802 1006188
rect 367940 1006176 367968 1006284
rect 369118 1006272 369124 1006324
rect 369176 1006312 369182 1006324
rect 380158 1006312 380164 1006324
rect 369176 1006284 380164 1006312
rect 369176 1006272 369182 1006284
rect 380158 1006272 380164 1006284
rect 380216 1006272 380222 1006324
rect 431678 1006312 431684 1006324
rect 412606 1006284 431684 1006312
rect 373258 1006176 373264 1006188
rect 367940 1006148 373264 1006176
rect 373258 1006136 373264 1006148
rect 373316 1006136 373322 1006188
rect 402238 1006136 402244 1006188
rect 402296 1006176 402302 1006188
rect 412606 1006176 412634 1006284
rect 431678 1006272 431684 1006284
rect 431736 1006272 431742 1006324
rect 431926 1006312 431954 1006420
rect 436738 1006408 436744 1006460
rect 436796 1006448 436802 1006460
rect 448514 1006448 448520 1006460
rect 436796 1006420 448520 1006448
rect 436796 1006408 436802 1006420
rect 448514 1006408 448520 1006420
rect 448572 1006408 448578 1006460
rect 513558 1006408 513564 1006460
rect 513616 1006448 513622 1006460
rect 519538 1006448 519544 1006460
rect 513616 1006420 519544 1006448
rect 513616 1006408 513622 1006420
rect 519538 1006408 519544 1006420
rect 519596 1006408 519602 1006460
rect 507854 1006340 507860 1006392
rect 507912 1006380 507918 1006392
rect 510522 1006380 510528 1006392
rect 507912 1006352 510528 1006380
rect 507912 1006340 507918 1006352
rect 510522 1006340 510528 1006352
rect 510580 1006340 510586 1006392
rect 555418 1006340 555424 1006392
rect 555476 1006380 555482 1006392
rect 558822 1006380 558828 1006392
rect 555476 1006352 558828 1006380
rect 555476 1006340 555482 1006352
rect 558822 1006340 558828 1006352
rect 558880 1006340 558886 1006392
rect 456794 1006312 456800 1006324
rect 431926 1006284 456800 1006312
rect 456794 1006272 456800 1006284
rect 456852 1006272 456858 1006324
rect 522298 1006312 522304 1006324
rect 514036 1006284 522304 1006312
rect 506198 1006204 506204 1006256
rect 506256 1006244 506262 1006256
rect 514036 1006244 514064 1006284
rect 522298 1006272 522304 1006284
rect 522356 1006272 522362 1006324
rect 571978 1006312 571984 1006324
rect 562336 1006284 571984 1006312
rect 506256 1006216 514064 1006244
rect 506256 1006204 506262 1006216
rect 553946 1006204 553952 1006256
rect 554004 1006244 554010 1006256
rect 562336 1006244 562364 1006284
rect 571978 1006272 571984 1006284
rect 572036 1006272 572042 1006324
rect 554004 1006216 562364 1006244
rect 554004 1006204 554010 1006216
rect 429194 1006176 429200 1006188
rect 402296 1006148 412634 1006176
rect 425348 1006148 429200 1006176
rect 402296 1006136 402302 1006148
rect 148870 1006068 148876 1006120
rect 148928 1006108 148934 1006120
rect 150066 1006108 150072 1006120
rect 148928 1006080 150072 1006108
rect 148928 1006068 148934 1006080
rect 150066 1006068 150072 1006080
rect 150124 1006068 150130 1006120
rect 93118 1006000 93124 1006052
rect 93176 1006040 93182 1006052
rect 96062 1006040 96068 1006052
rect 93176 1006012 96068 1006040
rect 93176 1006000 93182 1006012
rect 96062 1006000 96068 1006012
rect 96120 1006000 96126 1006052
rect 96246 1006000 96252 1006052
rect 96304 1006040 96310 1006052
rect 98270 1006040 98276 1006052
rect 96304 1006012 98276 1006040
rect 96304 1006000 96310 1006012
rect 98270 1006000 98276 1006012
rect 98328 1006000 98334 1006052
rect 101398 1006000 101404 1006052
rect 101456 1006040 101462 1006052
rect 103974 1006040 103980 1006052
rect 101456 1006012 103980 1006040
rect 101456 1006000 101462 1006012
rect 103974 1006000 103980 1006012
rect 104032 1006000 104038 1006052
rect 105998 1006000 106004 1006052
rect 106056 1006040 106062 1006052
rect 124858 1006040 124864 1006052
rect 106056 1006012 124864 1006040
rect 106056 1006000 106062 1006012
rect 124858 1006000 124864 1006012
rect 124916 1006000 124922 1006052
rect 158254 1006000 158260 1006052
rect 158312 1006040 158318 1006052
rect 171778 1006040 171784 1006052
rect 158312 1006012 171784 1006040
rect 158312 1006000 158318 1006012
rect 171778 1006000 171784 1006012
rect 171836 1006000 171842 1006052
rect 198182 1006000 198188 1006052
rect 198240 1006040 198246 1006052
rect 201034 1006040 201040 1006052
rect 198240 1006012 201040 1006040
rect 198240 1006000 198246 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 208394 1006000 208400 1006052
rect 208452 1006040 208458 1006052
rect 229738 1006040 229744 1006052
rect 208452 1006012 229744 1006040
rect 208452 1006000 208458 1006012
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 251082 1006000 251088 1006052
rect 251140 1006040 251146 1006052
rect 252462 1006040 252468 1006052
rect 251140 1006012 252468 1006040
rect 251140 1006000 251146 1006012
rect 252462 1006000 252468 1006012
rect 252520 1006000 252526 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 280798 1006040 280804 1006052
rect 261904 1006012 280804 1006040
rect 261904 1006000 261910 1006012
rect 280798 1006000 280804 1006012
rect 280856 1006000 280862 1006052
rect 298922 1006000 298928 1006052
rect 298980 1006040 298986 1006052
rect 311802 1006040 311808 1006052
rect 298980 1006012 311808 1006040
rect 298980 1006000 298986 1006012
rect 311802 1006000 311808 1006012
rect 311860 1006000 311866 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 320818 1006040 320824 1006052
rect 314712 1006012 320824 1006040
rect 314712 1006000 314718 1006012
rect 320818 1006000 320824 1006012
rect 320876 1006000 320882 1006052
rect 363414 1006000 363420 1006052
rect 363472 1006040 363478 1006052
rect 382918 1006040 382924 1006052
rect 363472 1006012 382924 1006040
rect 363472 1006000 363478 1006012
rect 382918 1006000 382924 1006012
rect 382976 1006000 382982 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 425348 1006040 425376 1006148
rect 429194 1006136 429200 1006148
rect 429252 1006136 429258 1006188
rect 434622 1006136 434628 1006188
rect 434680 1006176 434686 1006188
rect 471422 1006176 471428 1006188
rect 434680 1006148 471428 1006176
rect 434680 1006136 434686 1006148
rect 471422 1006136 471428 1006148
rect 471480 1006136 471486 1006188
rect 514202 1006136 514208 1006188
rect 514260 1006176 514266 1006188
rect 522482 1006176 522488 1006188
rect 514260 1006148 522488 1006176
rect 514260 1006136 514266 1006148
rect 522482 1006136 522488 1006148
rect 522540 1006136 522546 1006188
rect 562502 1006136 562508 1006188
rect 562560 1006176 562566 1006188
rect 570598 1006176 570604 1006188
rect 562560 1006148 570604 1006176
rect 562560 1006136 562566 1006148
rect 570598 1006136 570604 1006148
rect 570656 1006136 570662 1006188
rect 400916 1006012 425376 1006040
rect 400916 1006000 400922 1006012
rect 425514 1006000 425520 1006052
rect 425572 1006040 425578 1006052
rect 429194 1006040 429200 1006052
rect 425572 1006012 429200 1006040
rect 425572 1006000 425578 1006012
rect 429194 1006000 429200 1006012
rect 429252 1006000 429258 1006052
rect 430022 1006000 430028 1006052
rect 430080 1006040 430086 1006052
rect 471238 1006040 471244 1006052
rect 430080 1006012 471244 1006040
rect 430080 1006000 430086 1006012
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 496722 1006000 496728 1006052
rect 496780 1006040 496786 1006052
rect 498838 1006040 498844 1006052
rect 496780 1006012 498844 1006040
rect 496780 1006000 496786 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 500494 1006000 500500 1006052
rect 500552 1006040 500558 1006052
rect 513558 1006040 513564 1006052
rect 500552 1006012 513564 1006040
rect 500552 1006000 500558 1006012
rect 513558 1006000 513564 1006012
rect 513616 1006000 513622 1006052
rect 554314 1006000 554320 1006052
rect 554372 1006040 554378 1006052
rect 574738 1006040 574744 1006052
rect 554372 1006012 574744 1006040
rect 554372 1006000 554378 1006012
rect 574738 1006000 574744 1006012
rect 574796 1006000 574802 1006052
rect 509050 1005864 509056 1005916
rect 509108 1005904 509114 1005916
rect 514018 1005904 514024 1005916
rect 509108 1005876 514024 1005904
rect 509108 1005864 509114 1005876
rect 514018 1005864 514024 1005876
rect 514076 1005864 514082 1005916
rect 564434 1005864 564440 1005916
rect 564492 1005904 564498 1005916
rect 567838 1005904 567844 1005916
rect 564492 1005876 567844 1005904
rect 564492 1005864 564498 1005876
rect 567838 1005864 567844 1005876
rect 567896 1005864 567902 1005916
rect 427538 1005660 427544 1005712
rect 427596 1005700 427602 1005712
rect 440878 1005700 440884 1005712
rect 427596 1005672 440884 1005700
rect 427596 1005660 427602 1005672
rect 440878 1005660 440884 1005672
rect 440936 1005660 440942 1005712
rect 428366 1005524 428372 1005576
rect 428424 1005564 428430 1005576
rect 446398 1005564 446404 1005576
rect 428424 1005536 446404 1005564
rect 428424 1005524 428430 1005536
rect 446398 1005524 446404 1005536
rect 446456 1005524 446462 1005576
rect 360562 1005388 360568 1005440
rect 360620 1005428 360626 1005440
rect 378778 1005428 378784 1005440
rect 360620 1005400 378784 1005428
rect 360620 1005388 360626 1005400
rect 378778 1005388 378784 1005400
rect 378836 1005388 378842 1005440
rect 423490 1005388 423496 1005440
rect 423548 1005428 423554 1005440
rect 464338 1005428 464344 1005440
rect 423548 1005400 464344 1005428
rect 423548 1005388 423554 1005400
rect 464338 1005388 464344 1005400
rect 464396 1005388 464402 1005440
rect 555970 1005388 555976 1005440
rect 556028 1005428 556034 1005440
rect 573358 1005428 573364 1005440
rect 556028 1005400 573364 1005428
rect 556028 1005388 556034 1005400
rect 573358 1005388 573364 1005400
rect 573416 1005388 573422 1005440
rect 102778 1005252 102784 1005304
rect 102836 1005292 102842 1005304
rect 108850 1005292 108856 1005304
rect 102836 1005264 108856 1005292
rect 102836 1005252 102842 1005264
rect 108850 1005252 108856 1005264
rect 108908 1005252 108914 1005304
rect 204898 1005252 204904 1005304
rect 204956 1005292 204962 1005304
rect 212074 1005292 212080 1005304
rect 204956 1005264 212080 1005292
rect 204956 1005252 204962 1005264
rect 212074 1005252 212080 1005264
rect 212132 1005252 212138 1005304
rect 357710 1005252 357716 1005304
rect 357768 1005292 357774 1005304
rect 375374 1005292 375380 1005304
rect 357768 1005264 375380 1005292
rect 357768 1005252 357774 1005264
rect 375374 1005252 375380 1005264
rect 375432 1005252 375438 1005304
rect 424318 1005252 424324 1005304
rect 424376 1005292 424382 1005304
rect 465718 1005292 465724 1005304
rect 424376 1005264 465724 1005292
rect 424376 1005252 424382 1005264
rect 465718 1005252 465724 1005264
rect 465776 1005252 465782 1005304
rect 498838 1005252 498844 1005304
rect 498896 1005292 498902 1005304
rect 516778 1005292 516784 1005304
rect 498896 1005264 516784 1005292
rect 498896 1005252 498902 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 149698 1005048 149704 1005100
rect 149756 1005088 149762 1005100
rect 152918 1005088 152924 1005100
rect 149756 1005060 152924 1005088
rect 149756 1005048 149762 1005060
rect 152918 1005048 152924 1005060
rect 152976 1005048 152982 1005100
rect 354582 1005048 354588 1005100
rect 354640 1005088 354646 1005100
rect 356514 1005088 356520 1005100
rect 354640 1005060 356520 1005088
rect 354640 1005048 354646 1005060
rect 356514 1005048 356520 1005060
rect 356572 1005048 356578 1005100
rect 365070 1005048 365076 1005100
rect 365128 1005088 365134 1005100
rect 370498 1005088 370504 1005100
rect 365128 1005060 370504 1005088
rect 365128 1005048 365134 1005060
rect 370498 1005048 370504 1005060
rect 370556 1005048 370562 1005100
rect 551462 1005048 551468 1005100
rect 551520 1005088 551526 1005100
rect 569218 1005088 569224 1005100
rect 551520 1005060 569224 1005088
rect 551520 1005048 551526 1005060
rect 569218 1005048 569224 1005060
rect 569276 1005048 569282 1005100
rect 151078 1004912 151084 1004964
rect 151136 1004952 151142 1004964
rect 153746 1004952 153752 1004964
rect 151136 1004924 153752 1004952
rect 151136 1004912 151142 1004924
rect 153746 1004912 153752 1004924
rect 153804 1004912 153810 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 263042 1004912 263048 1004964
rect 263100 1004952 263106 1004964
rect 268378 1004952 268384 1004964
rect 263100 1004924 268384 1004952
rect 263100 1004912 263106 1004924
rect 268378 1004912 268384 1004924
rect 268436 1004912 268442 1004964
rect 353202 1004912 353208 1004964
rect 353260 1004952 353266 1004964
rect 355686 1004952 355692 1004964
rect 353260 1004924 355692 1004952
rect 353260 1004912 353266 1004924
rect 355686 1004912 355692 1004924
rect 355744 1004912 355750 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 364978 1004952 364984 1004964
rect 361448 1004924 364984 1004952
rect 361448 1004912 361454 1004924
rect 364978 1004912 364984 1004924
rect 365036 1004912 365042 1004964
rect 422018 1004912 422024 1004964
rect 422076 1004952 422082 1004964
rect 423490 1004952 423496 1004964
rect 422076 1004924 423496 1004952
rect 422076 1004912 422082 1004924
rect 423490 1004912 423496 1004924
rect 423548 1004912 423554 1004964
rect 433978 1004952 433984 1004964
rect 431926 1004924 433984 1004952
rect 149882 1004776 149888 1004828
rect 149940 1004816 149946 1004828
rect 152918 1004816 152924 1004828
rect 149940 1004788 152924 1004816
rect 149940 1004776 149946 1004788
rect 152918 1004776 152924 1004788
rect 152976 1004776 152982 1004828
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 211246 1004776 211252 1004828
rect 211304 1004816 211310 1004828
rect 215938 1004816 215944 1004828
rect 211304 1004788 215944 1004816
rect 211304 1004776 211310 1004788
rect 215938 1004776 215944 1004788
rect 215996 1004776 216002 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365162 1004816 365168 1004828
rect 362644 1004788 365168 1004816
rect 362644 1004776 362650 1004788
rect 365162 1004776 365168 1004788
rect 365220 1004776 365226 1004828
rect 420822 1004776 420828 1004828
rect 420880 1004816 420886 1004828
rect 422662 1004816 422668 1004828
rect 420880 1004788 422668 1004816
rect 420880 1004776 420886 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 430850 1004776 430856 1004828
rect 430908 1004816 430914 1004828
rect 431926 1004816 431954 1004924
rect 433978 1004912 433984 1004924
rect 434036 1004912 434042 1004964
rect 498102 1004912 498108 1004964
rect 498160 1004952 498166 1004964
rect 499666 1004952 499672 1004964
rect 498160 1004924 499672 1004952
rect 498160 1004912 498166 1004924
rect 499666 1004912 499672 1004924
rect 499724 1004912 499730 1004964
rect 508222 1004912 508228 1004964
rect 508280 1004952 508286 1004964
rect 511258 1004952 511264 1004964
rect 508280 1004924 511264 1004952
rect 508280 1004912 508286 1004924
rect 511258 1004912 511264 1004924
rect 511316 1004912 511322 1004964
rect 560846 1004912 560852 1004964
rect 560904 1004952 560910 1004964
rect 566458 1004952 566464 1004964
rect 560904 1004924 566464 1004952
rect 560904 1004912 560910 1004924
rect 566458 1004912 566464 1004924
rect 566516 1004912 566522 1004964
rect 430908 1004788 431954 1004816
rect 430908 1004776 430914 1004788
rect 432046 1004776 432052 1004828
rect 432104 1004816 432110 1004828
rect 436738 1004816 436744 1004828
rect 432104 1004788 436744 1004816
rect 432104 1004776 432110 1004788
rect 436738 1004776 436744 1004788
rect 436796 1004776 436802 1004828
rect 499298 1004776 499304 1004828
rect 499356 1004816 499362 1004828
rect 501322 1004816 501328 1004828
rect 499356 1004788 501328 1004816
rect 499356 1004776 499362 1004788
rect 501322 1004776 501328 1004788
rect 501380 1004776 501386 1004828
rect 507026 1004776 507032 1004828
rect 507084 1004816 507090 1004828
rect 509878 1004816 509884 1004828
rect 507084 1004788 509884 1004816
rect 507084 1004776 507090 1004788
rect 509878 1004776 509884 1004788
rect 509936 1004776 509942 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 151262 1004640 151268 1004692
rect 151320 1004680 151326 1004692
rect 154114 1004680 154120 1004692
rect 151320 1004652 154120 1004680
rect 151320 1004640 151326 1004652
rect 154114 1004640 154120 1004652
rect 154172 1004640 154178 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 430022 1004640 430028 1004692
rect 430080 1004680 430086 1004692
rect 431954 1004680 431960 1004692
rect 430080 1004652 431960 1004680
rect 430080 1004640 430086 1004652
rect 431954 1004640 431960 1004652
rect 432012 1004640 432018 1004692
rect 432874 1004640 432880 1004692
rect 432932 1004680 432938 1004692
rect 438118 1004680 438124 1004692
rect 432932 1004652 438124 1004680
rect 432932 1004640 432938 1004652
rect 438118 1004640 438124 1004652
rect 438176 1004640 438182 1004692
rect 503346 1004640 503352 1004692
rect 503404 1004680 503410 1004692
rect 507302 1004680 507308 1004692
rect 503404 1004652 507308 1004680
rect 503404 1004640 503410 1004652
rect 507302 1004640 507308 1004652
rect 507360 1004640 507366 1004692
rect 508222 1004640 508228 1004692
rect 508280 1004680 508286 1004692
rect 510614 1004680 510620 1004692
rect 508280 1004652 510620 1004680
rect 508280 1004640 508286 1004652
rect 510614 1004640 510620 1004652
rect 510672 1004640 510678 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559466 1004680 559472 1004692
rect 557684 1004652 559472 1004680
rect 557684 1004640 557690 1004652
rect 559466 1004640 559472 1004652
rect 559524 1004640 559530 1004692
rect 560846 1004640 560852 1004692
rect 560904 1004680 560910 1004692
rect 565078 1004680 565084 1004692
rect 560904 1004652 565084 1004680
rect 560904 1004640 560910 1004652
rect 565078 1004640 565084 1004652
rect 565136 1004640 565142 1004692
rect 422202 1004572 422208 1004624
rect 422260 1004612 422266 1004624
rect 424318 1004612 424324 1004624
rect 422260 1004584 424324 1004612
rect 422260 1004572 422266 1004584
rect 424318 1004572 424324 1004584
rect 424376 1004572 424382 1004624
rect 499482 1004572 499488 1004624
rect 499540 1004612 499546 1004624
rect 500494 1004612 500500 1004624
rect 499540 1004584 500500 1004612
rect 499540 1004572 499546 1004584
rect 500494 1004572 500500 1004584
rect 500552 1004572 500558 1004624
rect 510062 1004504 510068 1004556
rect 510120 1004544 510126 1004556
rect 515398 1004544 515404 1004556
rect 510120 1004516 515404 1004544
rect 510120 1004504 510126 1004516
rect 515398 1004504 515404 1004516
rect 515456 1004504 515462 1004556
rect 425514 1004164 425520 1004216
rect 425572 1004204 425578 1004216
rect 449158 1004204 449164 1004216
rect 425572 1004176 449164 1004204
rect 425572 1004164 425578 1004176
rect 449158 1004164 449164 1004176
rect 449216 1004164 449222 1004216
rect 451826 1004164 451832 1004216
rect 451884 1004204 451890 1004216
rect 467558 1004204 467564 1004216
rect 451884 1004176 467564 1004204
rect 451884 1004164 451890 1004176
rect 467558 1004164 467564 1004176
rect 467616 1004164 467622 1004216
rect 425146 1004028 425152 1004080
rect 425204 1004068 425210 1004080
rect 454862 1004068 454868 1004080
rect 425204 1004040 454868 1004068
rect 425204 1004028 425210 1004040
rect 454862 1004028 454868 1004040
rect 454920 1004028 454926 1004080
rect 456794 1004028 456800 1004080
rect 456852 1004068 456858 1004080
rect 456852 1004040 460934 1004068
rect 456852 1004028 456858 1004040
rect 422202 1003892 422208 1003944
rect 422260 1003932 422266 1003944
rect 458818 1003932 458824 1003944
rect 422260 1003904 458824 1003932
rect 422260 1003892 422266 1003904
rect 458818 1003892 458824 1003904
rect 458876 1003892 458882 1003944
rect 460906 1003932 460934 1004040
rect 502518 1004028 502524 1004080
rect 502576 1004068 502582 1004080
rect 514662 1004068 514668 1004080
rect 502576 1004040 514668 1004068
rect 502576 1004028 502582 1004040
rect 514662 1004028 514668 1004040
rect 514720 1004028 514726 1004080
rect 461578 1003932 461584 1003944
rect 460906 1003904 461584 1003932
rect 461578 1003892 461584 1003904
rect 461636 1003892 461642 1003944
rect 499482 1003892 499488 1003944
rect 499540 1003932 499546 1003944
rect 518342 1003932 518348 1003944
rect 499540 1003904 518348 1003932
rect 499540 1003892 499546 1003904
rect 518342 1003892 518348 1003904
rect 518400 1003892 518406 1003944
rect 422018 1003484 422024 1003536
rect 422076 1003524 422082 1003536
rect 423766 1003524 423772 1003536
rect 422076 1003496 423772 1003524
rect 422076 1003484 422082 1003496
rect 423766 1003484 423772 1003496
rect 423824 1003484 423830 1003536
rect 448514 1003280 448520 1003332
rect 448572 1003320 448578 1003332
rect 451642 1003320 451648 1003332
rect 448572 1003292 451648 1003320
rect 448572 1003280 448578 1003292
rect 451642 1003280 451648 1003292
rect 451700 1003280 451706 1003332
rect 97442 1002736 97448 1002788
rect 97500 1002776 97506 1002788
rect 102318 1002776 102324 1002788
rect 97500 1002748 102324 1002776
rect 97500 1002736 97506 1002748
rect 102318 1002736 102324 1002748
rect 102376 1002736 102382 1002788
rect 94498 1002600 94504 1002652
rect 94556 1002640 94562 1002652
rect 100294 1002640 100300 1002652
rect 94556 1002612 100300 1002640
rect 94556 1002600 94562 1002612
rect 100294 1002600 100300 1002612
rect 100352 1002600 100358 1002652
rect 253474 1002600 253480 1002652
rect 253532 1002640 253538 1002652
rect 256142 1002640 256148 1002652
rect 253532 1002612 256148 1002640
rect 253532 1002600 253538 1002612
rect 256142 1002600 256148 1002612
rect 256200 1002600 256206 1002652
rect 100018 1002464 100024 1002516
rect 100076 1002504 100082 1002516
rect 103146 1002504 103152 1002516
rect 100076 1002476 103152 1002504
rect 100076 1002464 100082 1002476
rect 103146 1002464 103152 1002476
rect 103204 1002464 103210 1002516
rect 252002 1002464 252008 1002516
rect 252060 1002504 252066 1002516
rect 255314 1002504 255320 1002516
rect 252060 1002476 255320 1002504
rect 252060 1002464 252066 1002476
rect 255314 1002464 255320 1002476
rect 255372 1002464 255378 1002516
rect 261018 1002464 261024 1002516
rect 261076 1002504 261082 1002516
rect 264238 1002504 264244 1002516
rect 261076 1002476 264244 1002504
rect 261076 1002464 261082 1002476
rect 264238 1002464 264244 1002476
rect 264296 1002464 264302 1002516
rect 557994 1002464 558000 1002516
rect 558052 1002504 558058 1002516
rect 560938 1002504 560944 1002516
rect 558052 1002476 560944 1002504
rect 558052 1002464 558058 1002476
rect 560938 1002464 560944 1002476
rect 560996 1002464 561002 1002516
rect 555142 1002396 555148 1002448
rect 555200 1002436 555206 1002448
rect 557534 1002436 557540 1002448
rect 555200 1002408 557540 1002436
rect 555200 1002396 555206 1002408
rect 557534 1002396 557540 1002408
rect 557592 1002396 557598 1002448
rect 97258 1002328 97264 1002380
rect 97316 1002368 97322 1002380
rect 100294 1002368 100300 1002380
rect 97316 1002340 100300 1002368
rect 97316 1002328 97322 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 107654 1002328 107660 1002380
rect 107712 1002368 107718 1002380
rect 109494 1002368 109500 1002380
rect 107712 1002340 109500 1002368
rect 107712 1002328 107718 1002340
rect 109494 1002328 109500 1002340
rect 109552 1002328 109558 1002380
rect 253014 1002328 253020 1002380
rect 253072 1002368 253078 1002380
rect 256142 1002368 256148 1002380
rect 253072 1002340 256148 1002368
rect 253072 1002328 253078 1002340
rect 256142 1002328 256148 1002340
rect 256200 1002328 256206 1002380
rect 558822 1002328 558828 1002380
rect 558880 1002368 558886 1002380
rect 562502 1002368 562508 1002380
rect 558880 1002340 562508 1002368
rect 558880 1002328 558886 1002340
rect 562502 1002328 562508 1002340
rect 562560 1002328 562566 1002380
rect 98638 1002192 98644 1002244
rect 98696 1002232 98702 1002244
rect 101950 1002232 101956 1002244
rect 98696 1002204 101956 1002232
rect 98696 1002192 98702 1002204
rect 101950 1002192 101956 1002204
rect 102008 1002192 102014 1002244
rect 105630 1002192 105636 1002244
rect 105688 1002232 105694 1002244
rect 107838 1002232 107844 1002244
rect 105688 1002204 107844 1002232
rect 105688 1002192 105694 1002204
rect 107838 1002192 107844 1002204
rect 107896 1002192 107902 1002244
rect 108022 1002192 108028 1002244
rect 108080 1002232 108086 1002244
rect 110414 1002232 110420 1002244
rect 108080 1002204 110420 1002232
rect 108080 1002192 108086 1002204
rect 110414 1002192 110420 1002204
rect 110472 1002192 110478 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 158714 1002232 158720 1002244
rect 155828 1002204 158720 1002232
rect 155828 1002192 155834 1002204
rect 158714 1002192 158720 1002204
rect 158772 1002192 158778 1002244
rect 203518 1002192 203524 1002244
rect 203576 1002232 203582 1002244
rect 206370 1002232 206376 1002244
rect 203576 1002204 206376 1002232
rect 203576 1002192 203582 1002204
rect 206370 1002192 206376 1002204
rect 206428 1002192 206434 1002244
rect 206738 1002192 206744 1002244
rect 206796 1002232 206802 1002244
rect 208394 1002232 208400 1002244
rect 206796 1002204 208400 1002232
rect 206796 1002192 206802 1002204
rect 208394 1002192 208400 1002204
rect 208452 1002192 208458 1002244
rect 210878 1002192 210884 1002244
rect 210936 1002232 210942 1002244
rect 213178 1002232 213184 1002244
rect 210936 1002204 213184 1002232
rect 210936 1002192 210942 1002204
rect 213178 1002192 213184 1002204
rect 213236 1002192 213242 1002244
rect 251818 1002192 251824 1002244
rect 251876 1002232 251882 1002244
rect 254486 1002232 254492 1002244
rect 251876 1002204 254492 1002232
rect 251876 1002192 251882 1002204
rect 254486 1002192 254492 1002204
rect 254544 1002192 254550 1002244
rect 358538 1002192 358544 1002244
rect 358596 1002232 358602 1002244
rect 360838 1002232 360844 1002244
rect 358596 1002204 360844 1002232
rect 358596 1002192 358602 1002204
rect 360838 1002192 360844 1002204
rect 360896 1002192 360902 1002244
rect 423582 1002192 423588 1002244
rect 423640 1002232 423646 1002244
rect 426342 1002232 426348 1002244
rect 423640 1002204 426348 1002232
rect 423640 1002192 423646 1002204
rect 426342 1002192 426348 1002204
rect 426400 1002192 426406 1002244
rect 501690 1002192 501696 1002244
rect 501748 1002232 501754 1002244
rect 504358 1002232 504364 1002244
rect 501748 1002204 504364 1002232
rect 501748 1002192 501754 1002204
rect 504358 1002192 504364 1002204
rect 504416 1002192 504422 1002244
rect 551922 1002192 551928 1002244
rect 551980 1002232 551986 1002244
rect 554314 1002232 554320 1002244
rect 551980 1002204 554320 1002232
rect 551980 1002192 551986 1002204
rect 554314 1002192 554320 1002204
rect 554372 1002192 554378 1002244
rect 557994 1002192 558000 1002244
rect 558052 1002232 558058 1002244
rect 560294 1002232 560300 1002244
rect 558052 1002204 560300 1002232
rect 558052 1002192 558058 1002204
rect 560294 1002192 560300 1002204
rect 560352 1002192 560358 1002244
rect 560478 1002192 560484 1002244
rect 560536 1002232 560542 1002244
rect 563054 1002232 563060 1002244
rect 560536 1002204 563060 1002232
rect 560536 1002192 560542 1002204
rect 563054 1002192 563060 1002204
rect 563112 1002192 563118 1002244
rect 96062 1002056 96068 1002108
rect 96120 1002096 96126 1002108
rect 99098 1002096 99104 1002108
rect 96120 1002068 99104 1002096
rect 96120 1002056 96126 1002068
rect 99098 1002056 99104 1002068
rect 99156 1002056 99162 1002108
rect 100202 1002056 100208 1002108
rect 100260 1002096 100266 1002108
rect 103146 1002096 103152 1002108
rect 100260 1002068 103152 1002096
rect 100260 1002056 100266 1002068
rect 103146 1002056 103152 1002068
rect 103204 1002056 103210 1002108
rect 103974 1002056 103980 1002108
rect 104032 1002096 104038 1002108
rect 106458 1002096 106464 1002108
rect 104032 1002068 106464 1002096
rect 104032 1002056 104038 1002068
rect 106458 1002056 106464 1002068
rect 106516 1002056 106522 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111794 1002096 111800 1002108
rect 109736 1002068 111800 1002096
rect 109736 1002056 109742 1002068
rect 111794 1002056 111800 1002068
rect 111852 1002056 111858 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 152458 1002056 152464 1002108
rect 152516 1002096 152522 1002108
rect 154574 1002096 154580 1002108
rect 152516 1002068 154580 1002096
rect 152516 1002056 152522 1002068
rect 154574 1002056 154580 1002068
rect 154632 1002056 154638 1002108
rect 205082 1002056 205088 1002108
rect 205140 1002096 205146 1002108
rect 207198 1002096 207204 1002108
rect 205140 1002068 207204 1002096
rect 205140 1002056 205146 1002068
rect 207198 1002056 207204 1002068
rect 207256 1002056 207262 1002108
rect 212534 1002056 212540 1002108
rect 212592 1002096 212598 1002108
rect 214558 1002096 214564 1002108
rect 212592 1002068 214564 1002096
rect 212592 1002056 212598 1002068
rect 214558 1002056 214564 1002068
rect 214616 1002056 214622 1002108
rect 263502 1002056 263508 1002108
rect 263560 1002096 263566 1002108
rect 265618 1002096 265624 1002108
rect 263560 1002068 265624 1002096
rect 263560 1002056 263566 1002068
rect 265618 1002056 265624 1002068
rect 265676 1002056 265682 1002108
rect 300302 1002056 300308 1002108
rect 300360 1002096 300366 1002108
rect 305270 1002096 305276 1002108
rect 300360 1002068 305276 1002096
rect 300360 1002056 300366 1002068
rect 305270 1002056 305276 1002068
rect 305328 1002056 305334 1002108
rect 310146 1002056 310152 1002108
rect 310204 1002096 310210 1002108
rect 311894 1002096 311900 1002108
rect 310204 1002068 311900 1002096
rect 310204 1002056 310210 1002068
rect 311894 1002056 311900 1002068
rect 311952 1002056 311958 1002108
rect 355778 1002056 355784 1002108
rect 355836 1002096 355842 1002108
rect 356514 1002096 356520 1002108
rect 355836 1002068 356520 1002096
rect 355836 1002056 355842 1002068
rect 356514 1002056 356520 1002068
rect 356572 1002056 356578 1002108
rect 504542 1002056 504548 1002108
rect 504600 1002096 504606 1002108
rect 507118 1002096 507124 1002108
rect 504600 1002068 507124 1002096
rect 504600 1002056 504606 1002068
rect 507118 1002056 507124 1002068
rect 507176 1002056 507182 1002108
rect 559650 1002056 559656 1002108
rect 559708 1002096 559714 1002108
rect 561490 1002096 561496 1002108
rect 559708 1002068 561496 1002096
rect 559708 1002056 559714 1002068
rect 561490 1002056 561496 1002068
rect 561548 1002056 561554 1002108
rect 561674 1002056 561680 1002108
rect 561732 1002096 561738 1002108
rect 563698 1002096 563704 1002108
rect 561732 1002068 563704 1002096
rect 561732 1002056 561738 1002068
rect 563698 1002056 563704 1002068
rect 563756 1002056 563762 1002108
rect 95878 1001920 95884 1001972
rect 95936 1001960 95942 1001972
rect 98270 1001960 98276 1001972
rect 95936 1001932 98276 1001960
rect 95936 1001920 95942 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 98822 1001920 98828 1001972
rect 98880 1001960 98886 1001972
rect 101122 1001960 101128 1001972
rect 98880 1001932 101128 1001960
rect 98880 1001920 98886 1001932
rect 101122 1001920 101128 1001932
rect 101180 1001920 101186 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 107746 1001960 107752 1001972
rect 106056 1001932 107752 1001960
rect 106056 1001920 106062 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 155770 1001920 155776 1001972
rect 155828 1001960 155834 1001972
rect 157334 1001960 157340 1001972
rect 155828 1001932 157340 1001960
rect 155828 1001920 155834 1001932
rect 157334 1001920 157340 1001932
rect 157392 1001920 157398 1001972
rect 157794 1001920 157800 1001972
rect 157852 1001960 157858 1001972
rect 160094 1001960 160100 1001972
rect 157852 1001932 160100 1001960
rect 157852 1001920 157858 1001932
rect 160094 1001920 160100 1001932
rect 160152 1001920 160158 1001972
rect 202966 1001920 202972 1001972
rect 203024 1001960 203030 1001972
rect 205542 1001960 205548 1001972
rect 203024 1001932 205548 1001960
rect 203024 1001920 203030 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 210878 1001920 210884 1001972
rect 210936 1001960 210942 1001972
rect 212534 1001960 212540 1001972
rect 210936 1001932 212540 1001960
rect 210936 1001920 210942 1001932
rect 212534 1001920 212540 1001932
rect 212592 1001920 212598 1001972
rect 261018 1001920 261024 1001972
rect 261076 1001960 261082 1001972
rect 263594 1001960 263600 1001972
rect 261076 1001932 263600 1001960
rect 261076 1001920 261082 1001932
rect 263594 1001920 263600 1001932
rect 263652 1001920 263658 1001972
rect 263870 1001920 263876 1001972
rect 263928 1001960 263934 1001972
rect 266998 1001960 267004 1001972
rect 263928 1001932 267004 1001960
rect 263928 1001920 263934 1001932
rect 266998 1001920 267004 1001932
rect 267056 1001920 267062 1001972
rect 310974 1001920 310980 1001972
rect 311032 1001960 311038 1001972
rect 313274 1001960 313280 1001972
rect 311032 1001932 313280 1001960
rect 311032 1001920 311038 1001932
rect 313274 1001920 313280 1001932
rect 313332 1001920 313338 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 360194 1001920 360200 1001972
rect 360252 1001960 360258 1001972
rect 362218 1001960 362224 1001972
rect 360252 1001932 362224 1001960
rect 360252 1001920 360258 1001932
rect 362218 1001920 362224 1001932
rect 362276 1001920 362282 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 425698 1001920 425704 1001972
rect 425756 1001960 425762 1001972
rect 427170 1001960 427176 1001972
rect 425756 1001932 427176 1001960
rect 425756 1001920 425762 1001932
rect 427170 1001920 427176 1001932
rect 427228 1001920 427234 1001972
rect 433334 1001920 433340 1001972
rect 433392 1001960 433398 1001972
rect 435358 1001960 435364 1001972
rect 433392 1001932 435364 1001960
rect 433392 1001920 433398 1001932
rect 435358 1001920 435364 1001932
rect 435416 1001920 435422 1001972
rect 500862 1001920 500868 1001972
rect 500920 1001960 500926 1001972
rect 501690 1001960 501696 1001972
rect 500920 1001932 501696 1001960
rect 500920 1001920 500926 1001932
rect 501690 1001920 501696 1001932
rect 501748 1001920 501754 1001972
rect 501874 1001920 501880 1001972
rect 501932 1001960 501938 1001972
rect 503346 1001960 503352 1001972
rect 501932 1001932 503352 1001960
rect 501932 1001920 501938 1001932
rect 503346 1001920 503352 1001932
rect 503404 1001920 503410 1001972
rect 504174 1001920 504180 1001972
rect 504232 1001960 504238 1001972
rect 505738 1001960 505744 1001972
rect 504232 1001932 505744 1001960
rect 504232 1001920 504238 1001932
rect 505738 1001920 505744 1001932
rect 505796 1001920 505802 1001972
rect 510338 1001920 510344 1001972
rect 510396 1001960 510402 1001972
rect 512638 1001960 512644 1001972
rect 510396 1001932 512644 1001960
rect 510396 1001920 510402 1001932
rect 512638 1001920 512644 1001932
rect 512696 1001920 512702 1001972
rect 560018 1001920 560024 1001972
rect 560076 1001960 560082 1001972
rect 562318 1001960 562324 1001972
rect 560076 1001932 562324 1001960
rect 560076 1001920 560082 1001932
rect 562318 1001920 562324 1001932
rect 562376 1001920 562382 1001972
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 423766 1001172 423772 1001224
rect 423824 1001212 423830 1001224
rect 456794 1001212 456800 1001224
rect 423824 1001184 456800 1001212
rect 423824 1001172 423830 1001184
rect 456794 1001172 456800 1001184
rect 456852 1001172 456858 1001224
rect 498102 1001172 498108 1001224
rect 498160 1001212 498166 1001224
rect 520366 1001212 520372 1001224
rect 498160 1001184 520372 1001212
rect 498160 1001172 498166 1001184
rect 520366 1001172 520372 1001184
rect 520424 1001172 520430 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 423582 1000900 423588 1000952
rect 423640 1000940 423646 1000952
rect 429378 1000940 429384 1000952
rect 423640 1000912 429384 1000940
rect 423640 1000900 423646 1000912
rect 429378 1000900 429384 1000912
rect 429436 1000900 429442 1000952
rect 298094 1000492 298100 1000544
rect 298152 1000532 298158 1000544
rect 308950 1000532 308956 1000544
rect 298152 1000504 308956 1000532
rect 298152 1000492 298158 1000504
rect 308950 1000492 308956 1000504
rect 309008 1000492 309014 1000544
rect 375374 1000492 375380 1000544
rect 375432 1000532 375438 1000544
rect 383286 1000532 383292 1000544
rect 375432 1000504 383292 1000532
rect 375432 1000492 375438 1000504
rect 383286 1000492 383292 1000504
rect 383344 1000492 383350 1000544
rect 92750 999744 92756 999796
rect 92808 999784 92814 999796
rect 102962 999784 102968 999796
rect 92808 999756 102968 999784
rect 92808 999744 92814 999756
rect 102962 999744 102968 999756
rect 103020 999744 103026 999796
rect 360838 999744 360844 999796
rect 360896 999784 360902 999796
rect 369854 999784 369860 999796
rect 360896 999756 369860 999784
rect 360896 999744 360902 999756
rect 369854 999744 369860 999756
rect 369912 999744 369918 999796
rect 373258 999064 373264 999116
rect 373316 999104 373322 999116
rect 374638 999104 374644 999116
rect 373316 999076 374644 999104
rect 373316 999064 373322 999076
rect 374638 999064 374644 999076
rect 374696 999064 374702 999116
rect 565262 999064 565268 999116
rect 565320 999104 565326 999116
rect 568206 999104 568212 999116
rect 565320 999076 568212 999104
rect 565320 999064 565326 999076
rect 568206 999064 568212 999076
rect 568264 999064 568270 999116
rect 196618 998996 196624 999048
rect 196676 999036 196682 999048
rect 204346 999036 204352 999048
rect 196676 999008 204352 999036
rect 196676 998996 196682 999008
rect 204346 998996 204352 999008
rect 204404 998996 204410 999048
rect 467558 998860 467564 998912
rect 467616 998900 467622 998912
rect 472618 998900 472624 998912
rect 467616 998872 472624 998900
rect 467616 998860 467622 998872
rect 472618 998860 472624 998872
rect 472676 998860 472682 998912
rect 200758 998724 200764 998776
rect 200816 998764 200822 998776
rect 203886 998764 203892 998776
rect 200816 998736 203892 998764
rect 200816 998724 200822 998736
rect 203886 998724 203892 998736
rect 203944 998724 203950 998776
rect 378778 998724 378784 998776
rect 378836 998764 378842 998776
rect 383562 998764 383568 998776
rect 378836 998736 383568 998764
rect 378836 998724 378842 998736
rect 383562 998724 383568 998736
rect 383620 998724 383626 998776
rect 426526 998656 426532 998708
rect 426584 998696 426590 998708
rect 466454 998696 466460 998708
rect 426584 998668 466460 998696
rect 426584 998656 426590 998668
rect 466454 998656 466460 998668
rect 466512 998656 466518 998708
rect 515582 998656 515588 998708
rect 515640 998696 515646 998708
rect 523862 998696 523868 998708
rect 515640 998668 523868 998696
rect 515640 998656 515646 998668
rect 523862 998656 523868 998668
rect 523920 998656 523926 998708
rect 197814 998588 197820 998640
rect 197872 998628 197878 998640
rect 202690 998628 202696 998640
rect 197872 998600 202696 998628
rect 197872 998588 197878 998600
rect 202690 998588 202696 998600
rect 202748 998588 202754 998640
rect 376754 998588 376760 998640
rect 376812 998628 376818 998640
rect 383470 998628 383476 998640
rect 376812 998600 383476 998628
rect 376812 998588 376818 998600
rect 383470 998588 383476 998600
rect 383528 998588 383534 998640
rect 247218 998520 247224 998572
rect 247276 998560 247282 998572
rect 256970 998560 256976 998572
rect 247276 998532 256976 998560
rect 247276 998520 247282 998532
rect 256970 998520 256976 998532
rect 257028 998520 257034 998572
rect 429378 998520 429384 998572
rect 429436 998560 429442 998572
rect 472434 998560 472440 998572
rect 429436 998532 472440 998560
rect 429436 998520 429442 998532
rect 472434 998520 472440 998532
rect 472492 998520 472498 998572
rect 514662 998520 514668 998572
rect 514720 998560 514726 998572
rect 524046 998560 524052 998572
rect 514720 998532 524052 998560
rect 514720 998520 514726 998532
rect 524046 998520 524052 998532
rect 524104 998520 524110 998572
rect 553118 998520 553124 998572
rect 553176 998560 553182 998572
rect 565814 998560 565820 998572
rect 553176 998532 565820 998560
rect 553176 998520 553182 998532
rect 565814 998520 565820 998532
rect 565872 998520 565878 998572
rect 200942 998452 200948 998504
rect 201000 998492 201006 998504
rect 203886 998492 203892 998504
rect 201000 998464 203892 998492
rect 201000 998452 201006 998464
rect 203886 998452 203892 998464
rect 203944 998452 203950 998504
rect 304258 998452 304264 998504
rect 304316 998492 304322 998504
rect 307294 998492 307300 998504
rect 304316 998464 307300 998492
rect 304316 998452 304322 998464
rect 307294 998452 307300 998464
rect 307352 998452 307358 998504
rect 92382 998384 92388 998436
rect 92440 998424 92446 998436
rect 100202 998424 100208 998436
rect 92440 998396 100208 998424
rect 92440 998384 92446 998396
rect 100202 998384 100208 998396
rect 100260 998384 100266 998436
rect 247402 998384 247408 998436
rect 247460 998424 247466 998436
rect 258994 998424 259000 998436
rect 247460 998396 259000 998424
rect 247460 998384 247466 998396
rect 258994 998384 259000 998396
rect 259052 998384 259058 998436
rect 351822 998384 351828 998436
rect 351880 998424 351886 998436
rect 382274 998424 382280 998436
rect 351880 998396 382280 998424
rect 351880 998384 351886 998396
rect 382274 998384 382280 998396
rect 382332 998384 382338 998436
rect 429194 998384 429200 998436
rect 429252 998424 429258 998436
rect 472250 998424 472256 998436
rect 429252 998396 472256 998424
rect 429252 998384 429258 998396
rect 472250 998384 472256 998396
rect 472308 998384 472314 998436
rect 499298 998384 499304 998436
rect 499356 998424 499362 998436
rect 517514 998424 517520 998436
rect 499356 998396 517520 998424
rect 499356 998384 499362 998396
rect 517514 998384 517520 998396
rect 517572 998384 517578 998436
rect 552290 998384 552296 998436
rect 552348 998424 552354 998436
rect 572714 998424 572720 998436
rect 552348 998396 572720 998424
rect 552348 998384 552354 998396
rect 572714 998384 572720 998396
rect 572772 998384 572778 998436
rect 200206 998316 200212 998368
rect 200264 998356 200270 998368
rect 202966 998356 202972 998368
rect 200264 998328 202972 998356
rect 200264 998316 200270 998328
rect 202966 998316 202972 998328
rect 203024 998316 203030 998368
rect 303062 998316 303068 998368
rect 303120 998356 303126 998368
rect 306098 998356 306104 998368
rect 303120 998328 306104 998356
rect 303120 998316 303126 998328
rect 306098 998316 306104 998328
rect 306156 998316 306162 998368
rect 247034 998248 247040 998300
rect 247092 998288 247098 998300
rect 253658 998288 253664 998300
rect 247092 998260 253664 998288
rect 247092 998248 247098 998260
rect 253658 998248 253664 998260
rect 253716 998248 253722 998300
rect 304442 998180 304448 998232
rect 304500 998220 304506 998232
rect 306926 998220 306932 998232
rect 304500 998192 306932 998220
rect 304500 998180 304506 998192
rect 306926 998180 306932 998192
rect 306984 998180 306990 998232
rect 568022 998180 568028 998232
rect 568080 998220 568086 998232
rect 572898 998220 572904 998232
rect 568080 998192 572904 998220
rect 568080 998180 568086 998192
rect 572898 998180 572904 998192
rect 572956 998180 572962 998232
rect 197998 998112 198004 998164
rect 198056 998152 198062 998164
rect 201862 998152 201868 998164
rect 198056 998124 201868 998152
rect 198056 998112 198062 998124
rect 201862 998112 201868 998124
rect 201920 998112 201926 998164
rect 202138 998112 202144 998164
rect 202196 998152 202202 998164
rect 205542 998152 205548 998164
rect 202196 998124 205548 998152
rect 202196 998112 202202 998124
rect 205542 998112 205548 998124
rect 205600 998112 205606 998164
rect 246758 998112 246764 998164
rect 246816 998152 246822 998164
rect 251082 998152 251088 998164
rect 246816 998124 251088 998152
rect 246816 998112 246822 998124
rect 251082 998112 251088 998124
rect 251140 998112 251146 998164
rect 258166 998112 258172 998164
rect 258224 998152 258230 998164
rect 259454 998152 259460 998164
rect 258224 998124 259460 998152
rect 258224 998112 258230 998124
rect 259454 998112 259460 998124
rect 259512 998112 259518 998164
rect 92566 998044 92572 998096
rect 92624 998084 92630 998096
rect 96246 998084 96252 998096
rect 92624 998056 96252 998084
rect 92624 998044 92630 998056
rect 96246 998044 96252 998056
rect 96304 998044 96310 998096
rect 260190 998044 260196 998096
rect 260248 998084 260254 998096
rect 262858 998084 262864 998096
rect 260248 998056 262864 998084
rect 260248 998044 260254 998056
rect 262858 998044 262864 998056
rect 262916 998044 262922 998096
rect 305638 998044 305644 998096
rect 305696 998084 305702 998096
rect 307754 998084 307760 998096
rect 305696 998056 307760 998084
rect 305696 998044 305702 998056
rect 307754 998044 307760 998056
rect 307812 998044 307818 998096
rect 308398 998044 308404 998096
rect 308456 998084 308462 998096
rect 310606 998084 310612 998096
rect 308456 998056 310612 998084
rect 308456 998044 308462 998056
rect 310606 998044 310612 998056
rect 310664 998044 310670 998096
rect 199378 997976 199384 998028
rect 199436 998016 199442 998028
rect 202690 998016 202696 998028
rect 199436 997988 202696 998016
rect 199436 997976 199442 997988
rect 202690 997976 202696 997988
rect 202748 997976 202754 998028
rect 250438 997976 250444 998028
rect 250496 998016 250502 998028
rect 253290 998016 253296 998028
rect 250496 997988 253296 998016
rect 250496 997976 250502 997988
rect 253290 997976 253296 997988
rect 253348 997976 253354 998028
rect 254578 997976 254584 998028
rect 254636 998016 254642 998028
rect 256510 998016 256516 998028
rect 254636 997988 256516 998016
rect 254636 997976 254642 997988
rect 256510 997976 256516 997988
rect 256568 997976 256574 998028
rect 259822 997908 259828 997960
rect 259880 997948 259886 997960
rect 262214 997948 262220 997960
rect 259880 997920 262220 997948
rect 259880 997908 259886 997920
rect 262214 997908 262220 997920
rect 262272 997908 262278 997960
rect 307202 997908 307208 997960
rect 307260 997948 307266 997960
rect 308950 997948 308956 997960
rect 307260 997920 308956 997948
rect 307260 997908 307266 997920
rect 308950 997908 308956 997920
rect 309008 997908 309014 997960
rect 591298 997908 591304 997960
rect 591356 997948 591362 997960
rect 625798 997948 625804 997960
rect 591356 997920 625804 997948
rect 591356 997908 591362 997920
rect 625798 997908 625804 997920
rect 625856 997908 625862 997960
rect 198366 997840 198372 997892
rect 198424 997880 198430 997892
rect 200666 997880 200672 997892
rect 198424 997852 200672 997880
rect 198424 997840 198430 997852
rect 200666 997840 200672 997852
rect 200724 997840 200730 997892
rect 247678 997840 247684 997892
rect 247736 997880 247742 997892
rect 252462 997880 252468 997892
rect 247736 997852 252468 997880
rect 247736 997840 247742 997852
rect 252462 997840 252468 997852
rect 252520 997840 252526 997892
rect 256326 997840 256332 997892
rect 256384 997880 256390 997892
rect 257338 997880 257344 997892
rect 256384 997852 257344 997880
rect 256384 997840 256390 997852
rect 257338 997840 257344 997852
rect 257396 997840 257402 997892
rect 202322 997772 202328 997824
rect 202380 997812 202386 997824
rect 204714 997812 204720 997824
rect 202380 997784 204720 997812
rect 202380 997772 202386 997784
rect 204714 997772 204720 997784
rect 204772 997772 204778 997824
rect 260190 997772 260196 997824
rect 260248 997812 260254 997824
rect 260926 997812 260932 997824
rect 260248 997784 260932 997812
rect 260248 997772 260254 997784
rect 260926 997772 260932 997784
rect 260984 997772 260990 997824
rect 302878 997772 302884 997824
rect 302936 997812 302942 997824
rect 306098 997812 306104 997824
rect 302936 997784 306104 997812
rect 302936 997772 302942 997784
rect 306098 997772 306104 997784
rect 306156 997772 306162 997824
rect 307018 997772 307024 997824
rect 307076 997812 307082 997824
rect 308122 997812 308128 997824
rect 307076 997784 308128 997812
rect 307076 997772 307082 997784
rect 308122 997772 308128 997784
rect 308180 997772 308186 997824
rect 549162 997772 549168 997824
rect 549220 997812 549226 997824
rect 551462 997812 551468 997824
rect 549220 997784 551468 997812
rect 549220 997772 549226 997784
rect 551462 997772 551468 997784
rect 551520 997772 551526 997824
rect 590838 997772 590844 997824
rect 590896 997812 590902 997824
rect 625614 997812 625620 997824
rect 590896 997784 625620 997812
rect 590896 997772 590902 997784
rect 625614 997772 625620 997784
rect 625672 997772 625678 997824
rect 93486 997704 93492 997756
rect 93544 997744 93550 997756
rect 106458 997744 106464 997756
rect 93544 997716 106464 997744
rect 93544 997704 93550 997716
rect 106458 997704 106464 997716
rect 106516 997704 106522 997756
rect 113818 997704 113824 997756
rect 113876 997744 113882 997756
rect 117130 997744 117136 997756
rect 113876 997716 117136 997744
rect 113876 997704 113882 997716
rect 117130 997704 117136 997716
rect 117188 997704 117194 997756
rect 143718 997704 143724 997756
rect 143776 997744 143782 997756
rect 160094 997744 160100 997756
rect 143776 997716 160100 997744
rect 143776 997704 143782 997716
rect 160094 997704 160100 997716
rect 160152 997704 160158 997756
rect 246574 997704 246580 997756
rect 246632 997744 246638 997756
rect 256326 997744 256332 997756
rect 246632 997716 256332 997744
rect 246632 997704 246638 997716
rect 256326 997704 256332 997716
rect 256384 997704 256390 997756
rect 359458 997704 359464 997756
rect 359516 997744 359522 997756
rect 372338 997744 372344 997756
rect 359516 997716 372344 997744
rect 359516 997704 359522 997716
rect 372338 997704 372344 997716
rect 372396 997704 372402 997756
rect 425698 997704 425704 997756
rect 425756 997744 425762 997756
rect 439682 997744 439688 997756
rect 425756 997716 439688 997744
rect 425756 997704 425762 997716
rect 439682 997704 439688 997716
rect 439740 997704 439746 997756
rect 507302 997704 507308 997756
rect 507360 997744 507366 997756
rect 516870 997744 516876 997756
rect 507360 997716 516876 997744
rect 507360 997704 507366 997716
rect 516870 997704 516876 997716
rect 516928 997704 516934 997756
rect 195238 997636 195244 997688
rect 195296 997676 195302 997688
rect 198366 997676 198372 997688
rect 195296 997648 198372 997676
rect 195296 997636 195302 997648
rect 198366 997636 198372 997648
rect 198424 997636 198430 997688
rect 540882 997636 540888 997688
rect 540940 997676 540946 997688
rect 555418 997676 555424 997688
rect 540940 997648 555424 997676
rect 540940 997636 540946 997648
rect 555418 997636 555424 997648
rect 555476 997636 555482 997688
rect 573358 997636 573364 997688
rect 573416 997676 573422 997688
rect 623682 997676 623688 997688
rect 573416 997648 623688 997676
rect 573416 997636 573422 997648
rect 623682 997636 623688 997648
rect 623740 997636 623746 997688
rect 109494 997568 109500 997620
rect 109552 997608 109558 997620
rect 116210 997608 116216 997620
rect 109552 997580 116216 997608
rect 109552 997568 109558 997580
rect 116210 997568 116216 997580
rect 116268 997568 116274 997620
rect 153930 997608 153936 997620
rect 147646 997580 153936 997608
rect 144178 997500 144184 997552
rect 144236 997540 144242 997552
rect 147646 997540 147674 997580
rect 153930 997568 153936 997580
rect 153988 997568 153994 997620
rect 369854 997568 369860 997620
rect 369912 997608 369918 997620
rect 372522 997608 372528 997620
rect 369912 997580 372528 997608
rect 369912 997568 369918 997580
rect 372522 997568 372528 997580
rect 372580 997568 372586 997620
rect 433978 997568 433984 997620
rect 434036 997608 434042 997620
rect 439866 997608 439872 997620
rect 434036 997580 439872 997608
rect 434036 997568 434042 997580
rect 439866 997568 439872 997580
rect 439924 997568 439930 997620
rect 509878 997568 509884 997620
rect 509936 997608 509942 997620
rect 517054 997608 517060 997620
rect 509936 997580 517060 997608
rect 509936 997568 509942 997580
rect 517054 997568 517060 997580
rect 517112 997568 517118 997620
rect 144236 997512 147674 997540
rect 144236 997500 144242 997512
rect 551922 997500 551928 997552
rect 551980 997540 551986 997552
rect 591298 997540 591304 997552
rect 551980 997512 591304 997540
rect 551980 997500 551986 997512
rect 591298 997500 591304 997512
rect 591356 997500 591362 997552
rect 502334 997432 502340 997484
rect 502392 997472 502398 997484
rect 516686 997472 516692 997484
rect 502392 997444 516692 997472
rect 502392 997432 502398 997444
rect 516686 997432 516692 997444
rect 516744 997432 516750 997484
rect 571978 997364 571984 997416
rect 572036 997404 572042 997416
rect 590562 997404 590568 997416
rect 572036 997376 590568 997404
rect 572036 997364 572042 997376
rect 590562 997364 590568 997376
rect 590620 997364 590626 997416
rect 488902 997296 488908 997348
rect 488960 997336 488966 997348
rect 510614 997336 510620 997348
rect 488960 997308 510620 997336
rect 488960 997296 488966 997308
rect 510614 997296 510620 997308
rect 510672 997296 510678 997348
rect 565814 997296 565820 997348
rect 565872 997336 565878 997348
rect 570230 997336 570236 997348
rect 565872 997308 570236 997336
rect 565872 997296 565878 997308
rect 570230 997296 570236 997308
rect 570288 997296 570294 997348
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 205082 997268 205088 997280
rect 200264 997240 205088 997268
rect 200264 997228 200270 997240
rect 205082 997228 205088 997240
rect 205140 997228 205146 997280
rect 574738 997228 574744 997280
rect 574796 997268 574802 997280
rect 590838 997268 590844 997280
rect 574796 997240 590844 997268
rect 574796 997228 574802 997240
rect 590838 997228 590844 997240
rect 590896 997228 590902 997280
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 557534 997160 557540 997212
rect 557592 997200 557598 997212
rect 570782 997200 570788 997212
rect 557592 997172 570788 997200
rect 557592 997160 557598 997172
rect 570782 997160 570788 997172
rect 570840 997160 570846 997212
rect 399938 997092 399944 997144
rect 399996 997132 400002 997144
rect 431954 997132 431960 997144
rect 399996 997104 431960 997132
rect 399996 997092 400002 997104
rect 431954 997092 431960 997104
rect 432012 997092 432018 997144
rect 144546 997024 144552 997076
rect 144604 997064 144610 997076
rect 158714 997064 158720 997076
rect 144604 997036 158720 997064
rect 144604 997024 144610 997036
rect 158714 997024 158720 997036
rect 158772 997024 158778 997076
rect 320818 997024 320824 997076
rect 320876 997064 320882 997076
rect 332594 997064 332600 997076
rect 320876 997036 332600 997064
rect 320876 997024 320882 997036
rect 332594 997024 332600 997036
rect 332652 997024 332658 997076
rect 505738 997024 505744 997076
rect 505796 997064 505802 997076
rect 517698 997064 517704 997076
rect 505796 997036 517704 997064
rect 505796 997024 505802 997036
rect 517698 997024 517704 997036
rect 517756 997024 517762 997076
rect 549162 997024 549168 997076
rect 549220 997064 549226 997076
rect 617150 997064 617156 997076
rect 549220 997036 617156 997064
rect 549220 997024 549226 997036
rect 617150 997024 617156 997036
rect 617208 997024 617214 997076
rect 365162 996956 365168 997008
rect 365220 996996 365226 997008
rect 372706 996996 372712 997008
rect 365220 996968 372712 996996
rect 365220 996956 365226 996968
rect 372706 996956 372712 996968
rect 372764 996956 372770 997008
rect 572714 996888 572720 996940
rect 572772 996928 572778 996940
rect 590378 996928 590384 996940
rect 572772 996900 590384 996928
rect 572772 996888 572778 996900
rect 590378 996888 590384 996900
rect 590436 996888 590442 996940
rect 558178 996752 558184 996804
rect 558236 996792 558242 996804
rect 558236 996764 586514 996792
rect 558236 996752 558242 996764
rect 586486 996724 586514 996764
rect 590562 996724 590568 996736
rect 586486 996696 590568 996724
rect 590562 996684 590568 996696
rect 590620 996684 590626 996736
rect 143718 996480 143724 996532
rect 143776 996520 143782 996532
rect 151262 996520 151268 996532
rect 143776 996492 151268 996520
rect 143776 996480 143782 996492
rect 151262 996480 151268 996492
rect 151320 996480 151326 996532
rect 92934 996344 92940 996396
rect 92992 996384 92998 996396
rect 121730 996384 121736 996396
rect 92992 996356 121736 996384
rect 92992 996344 92998 996356
rect 121730 996344 121736 996356
rect 121788 996344 121794 996396
rect 144178 996344 144184 996396
rect 144236 996384 144242 996396
rect 149882 996384 149888 996396
rect 144236 996356 149888 996384
rect 144236 996344 144242 996356
rect 149882 996344 149888 996356
rect 149940 996344 149946 996396
rect 549438 996344 549444 996396
rect 549496 996384 549502 996396
rect 550634 996384 550640 996396
rect 549496 996356 550640 996384
rect 549496 996344 549502 996356
rect 550634 996344 550640 996356
rect 550692 996344 550698 996396
rect 253198 996208 253204 996260
rect 253256 996248 253262 996260
rect 263594 996248 263600 996260
rect 253256 996220 263600 996248
rect 253256 996208 253262 996220
rect 263594 996208 263600 996220
rect 263652 996208 263658 996260
rect 368934 996208 368940 996260
rect 368992 996248 368998 996260
rect 377582 996248 377588 996260
rect 368992 996220 377588 996248
rect 368992 996208 368998 996220
rect 377582 996208 377588 996220
rect 377640 996208 377646 996260
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 211154 996112 211160 996124
rect 171836 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 211798 996072 211804 996124
rect 211856 996112 211862 996124
rect 260926 996112 260932 996124
rect 211856 996084 260932 996112
rect 211856 996072 211862 996084
rect 260926 996072 260932 996084
rect 260984 996072 260990 996124
rect 279418 996072 279424 996124
rect 279476 996112 279482 996124
rect 316034 996112 316040 996124
rect 279476 996084 316040 996112
rect 279476 996072 279482 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 354582 996072 354588 996124
rect 354640 996112 354646 996124
rect 354640 996072 354674 996112
rect 366358 996072 366364 996124
rect 366416 996112 366422 996124
rect 402238 996112 402244 996124
rect 366416 996084 386460 996112
rect 366416 996072 366422 996084
rect 144362 995976 144368 995988
rect 136468 995948 144368 995976
rect 136468 995852 136496 995948
rect 144362 995936 144368 995948
rect 144420 995936 144426 995988
rect 168742 995936 168748 995988
rect 168800 995976 168806 995988
rect 171502 995976 171508 995988
rect 168800 995948 171508 995976
rect 168800 995936 168806 995948
rect 171502 995936 171508 995948
rect 171560 995936 171566 995988
rect 177298 995936 177304 995988
rect 177356 995976 177362 995988
rect 212534 995976 212540 995988
rect 177356 995948 212540 995976
rect 177356 995936 177362 995948
rect 212534 995936 212540 995948
rect 212592 995936 212598 995988
rect 229738 995936 229744 995988
rect 229796 995976 229802 995988
rect 229796 995948 255636 995976
rect 229796 995936 229802 995948
rect 136450 995800 136456 995852
rect 136508 995800 136514 995852
rect 168558 995800 168564 995852
rect 168616 995840 168622 995852
rect 171226 995840 171232 995852
rect 168616 995812 171232 995840
rect 168616 995800 168622 995812
rect 171226 995800 171232 995812
rect 171284 995800 171290 995852
rect 213178 995800 213184 995852
rect 213236 995840 213242 995852
rect 255406 995840 255412 995852
rect 213236 995812 255412 995840
rect 213236 995800 213242 995812
rect 255406 995800 255412 995812
rect 255464 995800 255470 995852
rect 255608 995840 255636 995948
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 298922 995976 298928 995988
rect 264296 995948 298928 995976
rect 264296 995936 264302 995948
rect 298922 995936 298928 995948
rect 298980 995936 298986 995988
rect 354646 995976 354674 996072
rect 382734 995976 382740 995988
rect 354646 995948 382740 995976
rect 382734 995936 382740 995948
rect 382792 995936 382798 995988
rect 386432 995908 386460 996084
rect 391952 996084 402244 996112
rect 391952 995976 391980 996084
rect 402238 996072 402244 996084
rect 402296 996072 402302 996124
rect 511258 996072 511264 996124
rect 511316 996112 511322 996124
rect 563054 996112 563060 996124
rect 511316 996084 563060 996112
rect 511316 996072 511322 996084
rect 563054 996072 563060 996084
rect 563112 996072 563118 996124
rect 560294 995976 560300 995988
rect 386984 995948 391980 995976
rect 527376 995948 560300 995976
rect 386984 995908 387012 995948
rect 386432 995880 387012 995908
rect 522298 995868 522304 995920
rect 522356 995908 522362 995920
rect 527376 995908 527404 995948
rect 560294 995936 560300 995948
rect 560352 995936 560358 995988
rect 570598 995936 570604 995988
rect 570656 995976 570662 995988
rect 570656 995948 627914 995976
rect 570656 995936 570662 995948
rect 522356 995880 527404 995908
rect 522356 995868 522362 995880
rect 262214 995840 262220 995852
rect 255608 995812 262220 995840
rect 262214 995800 262220 995812
rect 262272 995800 262278 995852
rect 262858 995800 262864 995852
rect 262916 995840 262922 995852
rect 313274 995840 313280 995852
rect 262916 995812 313280 995840
rect 262916 995800 262922 995812
rect 313274 995800 313280 995812
rect 313332 995800 313338 995852
rect 355778 995800 355784 995852
rect 355836 995840 355842 995852
rect 368934 995840 368940 995852
rect 355836 995812 368940 995840
rect 355836 995800 355842 995812
rect 368934 995800 368940 995812
rect 368992 995800 368998 995852
rect 369302 995800 369308 995852
rect 369360 995840 369366 995852
rect 383102 995840 383108 995852
rect 369360 995812 383108 995840
rect 369360 995800 369366 995812
rect 383102 995800 383108 995812
rect 383160 995800 383166 995852
rect 506198 995800 506204 995852
rect 506256 995840 506262 995852
rect 509050 995840 509056 995852
rect 506256 995812 509056 995840
rect 506256 995800 506262 995812
rect 509050 995800 509056 995812
rect 509108 995800 509114 995852
rect 540238 995800 540244 995852
rect 540296 995840 540302 995852
rect 561674 995840 561680 995852
rect 540296 995812 561680 995840
rect 540296 995800 540302 995812
rect 561674 995800 561680 995812
rect 561732 995800 561738 995852
rect 562134 995800 562140 995852
rect 562192 995840 562198 995852
rect 625614 995840 625620 995852
rect 562192 995812 625620 995840
rect 562192 995800 562198 995812
rect 625614 995800 625620 995812
rect 625672 995800 625678 995852
rect 627886 995840 627914 995948
rect 642082 995908 642088 995920
rect 633406 995880 642088 995908
rect 633406 995840 633434 995880
rect 642082 995868 642088 995880
rect 642140 995868 642146 995920
rect 627886 995812 633434 995840
rect 92198 995528 92204 995580
rect 92256 995568 92262 995580
rect 92750 995568 92756 995580
rect 92256 995540 92756 995568
rect 92256 995528 92262 995540
rect 92750 995528 92756 995540
rect 92808 995528 92814 995580
rect 170674 995528 170680 995580
rect 170732 995568 170738 995580
rect 170732 995540 171916 995568
rect 170732 995528 170738 995540
rect 171888 995415 171916 995540
rect 194962 995528 194968 995580
rect 195020 995568 195026 995580
rect 201678 995568 201684 995580
rect 195020 995540 201684 995568
rect 195020 995528 195026 995540
rect 201678 995528 201684 995540
rect 201736 995528 201742 995580
rect 255406 995528 255412 995580
rect 255464 995568 255470 995580
rect 261846 995568 261852 995580
rect 255464 995540 261852 995568
rect 255464 995528 255470 995540
rect 261846 995528 261852 995540
rect 261904 995528 261910 995580
rect 299566 995528 299572 995580
rect 299624 995568 299630 995580
rect 301682 995568 301688 995580
rect 299624 995540 301688 995568
rect 299624 995528 299630 995540
rect 301682 995528 301688 995540
rect 301740 995528 301746 995580
rect 364978 995528 364984 995580
rect 365036 995568 365042 995580
rect 369302 995568 369308 995580
rect 365036 995540 369308 995568
rect 365036 995528 365042 995540
rect 369302 995528 369308 995540
rect 369360 995528 369366 995580
rect 377582 995528 377588 995580
rect 377640 995568 377646 995580
rect 377640 995540 379514 995568
rect 377640 995528 377646 995540
rect 246206 995460 246212 995512
rect 246264 995500 246270 995512
rect 247218 995500 247224 995512
rect 246264 995472 247224 995500
rect 246264 995460 246270 995472
rect 247218 995460 247224 995472
rect 247276 995460 247282 995512
rect 300118 995392 300124 995444
rect 300176 995432 300182 995444
rect 304074 995432 304080 995444
rect 300176 995404 304080 995432
rect 300176 995392 300182 995404
rect 304074 995392 304080 995404
rect 304132 995392 304138 995444
rect 379486 995432 379514 995540
rect 380158 995528 380164 995580
rect 380216 995568 380222 995580
rect 383286 995568 383292 995580
rect 380216 995540 383292 995568
rect 380216 995528 380222 995540
rect 383286 995528 383292 995540
rect 383344 995528 383350 995580
rect 383470 995528 383476 995580
rect 383528 995568 383534 995580
rect 385586 995568 385592 995580
rect 383528 995540 385592 995568
rect 383528 995528 383534 995540
rect 385586 995528 385592 995540
rect 385644 995528 385650 995580
rect 472618 995528 472624 995580
rect 472676 995568 472682 995580
rect 473354 995568 473360 995580
rect 472676 995540 473360 995568
rect 472676 995528 472682 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 524046 995528 524052 995580
rect 524104 995568 524110 995580
rect 525334 995568 525340 995580
rect 524104 995540 525340 995568
rect 524104 995528 524110 995540
rect 525334 995528 525340 995540
rect 525392 995528 525398 995580
rect 554682 995528 554688 995580
rect 554740 995568 554746 995580
rect 562134 995568 562140 995580
rect 554740 995540 562140 995568
rect 554740 995528 554746 995540
rect 562134 995528 562140 995540
rect 562192 995528 562198 995580
rect 623682 995528 623688 995580
rect 623740 995568 623746 995580
rect 626534 995568 626540 995580
rect 623740 995540 626540 995568
rect 623740 995528 623746 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 388806 995432 388812 995444
rect 379486 995404 388812 995432
rect 388806 995392 388812 995404
rect 388864 995392 388870 995444
rect 389818 995392 389824 995444
rect 389876 995432 389882 995444
rect 389876 995404 398834 995432
rect 389876 995392 389882 995404
rect 171686 995277 171692 995329
rect 171744 995277 171750 995329
rect 180702 995324 180708 995376
rect 180760 995364 180766 995376
rect 182634 995364 182640 995376
rect 180760 995336 182640 995364
rect 180760 995324 180766 995336
rect 182634 995324 182640 995336
rect 182692 995324 182698 995376
rect 185118 995324 185124 995376
rect 185176 995364 185182 995376
rect 186774 995364 186780 995376
rect 185176 995336 186780 995364
rect 185176 995324 185182 995336
rect 186774 995324 186780 995336
rect 186832 995324 186838 995376
rect 193122 995324 193128 995376
rect 193180 995364 193186 995376
rect 198182 995364 198188 995376
rect 193180 995336 198188 995364
rect 193180 995324 193186 995336
rect 198182 995324 198188 995336
rect 198240 995324 198246 995376
rect 228358 995324 228364 995376
rect 228416 995364 228422 995376
rect 253198 995364 253204 995376
rect 228416 995336 253204 995364
rect 228416 995324 228422 995336
rect 253198 995324 253204 995336
rect 253256 995324 253262 995376
rect 296162 995324 296168 995376
rect 296220 995364 296226 995376
rect 298278 995364 298284 995376
rect 296220 995336 298284 995364
rect 296220 995324 296226 995336
rect 298278 995324 298284 995336
rect 298336 995324 298342 995376
rect 398806 995364 398834 995404
rect 415394 995392 415400 995444
rect 415452 995432 415458 995444
rect 415452 995404 415716 995432
rect 415452 995392 415458 995404
rect 415688 995387 415716 995404
rect 398926 995364 398932 995376
rect 398806 995336 398932 995364
rect 398926 995324 398932 995336
rect 398984 995324 398990 995376
rect 415688 995359 415978 995387
rect 374638 995256 374644 995308
rect 374696 995296 374702 995308
rect 397638 995296 397644 995308
rect 374696 995268 389036 995296
rect 374696 995256 374702 995268
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 178862 995188 178868 995240
rect 178920 995228 178926 995240
rect 180334 995228 180340 995240
rect 178920 995200 180340 995228
rect 178920 995188 178926 995200
rect 180334 995188 180340 995200
rect 180392 995188 180398 995240
rect 180472 995188 180478 995240
rect 180530 995228 180536 995240
rect 202138 995228 202144 995240
rect 180530 995200 202144 995228
rect 180530 995188 180536 995200
rect 202138 995188 202144 995200
rect 202196 995188 202202 995240
rect 235580 995188 235586 995240
rect 235638 995228 235644 995240
rect 253014 995228 253020 995240
rect 235638 995200 253020 995228
rect 235638 995188 235644 995200
rect 253014 995188 253020 995200
rect 253072 995188 253078 995240
rect 389008 995228 389036 995268
rect 394666 995268 397644 995296
rect 394666 995228 394694 995268
rect 397638 995256 397644 995268
rect 397696 995256 397702 995308
rect 416130 995235 416136 995287
rect 416188 995235 416194 995287
rect 389008 995200 394694 995228
rect 362218 995120 362224 995172
rect 362276 995160 362282 995172
rect 387518 995160 387524 995172
rect 362276 995132 387524 995160
rect 362276 995120 362282 995132
rect 387518 995120 387524 995132
rect 387576 995120 387582 995172
rect 532142 995120 532148 995172
rect 532200 995160 532206 995172
rect 540238 995160 540244 995172
rect 532200 995132 540244 995160
rect 532200 995120 532206 995132
rect 540238 995120 540244 995132
rect 540296 995120 540302 995172
rect 171232 995105 171284 995111
rect 171232 995047 171284 995053
rect 180150 995052 180156 995104
rect 180208 995092 180214 995104
rect 206278 995092 206284 995104
rect 180208 995064 206284 995092
rect 180208 995052 180214 995064
rect 206278 995052 206284 995064
rect 206336 995052 206342 995104
rect 235258 995052 235264 995104
rect 235316 995092 235322 995104
rect 253474 995092 253480 995104
rect 235316 995064 253480 995092
rect 235316 995052 235322 995064
rect 253474 995052 253480 995064
rect 253532 995052 253538 995104
rect 282822 995052 282828 995104
rect 282880 995092 282886 995104
rect 311894 995092 311900 995104
rect 282880 995064 311900 995092
rect 282880 995052 282886 995064
rect 311894 995052 311900 995064
rect 311952 995052 311958 995104
rect 451642 995052 451648 995104
rect 451700 995092 451706 995104
rect 485958 995092 485964 995104
rect 451700 995064 485964 995092
rect 451700 995052 451706 995064
rect 485958 995052 485964 995064
rect 486016 995052 486022 995104
rect 507118 995052 507124 995104
rect 507176 995092 507182 995104
rect 528186 995092 528192 995104
rect 507176 995064 528192 995092
rect 507176 995052 507182 995064
rect 528186 995052 528192 995064
rect 528244 995052 528250 995104
rect 556614 995052 556620 995104
rect 556672 995092 556678 995104
rect 639506 995092 639512 995104
rect 556672 995064 639512 995092
rect 556672 995052 556678 995064
rect 639506 995052 639512 995064
rect 639564 995052 639570 995104
rect 357434 994984 357440 995036
rect 357492 995024 357498 995036
rect 395154 995024 395160 995036
rect 357492 994996 395160 995024
rect 357492 994984 357498 994996
rect 395154 994984 395160 994996
rect 395212 994984 395218 995036
rect 171244 994881 171272 994967
rect 180702 994916 180708 994968
rect 180760 994956 180766 994968
rect 208394 994956 208400 994968
rect 180760 994928 208400 994956
rect 180760 994916 180766 994928
rect 208394 994916 208400 994928
rect 208452 994916 208458 994968
rect 232866 994916 232872 994968
rect 232924 994956 232930 994968
rect 256050 994956 256056 994968
rect 232924 994928 256056 994956
rect 232924 994916 232930 994928
rect 256050 994916 256056 994928
rect 256108 994916 256114 994968
rect 283466 994916 283472 994968
rect 283524 994956 283530 994968
rect 307018 994956 307024 994968
rect 283524 994928 307024 994956
rect 283524 994916 283530 994928
rect 307018 994916 307024 994928
rect 307076 994916 307082 994968
rect 474550 994916 474556 994968
rect 474608 994956 474614 994968
rect 482922 994956 482928 994968
rect 474608 994928 482928 994956
rect 474608 994916 474614 994928
rect 482922 994916 482928 994928
rect 482980 994916 482986 994968
rect 486602 994916 486608 994968
rect 486660 994956 486666 994968
rect 489914 994956 489920 994968
rect 486660 994928 489920 994956
rect 486660 994916 486666 994928
rect 489914 994916 489920 994928
rect 489972 994916 489978 994968
rect 519814 994916 519820 994968
rect 519872 994956 519878 994968
rect 530210 994956 530216 994968
rect 519872 994928 530216 994956
rect 519872 994916 519878 994928
rect 530210 994916 530216 994928
rect 530268 994916 530274 994968
rect 534350 994916 534356 994968
rect 534408 994956 534414 994968
rect 538122 994956 538128 994968
rect 534408 994928 538128 994956
rect 534408 994916 534414 994928
rect 538122 994916 538128 994928
rect 538180 994916 538186 994968
rect 570782 994916 570788 994968
rect 570840 994956 570846 994968
rect 640702 994956 640708 994968
rect 570840 994928 640708 994956
rect 570840 994916 570846 994928
rect 640702 994916 640708 994928
rect 640760 994916 640766 994968
rect 78306 994780 78312 994832
rect 78364 994820 78370 994832
rect 104158 994820 104164 994832
rect 78364 994792 104164 994820
rect 78364 994780 78370 994792
rect 104158 994780 104164 994792
rect 104216 994780 104222 994832
rect 132126 994780 132132 994832
rect 132184 994820 132190 994832
rect 142982 994820 142988 994832
rect 132184 994792 142988 994820
rect 132184 994780 132190 994792
rect 142982 994780 142988 994792
rect 143040 994780 143046 994832
rect 143166 994780 143172 994832
rect 143224 994820 143230 994832
rect 155954 994820 155960 994832
rect 143224 994792 155960 994820
rect 143224 994780 143230 994792
rect 155954 994780 155960 994792
rect 156012 994780 156018 994832
rect 171042 994829 171048 994881
rect 171100 994829 171106 994881
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 371878 994848 371884 994900
rect 371936 994888 371942 994900
rect 396994 994888 397000 994900
rect 371936 994860 397000 994888
rect 371936 994848 371942 994860
rect 396994 994848 397000 994860
rect 397052 994848 397058 994900
rect 286502 994780 286508 994832
rect 286560 994820 286566 994832
rect 305638 994820 305644 994832
rect 286560 994792 305644 994820
rect 286560 994780 286566 994792
rect 305638 994780 305644 994792
rect 305696 994780 305702 994832
rect 458818 994780 458824 994832
rect 458876 994820 458882 994832
rect 482278 994820 482284 994832
rect 458876 994792 482284 994820
rect 458876 994780 458882 994792
rect 482278 994780 482284 994792
rect 482336 994780 482342 994832
rect 501874 994780 501880 994832
rect 501932 994820 501938 994832
rect 539226 994820 539232 994832
rect 501932 994792 539232 994820
rect 501932 994780 501938 994792
rect 539226 994780 539232 994792
rect 539284 994780 539290 994832
rect 567838 994780 567844 994832
rect 567896 994820 567902 994832
rect 639046 994820 639052 994832
rect 567896 994792 639052 994820
rect 567896 994780 567902 994792
rect 639046 994780 639052 994792
rect 639104 994780 639110 994832
rect 168558 994712 168564 994764
rect 168616 994752 168622 994764
rect 250438 994752 250444 994764
rect 168616 994724 250444 994752
rect 168616 994712 168622 994724
rect 250438 994712 250444 994724
rect 250496 994712 250502 994764
rect 363598 994712 363604 994764
rect 363656 994752 363662 994764
rect 393958 994752 393964 994764
rect 363656 994724 393964 994752
rect 363656 994712 363662 994724
rect 393958 994712 393964 994724
rect 394016 994712 394022 994764
rect 81342 994644 81348 994696
rect 81400 994684 81406 994696
rect 98638 994684 98644 994696
rect 81400 994656 98644 994684
rect 81400 994644 81406 994656
rect 98638 994644 98644 994656
rect 98696 994644 98702 994696
rect 129734 994644 129740 994696
rect 129792 994684 129798 994696
rect 134886 994684 134892 994696
rect 129792 994656 134892 994684
rect 129792 994644 129798 994656
rect 134886 994644 134892 994656
rect 134944 994644 134950 994696
rect 157334 994684 157340 994696
rect 135088 994656 157340 994684
rect 77662 994508 77668 994560
rect 77720 994548 77726 994560
rect 97442 994548 97448 994560
rect 77720 994520 97448 994548
rect 77720 994508 77726 994520
rect 97442 994508 97448 994520
rect 97500 994508 97506 994560
rect 128446 994508 128452 994560
rect 128504 994548 128510 994560
rect 135088 994548 135116 994656
rect 157334 994644 157340 994656
rect 157392 994644 157398 994696
rect 284110 994644 284116 994696
rect 284168 994684 284174 994696
rect 308398 994684 308404 994696
rect 284168 994656 308404 994684
rect 284168 994644 284174 994656
rect 308398 994644 308404 994656
rect 308456 994644 308462 994696
rect 419442 994644 419448 994696
rect 419500 994684 419506 994696
rect 660408 994684 660436 995121
rect 660574 994983 660580 995035
rect 660632 994983 660638 995035
rect 419500 994656 660436 994684
rect 419500 994644 419506 994656
rect 660776 994628 660804 994897
rect 168742 994576 168748 994628
rect 168800 994616 168806 994628
rect 243078 994616 243084 994628
rect 168800 994588 243084 994616
rect 168800 994576 168806 994588
rect 243078 994576 243084 994588
rect 243136 994576 243142 994628
rect 244182 994576 244188 994628
rect 244240 994616 244246 994628
rect 246758 994616 246764 994628
rect 244240 994588 246764 994616
rect 244240 994576 244246 994588
rect 246758 994576 246764 994588
rect 246816 994576 246822 994628
rect 356054 994576 356060 994628
rect 356112 994616 356118 994628
rect 393314 994616 393320 994628
rect 356112 994588 393320 994616
rect 356112 994576 356118 994588
rect 393314 994576 393320 994588
rect 393372 994576 393378 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 154574 994548 154580 994560
rect 128504 994520 135116 994548
rect 137204 994520 154580 994548
rect 128504 994508 128510 994520
rect 80698 994372 80704 994424
rect 80756 994412 80762 994424
rect 93118 994412 93124 994424
rect 80756 994384 93124 994412
rect 80756 994372 80762 994384
rect 93118 994372 93124 994384
rect 93176 994372 93182 994424
rect 131574 994372 131580 994424
rect 131632 994412 131638 994424
rect 137204 994412 137232 994520
rect 154574 994508 154580 994520
rect 154632 994508 154638 994560
rect 420822 994508 420828 994560
rect 420880 994548 420886 994560
rect 590562 994548 590568 994560
rect 420880 994520 590568 994548
rect 420880 994508 420886 994520
rect 590562 994508 590568 994520
rect 590620 994508 590626 994560
rect 625614 994508 625620 994560
rect 625672 994548 625678 994560
rect 633986 994548 633992 994560
rect 625672 994520 633992 994548
rect 625672 994508 625678 994520
rect 633986 994508 633992 994520
rect 634044 994508 634050 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 168926 994440 168932 994492
rect 168984 994480 168990 994492
rect 298738 994480 298744 994492
rect 168984 994452 298744 994480
rect 168984 994440 168990 994452
rect 298738 994440 298744 994452
rect 298796 994440 298802 994492
rect 383286 994440 383292 994492
rect 383344 994480 383350 994492
rect 389818 994480 389824 994492
rect 383344 994452 389824 994480
rect 383344 994440 383350 994452
rect 389818 994440 389824 994452
rect 389876 994440 389882 994492
rect 142798 994412 142804 994424
rect 131632 994384 137232 994412
rect 137296 994384 142804 994412
rect 131632 994372 131638 994384
rect 129090 994236 129096 994288
rect 129148 994276 129154 994288
rect 137296 994276 137324 994384
rect 142798 994372 142804 994384
rect 142856 994372 142862 994424
rect 142982 994372 142988 994424
rect 143040 994412 143046 994424
rect 148502 994412 148508 994424
rect 143040 994384 148508 994412
rect 143040 994372 143046 994384
rect 148502 994372 148508 994384
rect 148560 994372 148566 994424
rect 461578 994372 461584 994424
rect 461636 994412 461642 994424
rect 461636 994384 474780 994412
rect 461636 994372 461642 994384
rect 186774 994304 186780 994356
rect 186832 994344 186838 994356
rect 194962 994344 194968 994356
rect 186832 994316 194968 994344
rect 186832 994304 186838 994316
rect 194962 994304 194968 994316
rect 195020 994304 195026 994356
rect 232222 994304 232228 994356
rect 232280 994344 232286 994356
rect 254578 994344 254584 994356
rect 232280 994316 254584 994344
rect 232280 994304 232286 994316
rect 254578 994304 254584 994316
rect 254636 994304 254642 994356
rect 382734 994304 382740 994356
rect 382792 994344 382798 994356
rect 392670 994344 392676 994356
rect 382792 994316 392676 994344
rect 382792 994304 382798 994316
rect 392670 994304 392676 994316
rect 392728 994304 392734 994356
rect 143166 994276 143172 994288
rect 129148 994248 137324 994276
rect 137388 994248 143172 994276
rect 129148 994236 129154 994248
rect 134886 994100 134892 994152
rect 134944 994140 134950 994152
rect 137388 994140 137416 994248
rect 143166 994236 143172 994248
rect 143224 994236 143230 994288
rect 186498 994276 186504 994288
rect 171106 994248 186504 994276
rect 171106 994208 171134 994248
rect 186498 994236 186504 994248
rect 186556 994236 186562 994288
rect 295334 994236 295340 994288
rect 295392 994276 295398 994288
rect 381170 994276 381176 994288
rect 295392 994248 381176 994276
rect 295392 994236 295398 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 396350 994236 396356 994288
rect 396408 994276 396414 994288
rect 446122 994276 446128 994288
rect 396408 994248 446128 994276
rect 396408 994236 396414 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 456794 994236 456800 994288
rect 456852 994276 456858 994288
rect 474550 994276 474556 994288
rect 456852 994248 474556 994276
rect 456852 994236 456858 994248
rect 474550 994236 474556 994248
rect 474608 994236 474614 994288
rect 474752 994276 474780 994384
rect 475378 994372 475384 994424
rect 475436 994412 475442 994424
rect 487798 994412 487804 994424
rect 475436 994384 487804 994412
rect 475436 994372 475442 994384
rect 487798 994372 487804 994384
rect 487856 994372 487862 994424
rect 496722 994372 496728 994424
rect 496780 994412 496786 994424
rect 519814 994412 519820 994424
rect 496780 994384 519820 994412
rect 496780 994372 496786 994384
rect 519814 994372 519820 994384
rect 519872 994372 519878 994424
rect 523678 994372 523684 994424
rect 523736 994412 523742 994424
rect 538306 994412 538312 994424
rect 523736 994384 538312 994412
rect 523736 994372 523742 994384
rect 538306 994372 538312 994384
rect 538364 994372 538370 994424
rect 489914 994276 489920 994288
rect 474752 994248 489920 994276
rect 489914 994236 489920 994248
rect 489972 994236 489978 994288
rect 500862 994236 500868 994288
rect 500920 994276 500926 994288
rect 500920 994248 524414 994276
rect 500920 994236 500926 994248
rect 151786 994180 171134 994208
rect 134944 994112 137416 994140
rect 134944 994100 134950 994112
rect 144914 994100 144920 994152
rect 144972 994140 144978 994152
rect 151786 994140 151814 994180
rect 300118 994140 300124 994152
rect 144972 994112 151814 994140
rect 173452 994112 300124 994140
rect 144972 994100 144978 994112
rect 169386 994032 169392 994084
rect 169444 994072 169450 994084
rect 173452 994072 173480 994112
rect 300118 994100 300124 994112
rect 300176 994100 300182 994152
rect 466454 994100 466460 994152
rect 466512 994140 466518 994152
rect 475378 994140 475384 994152
rect 466512 994112 475384 994140
rect 466512 994100 466518 994112
rect 475378 994100 475384 994112
rect 475436 994100 475442 994152
rect 518342 994100 518348 994152
rect 518400 994140 518406 994152
rect 523678 994140 523684 994152
rect 518400 994112 523684 994140
rect 518400 994100 518406 994112
rect 523678 994100 523684 994112
rect 523736 994100 523742 994152
rect 524386 994140 524414 994248
rect 530210 994236 530216 994288
rect 530268 994276 530274 994288
rect 537662 994276 537668 994288
rect 530268 994248 537668 994276
rect 530268 994236 530274 994248
rect 537662 994236 537668 994248
rect 537720 994236 537726 994288
rect 550634 994236 550640 994288
rect 550692 994276 550698 994288
rect 572714 994276 572720 994288
rect 550692 994248 572720 994276
rect 550692 994236 550698 994248
rect 572714 994236 572720 994248
rect 572772 994236 572778 994288
rect 535546 994140 535552 994152
rect 524386 994112 535552 994140
rect 535546 994100 535552 994112
rect 535604 994100 535610 994152
rect 169444 994044 173480 994072
rect 169444 994032 169450 994044
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 142798 993964 142804 994016
rect 142856 994004 142862 994016
rect 151078 994004 151084 994016
rect 142856 993976 151084 994004
rect 142856 993964 142862 993976
rect 151078 993964 151084 993976
rect 151136 993964 151142 994016
rect 180334 993964 180340 994016
rect 180392 994004 180398 994016
rect 196618 994004 196624 994016
rect 180392 993976 196624 994004
rect 180392 993964 180398 993976
rect 196618 993964 196624 993976
rect 196676 993964 196682 994016
rect 243906 993964 243912 994016
rect 243964 994004 243970 994016
rect 247402 994004 247408 994016
rect 243964 993976 247408 994004
rect 243964 993964 243970 993976
rect 247402 993964 247408 993976
rect 247460 993964 247466 994016
rect 569218 993896 569224 993948
rect 569276 993936 569282 993948
rect 661328 993936 661356 994561
rect 569276 993908 661356 993936
rect 569276 993896 569282 993908
rect 243078 993828 243084 993880
rect 243136 993868 243142 993880
rect 247678 993868 247684 993880
rect 243136 993840 247684 993868
rect 243136 993828 243142 993840
rect 247678 993828 247684 993840
rect 247736 993828 247742 993880
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 195238 993800 195244 993812
rect 171284 993772 195244 993800
rect 171284 993760 171290 993772
rect 195238 993760 195244 993772
rect 195296 993760 195302 993812
rect 520366 993760 520372 993812
rect 520424 993800 520430 993812
rect 660942 993800 660948 993812
rect 520424 993772 660948 993800
rect 520424 993760 520430 993772
rect 660942 993760 660948 993772
rect 661000 993760 661006 993812
rect 171042 993624 171048 993676
rect 171100 993664 171106 993676
rect 197998 993664 198004 993676
rect 171100 993636 198004 993664
rect 171100 993624 171106 993636
rect 197998 993624 198004 993636
rect 198056 993624 198062 993676
rect 517238 993624 517244 993676
rect 517296 993664 517302 993676
rect 660758 993664 660764 993676
rect 517296 993636 660764 993664
rect 517296 993624 517302 993636
rect 660758 993624 660764 993636
rect 660816 993624 660822 993676
rect 164878 993420 164884 993472
rect 164936 993460 164942 993472
rect 169754 993460 169760 993472
rect 164936 993432 169760 993460
rect 164936 993420 164942 993432
rect 169754 993420 169760 993432
rect 169812 993420 169818 993472
rect 214558 993420 214564 993472
rect 214616 993460 214622 993472
rect 219434 993460 219440 993472
rect 214616 993432 219440 993460
rect 214616 993420 214622 993432
rect 219434 993420 219440 993432
rect 219492 993420 219498 993472
rect 50338 993148 50344 993200
rect 50396 993188 50402 993200
rect 107746 993188 107752 993200
rect 50396 993160 107752 993188
rect 50396 993148 50402 993160
rect 107746 993148 107752 993160
rect 107804 993148 107810 993200
rect 44818 993012 44824 993064
rect 44876 993052 44882 993064
rect 109034 993052 109040 993064
rect 44876 993024 109040 993052
rect 44876 993012 44882 993024
rect 109034 993012 109040 993024
rect 109092 993012 109098 993064
rect 138014 993012 138020 993064
rect 138072 993052 138078 993064
rect 163130 993052 163136 993064
rect 138072 993024 163136 993052
rect 138072 993012 138078 993024
rect 163130 993012 163136 993024
rect 163188 993012 163194 993064
rect 318058 993012 318064 993064
rect 318116 993052 318122 993064
rect 349154 993052 349160 993064
rect 318116 993024 349160 993052
rect 318116 993012 318122 993024
rect 349154 993012 349160 993024
rect 349212 993012 349218 993064
rect 562502 993012 562508 993064
rect 562560 993052 562566 993064
rect 660298 993052 660304 993064
rect 562560 993024 660304 993052
rect 562560 993012 562566 993024
rect 660298 993012 660304 993024
rect 660356 993012 660362 993064
rect 54478 992876 54484 992928
rect 54536 992916 54542 992928
rect 148318 992916 148324 992928
rect 54536 992888 148324 992916
rect 54536 992876 54542 992888
rect 148318 992876 148324 992888
rect 148376 992876 148382 992928
rect 319438 992876 319444 992928
rect 319496 992916 319502 992928
rect 364978 992916 364984 992928
rect 319496 992888 364984 992916
rect 319496 992876 319502 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 367738 992876 367744 992928
rect 367796 992916 367802 992928
rect 429930 992916 429936 992928
rect 367796 992888 429936 992916
rect 367796 992876 367802 992888
rect 429930 992876 429936 992888
rect 429988 992876 429994 992928
rect 435358 992876 435364 992928
rect 435416 992916 435422 992928
rect 478966 992916 478972 992928
rect 435416 992888 478972 992916
rect 435416 992876 435422 992888
rect 478966 992876 478972 992888
rect 479024 992876 479030 992928
rect 560938 992876 560944 992928
rect 560996 992916 561002 992928
rect 668578 992916 668584 992928
rect 560996 992888 668584 992916
rect 560996 992876 561002 992888
rect 668578 992876 668584 992888
rect 668636 992876 668642 992928
rect 638862 992264 638868 992316
rect 638920 992304 638926 992316
rect 640794 992304 640800 992316
rect 638920 992276 640800 992304
rect 638920 992264 638926 992276
rect 640794 992264 640800 992276
rect 640852 992264 640858 992316
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 51718 991584 51724 991636
rect 51776 991624 51782 991636
rect 110414 991624 110420 991636
rect 51776 991596 110420 991624
rect 51776 991584 51782 991596
rect 110414 991584 110420 991596
rect 110472 991584 110478 991636
rect 55858 991448 55864 991500
rect 55916 991488 55922 991500
rect 146938 991488 146944 991500
rect 55916 991460 146944 991488
rect 55916 991448 55922 991460
rect 146938 991448 146944 991460
rect 146996 991448 147002 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 369118 991448 369124 991500
rect 369176 991488 369182 991500
rect 414106 991488 414112 991500
rect 369176 991460 414112 991488
rect 369176 991448 369182 991460
rect 414106 991448 414112 991460
rect 414164 991448 414170 991500
rect 512638 991448 512644 991500
rect 512696 991488 512702 991500
rect 543826 991488 543832 991500
rect 512696 991460 543832 991488
rect 512696 991448 512702 991460
rect 543826 991448 543832 991460
rect 543884 991448 543890 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 53282 990224 53288 990276
rect 53340 990264 53346 990276
rect 95878 990264 95884 990276
rect 53340 990236 95884 990264
rect 53340 990224 53346 990236
rect 95878 990224 95884 990236
rect 95936 990224 95942 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 108114 990128 108120 990140
rect 49016 990100 108120 990128
rect 49016 990088 49022 990100
rect 108114 990088 108120 990100
rect 108172 990088 108178 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 669958 990128 669964 990140
rect 562376 990100 669964 990128
rect 562376 990088 562382 990100
rect 669958 990088 669964 990100
rect 670016 990088 670022 990140
rect 572714 989476 572720 989528
rect 572772 989516 572778 989528
rect 576302 989516 576308 989528
rect 572772 989488 576308 989516
rect 572772 989476 572778 989488
rect 576302 989476 576308 989488
rect 576360 989476 576366 989528
rect 89622 987368 89628 987420
rect 89680 987408 89686 987420
rect 111794 987408 111800 987420
rect 89680 987380 111800 987408
rect 89680 987368 89686 987380
rect 111794 987368 111800 987380
rect 111852 987368 111858 987420
rect 563698 987368 563704 987420
rect 563756 987408 563762 987420
rect 608778 987408 608784 987420
rect 563756 987380 608784 987408
rect 563756 987368 563762 987380
rect 608778 987368 608784 987380
rect 608836 987368 608842 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 204898 986660 204904 986672
rect 203208 986632 204904 986660
rect 203208 986620 203214 986632
rect 204898 986620 204904 986632
rect 204956 986620 204962 986672
rect 438118 986076 438124 986128
rect 438176 986116 438182 986128
rect 462774 986116 462780 986128
rect 438176 986088 462780 986116
rect 438176 986076 438182 986088
rect 462774 986076 462780 986088
rect 462832 986076 462838 986128
rect 515398 986076 515404 986128
rect 515456 986116 515462 986128
rect 527634 986116 527640 986128
rect 515456 986088 527640 986116
rect 515456 986076 515462 986088
rect 527634 986076 527640 986088
rect 527692 986076 527698 986128
rect 566458 986076 566464 986128
rect 566516 986116 566522 986128
rect 592494 986116 592500 986128
rect 566516 986088 592500 986116
rect 566516 986076 566522 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 370498 985940 370504 985992
rect 370556 985980 370562 985992
rect 397822 985980 397828 985992
rect 370556 985952 397828 985980
rect 370556 985940 370562 985952
rect 397822 985940 397828 985952
rect 397880 985940 397886 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 495158 985980 495164 985992
rect 436796 985952 495164 985980
rect 436796 985940 436802 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 672718 975712 672724 975724
rect 651708 975684 672724 975712
rect 651708 975672 651714 975684
rect 672718 975672 672724 975684
rect 672776 975672 672782 975724
rect 46198 961868 46204 961920
rect 46256 961908 46262 961920
rect 62114 961908 62120 961920
rect 46256 961880 62120 961908
rect 46256 961868 46262 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952348 36544 952400
rect 36596 952388 36602 952400
rect 41690 952388 41696 952400
rect 36596 952360 41696 952388
rect 36596 952348 36602 952360
rect 41690 952348 41696 952360
rect 41748 952348 41754 952400
rect 33778 951464 33784 951516
rect 33836 951504 33842 951516
rect 41506 951504 41512 951516
rect 33836 951476 41512 951504
rect 33836 951464 33842 951476
rect 41506 951464 41512 951476
rect 41564 951464 41570 951516
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 663058 948104 663064 948116
rect 652260 948076 663064 948104
rect 652260 948064 652266 948076
rect 663058 948064 663064 948076
rect 663116 948064 663122 948116
rect 45554 945956 45560 946008
rect 45612 945996 45618 946008
rect 62114 945996 62120 946008
rect 45612 945968 62120 945996
rect 45612 945956 45618 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 28718 945276 28724 945328
rect 28776 945316 28782 945328
rect 31754 945316 31760 945328
rect 28776 945288 31760 945316
rect 28776 945276 28782 945288
rect 31754 945276 31760 945288
rect 31812 945276 31818 945328
rect 35802 942556 35808 942608
rect 35860 942596 35866 942608
rect 41598 942596 41604 942608
rect 35860 942568 41604 942596
rect 35860 942556 35866 942568
rect 41598 942556 41604 942568
rect 41656 942556 41662 942608
rect 35802 941196 35808 941248
rect 35860 941236 35866 941248
rect 41414 941236 41420 941248
rect 35860 941208 41420 941236
rect 35860 941196 35866 941208
rect 41414 941196 41420 941208
rect 41472 941196 41478 941248
rect 35802 939768 35808 939820
rect 35860 939808 35866 939820
rect 41598 939808 41604 939820
rect 35860 939780 41604 939808
rect 35860 939768 35866 939780
rect 41598 939768 41604 939780
rect 41656 939768 41662 939820
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 663058 921856 663064 921868
rect 651524 921828 663064 921856
rect 651524 921816 651530 921828
rect 663058 921816 663064 921828
rect 663116 921816 663122 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 665818 909480 665824 909492
rect 652444 909452 665824 909480
rect 652444 909440 652450 909452
rect 665818 909440 665824 909452
rect 665876 909440 665882 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 671338 895676 671344 895688
rect 651524 895648 671344 895676
rect 651524 895636 651530 895648
rect 671338 895636 671344 895648
rect 671396 895636 671402 895688
rect 44082 892752 44088 892764
rect 42858 892724 44088 892752
rect 42858 892466 42886 892724
rect 44082 892712 44088 892724
rect 44140 892712 44146 892764
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43070 892202 43076 892254
rect 43128 892202 43134 892254
rect 43088 892058 43116 892202
rect 44082 891936 44088 891948
rect 43180 891908 44088 891936
rect 43180 891854 43208 891908
rect 44082 891896 44088 891908
rect 44140 891896 44146 891948
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 652386 855584 652392 855636
rect 652444 855624 652450 855636
rect 664438 855624 664444 855636
rect 652444 855596 664444 855624
rect 652444 855584 652450 855596
rect 664438 855584 664444 855596
rect 664496 855584 664502 855636
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651834 841780 651840 841832
rect 651892 841820 651898 841832
rect 669958 841820 669964 841832
rect 651892 841792 669964 841820
rect 651892 841780 651898 841792
rect 669958 841780 669964 841792
rect 670016 841780 670022 841832
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817028 35808 817080
rect 35860 817068 35866 817080
rect 41690 817068 41696 817080
rect 35860 817040 41696 817068
rect 35860 817028 35866 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 41414 815640 41420 815652
rect 35860 815612 41420 815640
rect 35860 815600 35866 815612
rect 41414 815600 41420 815612
rect 41472 815600 41478 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 661678 815640 661684 815652
rect 651524 815612 661684 815640
rect 651524 815600 651530 815612
rect 661678 815600 661684 815612
rect 661736 815600 661742 815652
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 41598 814280 41604 814292
rect 35860 814252 41604 814280
rect 35860 814240 35866 814252
rect 41598 814240 41604 814252
rect 41656 814240 41662 814292
rect 41322 811452 41328 811504
rect 41380 811492 41386 811504
rect 41690 811492 41696 811504
rect 41380 811464 41696 811492
rect 41380 811452 41386 811464
rect 41690 811452 41696 811464
rect 41748 811452 41754 811504
rect 40586 808528 40592 808580
rect 40644 808568 40650 808580
rect 41598 808568 41604 808580
rect 40644 808540 41604 808568
rect 40644 808528 40650 808540
rect 41598 808528 41604 808540
rect 41656 808528 41662 808580
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 35158 802408 35164 802460
rect 35216 802448 35222 802460
rect 41690 802448 41696 802460
rect 35216 802420 41696 802448
rect 35216 802408 35222 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 35894 802272 35900 802324
rect 35952 802312 35958 802324
rect 41690 802312 41696 802324
rect 35952 802284 41696 802312
rect 35952 802272 35958 802284
rect 41690 802272 41696 802284
rect 41748 802272 41754 802324
rect 53098 793568 53104 793620
rect 53156 793608 53162 793620
rect 62114 793608 62120 793620
rect 53156 793580 62120 793608
rect 53156 793568 53162 793580
rect 62114 793568 62120 793580
rect 62172 793568 62178 793620
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 652386 775548 652392 775600
rect 652444 775588 652450 775600
rect 668394 775588 668400 775600
rect 652444 775560 668400 775588
rect 652444 775548 652450 775560
rect 668394 775548 668400 775560
rect 668452 775548 668458 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35526 768952 35532 769004
rect 35584 768992 35590 769004
rect 40034 768992 40040 769004
rect 35584 768964 40040 768992
rect 35584 768952 35590 768964
rect 40034 768952 40040 768964
rect 40092 768952 40098 769004
rect 35342 768816 35348 768868
rect 35400 768856 35406 768868
rect 41690 768856 41696 768868
rect 35400 768828 41696 768856
rect 35400 768816 35406 768828
rect 41690 768816 41696 768828
rect 41748 768816 41754 768868
rect 35802 768680 35808 768732
rect 35860 768720 35866 768732
rect 41322 768720 41328 768732
rect 35860 768692 41328 768720
rect 35860 768680 35866 768692
rect 41322 768680 41328 768692
rect 41380 768680 41386 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 35526 767320 35532 767372
rect 35584 767360 35590 767372
rect 37918 767360 37924 767372
rect 35584 767332 37924 767360
rect 35584 767320 35590 767332
rect 37918 767320 37924 767332
rect 37976 767320 37982 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 37090 763240 37096 763292
rect 37148 763280 37154 763292
rect 39298 763280 39304 763292
rect 37148 763252 39304 763280
rect 37148 763240 37154 763252
rect 39298 763240 39304 763252
rect 39356 763240 39362 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 672166 761880 672172 761932
rect 672224 761920 672230 761932
rect 672718 761920 672724 761932
rect 672224 761892 672724 761920
rect 672224 761880 672230 761892
rect 672718 761880 672724 761892
rect 672776 761880 672782 761932
rect 31018 759636 31024 759688
rect 31076 759676 31082 759688
rect 39114 759676 39120 759688
rect 31076 759648 39120 759676
rect 31076 759636 31082 759648
rect 39114 759636 39120 759648
rect 39172 759636 39178 759688
rect 37918 759024 37924 759076
rect 37976 759064 37982 759076
rect 41506 759064 41512 759076
rect 37976 759036 41512 759064
rect 37976 759024 37982 759036
rect 41506 759024 41512 759036
rect 41564 759024 41570 759076
rect 35158 758276 35164 758328
rect 35216 758316 35222 758328
rect 41690 758316 41696 758328
rect 35216 758288 41696 758316
rect 35216 758276 35222 758288
rect 41690 758276 41696 758288
rect 41748 758276 41754 758328
rect 676030 757120 676036 757172
rect 676088 757160 676094 757172
rect 676582 757160 676588 757172
rect 676088 757132 676588 757160
rect 676088 757120 676094 757132
rect 676582 757120 676588 757132
rect 676640 757120 676646 757172
rect 675846 754264 675852 754316
rect 675904 754304 675910 754316
rect 683114 754304 683120 754316
rect 675904 754276 683120 754304
rect 675904 754264 675910 754276
rect 683114 754264 683120 754276
rect 683172 754264 683178 754316
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 35802 730056 35808 730108
rect 35860 730096 35866 730108
rect 41690 730096 41696 730108
rect 35860 730068 41696 730096
rect 35860 730056 35866 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 674208 728640 674406 728668
rect 673362 728560 673368 728612
rect 673420 728600 673426 728612
rect 674208 728600 674236 728640
rect 673420 728572 674236 728600
rect 673420 728560 673426 728572
rect 670694 728424 670700 728476
rect 670752 728464 670758 728476
rect 670752 728436 674268 728464
rect 670752 728424 670758 728436
rect 673362 728288 673368 728340
rect 673420 728328 673426 728340
rect 673420 728300 674176 728328
rect 673420 728288 673426 728300
rect 673362 728084 673368 728136
rect 673420 728124 673426 728136
rect 673420 728096 674058 728124
rect 673420 728084 673426 728096
rect 41322 725908 41328 725960
rect 41380 725948 41386 725960
rect 41690 725948 41696 725960
rect 41380 725920 41696 725948
rect 41380 725908 41386 725920
rect 41690 725908 41696 725920
rect 41748 725908 41754 725960
rect 41322 724480 41328 724532
rect 41380 724520 41386 724532
rect 41690 724520 41696 724532
rect 41380 724492 41696 724520
rect 41380 724480 41386 724492
rect 41690 724480 41696 724492
rect 41748 724480 41754 724532
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 33778 715776 33784 715828
rect 33836 715816 33842 715828
rect 41690 715816 41696 715828
rect 33836 715788 41696 715816
rect 33836 715776 33842 715788
rect 41690 715776 41696 715788
rect 41748 715776 41754 715828
rect 33042 715640 33048 715692
rect 33100 715680 33106 715692
rect 41138 715680 41144 715692
rect 33100 715652 41144 715680
rect 33100 715640 33106 715652
rect 41138 715640 41144 715652
rect 41196 715640 41202 715692
rect 31662 715504 31668 715556
rect 31720 715544 31726 715556
rect 41690 715544 41696 715556
rect 31720 715516 41696 715544
rect 31720 715504 31726 715516
rect 41690 715504 41696 715516
rect 41748 715504 41754 715556
rect 36538 714824 36544 714876
rect 36596 714864 36602 714876
rect 41690 714864 41696 714876
rect 36596 714836 41696 714864
rect 36596 714824 36602 714836
rect 41690 714824 41696 714836
rect 41748 714824 41754 714876
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 651466 709316 651472 709368
rect 651524 709356 651530 709368
rect 664438 709356 664444 709368
rect 651524 709328 664444 709356
rect 651524 709316 651530 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 651466 696940 651472 696992
rect 651524 696980 651530 696992
rect 661862 696980 661868 696992
rect 651524 696952 661868 696980
rect 651524 696940 651530 696952
rect 661862 696940 661868 696952
rect 661920 696940 661926 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 41322 687216 41328 687268
rect 41380 687256 41386 687268
rect 41690 687256 41696 687268
rect 41380 687228 41696 687256
rect 41380 687216 41386 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 41322 683136 41328 683188
rect 41380 683176 41386 683188
rect 41690 683176 41696 683188
rect 41380 683148 41696 683176
rect 41380 683136 41386 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 651650 683136 651656 683188
rect 651708 683176 651714 683188
rect 669958 683176 669964 683188
rect 651708 683148 669964 683176
rect 651708 683136 651714 683148
rect 669958 683136 669964 683148
rect 670016 683136 670022 683188
rect 41322 681844 41328 681896
rect 41380 681884 41386 681896
rect 41690 681884 41696 681896
rect 41380 681856 41696 681884
rect 41380 681844 41386 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 40034 677968 40040 678020
rect 40092 678008 40098 678020
rect 41690 678008 41696 678020
rect 40092 677980 41696 678008
rect 40092 677968 40098 677980
rect 41690 677968 41696 677980
rect 41748 677968 41754 678020
rect 51718 674840 51724 674892
rect 51776 674880 51782 674892
rect 62114 674880 62120 674892
rect 51776 674852 62120 674880
rect 51776 674840 51782 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 40126 672772 40132 672784
rect 35216 672744 40132 672772
rect 35216 672732 35222 672744
rect 40126 672732 40132 672744
rect 40184 672732 40190 672784
rect 36722 672052 36728 672104
rect 36780 672092 36786 672104
rect 41506 672092 41512 672104
rect 36780 672064 41512 672092
rect 36780 672052 36786 672064
rect 41506 672052 41512 672064
rect 41564 672052 41570 672104
rect 39942 671712 39948 671764
rect 40000 671752 40006 671764
rect 41690 671752 41696 671764
rect 40000 671724 41696 671752
rect 40000 671712 40006 671724
rect 41690 671712 41696 671724
rect 41748 671712 41754 671764
rect 651466 669332 651472 669384
rect 651524 669372 651530 669384
rect 661678 669372 661684 669384
rect 651524 669344 661684 669372
rect 651524 669332 651530 669344
rect 661678 669332 661684 669344
rect 661736 669332 661742 669384
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651466 656888 651472 656940
rect 651524 656928 651530 656940
rect 663058 656928 663064 656940
rect 651524 656900 663064 656928
rect 651524 656888 651530 656900
rect 663058 656888 663064 656900
rect 663116 656888 663122 656940
rect 46198 647844 46204 647896
rect 46256 647884 46262 647896
rect 62114 647884 62120 647896
rect 46256 647856 62120 647884
rect 46256 647844 46262 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639072 35808 639124
rect 35860 639112 35866 639124
rect 40034 639112 40040 639124
rect 35860 639084 40040 639112
rect 35860 639072 35866 639084
rect 40034 639072 40040 639084
rect 40092 639072 40098 639124
rect 35618 638936 35624 638988
rect 35676 638976 35682 638988
rect 41506 638976 41512 638988
rect 35676 638948 41512 638976
rect 35676 638936 35682 638948
rect 41506 638936 41512 638948
rect 41564 638936 41570 638988
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 40034 637616 40040 637628
rect 35860 637588 40040 637616
rect 35860 637576 35866 637588
rect 40034 637576 40040 637588
rect 40092 637576 40098 637628
rect 35802 636216 35808 636268
rect 35860 636256 35866 636268
rect 41690 636256 41696 636268
rect 35860 636228 41696 636256
rect 35860 636216 35866 636228
rect 41690 636216 41696 636228
rect 41748 636216 41754 636268
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 40034 635876 40040 635928
rect 40092 635916 40098 635928
rect 41690 635916 41696 635928
rect 40092 635888 41696 635916
rect 40092 635876 40098 635888
rect 41690 635876 41696 635888
rect 41748 635876 41754 635928
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651466 629280 651472 629332
rect 651524 629320 651530 629332
rect 667198 629320 667204 629332
rect 651524 629292 667204 629320
rect 651524 629280 651530 629292
rect 667198 629280 667204 629292
rect 667256 629280 667262 629332
rect 675846 626560 675852 626612
rect 675904 626600 675910 626612
rect 676490 626600 676496 626612
rect 675904 626572 676496 626600
rect 675904 626560 675910 626572
rect 676490 626560 676496 626572
rect 676548 626560 676554 626612
rect 673362 623976 673368 624028
rect 673420 623976 673426 624028
rect 673380 623892 673408 623976
rect 673362 623840 673368 623892
rect 673420 623840 673426 623892
rect 50338 623772 50344 623824
rect 50396 623812 50402 623824
rect 62114 623812 62120 623824
rect 50396 623784 62120 623812
rect 50396 623772 50402 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 672626 620984 672632 621036
rect 672684 621024 672690 621036
rect 672994 621024 673000 621036
rect 672684 620996 673000 621024
rect 672684 620984 672690 620996
rect 672994 620984 673000 620996
rect 673052 620984 673058 621036
rect 672258 618332 672264 618384
rect 672316 618372 672322 618384
rect 672902 618372 672908 618384
rect 672316 618344 672908 618372
rect 672316 618332 672322 618344
rect 672902 618332 672908 618344
rect 672960 618332 672966 618384
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 43806 612932 43812 612944
rect 43286 612904 43812 612932
rect 43806 612892 43812 612904
rect 43864 612892 43870 612944
rect 43714 612728 43720 612740
rect 43397 612700 43720 612728
rect 43714 612688 43720 612700
rect 43772 612688 43778 612740
rect 43990 612592 43996 612604
rect 43502 612564 43996 612592
rect 43502 612510 43530 612564
rect 43990 612552 43996 612564
rect 44048 612552 44054 612604
rect 43582 612332 43634 612338
rect 43714 612280 43720 612332
rect 43772 612280 43778 612332
rect 43582 612274 43634 612280
rect 43732 612102 43760 612280
rect 46014 611912 46020 611924
rect 43838 611884 46020 611912
rect 46014 611872 46020 611884
rect 46072 611872 46078 611924
rect 47946 611708 47952 611720
rect 43957 611680 47952 611708
rect 47946 611668 47952 611680
rect 48004 611668 48010 611720
rect 46934 611504 46940 611516
rect 44068 611476 46940 611504
rect 46934 611464 46940 611476
rect 46992 611464 46998 611516
rect 44155 611312 44207 611318
rect 44155 611254 44207 611260
rect 44373 611056 44379 611108
rect 44431 611056 44437 611108
rect 44272 610972 44324 610978
rect 44391 610946 44419 611056
rect 44272 610914 44324 610920
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 664622 603140 664628 603152
rect 651524 603112 664628 603140
rect 651524 603100 651530 603112
rect 664622 603100 664628 603112
rect 664680 603100 664686 603152
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 41230 594668 41236 594720
rect 41288 594708 41294 594720
rect 41506 594708 41512 594720
rect 41288 594680 41512 594708
rect 41288 594668 41294 594680
rect 41506 594668 41512 594680
rect 41564 594668 41570 594720
rect 676030 591336 676036 591388
rect 676088 591376 676094 591388
rect 682378 591376 682384 591388
rect 676088 591348 682384 591376
rect 676088 591336 676094 591348
rect 682378 591336 682384 591348
rect 682436 591336 682442 591388
rect 652386 590656 652392 590708
rect 652444 590696 652450 590708
rect 658918 590696 658924 590708
rect 652444 590668 658924 590696
rect 652444 590656 652450 590668
rect 658918 590656 658924 590668
rect 658976 590656 658982 590708
rect 40494 589636 40500 589688
rect 40552 589676 40558 589688
rect 41690 589676 41696 589688
rect 40552 589648 41696 589676
rect 40552 589636 40558 589648
rect 41690 589636 41696 589648
rect 41748 589636 41754 589688
rect 33778 585760 33784 585812
rect 33836 585800 33842 585812
rect 39666 585800 39672 585812
rect 33836 585772 39672 585800
rect 33836 585760 33842 585772
rect 39666 585760 39672 585772
rect 39724 585760 39730 585812
rect 37918 585284 37924 585336
rect 37976 585324 37982 585336
rect 41414 585324 41420 585336
rect 37976 585296 41420 585324
rect 37976 585284 37982 585296
rect 41414 585284 41420 585296
rect 41472 585284 41478 585336
rect 36538 585148 36544 585200
rect 36596 585188 36602 585200
rect 40218 585188 40224 585200
rect 36596 585160 40224 585188
rect 36596 585148 36602 585160
rect 40218 585148 40224 585160
rect 40276 585148 40282 585200
rect 51718 583720 51724 583772
rect 51776 583760 51782 583772
rect 62114 583760 62120 583772
rect 51776 583732 62120 583760
rect 51776 583720 51782 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 666002 576892 666008 576904
rect 651524 576864 666008 576892
rect 651524 576852 651530 576864
rect 666002 576852 666008 576864
rect 666060 576852 666066 576904
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 659102 563088 659108 563100
rect 651708 563060 659108 563088
rect 651708 563048 651714 563060
rect 659102 563048 659108 563060
rect 659160 563048 659166 563100
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 41506 557580 41512 557592
rect 35860 557552 41512 557580
rect 35860 557540 35866 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 41690 554792 41696 554804
rect 35860 554764 41696 554792
rect 35860 554752 35866 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 35802 553528 35808 553580
rect 35860 553568 35866 553580
rect 41414 553568 41420 553580
rect 35860 553540 41420 553568
rect 35860 553528 35866 553540
rect 41414 553528 41420 553540
rect 41472 553528 41478 553580
rect 35618 553392 35624 553444
rect 35676 553432 35682 553444
rect 41690 553432 41696 553444
rect 35676 553404 41696 553432
rect 35676 553392 35682 553404
rect 41690 553392 41696 553404
rect 41748 553392 41754 553444
rect 41230 550740 41236 550792
rect 41288 550780 41294 550792
rect 41690 550780 41696 550792
rect 41288 550752 41696 550780
rect 41288 550740 41294 550752
rect 41690 550740 41696 550752
rect 41748 550740 41754 550792
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 41690 549352 41696 549364
rect 41386 549324 41696 549352
rect 41230 549244 41236 549296
rect 41288 549284 41294 549296
rect 41386 549284 41414 549324
rect 41690 549312 41696 549324
rect 41748 549312 41754 549364
rect 41288 549256 41414 549284
rect 41288 549244 41294 549256
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 675938 547612 675944 547664
rect 675996 547652 676002 547664
rect 678238 547652 678244 547664
rect 675996 547624 678244 547652
rect 675996 547612 676002 547624
rect 678238 547612 678244 547624
rect 678296 547612 678302 547664
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 37182 547448 37188 547460
rect 31812 547420 37188 547448
rect 31812 547408 31818 547420
rect 37182 547408 37188 547420
rect 37240 547408 37246 547460
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 41506 543028 41512 543040
rect 33836 543000 41512 543028
rect 33836 542988 33842 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 37182 542308 37188 542360
rect 37240 542348 37246 542360
rect 41690 542348 41696 542360
rect 37240 542320 41696 542348
rect 37240 542308 37246 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669958 536840 669964 536852
rect 651524 536812 669964 536840
rect 651524 536800 651530 536812
rect 669958 536800 669964 536812
rect 670016 536800 670022 536852
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 672718 532108 672724 532160
rect 672776 532148 672782 532160
rect 674006 532148 674012 532160
rect 672776 532120 674012 532148
rect 672776 532108 672782 532120
rect 674006 532108 674012 532120
rect 674064 532108 674070 532160
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 676030 518780 676036 518832
rect 676088 518820 676094 518832
rect 677870 518820 677876 518832
rect 676088 518792 677876 518820
rect 676088 518780 676094 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675846 503616 675852 503668
rect 675904 503656 675910 503668
rect 680998 503656 681004 503668
rect 675904 503628 681004 503656
rect 675904 503616 675910 503628
rect 680998 503616 681004 503628
rect 681056 503616 681062 503668
rect 675846 499536 675852 499588
rect 675904 499576 675910 499588
rect 679618 499576 679624 499588
rect 675904 499548 679624 499576
rect 675904 499536 675910 499548
rect 679618 499536 679624 499548
rect 679676 499536 679682 499588
rect 652570 494708 652576 494760
rect 652628 494748 652634 494760
rect 665818 494748 665824 494760
rect 652628 494720 665824 494748
rect 652628 494708 652634 494720
rect 665818 494708 665824 494720
rect 665876 494708 665882 494760
rect 675846 492668 675852 492720
rect 675904 492708 675910 492720
rect 683114 492708 683120 492720
rect 675904 492680 683120 492708
rect 675904 492668 675910 492680
rect 683114 492668 683120 492680
rect 683172 492668 683178 492720
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 670142 484412 670148 484424
rect 654106 484384 670148 484412
rect 670142 484372 670148 484384
rect 670200 484372 670206 484424
rect 675846 480360 675852 480412
rect 675904 480400 675910 480412
rect 683114 480400 683120 480412
rect 675904 480372 683120 480400
rect 675904 480360 675910 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 675846 476076 675852 476128
rect 675904 476116 675910 476128
rect 680354 476116 680360 476128
rect 675904 476088 680360 476116
rect 675904 476076 675910 476088
rect 680354 476076 680360 476088
rect 680412 476076 680418 476128
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 663058 470608 663064 470620
rect 651524 470580 663064 470608
rect 651524 470568 651530 470580
rect 663058 470568 663064 470580
rect 663116 470568 663122 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 676122 457444 676128 457496
rect 676180 457444 676186 457496
rect 676306 457444 676312 457496
rect 676364 457484 676370 457496
rect 676858 457484 676864 457496
rect 676364 457456 676864 457484
rect 676364 457444 676370 457456
rect 676858 457444 676864 457456
rect 676916 457444 676922 457496
rect 676140 457224 676168 457444
rect 676122 457172 676128 457224
rect 676180 457172 676186 457224
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 667198 456804 667204 456816
rect 652444 456776 667204 456804
rect 652444 456764 652450 456776
rect 667198 456764 667204 456776
rect 667256 456764 667262 456816
rect 673178 456764 673184 456816
rect 673236 456804 673242 456816
rect 673236 456776 673454 456804
rect 673236 456764 673242 456776
rect 673426 456668 673454 456776
rect 673426 456640 673988 456668
rect 673960 456246 673988 456640
rect 675846 456084 675852 456136
rect 675904 456124 675910 456136
rect 677134 456124 677140 456136
rect 675904 456096 677140 456124
rect 675904 456084 675910 456096
rect 677134 456084 677140 456096
rect 677192 456084 677198 456136
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673736 455864 673788 455870
rect 673736 455806 673788 455812
rect 673454 455540 673460 455592
rect 673512 455580 673518 455592
rect 673512 455552 673624 455580
rect 673512 455540 673518 455552
rect 673506 455388 673558 455394
rect 673506 455330 673558 455336
rect 672074 455200 672080 455252
rect 672132 455240 672138 455252
rect 672132 455212 673316 455240
rect 672132 455200 672138 455212
rect 673288 455022 673316 455212
rect 673388 455184 673440 455190
rect 673388 455126 673440 455132
rect 673158 454928 673164 454980
rect 673216 454928 673222 454980
rect 673040 454792 673046 454844
rect 673098 454792 673104 454844
rect 673176 454818 673204 454928
rect 673058 454614 673086 454792
rect 672810 454384 672816 454436
rect 672868 454384 672874 454436
rect 672828 454206 672856 454384
rect 672954 454232 673006 454238
rect 672954 454174 673006 454180
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 671338 430624 671344 430636
rect 651524 430596 671344 430624
rect 651524 430584 651530 430596
rect 671338 430584 671344 430596
rect 671396 430584 671402 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41322 423784 41328 423836
rect 41380 423824 41386 423836
rect 41690 423824 41696 423836
rect 41380 423796 41696 423824
rect 41380 423784 41386 423796
rect 41690 423784 41696 423796
rect 41748 423784 41754 423836
rect 40954 423172 40960 423224
rect 41012 423212 41018 423224
rect 41598 423212 41604 423224
rect 41012 423184 41604 423212
rect 41012 423172 41018 423184
rect 41598 423172 41604 423184
rect 41656 423172 41662 423224
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 661678 416820 661684 416832
rect 651892 416792 661684 416820
rect 651892 416780 651898 416792
rect 661678 416780 661684 416792
rect 661736 416780 661742 416832
rect 49142 415420 49148 415472
rect 49200 415460 49206 415472
rect 62114 415460 62120 415472
rect 49200 415432 62120 415460
rect 49200 415420 49206 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 36538 415352 36544 415404
rect 36596 415392 36602 415404
rect 41690 415392 41696 415404
rect 36596 415364 41696 415392
rect 36596 415352 36602 415364
rect 41690 415352 41696 415364
rect 41748 415352 41754 415404
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 41138 387064 41144 387116
rect 41196 387104 41202 387116
rect 41690 387104 41696 387116
rect 41196 387076 41696 387104
rect 41196 387064 41202 387076
rect 41690 387064 41696 387076
rect 41748 387064 41754 387116
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41690 382412 41696 382424
rect 41380 382384 41696 382412
rect 41380 382372 41386 382384
rect 41690 382372 41696 382384
rect 41748 382372 41754 382424
rect 41138 382236 41144 382288
rect 41196 382276 41202 382288
rect 41690 382276 41696 382288
rect 41196 382248 41696 382276
rect 41196 382236 41202 382248
rect 41690 382236 41696 382248
rect 41748 382236 41754 382288
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 41690 379556 41696 379568
rect 35860 379528 41696 379556
rect 35860 379516 35866 379528
rect 41690 379516 41696 379528
rect 41748 379516 41754 379568
rect 35802 375980 35808 376032
rect 35860 376020 35866 376032
rect 39482 376020 39488 376032
rect 35860 375992 39488 376020
rect 35860 375980 35866 375992
rect 39482 375980 39488 375992
rect 39540 375980 39546 376032
rect 51718 375368 51724 375420
rect 51776 375408 51782 375420
rect 62114 375408 62120 375420
rect 51776 375380 62120 375408
rect 51776 375368 51782 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 28902 371832 28908 371884
rect 28960 371872 28966 371884
rect 41690 371872 41696 371884
rect 28960 371844 41696 371872
rect 28960 371832 28966 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 651650 364352 651656 364404
rect 651708 364392 651714 364404
rect 663242 364392 663248 364404
rect 651708 364364 663248 364392
rect 651708 364352 651714 364364
rect 663242 364352 663248 364364
rect 663300 364352 663306 364404
rect 46382 362924 46388 362976
rect 46440 362964 46446 362976
rect 62114 362964 62120 362976
rect 46440 362936 62120 362964
rect 46440 362924 46446 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 45002 355784 45008 355836
rect 45060 355824 45066 355836
rect 45646 355824 45652 355836
rect 45060 355796 45652 355824
rect 45060 355784 45066 355796
rect 45646 355784 45652 355796
rect 45704 355784 45710 355836
rect 44634 355648 44640 355700
rect 44692 355688 44698 355700
rect 44692 355660 45048 355688
rect 44692 355648 44698 355660
rect 44569 354832 44575 354884
rect 44627 354872 44633 354884
rect 44627 354844 44839 354872
rect 44627 354832 44633 354844
rect 44575 354680 44627 354686
rect 44575 354622 44627 354628
rect 44811 354600 44839 354844
rect 44811 354572 44956 354600
rect 44793 354424 44799 354476
rect 44851 354424 44857 354476
rect 44686 354340 44738 354346
rect 44811 354314 44839 354424
rect 44686 354282 44738 354288
rect 44928 354110 44956 354572
rect 45020 354532 45048 355660
rect 45020 354504 45063 354532
rect 45035 353906 45063 354504
rect 45646 354056 45652 354068
rect 45158 354028 45652 354056
rect 45158 353702 45186 354028
rect 45646 354016 45652 354028
rect 45704 354016 45710 354068
rect 45922 353784 45928 353796
rect 45250 353756 45928 353784
rect 45250 353498 45278 353756
rect 45922 353744 45928 353756
rect 45980 353744 45986 353796
rect 45554 353240 45560 353252
rect 45385 353212 45560 353240
rect 45554 353200 45560 353212
rect 45612 353200 45618 353252
rect 651466 350548 651472 350600
rect 651524 350588 651530 350600
rect 667382 350588 667388 350600
rect 651524 350560 667388 350588
rect 651524 350548 651530 350560
rect 667382 350548 667388 350560
rect 667440 350548 667446 350600
rect 28902 345040 28908 345092
rect 28960 345080 28966 345092
rect 38286 345080 38292 345092
rect 28960 345052 38292 345080
rect 28960 345040 28966 345052
rect 38286 345040 38292 345052
rect 38344 345040 38350 345092
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 37918 339504 37924 339516
rect 35860 339476 37924 339504
rect 35860 339464 35866 339476
rect 37918 339464 37924 339476
rect 37976 339464 37982 339516
rect 651466 338104 651472 338156
rect 651524 338144 651530 338156
rect 666370 338144 666376 338156
rect 651524 338116 666376 338144
rect 651524 338104 651530 338116
rect 666370 338104 666376 338116
rect 666428 338104 666434 338156
rect 50338 336744 50344 336796
rect 50396 336784 50402 336796
rect 62114 336784 62120 336796
rect 50396 336756 62120 336784
rect 50396 336744 50402 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 666646 324340 666652 324352
rect 651524 324312 666652 324340
rect 651524 324300 651530 324312
rect 666646 324300 666652 324312
rect 666704 324300 666710 324352
rect 53098 310496 53104 310548
rect 53156 310536 53162 310548
rect 62114 310536 62120 310548
rect 53156 310508 62120 310536
rect 53156 310496 53162 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667198 310536 667204 310548
rect 651524 310508 667204 310536
rect 651524 310496 651530 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 676030 304852 676036 304904
rect 676088 304892 676094 304904
rect 676306 304892 676312 304904
rect 676088 304864 676312 304892
rect 676088 304852 676094 304864
rect 676306 304852 676312 304864
rect 676364 304852 676370 304904
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 678974 298092 678980 298104
rect 675904 298064 678980 298092
rect 675904 298052 675910 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676030 297032 676036 297084
rect 676088 297072 676094 297084
rect 680998 297072 681004 297084
rect 676088 297044 681004 297072
rect 676088 297032 676094 297044
rect 680998 297032 681004 297044
rect 681056 297032 681062 297084
rect 41322 285064 41328 285116
rect 41380 285104 41386 285116
rect 41690 285104 41696 285116
rect 41380 285076 41696 285104
rect 41380 285064 41386 285076
rect 41690 285064 41696 285076
rect 41748 285064 41754 285116
rect 32398 284928 32404 284980
rect 32456 284968 32462 284980
rect 41690 284968 41696 284980
rect 32456 284940 41696 284968
rect 32456 284928 32462 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667566 284356 667572 284368
rect 651524 284328 667572 284356
rect 651524 284316 651530 284328
rect 667566 284316 667572 284328
rect 667624 284316 667630 284368
rect 88334 275952 88340 276004
rect 88392 275992 88398 276004
rect 143350 275992 143356 276004
rect 88392 275964 143356 275992
rect 88392 275952 88398 275964
rect 143350 275952 143356 275964
rect 143408 275952 143414 276004
rect 156874 275952 156880 276004
rect 156932 275992 156938 276004
rect 193858 275992 193864 276004
rect 156932 275964 193864 275992
rect 156932 275952 156938 275964
rect 193858 275952 193864 275964
rect 193916 275952 193922 276004
rect 201770 275952 201776 276004
rect 201828 275992 201834 276004
rect 222102 275992 222108 276004
rect 201828 275964 222108 275992
rect 201828 275952 201834 275964
rect 222102 275952 222108 275964
rect 222160 275952 222166 276004
rect 389174 275952 389180 276004
rect 389232 275992 389238 276004
rect 393314 275992 393320 276004
rect 389232 275964 393320 275992
rect 389232 275952 389238 275964
rect 393314 275952 393320 275964
rect 393372 275952 393378 276004
rect 413094 275952 413100 276004
rect 413152 275992 413158 276004
rect 434714 275992 434720 276004
rect 413152 275964 434720 275992
rect 413152 275952 413158 275964
rect 434714 275952 434720 275964
rect 434772 275952 434778 276004
rect 437474 275952 437480 276004
rect 437532 275992 437538 276004
rect 450078 275992 450084 276004
rect 437532 275964 450084 275992
rect 437532 275952 437538 275964
rect 450078 275952 450084 275964
rect 450136 275952 450142 276004
rect 456794 275952 456800 276004
rect 456852 275992 456858 276004
rect 460658 275992 460664 276004
rect 456852 275964 460664 275992
rect 456852 275952 456858 275964
rect 460658 275952 460664 275964
rect 460716 275952 460722 276004
rect 460842 275952 460848 276004
rect 460900 275992 460906 276004
rect 502058 275992 502064 276004
rect 460900 275964 502064 275992
rect 460900 275952 460906 275964
rect 502058 275952 502064 275964
rect 502116 275952 502122 276004
rect 510246 275952 510252 276004
rect 510304 275992 510310 276004
rect 597830 275992 597836 276004
rect 510304 275964 597836 275992
rect 510304 275952 510310 275964
rect 597830 275952 597836 275964
rect 597888 275952 597894 276004
rect 95418 275816 95424 275868
rect 95476 275856 95482 275868
rect 104802 275856 104808 275868
rect 95476 275828 104808 275856
rect 95476 275816 95482 275828
rect 104802 275816 104808 275828
rect 104860 275816 104866 275868
rect 113174 275816 113180 275868
rect 113232 275856 113238 275868
rect 169938 275856 169944 275868
rect 113232 275828 169944 275856
rect 113232 275816 113238 275828
rect 169938 275816 169944 275828
rect 169996 275816 170002 275868
rect 181714 275816 181720 275868
rect 181772 275856 181778 275868
rect 218882 275856 218888 275868
rect 181772 275828 218888 275856
rect 181772 275816 181778 275828
rect 218882 275816 218888 275828
rect 218940 275816 218946 275868
rect 396350 275816 396356 275868
rect 396408 275856 396414 275868
rect 412266 275856 412272 275868
rect 396408 275828 412272 275856
rect 396408 275816 396414 275828
rect 412266 275816 412272 275828
rect 412324 275816 412330 275868
rect 416406 275816 416412 275868
rect 416464 275856 416470 275868
rect 463050 275856 463056 275868
rect 416464 275828 463056 275856
rect 416464 275816 416470 275828
rect 463050 275816 463056 275828
rect 463108 275816 463114 275868
rect 471146 275816 471152 275868
rect 471204 275856 471210 275868
rect 493778 275856 493784 275868
rect 471204 275828 493784 275856
rect 471204 275816 471210 275828
rect 493778 275816 493784 275828
rect 493836 275816 493842 275868
rect 493962 275816 493968 275868
rect 494020 275856 494026 275868
rect 497366 275856 497372 275868
rect 494020 275828 497372 275856
rect 494020 275816 494026 275828
rect 497366 275816 497372 275828
rect 497424 275816 497430 275868
rect 498194 275816 498200 275868
rect 498252 275856 498258 275868
rect 498252 275828 499574 275856
rect 498252 275816 498258 275828
rect 81250 275680 81256 275732
rect 81308 275720 81314 275732
rect 88978 275720 88984 275732
rect 81308 275692 88984 275720
rect 81308 275680 81314 275692
rect 88978 275680 88984 275692
rect 89036 275680 89042 275732
rect 103698 275680 103704 275732
rect 103756 275720 103762 275732
rect 160094 275720 160100 275732
rect 103756 275692 160100 275720
rect 103756 275680 103762 275692
rect 160094 275680 160100 275692
rect 160152 275680 160158 275732
rect 178126 275680 178132 275732
rect 178184 275720 178190 275732
rect 216858 275720 216864 275732
rect 178184 275692 216864 275720
rect 178184 275680 178190 275692
rect 216858 275680 216864 275692
rect 216916 275680 216922 275732
rect 370498 275680 370504 275732
rect 370556 275720 370562 275732
rect 388622 275720 388628 275732
rect 370556 275692 388628 275720
rect 370556 275680 370562 275692
rect 388622 275680 388628 275692
rect 388680 275680 388686 275732
rect 410058 275680 410064 275732
rect 410116 275720 410122 275732
rect 428826 275720 428832 275732
rect 410116 275692 428832 275720
rect 410116 275680 410122 275692
rect 428826 275680 428832 275692
rect 428884 275680 428890 275732
rect 433150 275680 433156 275732
rect 433208 275720 433214 275732
rect 487890 275720 487896 275732
rect 433208 275692 487896 275720
rect 433208 275680 433214 275692
rect 487890 275680 487896 275692
rect 487948 275680 487954 275732
rect 488074 275680 488080 275732
rect 488132 275720 488138 275732
rect 498746 275720 498752 275732
rect 488132 275692 498752 275720
rect 488132 275680 488138 275692
rect 498746 275680 498752 275692
rect 498804 275680 498810 275732
rect 499546 275720 499574 275828
rect 504174 275816 504180 275868
rect 504232 275856 504238 275868
rect 509142 275856 509148 275868
rect 504232 275828 509148 275856
rect 504232 275816 504238 275828
rect 509142 275816 509148 275828
rect 509200 275816 509206 275868
rect 512178 275816 512184 275868
rect 512236 275856 512242 275868
rect 519814 275856 519820 275868
rect 512236 275828 519820 275856
rect 512236 275816 512242 275828
rect 519814 275816 519820 275828
rect 519872 275816 519878 275868
rect 604914 275856 604920 275868
rect 520016 275828 604920 275856
rect 505646 275720 505652 275732
rect 499546 275692 505652 275720
rect 505646 275680 505652 275692
rect 505704 275680 505710 275732
rect 507118 275680 507124 275732
rect 507176 275720 507182 275732
rect 512730 275720 512736 275732
rect 507176 275692 512736 275720
rect 507176 275680 507182 275692
rect 512730 275680 512736 275692
rect 512788 275680 512794 275732
rect 512914 275680 512920 275732
rect 512972 275720 512978 275732
rect 516226 275720 516232 275732
rect 512972 275692 516232 275720
rect 512972 275680 512978 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 516778 275680 516784 275732
rect 516836 275720 516842 275732
rect 520016 275720 520044 275828
rect 604914 275816 604920 275828
rect 604972 275816 604978 275868
rect 516836 275692 520044 275720
rect 516836 275680 516842 275692
rect 520182 275680 520188 275732
rect 520240 275720 520246 275732
rect 525518 275720 525524 275732
rect 520240 275692 525524 275720
rect 520240 275680 520246 275692
rect 525518 275680 525524 275692
rect 525576 275680 525582 275732
rect 525886 275680 525892 275732
rect 525944 275720 525950 275732
rect 527266 275720 527272 275732
rect 525944 275692 527272 275720
rect 525944 275680 525950 275692
rect 527266 275680 527272 275692
rect 527324 275680 527330 275732
rect 527726 275680 527732 275732
rect 527784 275720 527790 275732
rect 611998 275720 612004 275732
rect 527784 275692 612004 275720
rect 527784 275680 527790 275692
rect 611998 275680 612004 275692
rect 612056 275680 612062 275732
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86862 275584 86868 275596
rect 76524 275556 86868 275584
rect 76524 275544 76530 275556
rect 86862 275544 86868 275556
rect 86920 275544 86926 275596
rect 96614 275544 96620 275596
rect 96672 275584 96678 275596
rect 156598 275584 156604 275596
rect 96672 275556 156604 275584
rect 96672 275544 96678 275556
rect 156598 275544 156604 275556
rect 156656 275544 156662 275596
rect 163958 275544 163964 275596
rect 164016 275584 164022 275596
rect 202138 275584 202144 275596
rect 164016 275556 202144 275584
rect 164016 275544 164022 275556
rect 202138 275544 202144 275556
rect 202196 275544 202202 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 233878 275584 233884 275596
rect 221976 275556 233884 275584
rect 221976 275544 221982 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 236086 275544 236092 275596
rect 236144 275584 236150 275596
rect 255498 275584 255504 275596
rect 236144 275556 255504 275584
rect 236144 275544 236150 275556
rect 255498 275544 255504 275556
rect 255556 275544 255562 275596
rect 350718 275544 350724 275596
rect 350776 275584 350782 275596
rect 361390 275584 361396 275596
rect 350776 275556 361396 275584
rect 350776 275544 350782 275556
rect 361390 275544 361396 275556
rect 361448 275544 361454 275596
rect 361574 275544 361580 275596
rect 361632 275584 361638 275596
rect 385034 275584 385040 275596
rect 361632 275556 385040 275584
rect 361632 275544 361638 275556
rect 385034 275544 385040 275556
rect 385092 275544 385098 275596
rect 388070 275544 388076 275596
rect 388128 275584 388134 275596
rect 418154 275584 418160 275596
rect 388128 275556 418160 275584
rect 388128 275544 388134 275556
rect 418154 275544 418160 275556
rect 418212 275544 418218 275596
rect 418338 275544 418344 275596
rect 418396 275584 418402 275596
rect 435910 275584 435916 275596
rect 418396 275556 435916 275584
rect 418396 275544 418402 275556
rect 435910 275544 435916 275556
rect 435968 275544 435974 275596
rect 439498 275544 439504 275596
rect 439556 275584 439562 275596
rect 494974 275584 494980 275596
rect 439556 275556 494980 275584
rect 439556 275544 439562 275556
rect 494974 275544 494980 275556
rect 495032 275544 495038 275596
rect 496814 275544 496820 275596
rect 496872 275584 496878 275596
rect 538214 275584 538220 275596
rect 496872 275556 538220 275584
rect 496872 275544 496878 275556
rect 538214 275544 538220 275556
rect 538272 275544 538278 275596
rect 542998 275584 543004 275596
rect 538416 275556 543004 275584
rect 85942 275408 85948 275460
rect 86000 275448 86006 275460
rect 146754 275448 146760 275460
rect 86000 275420 146760 275448
rect 86000 275408 86006 275420
rect 146754 275408 146760 275420
rect 146812 275408 146818 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 167730 275448 167736 275460
rect 160520 275420 167736 275448
rect 160520 275408 160526 275420
rect 167730 275408 167736 275420
rect 167788 275408 167794 275460
rect 171042 275408 171048 275460
rect 171100 275448 171106 275460
rect 210418 275448 210424 275460
rect 171100 275420 210424 275448
rect 171100 275408 171106 275420
rect 210418 275408 210424 275420
rect 210476 275408 210482 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 237374 275448 237380 275460
rect 218388 275420 237380 275448
rect 218388 275408 218394 275420
rect 237374 275408 237380 275420
rect 237432 275408 237438 275460
rect 260926 275408 260932 275460
rect 260984 275448 260990 275460
rect 273530 275448 273536 275460
rect 260984 275420 273536 275448
rect 260984 275408 260990 275420
rect 273530 275408 273536 275420
rect 273588 275408 273594 275460
rect 284570 275408 284576 275460
rect 284628 275448 284634 275460
rect 290090 275448 290096 275460
rect 284628 275420 290096 275448
rect 284628 275408 284634 275420
rect 290090 275408 290096 275420
rect 290148 275408 290154 275460
rect 341518 275408 341524 275460
rect 341576 275448 341582 275460
rect 354306 275448 354312 275460
rect 341576 275420 354312 275448
rect 341576 275408 341582 275420
rect 354306 275408 354312 275420
rect 354364 275408 354370 275460
rect 360194 275448 360200 275460
rect 354646 275420 360200 275448
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 142706 275272 142712 275324
rect 142764 275312 142770 275324
rect 183462 275312 183468 275324
rect 142764 275284 183468 275312
rect 142764 275272 142770 275284
rect 183462 275272 183468 275284
rect 183520 275272 183526 275324
rect 186406 275272 186412 275324
rect 186464 275312 186470 275324
rect 187786 275312 187792 275324
rect 186464 275284 187792 275312
rect 186464 275272 186470 275284
rect 187786 275272 187792 275284
rect 187844 275272 187850 275324
rect 188798 275272 188804 275324
rect 188856 275312 188862 275324
rect 222838 275312 222844 275324
rect 188856 275284 222844 275312
rect 188856 275272 188862 275284
rect 222838 275272 222844 275284
rect 222896 275272 222902 275324
rect 225414 275272 225420 275324
rect 225472 275312 225478 275324
rect 245102 275312 245108 275324
rect 225472 275284 245108 275312
rect 225472 275272 225478 275284
rect 245102 275272 245108 275284
rect 245160 275272 245166 275324
rect 250254 275272 250260 275324
rect 250312 275312 250318 275324
rect 266630 275312 266636 275324
rect 250312 275284 266636 275312
rect 250312 275272 250318 275284
rect 266630 275272 266636 275284
rect 266688 275272 266694 275324
rect 273898 275272 273904 275324
rect 273956 275312 273962 275324
rect 282914 275312 282920 275324
rect 273956 275284 282920 275312
rect 273956 275272 273962 275284
rect 282914 275272 282920 275284
rect 282972 275272 282978 275324
rect 334342 275272 334348 275324
rect 334400 275312 334406 275324
rect 338942 275312 338948 275324
rect 334400 275284 338948 275312
rect 334400 275272 334406 275284
rect 338942 275272 338948 275284
rect 339000 275272 339006 275324
rect 353110 275312 353116 275324
rect 344986 275284 353116 275312
rect 290458 275204 290464 275256
rect 290516 275244 290522 275256
rect 294322 275244 294328 275256
rect 290516 275216 294328 275244
rect 290516 275204 290522 275216
rect 294322 275204 294328 275216
rect 294380 275204 294386 275256
rect 74074 275136 74080 275188
rect 74132 275176 74138 275188
rect 77202 275176 77208 275188
rect 74132 275148 77208 275176
rect 74132 275136 74138 275148
rect 77202 275136 77208 275148
rect 77260 275136 77266 275188
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 162118 275176 162124 275188
rect 110840 275148 162124 275176
rect 110840 275136 110846 275148
rect 162118 275136 162124 275148
rect 162176 275136 162182 275188
rect 338942 275136 338948 275188
rect 339000 275176 339006 275188
rect 344986 275176 345014 275284
rect 353110 275272 353116 275284
rect 353168 275272 353174 275324
rect 353938 275272 353944 275324
rect 353996 275312 354002 275324
rect 354646 275312 354674 275420
rect 360194 275408 360200 275420
rect 360252 275408 360258 275460
rect 363046 275408 363052 275460
rect 363104 275448 363110 275460
rect 367278 275448 367284 275460
rect 363104 275420 367284 275448
rect 363104 275408 363110 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 369118 275408 369124 275460
rect 369176 275448 369182 275460
rect 377950 275448 377956 275460
rect 369176 275420 377956 275448
rect 369176 275408 369182 275420
rect 377950 275408 377956 275420
rect 378008 275408 378014 275460
rect 382274 275408 382280 275460
rect 382332 275448 382338 275460
rect 414566 275448 414572 275460
rect 382332 275420 414572 275448
rect 382332 275408 382338 275420
rect 414566 275408 414572 275420
rect 414624 275408 414630 275460
rect 415302 275408 415308 275460
rect 415360 275448 415366 275460
rect 425238 275448 425244 275460
rect 415360 275420 425244 275448
rect 415360 275408 415366 275420
rect 425238 275408 425244 275420
rect 425296 275408 425302 275460
rect 429194 275408 429200 275460
rect 429252 275448 429258 275460
rect 446490 275448 446496 275460
rect 429252 275420 446496 275448
rect 429252 275408 429258 275420
rect 446490 275408 446496 275420
rect 446548 275408 446554 275460
rect 449894 275408 449900 275460
rect 449952 275448 449958 275460
rect 504174 275448 504180 275460
rect 449952 275420 504180 275448
rect 449952 275408 449958 275420
rect 504174 275408 504180 275420
rect 504232 275408 504238 275460
rect 504358 275408 504364 275460
rect 504416 275448 504422 275460
rect 504416 275420 514064 275448
rect 504416 275408 504422 275420
rect 353996 275284 354674 275312
rect 353996 275272 354002 275284
rect 356330 275272 356336 275324
rect 356388 275312 356394 275324
rect 368474 275312 368480 275324
rect 356388 275284 368480 275312
rect 356388 275272 356394 275284
rect 368474 275272 368480 275284
rect 368532 275272 368538 275324
rect 375098 275272 375104 275324
rect 375156 275312 375162 275324
rect 403986 275312 403992 275324
rect 375156 275284 403992 275312
rect 375156 275272 375162 275284
rect 403986 275272 403992 275284
rect 404044 275272 404050 275324
rect 411254 275272 411260 275324
rect 411312 275312 411318 275324
rect 455966 275312 455972 275324
rect 411312 275284 455972 275312
rect 411312 275272 411318 275284
rect 455966 275272 455972 275284
rect 456024 275272 456030 275324
rect 456150 275272 456156 275324
rect 456208 275312 456214 275324
rect 512914 275312 512920 275324
rect 456208 275284 512920 275312
rect 456208 275272 456214 275284
rect 512914 275272 512920 275284
rect 512972 275272 512978 275324
rect 514036 275312 514064 275420
rect 517514 275408 517520 275460
rect 517572 275448 517578 275460
rect 521010 275448 521016 275460
rect 517572 275420 521016 275448
rect 517572 275408 517578 275420
rect 521010 275408 521016 275420
rect 521068 275408 521074 275460
rect 521194 275408 521200 275460
rect 521252 275448 521258 275460
rect 523402 275448 523408 275460
rect 521252 275420 523408 275448
rect 521252 275408 521258 275420
rect 523402 275408 523408 275420
rect 523460 275408 523466 275460
rect 530118 275448 530124 275460
rect 523696 275420 530124 275448
rect 523696 275312 523724 275420
rect 530118 275408 530124 275420
rect 530176 275408 530182 275460
rect 531314 275408 531320 275460
rect 531372 275448 531378 275460
rect 537570 275448 537576 275460
rect 531372 275420 537576 275448
rect 531372 275408 531378 275420
rect 537570 275408 537576 275420
rect 537628 275408 537634 275460
rect 538416 275448 538444 275556
rect 542998 275544 543004 275556
rect 543056 275544 543062 275596
rect 545114 275544 545120 275596
rect 545172 275584 545178 275596
rect 552658 275584 552664 275596
rect 545172 275556 552664 275584
rect 545172 275544 545178 275556
rect 552658 275544 552664 275556
rect 552716 275544 552722 275596
rect 552842 275544 552848 275596
rect 552900 275584 552906 275596
rect 552900 275556 586514 275584
rect 552900 275544 552906 275556
rect 577222 275448 577228 275460
rect 537772 275420 538444 275448
rect 538692 275420 577228 275448
rect 514036 275284 523724 275312
rect 525518 275272 525524 275324
rect 525576 275312 525582 275324
rect 527082 275312 527088 275324
rect 525576 275284 527088 275312
rect 525576 275272 525582 275284
rect 527082 275272 527088 275284
rect 527140 275272 527146 275324
rect 527266 275272 527272 275324
rect 527324 275312 527330 275324
rect 532786 275312 532792 275324
rect 527324 275284 532792 275312
rect 527324 275272 527330 275284
rect 532786 275272 532792 275284
rect 532844 275272 532850 275324
rect 532970 275272 532976 275324
rect 533028 275312 533034 275324
rect 535270 275312 535276 275324
rect 533028 275284 535276 275312
rect 533028 275272 533034 275284
rect 535270 275272 535276 275284
rect 535328 275272 535334 275324
rect 535454 275272 535460 275324
rect 535512 275312 535518 275324
rect 537772 275312 537800 275420
rect 535512 275284 537800 275312
rect 535512 275272 535518 275284
rect 537938 275272 537944 275324
rect 537996 275312 538002 275324
rect 538692 275312 538720 275420
rect 577222 275408 577228 275420
rect 577280 275408 577286 275460
rect 586486 275448 586514 275556
rect 599118 275448 599124 275460
rect 586486 275420 599124 275448
rect 599118 275408 599124 275420
rect 599176 275408 599182 275460
rect 611354 275408 611360 275460
rect 611412 275448 611418 275460
rect 616782 275448 616788 275460
rect 611412 275420 616788 275448
rect 611412 275408 611418 275420
rect 616782 275408 616788 275420
rect 616840 275408 616846 275460
rect 626166 275448 626172 275460
rect 620296 275420 626172 275448
rect 537996 275284 538720 275312
rect 537996 275272 538002 275284
rect 538858 275272 538864 275324
rect 538916 275312 538922 275324
rect 590746 275312 590752 275324
rect 538916 275284 590752 275312
rect 538916 275272 538922 275284
rect 590746 275272 590752 275284
rect 590804 275272 590810 275324
rect 620296 275312 620324 275420
rect 626166 275408 626172 275420
rect 626224 275408 626230 275460
rect 626442 275408 626448 275460
rect 626500 275448 626506 275460
rect 641622 275448 641628 275460
rect 626500 275420 641628 275448
rect 626500 275408 626506 275420
rect 641622 275408 641628 275420
rect 641680 275408 641686 275460
rect 596146 275284 620324 275312
rect 339000 275148 345014 275176
rect 339000 275136 339006 275148
rect 400582 275136 400588 275188
rect 400640 275176 400646 275188
rect 415762 275176 415768 275188
rect 400640 275148 415768 275176
rect 400640 275136 400646 275148
rect 415762 275136 415768 275148
rect 415820 275136 415826 275188
rect 427814 275136 427820 275188
rect 427872 275176 427878 275188
rect 442994 275176 443000 275188
rect 427872 275148 443000 275176
rect 427872 275136 427878 275148
rect 442994 275136 443000 275148
rect 443052 275136 443058 275188
rect 445938 275136 445944 275188
rect 445996 275176 446002 275188
rect 471330 275176 471336 275188
rect 445996 275148 471336 275176
rect 445996 275136 446002 275148
rect 471330 275136 471336 275148
rect 471388 275136 471394 275188
rect 484578 275136 484584 275188
rect 484636 275176 484642 275188
rect 488074 275176 488080 275188
rect 484636 275148 488080 275176
rect 484636 275136 484642 275148
rect 488074 275136 488080 275148
rect 488132 275136 488138 275188
rect 492490 275136 492496 275188
rect 492548 275176 492554 275188
rect 504358 275176 504364 275188
rect 492548 275148 504364 275176
rect 492548 275136 492554 275148
rect 504358 275136 504364 275148
rect 504416 275136 504422 275188
rect 505186 275136 505192 275188
rect 505244 275176 505250 275188
rect 506842 275176 506848 275188
rect 505244 275148 506848 275176
rect 505244 275136 505250 275148
rect 506842 275136 506848 275148
rect 506900 275136 506906 275188
rect 508038 275136 508044 275188
rect 508096 275176 508102 275188
rect 577038 275176 577044 275188
rect 508096 275148 577044 275176
rect 508096 275136 508102 275148
rect 577038 275136 577044 275148
rect 577096 275136 577102 275188
rect 577222 275136 577228 275188
rect 577280 275176 577286 275188
rect 596146 275176 596174 275284
rect 577280 275148 596174 275176
rect 577280 275136 577286 275148
rect 599118 275136 599124 275188
rect 599176 275176 599182 275188
rect 633342 275176 633348 275188
rect 599176 275148 633348 275176
rect 599176 275136 599182 275148
rect 633342 275136 633348 275148
rect 633400 275136 633406 275188
rect 224218 275068 224224 275120
rect 224276 275108 224282 275120
rect 226150 275108 226156 275120
rect 224276 275080 226156 275108
rect 224276 275068 224282 275080
rect 226150 275068 226156 275080
rect 226208 275068 226214 275120
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 182082 275040 182088 275052
rect 135680 275012 182088 275040
rect 135680 275000 135686 275012
rect 182082 275000 182088 275012
rect 182140 275000 182146 275052
rect 443362 275000 443368 275052
rect 443420 275040 443426 275052
rect 453574 275040 453580 275052
rect 443420 275012 453580 275040
rect 443420 275000 443426 275012
rect 453574 275000 453580 275012
rect 453632 275000 453638 275052
rect 462958 275000 462964 275052
rect 463016 275040 463022 275052
rect 467834 275040 467840 275052
rect 463016 275012 467840 275040
rect 463016 275000 463022 275012
rect 467834 275000 467840 275012
rect 467892 275000 467898 275052
rect 473078 275000 473084 275052
rect 473136 275040 473142 275052
rect 538030 275040 538036 275052
rect 473136 275012 538036 275040
rect 473136 275000 473142 275012
rect 538030 275000 538036 275012
rect 538088 275000 538094 275052
rect 540974 275040 540980 275052
rect 538324 275012 540980 275040
rect 71774 274932 71780 274984
rect 71832 274972 71838 274984
rect 73798 274972 73804 274984
rect 71832 274944 73804 274972
rect 71832 274932 71838 274944
rect 73798 274932 73804 274944
rect 73856 274932 73862 274984
rect 277486 274932 277492 274984
rect 277544 274972 277550 274984
rect 284294 274972 284300 274984
rect 277544 274944 284300 274972
rect 277544 274932 277550 274944
rect 284294 274932 284300 274944
rect 284352 274932 284358 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136542 274904 136548 274916
rect 129700 274876 136548 274904
rect 129700 274864 129706 274876
rect 136542 274864 136548 274876
rect 136600 274864 136606 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 185578 274904 185584 274916
rect 149848 274876 185584 274904
rect 149848 274864 149854 274876
rect 185578 274864 185584 274876
rect 185636 274864 185642 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 293402 274904 293408 274916
rect 289320 274876 293408 274904
rect 289320 274864 289326 274876
rect 293402 274864 293408 274876
rect 293460 274864 293466 274916
rect 453390 274864 453396 274916
rect 453448 274904 453454 274916
rect 457162 274904 457168 274916
rect 453448 274876 457168 274904
rect 453448 274864 453454 274876
rect 457162 274864 457168 274876
rect 457220 274864 457226 274916
rect 467742 274864 467748 274916
rect 467800 274904 467806 274916
rect 531314 274904 531320 274916
rect 467800 274876 531320 274904
rect 467800 274864 467806 274876
rect 531314 274864 531320 274876
rect 531372 274864 531378 274916
rect 531498 274864 531504 274916
rect 531556 274904 531562 274916
rect 533982 274904 533988 274916
rect 531556 274876 533988 274904
rect 531556 274864 531562 274876
rect 533982 274864 533988 274876
rect 534040 274864 534046 274916
rect 534166 274864 534172 274916
rect 534224 274904 534230 274916
rect 537202 274904 537208 274916
rect 534224 274876 537208 274904
rect 534224 274864 534230 274876
rect 537202 274864 537208 274876
rect 537260 274864 537266 274916
rect 537386 274864 537392 274916
rect 537444 274904 537450 274916
rect 538324 274904 538352 275012
rect 540974 275000 540980 275012
rect 541032 275000 541038 275052
rect 542998 275000 543004 275052
rect 543056 275040 543062 275052
rect 543056 275012 552520 275040
rect 543056 275000 543062 275012
rect 537444 274876 538352 274904
rect 537444 274864 537450 274876
rect 538490 274864 538496 274916
rect 538548 274904 538554 274916
rect 545850 274904 545856 274916
rect 538548 274876 545856 274904
rect 538548 274864 538554 274876
rect 545850 274864 545856 274876
rect 545908 274864 545914 274916
rect 546034 274864 546040 274916
rect 546092 274904 546098 274916
rect 550542 274904 550548 274916
rect 546092 274876 550548 274904
rect 546092 274864 546098 274876
rect 550542 274864 550548 274876
rect 550600 274864 550606 274916
rect 552492 274904 552520 275012
rect 552658 275000 552664 275052
rect 552716 275040 552722 275052
rect 578878 275040 578884 275052
rect 552716 275012 578884 275040
rect 552716 275000 552722 275012
rect 578878 275000 578884 275012
rect 578936 275000 578942 275052
rect 552842 274904 552848 274916
rect 552492 274876 552848 274904
rect 552842 274864 552848 274876
rect 552900 274864 552906 274916
rect 577038 274864 577044 274916
rect 577096 274904 577102 274916
rect 583662 274904 583668 274916
rect 577096 274876 583668 274904
rect 577096 274864 577102 274876
rect 583662 274864 583668 274876
rect 583720 274864 583726 274916
rect 604454 274864 604460 274916
rect 604512 274904 604518 274916
rect 607306 274904 607312 274916
rect 604512 274876 607312 274904
rect 604512 274864 604518 274876
rect 607306 274864 607312 274876
rect 607364 274864 607370 274916
rect 283374 274796 283380 274848
rect 283432 274836 283438 274848
rect 289078 274836 289084 274848
rect 283432 274808 289084 274836
rect 283432 274796 283438 274808
rect 289078 274796 289084 274808
rect 289136 274796 289142 274848
rect 407114 274796 407120 274848
rect 407172 274836 407178 274848
rect 411070 274836 411076 274848
rect 407172 274808 411076 274836
rect 407172 274796 407178 274808
rect 411070 274796 411076 274808
rect 411128 274796 411134 274848
rect 105998 274728 106004 274780
rect 106056 274768 106062 274780
rect 110414 274768 110420 274780
rect 106056 274740 110420 274768
rect 106056 274728 106062 274740
rect 110414 274728 110420 274740
rect 110472 274728 110478 274780
rect 140314 274728 140320 274780
rect 140372 274768 140378 274780
rect 144638 274768 144644 274780
rect 140372 274740 144644 274768
rect 140372 274728 140378 274740
rect 144638 274728 144644 274740
rect 144696 274728 144702 274780
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149882 274768 149888 274780
rect 146260 274740 149888 274768
rect 146260 274728 146266 274740
rect 149882 274728 149888 274740
rect 149940 274728 149946 274780
rect 425330 274728 425336 274780
rect 425388 274768 425394 274780
rect 432322 274768 432328 274780
rect 425388 274740 432328 274768
rect 425388 274728 425394 274740
rect 432322 274728 432328 274740
rect 432380 274728 432386 274780
rect 435542 274728 435548 274780
rect 435600 274768 435606 274780
rect 439038 274768 439044 274780
rect 435600 274740 439044 274768
rect 435600 274728 435606 274740
rect 439038 274728 439044 274740
rect 439096 274728 439102 274780
rect 462222 274728 462228 274780
rect 462280 274768 462286 274780
rect 466638 274768 466644 274780
rect 462280 274740 466644 274768
rect 462280 274728 462286 274740
rect 466638 274728 466644 274740
rect 466696 274728 466702 274780
rect 498746 274728 498752 274780
rect 498804 274768 498810 274780
rect 521194 274768 521200 274780
rect 498804 274740 521200 274768
rect 498804 274728 498810 274740
rect 521194 274728 521200 274740
rect 521252 274728 521258 274780
rect 521654 274728 521660 274780
rect 521712 274768 521718 274780
rect 526898 274768 526904 274780
rect 521712 274740 526904 274768
rect 521712 274728 521718 274740
rect 526898 274728 526904 274740
rect 526956 274728 526962 274780
rect 527082 274728 527088 274780
rect 527140 274768 527146 274780
rect 619082 274768 619088 274780
rect 527140 274740 619088 274768
rect 527140 274728 527146 274740
rect 619082 274728 619088 274740
rect 619140 274728 619146 274780
rect 66990 274660 66996 274712
rect 67048 274700 67054 274712
rect 71038 274700 71044 274712
rect 67048 274672 71044 274700
rect 67048 274660 67054 274672
rect 71038 274660 71044 274672
rect 71096 274660 71102 274712
rect 90634 274660 90640 274712
rect 90692 274700 90698 274712
rect 95878 274700 95884 274712
rect 90692 274672 95884 274700
rect 90692 274660 90698 274672
rect 95878 274660 95884 274672
rect 95936 274660 95942 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163130 274700 163136 274712
rect 161624 274672 163136 274700
rect 161624 274660 161630 274672
rect 163130 274660 163136 274672
rect 163188 274660 163194 274712
rect 170122 274660 170128 274712
rect 170180 274700 170186 274712
rect 173066 274700 173072 274712
rect 170180 274672 173072 274700
rect 170180 274660 170186 274672
rect 173066 274660 173072 274672
rect 173124 274660 173130 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 187142 274700 187148 274712
rect 185268 274672 187148 274700
rect 185268 274660 185274 274672
rect 187142 274660 187148 274672
rect 187200 274660 187206 274712
rect 210050 274660 210056 274712
rect 210108 274700 210114 274712
rect 210108 274672 212580 274700
rect 210108 274660 210114 274672
rect 104802 274592 104808 274644
rect 104860 274632 104866 274644
rect 157610 274632 157616 274644
rect 104860 274604 157616 274632
rect 104860 274592 104866 274604
rect 157610 274592 157616 274604
rect 157668 274592 157674 274644
rect 195882 274592 195888 274644
rect 195940 274632 195946 274644
rect 206278 274632 206284 274644
rect 195940 274604 206284 274632
rect 195940 274592 195946 274604
rect 206278 274592 206284 274604
rect 206336 274592 206342 274644
rect 212552 274564 212580 274672
rect 238478 274660 238484 274712
rect 238536 274700 238542 274712
rect 239766 274700 239772 274712
rect 238536 274672 239772 274700
rect 238536 274660 238542 274672
rect 239766 274660 239772 274672
rect 239824 274660 239830 274712
rect 244366 274660 244372 274712
rect 244424 274700 244430 274712
rect 251082 274700 251088 274712
rect 244424 274672 251088 274700
rect 244424 274660 244430 274672
rect 251082 274660 251088 274672
rect 251140 274660 251146 274712
rect 270402 274660 270408 274712
rect 270460 274700 270466 274712
rect 271138 274700 271144 274712
rect 270460 274672 271144 274700
rect 270460 274660 270466 274672
rect 271138 274660 271144 274672
rect 271196 274660 271202 274712
rect 285766 274660 285772 274712
rect 285824 274700 285830 274712
rect 286962 274700 286968 274712
rect 285824 274672 286968 274700
rect 285824 274660 285830 274672
rect 286962 274660 286968 274672
rect 287020 274660 287026 274712
rect 292850 274660 292856 274712
rect 292908 274700 292914 274712
rect 293862 274700 293868 274712
rect 292908 274672 293868 274700
rect 292908 274660 292914 274672
rect 293862 274660 293868 274672
rect 293920 274660 293926 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 298738 274660 298744 274712
rect 298796 274700 298802 274712
rect 300118 274700 300124 274712
rect 298796 274672 300124 274700
rect 298796 274660 298802 274672
rect 300118 274660 300124 274672
rect 300176 274660 300182 274712
rect 321370 274660 321376 274712
rect 321428 274700 321434 274712
rect 328270 274700 328276 274712
rect 321428 274672 328276 274700
rect 321428 274660 321434 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 331398 274660 331404 274712
rect 331456 274700 331462 274712
rect 335354 274700 335360 274712
rect 331456 274672 335360 274700
rect 331456 274660 331462 274672
rect 335354 274660 335360 274672
rect 335412 274660 335418 274712
rect 360286 274660 360292 274712
rect 360344 274700 360350 274712
rect 363782 274700 363788 274712
rect 360344 274672 363788 274700
rect 360344 274660 360350 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 367094 274660 367100 274712
rect 367152 274700 367158 274712
rect 369670 274700 369676 274712
rect 367152 274672 369676 274700
rect 367152 274660 367158 274672
rect 369670 274660 369676 274672
rect 369728 274660 369734 274712
rect 386046 274660 386052 274712
rect 386104 274700 386110 274712
rect 389726 274700 389732 274712
rect 386104 274672 389732 274700
rect 386104 274660 386110 274672
rect 389726 274660 389732 274672
rect 389784 274660 389790 274712
rect 404262 274660 404268 274712
rect 404320 274700 404326 274712
rect 407482 274700 407488 274712
rect 404320 274672 407488 274700
rect 404320 274660 404326 274672
rect 407482 274660 407488 274672
rect 407540 274660 407546 274712
rect 409138 274660 409144 274712
rect 409196 274700 409202 274712
rect 409874 274700 409880 274712
rect 409196 274672 409880 274700
rect 409196 274660 409202 274672
rect 409874 274660 409880 274672
rect 409932 274660 409938 274712
rect 488534 274660 488540 274712
rect 488592 274700 488598 274712
rect 492214 274700 492220 274712
rect 488592 274672 492220 274700
rect 488592 274660 488598 274672
rect 492214 274660 492220 274672
rect 492272 274660 492278 274712
rect 494054 274660 494060 274712
rect 494112 274700 494118 274712
rect 498562 274700 498568 274712
rect 494112 274672 498568 274700
rect 494112 274660 494118 274672
rect 498562 274660 498568 274672
rect 498620 274660 498626 274712
rect 619542 274660 619548 274712
rect 619600 274700 619606 274712
rect 623866 274700 623872 274712
rect 619600 274672 623872 274700
rect 619600 274660 619606 274672
rect 623866 274660 623872 274672
rect 623924 274660 623930 274712
rect 410242 274592 410248 274644
rect 410300 274632 410306 274644
rect 437474 274632 437480 274644
rect 410300 274604 437480 274632
rect 410300 274592 410306 274604
rect 437474 274592 437480 274604
rect 437532 274592 437538 274644
rect 440878 274592 440884 274644
rect 440936 274632 440942 274644
rect 486694 274632 486700 274644
rect 440936 274604 486700 274632
rect 440936 274592 440942 274604
rect 486694 274592 486700 274604
rect 486752 274592 486758 274644
rect 498746 274592 498752 274644
rect 498804 274632 498810 274644
rect 571794 274632 571800 274644
rect 498804 274604 571800 274632
rect 498804 274592 498810 274604
rect 571794 274592 571800 274604
rect 571852 274592 571858 274644
rect 212552 274536 219434 274564
rect 121362 274456 121368 274508
rect 121420 274496 121426 274508
rect 176746 274496 176752 274508
rect 121420 274468 176752 274496
rect 121420 274456 121426 274468
rect 176746 274456 176752 274468
rect 176804 274456 176810 274508
rect 182910 274456 182916 274508
rect 182968 274496 182974 274508
rect 199654 274496 199660 274508
rect 182968 274468 199660 274496
rect 182968 274456 182974 274468
rect 199654 274456 199660 274468
rect 199712 274456 199718 274508
rect 219406 274496 219434 274536
rect 237834 274496 237840 274508
rect 219406 274468 237840 274496
rect 237834 274456 237840 274468
rect 237892 274456 237898 274508
rect 362862 274456 362868 274508
rect 362920 274496 362926 274508
rect 386230 274496 386236 274508
rect 362920 274468 386236 274496
rect 362920 274456 362926 274468
rect 386230 274456 386236 274468
rect 386288 274456 386294 274508
rect 395890 274456 395896 274508
rect 395948 274496 395954 274508
rect 413094 274496 413100 274508
rect 395948 274468 413100 274496
rect 395948 274456 395954 274468
rect 413094 274456 413100 274468
rect 413152 274456 413158 274508
rect 427078 274456 427084 274508
rect 427136 274496 427142 274508
rect 477218 274496 477224 274508
rect 427136 274468 477224 274496
rect 427136 274456 427142 274468
rect 477218 274456 477224 274468
rect 477276 274456 477282 274508
rect 491478 274496 491484 274508
rect 477512 274468 491484 274496
rect 101306 274320 101312 274372
rect 101364 274360 101370 274372
rect 160922 274360 160928 274372
rect 101364 274332 160928 274360
rect 101364 274320 101370 274332
rect 160922 274320 160928 274332
rect 160980 274320 160986 274372
rect 187786 274320 187792 274372
rect 187844 274360 187850 274372
rect 220906 274360 220912 274372
rect 187844 274332 220912 274360
rect 187844 274320 187850 274332
rect 220906 274320 220912 274332
rect 220964 274320 220970 274372
rect 237374 274320 237380 274372
rect 237432 274360 237438 274372
rect 243722 274360 243728 274372
rect 237432 274332 243728 274360
rect 237432 274320 237438 274332
rect 243722 274320 243728 274332
rect 243780 274320 243786 274372
rect 384942 274320 384948 274372
rect 385000 274360 385006 274372
rect 419350 274360 419356 274372
rect 385000 274332 419356 274360
rect 385000 274320 385006 274332
rect 419350 274320 419356 274332
rect 419408 274320 419414 274372
rect 424962 274320 424968 274372
rect 425020 274360 425026 274372
rect 474918 274360 474924 274372
rect 425020 274332 474924 274360
rect 425020 274320 425026 274332
rect 474918 274320 474924 274332
rect 474976 274320 474982 274372
rect 476574 274320 476580 274372
rect 476632 274360 476638 274372
rect 477512 274360 477540 274468
rect 491478 274456 491484 274468
rect 491536 274456 491542 274508
rect 492306 274456 492312 274508
rect 492364 274496 492370 274508
rect 496354 274496 496360 274508
rect 492364 274468 496360 274496
rect 492364 274456 492370 274468
rect 496354 274456 496360 274468
rect 496412 274456 496418 274508
rect 496630 274456 496636 274508
rect 496688 274496 496694 274508
rect 577774 274496 577780 274508
rect 496688 274468 577780 274496
rect 496688 274456 496694 274468
rect 577774 274456 577780 274468
rect 577832 274456 577838 274508
rect 585778 274456 585784 274508
rect 585836 274496 585842 274508
rect 585836 274468 586514 274496
rect 585836 274456 585842 274468
rect 476632 274332 477540 274360
rect 476632 274320 476638 274332
rect 477678 274320 477684 274372
rect 477736 274360 477742 274372
rect 528508 274360 528514 274372
rect 477736 274332 528514 274360
rect 477736 274320 477742 274332
rect 528508 274320 528514 274332
rect 528566 274320 528572 274372
rect 528646 274320 528652 274372
rect 528704 274360 528710 274372
rect 538122 274360 538128 274372
rect 528704 274332 538128 274360
rect 528704 274320 528710 274332
rect 538122 274320 538128 274332
rect 538180 274320 538186 274372
rect 538306 274320 538312 274372
rect 538364 274360 538370 274372
rect 586054 274360 586060 274372
rect 538364 274332 586060 274360
rect 538364 274320 538370 274332
rect 586054 274320 586060 274332
rect 586112 274320 586118 274372
rect 586486 274360 586514 274468
rect 601418 274360 601424 274372
rect 586486 274332 601424 274360
rect 601418 274320 601424 274332
rect 601476 274320 601482 274372
rect 82354 274184 82360 274236
rect 82412 274224 82418 274236
rect 145558 274224 145564 274236
rect 82412 274196 145564 274224
rect 82412 274184 82418 274196
rect 145558 274184 145564 274196
rect 145616 274184 145622 274236
rect 160094 274184 160100 274236
rect 160152 274224 160158 274236
rect 164234 274224 164240 274236
rect 160152 274196 164240 274224
rect 160152 274184 160158 274196
rect 164234 274184 164240 274196
rect 164292 274184 164298 274236
rect 176930 274184 176936 274236
rect 176988 274224 176994 274236
rect 214650 274224 214656 274236
rect 176988 274196 214656 274224
rect 176988 274184 176994 274196
rect 214650 274184 214656 274196
rect 214708 274184 214714 274236
rect 220538 274184 220544 274236
rect 220596 274224 220602 274236
rect 240594 274224 240600 274236
rect 220596 274196 240600 274224
rect 220596 274184 220602 274196
rect 240594 274184 240600 274196
rect 240652 274184 240658 274236
rect 342898 274184 342904 274236
rect 342956 274224 342962 274236
rect 347222 274224 347228 274236
rect 342956 274196 347228 274224
rect 342956 274184 342962 274196
rect 347222 274184 347228 274196
rect 347280 274184 347286 274236
rect 366910 274184 366916 274236
rect 366968 274224 366974 274236
rect 389174 274224 389180 274236
rect 366968 274196 389180 274224
rect 366968 274184 366974 274196
rect 389174 274184 389180 274196
rect 389232 274184 389238 274236
rect 390278 274184 390284 274236
rect 390336 274224 390342 274236
rect 426434 274224 426440 274236
rect 390336 274196 426440 274224
rect 390336 274184 390342 274196
rect 426434 274184 426440 274196
rect 426492 274184 426498 274236
rect 438762 274184 438768 274236
rect 438820 274224 438826 274236
rect 496170 274224 496176 274236
rect 438820 274196 496176 274224
rect 438820 274184 438826 274196
rect 496170 274184 496176 274196
rect 496228 274184 496234 274236
rect 496354 274184 496360 274236
rect 496412 274224 496418 274236
rect 498746 274224 498752 274236
rect 496412 274196 498752 274224
rect 496412 274184 496418 274196
rect 498746 274184 498752 274196
rect 498804 274184 498810 274236
rect 501966 274184 501972 274236
rect 502024 274224 502030 274236
rect 502024 274196 523724 274224
rect 502024 274184 502030 274196
rect 84746 274048 84752 274100
rect 84804 274088 84810 274100
rect 148318 274088 148324 274100
rect 84804 274060 148324 274088
rect 84804 274048 84810 274060
rect 148318 274048 148324 274060
rect 148376 274048 148382 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 200666 274088 200672 274100
rect 158128 274060 200672 274088
rect 158128 274048 158134 274060
rect 200666 274048 200672 274060
rect 200724 274048 200730 274100
rect 206554 274048 206560 274100
rect 206612 274088 206618 274100
rect 235442 274088 235448 274100
rect 206612 274060 235448 274088
rect 206612 274048 206618 274060
rect 235442 274048 235448 274060
rect 235500 274048 235506 274100
rect 239582 274048 239588 274100
rect 239640 274088 239646 274100
rect 258626 274088 258632 274100
rect 239640 274060 258632 274088
rect 239640 274048 239646 274060
rect 258626 274048 258632 274060
rect 258684 274048 258690 274100
rect 346118 274048 346124 274100
rect 346176 274088 346182 274100
rect 362586 274088 362592 274100
rect 346176 274060 362592 274088
rect 346176 274048 346182 274060
rect 362586 274048 362592 274060
rect 362644 274048 362650 274100
rect 377766 274048 377772 274100
rect 377824 274088 377830 274100
rect 408678 274088 408684 274100
rect 377824 274060 408684 274088
rect 377824 274048 377830 274060
rect 408678 274048 408684 274060
rect 408736 274048 408742 274100
rect 413922 274048 413928 274100
rect 413980 274088 413986 274100
rect 456794 274088 456800 274100
rect 413980 274060 456800 274088
rect 413980 274048 413986 274060
rect 456794 274048 456800 274060
rect 456852 274048 456858 274100
rect 459370 274048 459376 274100
rect 459428 274088 459434 274100
rect 523494 274088 523500 274100
rect 459428 274060 523500 274088
rect 459428 274048 459434 274060
rect 523494 274048 523500 274060
rect 523552 274048 523558 274100
rect 523696 274088 523724 274196
rect 523862 274184 523868 274236
rect 523920 274224 523926 274236
rect 602154 274224 602160 274236
rect 523920 274196 602160 274224
rect 523920 274184 523926 274196
rect 602154 274184 602160 274196
rect 602212 274184 602218 274236
rect 602338 274184 602344 274236
rect 602396 274224 602402 274236
rect 608502 274224 608508 274236
rect 602396 274196 608508 274224
rect 602396 274184 602402 274196
rect 608502 274184 608508 274196
rect 608560 274184 608566 274236
rect 528508 274088 528514 274100
rect 523696 274060 528514 274088
rect 528508 274048 528514 274060
rect 528566 274048 528572 274100
rect 528646 274048 528652 274100
rect 528704 274088 528710 274100
rect 619542 274088 619548 274100
rect 528704 274060 619548 274088
rect 528704 274048 528710 274060
rect 619542 274048 619548 274060
rect 619600 274048 619606 274100
rect 77202 273912 77208 273964
rect 77260 273952 77266 273964
rect 143534 273952 143540 273964
rect 77260 273924 143540 273952
rect 77260 273912 77266 273924
rect 143534 273912 143540 273924
rect 143592 273912 143598 273964
rect 145006 273912 145012 273964
rect 145064 273952 145070 273964
rect 192478 273952 192484 273964
rect 145064 273924 192484 273952
rect 145064 273912 145070 273924
rect 192478 273912 192484 273924
rect 192536 273912 192542 273964
rect 193490 273912 193496 273964
rect 193548 273952 193554 273964
rect 226334 273952 226340 273964
rect 193548 273924 226340 273952
rect 193548 273912 193554 273924
rect 226334 273912 226340 273924
rect 226392 273912 226398 273964
rect 234890 273912 234896 273964
rect 234948 273952 234954 273964
rect 255682 273952 255688 273964
rect 234948 273924 255688 273952
rect 234948 273912 234954 273924
rect 255682 273912 255688 273924
rect 255740 273912 255746 273964
rect 256142 273912 256148 273964
rect 256200 273952 256206 273964
rect 270586 273952 270592 273964
rect 256200 273924 270592 273952
rect 256200 273912 256206 273924
rect 270586 273912 270592 273924
rect 270644 273912 270650 273964
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280798 273952 280804 273964
rect 271564 273924 280804 273952
rect 271564 273912 271570 273924
rect 280798 273912 280804 273924
rect 280856 273912 280862 273964
rect 331030 273912 331036 273964
rect 331088 273952 331094 273964
rect 342438 273952 342444 273964
rect 331088 273924 342444 273952
rect 331088 273912 331094 273924
rect 342438 273912 342444 273924
rect 342496 273912 342502 273964
rect 360102 273912 360108 273964
rect 360160 273952 360166 273964
rect 383838 273952 383844 273964
rect 360160 273924 383844 273952
rect 360160 273912 360166 273924
rect 383838 273912 383844 273924
rect 383896 273912 383902 273964
rect 385494 273912 385500 273964
rect 385552 273952 385558 273964
rect 395706 273952 395712 273964
rect 385552 273924 395712 273952
rect 385552 273912 385558 273924
rect 395706 273912 395712 273924
rect 395764 273912 395770 273964
rect 404998 273912 405004 273964
rect 405056 273952 405062 273964
rect 444190 273952 444196 273964
rect 405056 273924 444196 273952
rect 405056 273912 405062 273924
rect 444190 273912 444196 273924
rect 444248 273912 444254 273964
rect 451182 273912 451188 273964
rect 451240 273952 451246 273964
rect 513926 273952 513932 273964
rect 451240 273924 513932 273952
rect 451240 273912 451246 273924
rect 513926 273912 513932 273924
rect 513984 273912 513990 273964
rect 514110 273912 514116 273964
rect 514168 273952 514174 273964
rect 523862 273952 523868 273964
rect 514168 273924 523868 273952
rect 514168 273912 514174 273924
rect 523862 273912 523868 273924
rect 523920 273912 523926 273964
rect 524046 273912 524052 273964
rect 524104 273952 524110 273964
rect 613194 273952 613200 273964
rect 524104 273924 613200 273952
rect 524104 273912 524110 273924
rect 613194 273912 613200 273924
rect 613252 273912 613258 273964
rect 123754 273776 123760 273828
rect 123812 273816 123818 273828
rect 177482 273816 177488 273828
rect 123812 273788 177488 273816
rect 123812 273776 123818 273788
rect 177482 273776 177488 273788
rect 177540 273776 177546 273828
rect 406838 273776 406844 273828
rect 406896 273816 406902 273828
rect 410242 273816 410248 273828
rect 406896 273788 410248 273816
rect 406896 273776 406902 273788
rect 410242 273776 410248 273788
rect 410300 273776 410306 273828
rect 428458 273776 428464 273828
rect 428516 273816 428522 273828
rect 458358 273816 458364 273828
rect 428516 273788 458364 273816
rect 428516 273776 428522 273788
rect 458358 273776 458364 273788
rect 458416 273776 458422 273828
rect 465718 273776 465724 273828
rect 465776 273816 465782 273828
rect 482002 273816 482008 273828
rect 465776 273788 482008 273816
rect 465776 273776 465782 273788
rect 482002 273776 482008 273788
rect 482060 273776 482066 273828
rect 491202 273776 491208 273828
rect 491260 273816 491266 273828
rect 570690 273816 570696 273828
rect 491260 273788 570696 273816
rect 491260 273776 491266 273788
rect 570690 273776 570696 273788
rect 570748 273776 570754 273828
rect 587158 273816 587164 273828
rect 576826 273788 587164 273816
rect 280982 273708 280988 273760
rect 281040 273748 281046 273760
rect 287514 273748 287520 273760
rect 281040 273720 287520 273748
rect 281040 273708 281046 273720
rect 287514 273708 287520 273720
rect 287572 273708 287578 273760
rect 134426 273640 134432 273692
rect 134484 273680 134490 273692
rect 185026 273680 185032 273692
rect 134484 273652 185032 273680
rect 134484 273640 134490 273652
rect 185026 273640 185032 273652
rect 185084 273640 185090 273692
rect 457438 273640 457444 273692
rect 457496 273680 457502 273692
rect 484302 273680 484308 273692
rect 457496 273652 484308 273680
rect 457496 273640 457502 273652
rect 484302 273640 484308 273652
rect 484360 273640 484366 273692
rect 487062 273640 487068 273692
rect 487120 273680 487126 273692
rect 563514 273680 563520 273692
rect 487120 273652 563520 273680
rect 487120 273640 487126 273652
rect 563514 273640 563520 273652
rect 563572 273640 563578 273692
rect 570598 273640 570604 273692
rect 570656 273680 570662 273692
rect 576826 273680 576854 273788
rect 587158 273776 587164 273788
rect 587216 273776 587222 273828
rect 613378 273708 613384 273760
rect 613436 273748 613442 273760
rect 615586 273748 615592 273760
rect 613436 273720 615592 273748
rect 613436 273708 613442 273720
rect 615586 273708 615592 273720
rect 615644 273708 615650 273760
rect 570656 273652 576854 273680
rect 570656 273640 570662 273652
rect 144638 273504 144644 273556
rect 144696 273544 144702 273556
rect 187786 273544 187792 273556
rect 144696 273516 187792 273544
rect 144696 273504 144702 273516
rect 187786 273504 187792 273516
rect 187844 273504 187850 273556
rect 475562 273504 475568 273556
rect 475620 273544 475626 273556
rect 477678 273544 477684 273556
rect 475620 273516 477684 273544
rect 475620 273504 475626 273516
rect 477678 273504 477684 273516
rect 477736 273504 477742 273556
rect 482462 273504 482468 273556
rect 482520 273544 482526 273556
rect 558822 273544 558828 273556
rect 482520 273516 558828 273544
rect 482520 273504 482526 273516
rect 558822 273504 558828 273516
rect 558880 273504 558886 273556
rect 481358 273368 481364 273420
rect 481416 273408 481422 273420
rect 556430 273408 556436 273420
rect 481416 273380 556436 273408
rect 481416 273368 481422 273380
rect 556430 273368 556436 273380
rect 556488 273368 556494 273420
rect 347038 273232 347044 273284
rect 347096 273272 347102 273284
rect 349614 273272 349620 273284
rect 347096 273244 349620 273272
rect 347096 273232 347102 273244
rect 349614 273232 349620 273244
rect 349672 273232 349678 273284
rect 350258 273232 350264 273284
rect 350316 273272 350322 273284
rect 356330 273272 356336 273284
rect 350316 273244 356336 273272
rect 350316 273232 350322 273244
rect 356330 273232 356336 273244
rect 356388 273232 356394 273284
rect 114278 273164 114284 273216
rect 114336 273204 114342 273216
rect 169018 273204 169024 273216
rect 114336 273176 169024 273204
rect 114336 273164 114342 273176
rect 169018 273164 169024 273176
rect 169076 273164 169082 273216
rect 211798 273204 211804 273216
rect 200086 273176 211804 273204
rect 104986 273028 104992 273080
rect 105044 273068 105050 273080
rect 163314 273068 163320 273080
rect 105044 273040 163320 273068
rect 105044 273028 105050 273040
rect 163314 273028 163320 273040
rect 163372 273028 163378 273080
rect 167546 273028 167552 273080
rect 167604 273068 167610 273080
rect 184198 273068 184204 273080
rect 167604 273040 184204 273068
rect 167604 273028 167610 273040
rect 184198 273028 184204 273040
rect 184256 273028 184262 273080
rect 187602 273028 187608 273080
rect 187660 273068 187666 273080
rect 200086 273068 200114 273176
rect 211798 273164 211804 273176
rect 211856 273164 211862 273216
rect 419166 273164 419172 273216
rect 419224 273204 419230 273216
rect 462958 273204 462964 273216
rect 419224 273176 462964 273204
rect 419224 273164 419230 273176
rect 462958 273164 462964 273176
rect 463016 273164 463022 273216
rect 473446 273164 473452 273216
rect 473504 273204 473510 273216
rect 496814 273204 496820 273216
rect 473504 273176 496820 273204
rect 473504 273164 473510 273176
rect 496814 273164 496820 273176
rect 496872 273164 496878 273216
rect 500954 273164 500960 273216
rect 501012 273204 501018 273216
rect 581270 273204 581276 273216
rect 501012 273176 581276 273204
rect 501012 273164 501018 273176
rect 581270 273164 581276 273176
rect 581328 273164 581334 273216
rect 187660 273040 200114 273068
rect 187660 273028 187666 273040
rect 211246 273028 211252 273080
rect 211304 273068 211310 273080
rect 220078 273068 220084 273080
rect 211304 273040 220084 273068
rect 211304 273028 211310 273040
rect 220078 273028 220084 273040
rect 220136 273028 220142 273080
rect 397270 273028 397276 273080
rect 397328 273068 397334 273080
rect 418338 273068 418344 273080
rect 397328 273040 418344 273068
rect 397328 273028 397334 273040
rect 418338 273028 418344 273040
rect 418396 273028 418402 273080
rect 426342 273028 426348 273080
rect 426400 273068 426406 273080
rect 478414 273068 478420 273080
rect 426400 273040 478420 273068
rect 426400 273028 426406 273040
rect 478414 273028 478420 273040
rect 478472 273028 478478 273080
rect 485038 273028 485044 273080
rect 485096 273068 485102 273080
rect 492490 273068 492496 273080
rect 485096 273040 492496 273068
rect 485096 273028 485102 273040
rect 492490 273028 492496 273040
rect 492548 273028 492554 273080
rect 493594 273028 493600 273080
rect 493652 273068 493658 273080
rect 574186 273068 574192 273080
rect 493652 273040 574192 273068
rect 493652 273028 493658 273040
rect 574186 273028 574192 273040
rect 574244 273028 574250 273080
rect 580258 273028 580264 273080
rect 580316 273068 580322 273080
rect 640426 273068 640432 273080
rect 580316 273040 640432 273068
rect 580316 273028 580322 273040
rect 640426 273028 640432 273040
rect 640484 273028 640490 273080
rect 78858 272892 78864 272944
rect 78916 272932 78922 272944
rect 138658 272932 138664 272944
rect 78916 272904 138664 272932
rect 78916 272892 78922 272904
rect 138658 272892 138664 272904
rect 138716 272892 138722 272944
rect 141786 272892 141792 272944
rect 141844 272932 141850 272944
rect 189810 272932 189816 272944
rect 141844 272904 189816 272932
rect 141844 272892 141850 272904
rect 189810 272892 189816 272904
rect 189868 272892 189874 272944
rect 191190 272892 191196 272944
rect 191248 272932 191254 272944
rect 224862 272932 224868 272944
rect 191248 272904 224868 272932
rect 191248 272892 191254 272904
rect 224862 272892 224868 272904
rect 224920 272892 224926 272944
rect 288066 272892 288072 272944
rect 288124 272932 288130 272944
rect 290458 272932 290464 272944
rect 288124 272904 290464 272932
rect 288124 272892 288130 272904
rect 290458 272892 290464 272904
rect 290516 272892 290522 272944
rect 373166 272892 373172 272944
rect 373224 272932 373230 272944
rect 382642 272932 382648 272944
rect 373224 272904 382648 272932
rect 373224 272892 373230 272904
rect 382642 272892 382648 272904
rect 382700 272892 382706 272944
rect 391750 272892 391756 272944
rect 391808 272932 391814 272944
rect 410058 272932 410064 272944
rect 391808 272904 410064 272932
rect 391808 272892 391814 272904
rect 410058 272892 410064 272904
rect 410116 272892 410122 272944
rect 412450 272892 412456 272944
rect 412508 272932 412514 272944
rect 453390 272932 453396 272944
rect 412508 272904 453396 272932
rect 412508 272892 412514 272904
rect 453390 272892 453396 272904
rect 453448 272892 453454 272944
rect 458082 272892 458088 272944
rect 458140 272932 458146 272944
rect 521838 272932 521844 272944
rect 458140 272904 521844 272932
rect 458140 272892 458146 272904
rect 521838 272892 521844 272904
rect 521896 272892 521902 272944
rect 528508 272932 528514 272944
rect 523604 272904 528514 272932
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 156046 272796 156052 272808
rect 94280 272768 156052 272796
rect 94280 272756 94286 272768
rect 156046 272756 156052 272768
rect 156104 272756 156110 272808
rect 180518 272756 180524 272808
rect 180576 272796 180582 272808
rect 217226 272796 217232 272808
rect 180576 272768 217232 272796
rect 180576 272756 180582 272768
rect 217226 272756 217232 272768
rect 217284 272756 217290 272808
rect 228818 272756 228824 272808
rect 228876 272796 228882 272808
rect 249058 272796 249064 272808
rect 228876 272768 249064 272796
rect 228876 272756 228882 272768
rect 249058 272756 249064 272768
rect 249116 272756 249122 272808
rect 352926 272756 352932 272808
rect 352984 272796 352990 272808
rect 372982 272796 372988 272808
rect 352984 272768 372988 272796
rect 352984 272756 352990 272768
rect 372982 272756 372988 272768
rect 373040 272756 373046 272808
rect 380710 272756 380716 272808
rect 380768 272796 380774 272808
rect 396350 272796 396356 272808
rect 380768 272768 396356 272796
rect 380768 272756 380774 272768
rect 396350 272756 396356 272768
rect 396408 272756 396414 272808
rect 403986 272756 403992 272808
rect 404044 272796 404050 272808
rect 429194 272796 429200 272808
rect 404044 272768 429200 272796
rect 404044 272756 404050 272768
rect 429194 272756 429200 272768
rect 429252 272756 429258 272808
rect 434622 272756 434628 272808
rect 434680 272796 434686 272808
rect 488718 272796 488724 272808
rect 434680 272768 488724 272796
rect 434680 272756 434686 272768
rect 488718 272756 488724 272768
rect 488776 272756 488782 272808
rect 496262 272756 496268 272808
rect 496320 272796 496326 272808
rect 523604 272796 523632 272904
rect 528508 272892 528514 272904
rect 528566 272892 528572 272944
rect 528646 272892 528652 272944
rect 528704 272932 528710 272944
rect 611354 272932 611360 272944
rect 528704 272904 611360 272932
rect 528704 272892 528710 272904
rect 611354 272892 611360 272904
rect 611412 272892 611418 272944
rect 606110 272796 606116 272808
rect 496320 272768 523632 272796
rect 523696 272768 606116 272796
rect 496320 272756 496326 272768
rect 87138 272620 87144 272672
rect 87196 272660 87202 272672
rect 151998 272660 152004 272672
rect 87196 272632 152004 272660
rect 87196 272620 87202 272632
rect 151998 272620 152004 272632
rect 152056 272620 152062 272672
rect 168650 272620 168656 272672
rect 168708 272660 168714 272672
rect 208486 272660 208492 272672
rect 168708 272632 208492 272660
rect 168708 272620 168714 272632
rect 208486 272620 208492 272632
rect 208544 272620 208550 272672
rect 217410 272620 217416 272672
rect 217468 272660 217474 272672
rect 242158 272660 242164 272672
rect 217468 272632 242164 272660
rect 217468 272620 217474 272632
rect 242158 272620 242164 272632
rect 242216 272620 242222 272672
rect 242342 272620 242348 272672
rect 242400 272660 242406 272672
rect 259546 272660 259552 272672
rect 242400 272632 259552 272660
rect 242400 272620 242406 272632
rect 259546 272620 259552 272632
rect 259604 272620 259610 272672
rect 333606 272620 333612 272672
rect 333664 272660 333670 272672
rect 344830 272660 344836 272672
rect 333664 272632 344836 272660
rect 333664 272620 333670 272632
rect 344830 272620 344836 272632
rect 344888 272620 344894 272672
rect 368382 272620 368388 272672
rect 368440 272660 368446 272672
rect 393774 272660 393780 272672
rect 368440 272632 393780 272660
rect 368440 272620 368446 272632
rect 393774 272620 393780 272632
rect 393832 272620 393838 272672
rect 393958 272620 393964 272672
rect 394016 272660 394022 272672
rect 406286 272660 406292 272672
rect 394016 272632 406292 272660
rect 394016 272620 394022 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 408402 272620 408408 272672
rect 408460 272660 408466 272672
rect 452470 272660 452476 272672
rect 408460 272632 452476 272660
rect 408460 272620 408466 272632
rect 452470 272620 452476 272632
rect 452528 272620 452534 272672
rect 453850 272620 453856 272672
rect 453908 272660 453914 272672
rect 516410 272660 516416 272672
rect 453908 272632 516416 272660
rect 453908 272620 453914 272632
rect 516410 272620 516416 272632
rect 516468 272620 516474 272672
rect 516594 272620 516600 272672
rect 516652 272660 516658 272672
rect 523696 272660 523724 272768
rect 606110 272756 606116 272768
rect 606168 272756 606174 272808
rect 516652 272632 523724 272660
rect 516652 272620 516658 272632
rect 524322 272620 524328 272672
rect 524380 272660 524386 272672
rect 527910 272660 527916 272672
rect 524380 272632 527916 272660
rect 524380 272620 524386 272632
rect 527910 272620 527916 272632
rect 527968 272620 527974 272672
rect 528370 272620 528376 272672
rect 528428 272660 528434 272672
rect 614390 272660 614396 272672
rect 528428 272632 614396 272660
rect 528428 272620 528434 272632
rect 614390 272620 614396 272632
rect 614448 272620 614454 272672
rect 77662 272484 77668 272536
rect 77720 272524 77726 272536
rect 145098 272524 145104 272536
rect 77720 272496 145104 272524
rect 77720 272484 77726 272496
rect 145098 272484 145104 272496
rect 145156 272484 145162 272536
rect 152182 272484 152188 272536
rect 152240 272524 152246 272536
rect 197538 272524 197544 272536
rect 152240 272496 197544 272524
rect 152240 272484 152246 272496
rect 197538 272484 197544 272496
rect 197596 272484 197602 272536
rect 199470 272484 199476 272536
rect 199528 272524 199534 272536
rect 230566 272524 230572 272536
rect 199528 272496 230572 272524
rect 199528 272484 199534 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 252738 272524 252744 272536
rect 231452 272496 252744 272524
rect 231452 272484 231458 272496
rect 252738 272484 252744 272496
rect 252796 272484 252802 272536
rect 252922 272484 252928 272536
rect 252980 272524 252986 272536
rect 267826 272524 267832 272536
rect 252980 272496 267832 272524
rect 252980 272484 252986 272496
rect 267826 272484 267832 272496
rect 267884 272484 267890 272536
rect 268010 272484 268016 272536
rect 268068 272524 268074 272536
rect 278774 272524 278780 272536
rect 268068 272496 278780 272524
rect 268068 272484 268074 272496
rect 278774 272484 278780 272496
rect 278832 272484 278838 272536
rect 279786 272484 279792 272536
rect 279844 272524 279850 272536
rect 287146 272524 287152 272536
rect 279844 272496 287152 272524
rect 279844 272484 279850 272496
rect 287146 272484 287152 272496
rect 287204 272484 287210 272536
rect 322566 272484 322572 272536
rect 322624 272524 322630 272536
rect 330662 272524 330668 272536
rect 322624 272496 330668 272524
rect 322624 272484 322630 272496
rect 330662 272484 330668 272496
rect 330720 272484 330726 272536
rect 338022 272484 338028 272536
rect 338080 272524 338086 272536
rect 351914 272524 351920 272536
rect 338080 272496 351920 272524
rect 338080 272484 338086 272496
rect 351914 272484 351920 272496
rect 351972 272484 351978 272536
rect 358630 272484 358636 272536
rect 358688 272524 358694 272536
rect 380342 272524 380348 272536
rect 358688 272496 380348 272524
rect 358688 272484 358694 272496
rect 380342 272484 380348 272496
rect 380400 272484 380406 272536
rect 382918 272484 382924 272536
rect 382976 272524 382982 272536
rect 413370 272524 413376 272536
rect 382976 272496 413376 272524
rect 382976 272484 382982 272496
rect 413370 272484 413376 272496
rect 413428 272484 413434 272536
rect 415118 272484 415124 272536
rect 415176 272524 415182 272536
rect 461854 272524 461860 272536
rect 415176 272496 461860 272524
rect 415176 272484 415182 272496
rect 461854 272484 461860 272496
rect 461912 272484 461918 272536
rect 463510 272484 463516 272536
rect 463568 272524 463574 272536
rect 528554 272524 528560 272536
rect 463568 272496 528560 272524
rect 463568 272484 463574 272496
rect 528554 272484 528560 272496
rect 528612 272484 528618 272536
rect 529014 272484 529020 272536
rect 529072 272524 529078 272536
rect 538122 272524 538128 272536
rect 529072 272496 538128 272524
rect 529072 272484 529078 272496
rect 538122 272484 538128 272496
rect 538180 272484 538186 272536
rect 538306 272484 538312 272536
rect 538364 272524 538370 272536
rect 632146 272524 632152 272536
rect 538364 272496 632152 272524
rect 538364 272484 538370 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 127342 272348 127348 272400
rect 127400 272388 127406 272400
rect 179874 272388 179880 272400
rect 127400 272360 179880 272388
rect 127400 272348 127406 272360
rect 179874 272348 179880 272360
rect 179932 272348 179938 272400
rect 451734 272348 451740 272400
rect 451792 272388 451798 272400
rect 451792 272360 471284 272388
rect 451792 272348 451798 272360
rect 139118 272212 139124 272264
rect 139176 272252 139182 272264
rect 141602 272252 141608 272264
rect 139176 272224 141608 272252
rect 139176 272212 139182 272224
rect 141602 272212 141608 272224
rect 141660 272212 141666 272264
rect 143902 272212 143908 272264
rect 143960 272252 143966 272264
rect 190730 272252 190736 272264
rect 143960 272224 190736 272252
rect 143960 272212 143966 272224
rect 190730 272212 190736 272224
rect 190788 272212 190794 272264
rect 447594 272212 447600 272264
rect 447652 272252 447658 272264
rect 470042 272252 470048 272264
rect 447652 272224 470048 272252
rect 447652 272212 447658 272224
rect 470042 272212 470048 272224
rect 470100 272212 470106 272264
rect 471256 272252 471284 272360
rect 471422 272348 471428 272400
rect 471480 272388 471486 272400
rect 485038 272388 485044 272400
rect 471480 272360 485044 272388
rect 471480 272348 471486 272360
rect 485038 272348 485044 272360
rect 485096 272348 485102 272400
rect 488350 272348 488356 272400
rect 488408 272388 488414 272400
rect 567102 272388 567108 272400
rect 488408 272360 567108 272388
rect 488408 272348 488414 272360
rect 567102 272348 567108 272360
rect 567160 272348 567166 272400
rect 578878 272348 578884 272400
rect 578936 272388 578942 272400
rect 594334 272388 594340 272400
rect 578936 272360 594340 272388
rect 578936 272348 578942 272360
rect 594334 272348 594340 272360
rect 594392 272348 594398 272400
rect 471256 272224 480254 272252
rect 153286 272076 153292 272128
rect 153344 272116 153350 272128
rect 171778 272116 171784 272128
rect 153344 272088 171784 272116
rect 153344 272076 153350 272088
rect 171778 272076 171784 272088
rect 171836 272076 171842 272128
rect 463142 272076 463148 272128
rect 463200 272116 463206 272128
rect 471422 272116 471428 272128
rect 463200 272088 471428 272116
rect 463200 272076 463206 272088
rect 471422 272076 471428 272088
rect 471480 272076 471486 272128
rect 480226 272116 480254 272224
rect 487982 272212 487988 272264
rect 488040 272252 488046 272264
rect 565906 272252 565912 272264
rect 488040 272224 565912 272252
rect 488040 272212 488046 272224
rect 565906 272212 565912 272224
rect 565964 272212 565970 272264
rect 480806 272116 480812 272128
rect 480226 272088 480812 272116
rect 480806 272076 480812 272088
rect 480864 272076 480870 272128
rect 483750 272076 483756 272128
rect 483808 272116 483814 272128
rect 560018 272116 560024 272128
rect 483808 272088 560024 272116
rect 483808 272076 483814 272088
rect 560018 272076 560024 272088
rect 560076 272076 560082 272128
rect 470042 271940 470048 271992
rect 470100 271980 470106 271992
rect 473722 271980 473728 271992
rect 470100 271952 473728 271980
rect 470100 271940 470106 271952
rect 473722 271940 473728 271952
rect 473780 271940 473786 271992
rect 478690 271940 478696 271992
rect 478748 271980 478754 271992
rect 552474 271980 552480 271992
rect 478748 271952 552480 271980
rect 478748 271940 478754 271952
rect 552474 271940 552480 271952
rect 552532 271940 552538 271992
rect 552658 271940 552664 271992
rect 552716 271980 552722 271992
rect 580074 271980 580080 271992
rect 552716 271952 580080 271980
rect 552716 271940 552722 271952
rect 580074 271940 580080 271952
rect 580132 271940 580138 271992
rect 110414 271804 110420 271856
rect 110472 271844 110478 271856
rect 164970 271844 164976 271856
rect 110472 271816 164976 271844
rect 110472 271804 110478 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 175826 271804 175832 271856
rect 175884 271844 175890 271856
rect 207658 271844 207664 271856
rect 175884 271816 207664 271844
rect 175884 271804 175890 271816
rect 207658 271804 207664 271816
rect 207716 271804 207722 271856
rect 214834 271804 214840 271856
rect 214892 271844 214898 271856
rect 221458 271844 221464 271856
rect 214892 271816 221464 271844
rect 214892 271804 214898 271816
rect 221458 271804 221464 271816
rect 221516 271804 221522 271856
rect 222102 271804 222108 271856
rect 222160 271844 222166 271856
rect 232130 271844 232136 271856
rect 222160 271816 232136 271844
rect 222160 271804 222166 271816
rect 232130 271804 232136 271816
rect 232188 271804 232194 271856
rect 381354 271804 381360 271856
rect 381412 271844 381418 271856
rect 399202 271844 399208 271856
rect 381412 271816 399208 271844
rect 381412 271804 381418 271816
rect 399202 271804 399208 271816
rect 399260 271804 399266 271856
rect 411898 271804 411904 271856
rect 411956 271844 411962 271856
rect 438210 271844 438216 271856
rect 411956 271816 438216 271844
rect 411956 271804 411962 271816
rect 438210 271804 438216 271816
rect 438268 271804 438274 271856
rect 443638 271804 443644 271856
rect 443696 271844 443702 271856
rect 500494 271844 500500 271856
rect 443696 271816 500500 271844
rect 443696 271804 443702 271816
rect 500494 271804 500500 271816
rect 500552 271804 500558 271856
rect 500678 271804 500684 271856
rect 500736 271844 500742 271856
rect 508038 271844 508044 271856
rect 500736 271816 508044 271844
rect 500736 271804 500742 271816
rect 508038 271804 508044 271816
rect 508096 271804 508102 271856
rect 508958 271804 508964 271856
rect 509016 271844 509022 271856
rect 596634 271844 596640 271856
rect 509016 271816 596640 271844
rect 509016 271804 509022 271816
rect 596634 271804 596640 271816
rect 596692 271804 596698 271856
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 93026 271668 93032 271720
rect 93084 271708 93090 271720
rect 120718 271708 120724 271720
rect 93084 271680 120724 271708
rect 93084 271668 93090 271680
rect 120718 271668 120724 271680
rect 120776 271668 120782 271720
rect 120902 271668 120908 271720
rect 120960 271708 120966 271720
rect 175274 271708 175280 271720
rect 120960 271680 175280 271708
rect 120960 271668 120966 271680
rect 175274 271668 175280 271680
rect 175332 271668 175338 271720
rect 192294 271668 192300 271720
rect 192352 271708 192358 271720
rect 225506 271708 225512 271720
rect 192352 271680 225512 271708
rect 192352 271668 192358 271680
rect 225506 271668 225512 271680
rect 225564 271668 225570 271720
rect 372522 271668 372528 271720
rect 372580 271708 372586 271720
rect 400398 271708 400404 271720
rect 372580 271680 400404 271708
rect 372580 271668 372586 271680
rect 400398 271668 400404 271680
rect 400456 271668 400462 271720
rect 401318 271668 401324 271720
rect 401376 271708 401382 271720
rect 427814 271708 427820 271720
rect 401376 271680 427820 271708
rect 401376 271668 401382 271680
rect 427814 271668 427820 271680
rect 427872 271668 427878 271720
rect 453298 271668 453304 271720
rect 453356 271708 453362 271720
rect 511534 271708 511540 271720
rect 453356 271680 511540 271708
rect 453356 271668 453362 271680
rect 511534 271668 511540 271680
rect 511592 271668 511598 271720
rect 511902 271668 511908 271720
rect 511960 271708 511966 271720
rect 600222 271708 600228 271720
rect 511960 271680 600228 271708
rect 511960 271668 511966 271680
rect 600222 271668 600228 271680
rect 600280 271668 600286 271720
rect 111978 271532 111984 271584
rect 112036 271572 112042 271584
rect 168374 271572 168380 271584
rect 112036 271544 168380 271572
rect 112036 271532 112042 271544
rect 168374 271532 168380 271544
rect 168432 271532 168438 271584
rect 173434 271532 173440 271584
rect 173492 271572 173498 271584
rect 212626 271572 212632 271584
rect 173492 271544 212632 271572
rect 173492 271532 173498 271544
rect 212626 271532 212632 271544
rect 212684 271532 212690 271584
rect 226150 271532 226156 271584
rect 226208 271572 226214 271584
rect 247218 271572 247224 271584
rect 226208 271544 247224 271572
rect 226208 271532 226214 271544
rect 247218 271532 247224 271544
rect 247276 271532 247282 271584
rect 259730 271532 259736 271584
rect 259788 271572 259794 271584
rect 268378 271572 268384 271584
rect 259788 271544 268384 271572
rect 259788 271532 259794 271544
rect 268378 271532 268384 271544
rect 268436 271532 268442 271584
rect 362218 271532 362224 271584
rect 362276 271572 362282 271584
rect 381170 271572 381176 271584
rect 362276 271544 381176 271572
rect 362276 271532 362282 271544
rect 381170 271532 381176 271544
rect 381228 271532 381234 271584
rect 394326 271532 394332 271584
rect 394384 271572 394390 271584
rect 425330 271572 425336 271584
rect 394384 271544 425336 271572
rect 394384 271532 394390 271544
rect 425330 271532 425336 271544
rect 425388 271532 425394 271584
rect 443362 271572 443368 271584
rect 431926 271544 443368 271572
rect 89714 271396 89720 271448
rect 89772 271436 89778 271448
rect 152642 271436 152648 271448
rect 89772 271408 152648 271436
rect 89772 271396 89778 271408
rect 152642 271396 152648 271408
rect 152700 271396 152706 271448
rect 165154 271396 165160 271448
rect 165212 271436 165218 271448
rect 205726 271436 205732 271448
rect 165212 271408 205732 271436
rect 165212 271396 165218 271408
rect 205726 271396 205732 271408
rect 205784 271396 205790 271448
rect 223574 271396 223580 271448
rect 223632 271436 223638 271448
rect 247402 271436 247408 271448
rect 223632 271408 247408 271436
rect 223632 271396 223638 271408
rect 247402 271396 247408 271408
rect 247460 271396 247466 271448
rect 247862 271396 247868 271448
rect 247920 271436 247926 271448
rect 264330 271436 264336 271448
rect 247920 271408 264336 271436
rect 247920 271396 247926 271408
rect 264330 271396 264336 271408
rect 264388 271396 264394 271448
rect 275094 271396 275100 271448
rect 275152 271436 275158 271448
rect 283466 271436 283472 271448
rect 275152 271408 283472 271436
rect 275152 271396 275158 271408
rect 283466 271396 283472 271408
rect 283524 271396 283530 271448
rect 340598 271396 340604 271448
rect 340656 271436 340662 271448
rect 355134 271436 355140 271448
rect 340656 271408 355140 271436
rect 340656 271396 340662 271408
rect 355134 271396 355140 271408
rect 355192 271396 355198 271448
rect 355318 271396 355324 271448
rect 355376 271436 355382 271448
rect 374362 271436 374368 271448
rect 355376 271408 374368 271436
rect 355376 271396 355382 271408
rect 374362 271396 374368 271408
rect 374420 271396 374426 271448
rect 379422 271396 379428 271448
rect 379480 271436 379486 271448
rect 407114 271436 407120 271448
rect 379480 271408 407120 271436
rect 379480 271396 379486 271408
rect 407114 271396 407120 271408
rect 407172 271396 407178 271448
rect 409782 271396 409788 271448
rect 409840 271436 409846 271448
rect 431926 271436 431954 271544
rect 443362 271532 443368 271544
rect 443420 271532 443426 271584
rect 445662 271532 445668 271584
rect 445720 271572 445726 271584
rect 504542 271572 504548 271584
rect 445720 271544 504548 271572
rect 445720 271532 445726 271544
rect 504542 271532 504548 271544
rect 504600 271532 504606 271584
rect 504726 271532 504732 271584
rect 504784 271572 504790 271584
rect 589366 271572 589372 271584
rect 504784 271544 589372 271572
rect 504784 271532 504790 271544
rect 589366 271532 589372 271544
rect 589424 271532 589430 271584
rect 591298 271532 591304 271584
rect 591356 271572 591362 271584
rect 603718 271572 603724 271584
rect 591356 271544 603724 271572
rect 591356 271532 591362 271544
rect 603718 271532 603724 271544
rect 603776 271532 603782 271584
rect 607858 271532 607864 271584
rect 607916 271572 607922 271584
rect 643922 271572 643928 271584
rect 607916 271544 643928 271572
rect 607916 271532 607922 271544
rect 643922 271532 643928 271544
rect 643980 271532 643986 271584
rect 409840 271408 431954 271436
rect 409840 271396 409846 271408
rect 435358 271396 435364 271448
rect 435416 271436 435422 271448
rect 454494 271436 454500 271448
rect 435416 271408 454500 271436
rect 435416 271396 435422 271408
rect 454494 271396 454500 271408
rect 454552 271396 454558 271448
rect 454678 271396 454684 271448
rect 454736 271436 454742 271448
rect 515122 271436 515128 271448
rect 454736 271408 515128 271436
rect 454736 271396 454742 271408
rect 515122 271396 515128 271408
rect 515180 271396 515186 271448
rect 517330 271396 517336 271448
rect 517388 271436 517394 271448
rect 604454 271436 604460 271448
rect 517388 271408 604460 271436
rect 517388 271396 517394 271408
rect 604454 271396 604460 271408
rect 604512 271396 604518 271448
rect 68186 271260 68192 271312
rect 68244 271300 68250 271312
rect 138474 271300 138480 271312
rect 68244 271272 138480 271300
rect 68244 271260 68250 271272
rect 138474 271260 138480 271272
rect 138532 271260 138538 271312
rect 150986 271260 150992 271312
rect 151044 271300 151050 271312
rect 195974 271300 195980 271312
rect 151044 271272 195980 271300
rect 151044 271260 151050 271272
rect 195974 271260 195980 271272
rect 196032 271260 196038 271312
rect 215938 271260 215944 271312
rect 215996 271300 216002 271312
rect 242066 271300 242072 271312
rect 215996 271272 242072 271300
rect 215996 271260 216002 271272
rect 242066 271260 242072 271272
rect 242124 271260 242130 271312
rect 243170 271260 243176 271312
rect 243228 271300 243234 271312
rect 261018 271300 261024 271312
rect 243228 271272 261024 271300
rect 243228 271260 243234 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 266814 271260 266820 271312
rect 266872 271300 266878 271312
rect 276658 271300 276664 271312
rect 266872 271272 276664 271300
rect 266872 271260 266878 271272
rect 276658 271260 276664 271272
rect 276716 271260 276722 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 325510 271260 325516 271312
rect 325568 271300 325574 271312
rect 334158 271300 334164 271312
rect 325568 271272 334164 271300
rect 325568 271260 325574 271272
rect 334158 271260 334164 271272
rect 334216 271260 334222 271312
rect 334802 271260 334808 271312
rect 334860 271300 334866 271312
rect 341334 271300 341340 271312
rect 334860 271272 341340 271300
rect 334860 271260 334866 271272
rect 341334 271260 341340 271272
rect 341392 271260 341398 271312
rect 344646 271260 344652 271312
rect 344704 271300 344710 271312
rect 350718 271300 350724 271312
rect 344704 271272 350724 271300
rect 344704 271260 344710 271272
rect 350718 271260 350724 271272
rect 350776 271260 350782 271312
rect 351822 271260 351828 271312
rect 351880 271300 351886 271312
rect 372062 271300 372068 271312
rect 351880 271272 372068 271300
rect 351880 271260 351886 271272
rect 372062 271260 372068 271272
rect 372120 271260 372126 271312
rect 387702 271260 387708 271312
rect 387760 271300 387766 271312
rect 421650 271300 421656 271312
rect 387760 271272 421656 271300
rect 387760 271260 387766 271272
rect 421650 271260 421656 271272
rect 421708 271260 421714 271312
rect 422110 271260 422116 271312
rect 422168 271300 422174 271312
rect 445938 271300 445944 271312
rect 422168 271272 445944 271300
rect 422168 271260 422174 271272
rect 445938 271260 445944 271272
rect 445996 271260 446002 271312
rect 461578 271260 461584 271312
rect 461636 271300 461642 271312
rect 514294 271300 514300 271312
rect 461636 271272 514300 271300
rect 461636 271260 461642 271272
rect 514294 271260 514300 271272
rect 514352 271260 514358 271312
rect 514478 271260 514484 271312
rect 514536 271300 514542 271312
rect 514536 271272 523724 271300
rect 514536 271260 514542 271272
rect 72970 271124 72976 271176
rect 73028 271164 73034 271176
rect 142154 271164 142160 271176
rect 73028 271136 142160 271164
rect 73028 271124 73034 271136
rect 142154 271124 142160 271136
rect 142212 271124 142218 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 208854 271124 208860 271176
rect 208912 271164 208918 271176
rect 237466 271164 237472 271176
rect 208912 271136 237472 271164
rect 208912 271124 208918 271136
rect 237466 271124 237472 271136
rect 237524 271124 237530 271176
rect 240778 271124 240784 271176
rect 240836 271164 240842 271176
rect 259822 271164 259828 271176
rect 240836 271136 259828 271164
rect 240836 271124 240842 271136
rect 259822 271124 259828 271136
rect 259880 271124 259886 271176
rect 262122 271124 262128 271176
rect 262180 271164 262186 271176
rect 274634 271164 274640 271176
rect 262180 271136 274640 271164
rect 262180 271124 262186 271136
rect 274634 271124 274640 271136
rect 274692 271124 274698 271176
rect 276290 271124 276296 271176
rect 276348 271164 276354 271176
rect 284478 271164 284484 271176
rect 276348 271136 284484 271164
rect 276348 271124 276354 271136
rect 284478 271124 284484 271136
rect 284536 271124 284542 271176
rect 328086 271124 328092 271176
rect 328144 271164 328150 271176
rect 337746 271164 337752 271176
rect 328144 271136 337752 271164
rect 328144 271124 328150 271136
rect 337746 271124 337752 271136
rect 337804 271124 337810 271176
rect 342162 271124 342168 271176
rect 342220 271164 342226 271176
rect 356146 271164 356152 271176
rect 342220 271136 356152 271164
rect 342220 271124 342226 271136
rect 356146 271124 356152 271136
rect 356204 271124 356210 271176
rect 364150 271124 364156 271176
rect 364208 271164 364214 271176
rect 386046 271164 386052 271176
rect 364208 271136 386052 271164
rect 364208 271124 364214 271136
rect 386046 271124 386052 271136
rect 386104 271124 386110 271176
rect 431678 271124 431684 271176
rect 431736 271164 431742 271176
rect 484026 271164 484032 271176
rect 431736 271136 484032 271164
rect 431736 271124 431742 271136
rect 484026 271124 484032 271136
rect 484084 271124 484090 271176
rect 484210 271124 484216 271176
rect 484268 271164 484274 271176
rect 519722 271164 519728 271176
rect 484268 271136 519728 271164
rect 484268 271124 484274 271136
rect 519722 271124 519728 271136
rect 519780 271124 519786 271176
rect 519906 271124 519912 271176
rect 519964 271164 519970 271176
rect 523494 271164 523500 271176
rect 519964 271136 523500 271164
rect 519964 271124 519970 271136
rect 523494 271124 523500 271136
rect 523552 271124 523558 271176
rect 523696 271164 523724 271272
rect 523862 271260 523868 271312
rect 523920 271300 523926 271312
rect 610802 271300 610808 271312
rect 523920 271272 610808 271300
rect 523920 271260 523926 271272
rect 610802 271260 610808 271272
rect 610860 271260 610866 271312
rect 621658 271260 621664 271312
rect 621716 271300 621722 271312
rect 636838 271300 636844 271312
rect 621716 271272 636844 271300
rect 621716 271260 621722 271272
rect 636838 271260 636844 271272
rect 636896 271260 636902 271312
rect 538030 271164 538036 271176
rect 523696 271136 538036 271164
rect 538030 271124 538036 271136
rect 538088 271124 538094 271176
rect 538168 271124 538174 271176
rect 538226 271164 538232 271176
rect 625062 271164 625068 271176
rect 538226 271136 625068 271164
rect 538226 271124 538232 271136
rect 625062 271124 625068 271136
rect 625120 271124 625126 271176
rect 356514 271056 356520 271108
rect 356572 271096 356578 271108
rect 358998 271096 359004 271108
rect 356572 271068 359004 271096
rect 356572 271056 356578 271068
rect 358998 271056 359004 271068
rect 359056 271056 359062 271108
rect 128538 270988 128544 271040
rect 128596 271028 128602 271040
rect 181346 271028 181352 271040
rect 128596 271000 181352 271028
rect 128596 270988 128602 271000
rect 181346 270988 181352 271000
rect 181404 270988 181410 271040
rect 189994 270988 190000 271040
rect 190052 271028 190058 271040
rect 216122 271028 216128 271040
rect 190052 271000 216128 271028
rect 190052 270988 190058 271000
rect 216122 270988 216128 271000
rect 216180 270988 216186 271040
rect 389082 270988 389088 271040
rect 389140 271028 389146 271040
rect 415302 271028 415308 271040
rect 389140 271000 415308 271028
rect 389140 270988 389146 271000
rect 415302 270988 415308 271000
rect 415360 270988 415366 271040
rect 439958 270988 439964 271040
rect 440016 271028 440022 271040
rect 493778 271028 493784 271040
rect 440016 271000 493784 271028
rect 440016 270988 440022 271000
rect 493778 270988 493784 271000
rect 493836 270988 493842 271040
rect 499942 270988 499948 271040
rect 500000 271028 500006 271040
rect 500678 271028 500684 271040
rect 500000 271000 500684 271028
rect 500000 270988 500006 271000
rect 500678 270988 500684 271000
rect 500736 270988 500742 271040
rect 507670 270988 507676 271040
rect 507728 271028 507734 271040
rect 593138 271028 593144 271040
rect 507728 271000 593144 271028
rect 507728 270988 507734 271000
rect 593138 270988 593144 271000
rect 593196 270988 593202 271040
rect 130838 270852 130844 270904
rect 130896 270892 130902 270904
rect 182450 270892 182456 270904
rect 130896 270864 182456 270892
rect 130896 270852 130902 270864
rect 182450 270852 182456 270864
rect 182508 270852 182514 270904
rect 200482 270852 200488 270904
rect 200540 270892 200546 270904
rect 224218 270892 224224 270904
rect 200540 270864 224224 270892
rect 200540 270852 200546 270864
rect 224218 270852 224224 270864
rect 224276 270852 224282 270904
rect 416590 270852 416596 270904
rect 416648 270892 416654 270904
rect 463970 270892 463976 270904
rect 416648 270864 463976 270892
rect 416648 270852 416654 270864
rect 463970 270852 463976 270864
rect 464028 270852 464034 270904
rect 464338 270852 464344 270904
rect 464396 270892 464402 270904
rect 519630 270892 519636 270904
rect 464396 270864 519636 270892
rect 464396 270852 464402 270864
rect 519630 270852 519636 270864
rect 519688 270852 519694 270904
rect 520182 270852 520188 270904
rect 520240 270892 520246 270904
rect 523862 270892 523868 270904
rect 520240 270864 523868 270892
rect 520240 270852 520246 270864
rect 523862 270852 523868 270864
rect 523920 270852 523926 270904
rect 526806 270852 526812 270904
rect 526864 270892 526870 270904
rect 621474 270892 621480 270904
rect 526864 270864 621480 270892
rect 526864 270852 526870 270864
rect 621474 270852 621480 270864
rect 621532 270852 621538 270904
rect 137922 270716 137928 270768
rect 137980 270756 137986 270768
rect 187878 270756 187884 270768
rect 137980 270728 187884 270756
rect 137980 270716 137986 270728
rect 187878 270716 187884 270728
rect 187936 270716 187942 270768
rect 418062 270716 418068 270768
rect 418120 270756 418126 270768
rect 462222 270756 462228 270768
rect 418120 270728 462228 270756
rect 418120 270716 418126 270728
rect 462222 270716 462228 270728
rect 462280 270716 462286 270768
rect 464798 270716 464804 270768
rect 464856 270756 464862 270768
rect 484210 270756 484216 270768
rect 464856 270728 484216 270756
rect 464856 270716 464862 270728
rect 484210 270716 484216 270728
rect 484268 270716 484274 270768
rect 484394 270716 484400 270768
rect 484452 270756 484458 270768
rect 485498 270756 485504 270768
rect 484452 270728 485504 270756
rect 484452 270716 484458 270728
rect 485498 270716 485504 270728
rect 485556 270716 485562 270768
rect 489362 270716 489368 270768
rect 489420 270756 489426 270768
rect 551738 270756 551744 270768
rect 489420 270728 551744 270756
rect 489420 270716 489426 270728
rect 551738 270716 551744 270728
rect 551796 270716 551802 270768
rect 591298 270756 591304 270768
rect 557506 270728 591304 270756
rect 116670 270580 116676 270632
rect 116728 270620 116734 270632
rect 151078 270620 151084 270632
rect 116728 270592 151084 270620
rect 116728 270580 116734 270592
rect 151078 270580 151084 270592
rect 151136 270580 151142 270632
rect 237190 270580 237196 270632
rect 237248 270620 237254 270632
rect 237248 270592 237512 270620
rect 237248 270580 237254 270592
rect 115842 270444 115848 270496
rect 115900 270484 115906 270496
rect 171226 270484 171232 270496
rect 115900 270456 171232 270484
rect 115900 270444 115906 270456
rect 171226 270444 171232 270456
rect 171284 270444 171290 270496
rect 172422 270444 172428 270496
rect 172480 270484 172486 270496
rect 209498 270484 209504 270496
rect 172480 270456 209504 270484
rect 172480 270444 172486 270456
rect 209498 270444 209504 270456
rect 209556 270444 209562 270496
rect 233142 270444 233148 270496
rect 233200 270484 233206 270496
rect 237282 270484 237288 270496
rect 233200 270456 237288 270484
rect 233200 270444 233206 270456
rect 237282 270444 237288 270456
rect 237340 270444 237346 270496
rect 237484 270484 237512 270592
rect 400122 270580 400128 270632
rect 400180 270620 400186 270632
rect 435542 270620 435548 270632
rect 400180 270592 435548 270620
rect 400180 270580 400186 270592
rect 435542 270580 435548 270592
rect 435600 270580 435606 270632
rect 437382 270580 437388 270632
rect 437440 270620 437446 270632
rect 471146 270620 471152 270632
rect 437440 270592 471152 270620
rect 437440 270580 437446 270592
rect 471146 270580 471152 270592
rect 471204 270580 471210 270632
rect 474734 270580 474740 270632
rect 474792 270620 474798 270632
rect 538030 270620 538036 270632
rect 474792 270592 538036 270620
rect 474792 270580 474798 270592
rect 538030 270580 538036 270592
rect 538088 270580 538094 270632
rect 538168 270580 538174 270632
rect 538226 270620 538232 270632
rect 557506 270620 557534 270728
rect 591298 270716 591304 270728
rect 591356 270716 591362 270768
rect 538226 270592 557534 270620
rect 538226 270580 538232 270592
rect 237484 270456 248414 270484
rect 110230 270308 110236 270360
rect 110288 270348 110294 270360
rect 167914 270348 167920 270360
rect 110288 270320 167920 270348
rect 110288 270308 110294 270320
rect 167914 270308 167920 270320
rect 167972 270308 167978 270360
rect 173066 270308 173072 270360
rect 173124 270348 173130 270360
rect 210142 270348 210148 270360
rect 173124 270320 210148 270348
rect 173124 270308 173130 270320
rect 210142 270308 210148 270320
rect 210200 270308 210206 270360
rect 213822 270308 213828 270360
rect 213880 270348 213886 270360
rect 240502 270348 240508 270360
rect 213880 270320 240508 270348
rect 213880 270308 213886 270320
rect 240502 270308 240508 270320
rect 240560 270308 240566 270360
rect 248386 270348 248414 270456
rect 249610 270444 249616 270496
rect 249668 270484 249674 270496
rect 253658 270484 253664 270496
rect 249668 270456 253664 270484
rect 249668 270444 249674 270456
rect 253658 270444 253664 270456
rect 253716 270444 253722 270496
rect 291654 270444 291660 270496
rect 291712 270484 291718 270496
rect 295518 270484 295524 270496
rect 291712 270456 295524 270484
rect 291712 270444 291718 270456
rect 295518 270444 295524 270456
rect 295576 270444 295582 270496
rect 297910 270444 297916 270496
rect 297968 270484 297974 270496
rect 299566 270484 299572 270496
rect 297968 270456 299572 270484
rect 297968 270444 297974 270456
rect 299566 270444 299572 270456
rect 299624 270444 299630 270496
rect 299934 270444 299940 270496
rect 299992 270484 299998 270496
rect 300854 270484 300860 270496
rect 299992 270456 300860 270484
rect 299992 270444 299998 270456
rect 300854 270444 300860 270456
rect 300912 270444 300918 270496
rect 359918 270444 359924 270496
rect 359976 270484 359982 270496
rect 376754 270484 376760 270496
rect 359976 270456 376760 270484
rect 359976 270444 359982 270456
rect 376754 270444 376760 270456
rect 376812 270444 376818 270496
rect 377582 270444 377588 270496
rect 377640 270484 377646 270496
rect 391934 270484 391940 270496
rect 377640 270456 391940 270484
rect 377640 270444 377646 270456
rect 391934 270444 391940 270456
rect 391992 270444 391998 270496
rect 396258 270444 396264 270496
rect 396316 270484 396322 270496
rect 423674 270484 423680 270496
rect 396316 270456 423680 270484
rect 396316 270444 396322 270456
rect 423674 270444 423680 270456
rect 423732 270444 423738 270496
rect 429562 270444 429568 270496
rect 429620 270484 429626 270496
rect 480162 270484 480168 270496
rect 429620 270456 480168 270484
rect 429620 270444 429626 270456
rect 480162 270444 480168 270456
rect 480220 270444 480226 270496
rect 480346 270444 480352 270496
rect 480404 270484 480410 270496
rect 485038 270484 485044 270496
rect 480404 270456 485044 270484
rect 480404 270444 480410 270456
rect 485038 270444 485044 270456
rect 485096 270444 485102 270496
rect 486694 270444 486700 270496
rect 486752 270484 486758 270496
rect 494698 270484 494704 270496
rect 486752 270456 494704 270484
rect 486752 270444 486758 270456
rect 494698 270444 494704 270456
rect 494756 270444 494762 270496
rect 494882 270444 494888 270496
rect 494940 270484 494946 270496
rect 560846 270484 560852 270496
rect 494940 270456 560852 270484
rect 494940 270444 494946 270456
rect 560846 270444 560852 270456
rect 560904 270444 560910 270496
rect 252002 270348 252008 270360
rect 248386 270320 252008 270348
rect 252002 270308 252008 270320
rect 252060 270308 252066 270360
rect 262306 270348 262312 270360
rect 253216 270320 262312 270348
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 166902 270172 166908 270224
rect 166960 270212 166966 270224
rect 207382 270212 207388 270224
rect 166960 270184 207388 270212
rect 166960 270172 166966 270184
rect 207382 270172 207388 270184
rect 207440 270172 207446 270224
rect 212442 270172 212448 270224
rect 212500 270212 212506 270224
rect 239950 270212 239956 270224
rect 212500 270184 239956 270212
rect 212500 270172 212506 270184
rect 239950 270172 239956 270184
rect 240008 270172 240014 270224
rect 251082 270172 251088 270224
rect 251140 270212 251146 270224
rect 253216 270212 253244 270320
rect 262306 270308 262312 270320
rect 262364 270308 262370 270360
rect 348418 270308 348424 270360
rect 348476 270348 348482 270360
rect 363046 270348 363052 270360
rect 348476 270320 363052 270348
rect 348476 270308 348482 270320
rect 363046 270308 363052 270320
rect 363104 270308 363110 270360
rect 369394 270308 369400 270360
rect 369452 270348 369458 270360
rect 396074 270348 396080 270360
rect 369452 270320 396080 270348
rect 369452 270308 369458 270320
rect 396074 270308 396080 270320
rect 396132 270308 396138 270360
rect 402054 270308 402060 270360
rect 402112 270348 402118 270360
rect 430574 270348 430580 270360
rect 402112 270320 430580 270348
rect 402112 270308 402118 270320
rect 430574 270308 430580 270320
rect 430632 270308 430638 270360
rect 446950 270308 446956 270360
rect 447008 270348 447014 270360
rect 504910 270348 504916 270360
rect 447008 270320 504916 270348
rect 447008 270308 447014 270320
rect 504910 270308 504916 270320
rect 504968 270308 504974 270360
rect 505048 270308 505054 270360
rect 505106 270348 505112 270360
rect 543182 270348 543188 270360
rect 505106 270320 543188 270348
rect 505106 270308 505112 270320
rect 543182 270308 543188 270320
rect 543240 270308 543246 270360
rect 543366 270308 543372 270360
rect 543424 270348 543430 270360
rect 627914 270348 627920 270360
rect 543424 270320 627920 270348
rect 543424 270308 543430 270320
rect 627914 270308 627920 270320
rect 627972 270308 627978 270360
rect 316954 270240 316960 270292
rect 317012 270280 317018 270292
rect 321554 270280 321560 270292
rect 317012 270252 321560 270280
rect 317012 270240 317018 270252
rect 321554 270240 321560 270252
rect 321612 270240 321618 270292
rect 339310 270240 339316 270292
rect 339368 270280 339374 270292
rect 341518 270280 341524 270292
rect 339368 270252 341524 270280
rect 339368 270240 339374 270252
rect 341518 270240 341524 270252
rect 341576 270240 341582 270292
rect 251140 270184 253244 270212
rect 251140 270172 251146 270184
rect 253842 270172 253848 270224
rect 253900 270212 253906 270224
rect 265066 270212 265072 270224
rect 253900 270184 265072 270212
rect 253900 270172 253906 270184
rect 265066 270172 265072 270184
rect 265124 270172 265130 270224
rect 356698 270172 356704 270224
rect 356756 270212 356762 270224
rect 378134 270212 378140 270224
rect 356756 270184 378140 270212
rect 356756 270172 356762 270184
rect 378134 270172 378140 270184
rect 378192 270172 378198 270224
rect 381538 270172 381544 270224
rect 381596 270212 381602 270224
rect 382274 270212 382280 270224
rect 381596 270184 382280 270212
rect 381596 270172 381602 270184
rect 382274 270172 382280 270184
rect 382332 270172 382338 270224
rect 385678 270172 385684 270224
rect 385736 270212 385742 270224
rect 419534 270212 419540 270224
rect 385736 270184 419540 270212
rect 385736 270172 385742 270184
rect 419534 270172 419540 270184
rect 419592 270172 419598 270224
rect 428274 270172 428280 270224
rect 428332 270212 428338 270224
rect 459554 270212 459560 270224
rect 428332 270184 459560 270212
rect 428332 270172 428338 270184
rect 459554 270172 459560 270184
rect 459612 270172 459618 270224
rect 461854 270172 461860 270224
rect 461912 270212 461918 270224
rect 529198 270212 529204 270224
rect 461912 270184 529204 270212
rect 461912 270172 461918 270184
rect 529198 270172 529204 270184
rect 529256 270172 529262 270224
rect 529658 270172 529664 270224
rect 529716 270212 529722 270224
rect 530762 270212 530768 270224
rect 529716 270184 530768 270212
rect 529716 270172 529722 270184
rect 530762 270172 530768 270184
rect 530820 270172 530826 270224
rect 530946 270172 530952 270224
rect 531004 270212 531010 270224
rect 536098 270212 536104 270224
rect 531004 270184 536104 270212
rect 531004 270172 531010 270184
rect 536098 270172 536104 270184
rect 536156 270172 536162 270224
rect 536282 270172 536288 270224
rect 536340 270212 536346 270224
rect 538030 270212 538036 270224
rect 536340 270184 538036 270212
rect 536340 270172 536346 270184
rect 538030 270172 538036 270184
rect 538088 270172 538094 270224
rect 538168 270172 538174 270224
rect 538226 270212 538232 270224
rect 626626 270212 626632 270224
rect 538226 270184 626632 270212
rect 538226 270172 538232 270184
rect 626626 270172 626632 270184
rect 626684 270172 626690 270224
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 146754 270036 146760 270088
rect 146812 270076 146818 270088
rect 151354 270076 151360 270088
rect 146812 270048 151360 270076
rect 146812 270036 146818 270048
rect 151354 270036 151360 270048
rect 151412 270036 151418 270088
rect 153838 270076 153844 270088
rect 151786 270048 153844 270076
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 142614 269940 142620 269952
rect 75880 269912 142620 269940
rect 75880 269900 75886 269912
rect 142614 269900 142620 269912
rect 142672 269900 142678 269952
rect 143350 269900 143356 269952
rect 143408 269940 143414 269952
rect 151786 269940 151814 270048
rect 153838 270036 153844 270048
rect 153896 270036 153902 270088
rect 159910 270036 159916 270088
rect 159968 270076 159974 270088
rect 202690 270076 202696 270088
rect 159968 270048 202696 270076
rect 159968 270036 159974 270048
rect 202690 270036 202696 270048
rect 202748 270036 202754 270088
rect 205542 270036 205548 270088
rect 205600 270076 205606 270088
rect 234982 270076 234988 270088
rect 205600 270048 234988 270076
rect 205600 270036 205606 270048
rect 234982 270036 234988 270048
rect 235040 270036 235046 270088
rect 239766 270036 239772 270088
rect 239824 270076 239830 270088
rect 250898 270076 250904 270088
rect 239824 270048 250904 270076
rect 239824 270036 239830 270048
rect 250898 270036 250904 270048
rect 250956 270036 250962 270088
rect 266262 270036 266268 270088
rect 266320 270076 266326 270088
rect 277210 270076 277216 270088
rect 266320 270048 277216 270076
rect 266320 270036 266326 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 326890 270036 326896 270088
rect 326948 270076 326954 270088
rect 335538 270076 335544 270088
rect 326948 270048 335544 270076
rect 326948 270036 326954 270048
rect 335538 270036 335544 270048
rect 335596 270036 335602 270088
rect 336826 270036 336832 270088
rect 336884 270076 336890 270088
rect 350534 270076 350540 270088
rect 336884 270048 350540 270076
rect 336884 270036 336890 270048
rect 350534 270036 350540 270048
rect 350592 270036 350598 270088
rect 354214 270036 354220 270088
rect 354272 270076 354278 270088
rect 375374 270076 375380 270088
rect 354272 270048 375380 270076
rect 354272 270036 354278 270048
rect 375374 270036 375380 270048
rect 375432 270036 375438 270088
rect 376570 270036 376576 270088
rect 376628 270076 376634 270088
rect 376628 270048 402974 270076
rect 376628 270036 376634 270048
rect 143408 269912 151814 269940
rect 143408 269900 143414 269912
rect 154482 269900 154488 269952
rect 154540 269940 154546 269952
rect 198182 269940 198188 269952
rect 154540 269912 198188 269940
rect 154540 269900 154546 269912
rect 198182 269900 198188 269912
rect 198240 269900 198246 269952
rect 198642 269900 198648 269952
rect 198700 269940 198706 269952
rect 230014 269940 230020 269952
rect 198700 269912 230020 269940
rect 198700 269900 198706 269912
rect 230014 269900 230020 269912
rect 230072 269900 230078 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 252370 269940 252376 269952
rect 230440 269912 252376 269940
rect 230440 269900 230446 269912
rect 252370 269900 252376 269912
rect 252428 269900 252434 269952
rect 258442 269900 258448 269952
rect 258500 269940 258506 269952
rect 272242 269940 272248 269952
rect 258500 269912 272248 269940
rect 258500 269900 258506 269912
rect 272242 269900 272248 269912
rect 272300 269900 272306 269952
rect 273070 269900 273076 269952
rect 273128 269940 273134 269952
rect 282178 269940 282184 269952
rect 273128 269912 282184 269940
rect 273128 269900 273134 269912
rect 282178 269900 282184 269912
rect 282236 269900 282242 269952
rect 286778 269900 286784 269952
rect 286836 269940 286842 269952
rect 292114 269940 292120 269952
rect 286836 269912 292120 269940
rect 286836 269900 286842 269912
rect 292114 269900 292120 269912
rect 292172 269900 292178 269952
rect 323578 269900 323584 269952
rect 323636 269940 323642 269952
rect 331214 269940 331220 269952
rect 323636 269912 331220 269940
rect 323636 269900 323642 269912
rect 331214 269900 331220 269912
rect 331272 269900 331278 269952
rect 333882 269900 333888 269952
rect 333940 269940 333946 269952
rect 345106 269940 345112 269952
rect 333940 269912 345112 269940
rect 333940 269900 333946 269912
rect 345106 269900 345112 269912
rect 345164 269900 345170 269952
rect 347590 269900 347596 269952
rect 347648 269940 347654 269952
rect 365714 269940 365720 269952
rect 347648 269912 365720 269940
rect 347648 269900 347654 269912
rect 365714 269900 365720 269912
rect 365772 269900 365778 269952
rect 372338 269900 372344 269952
rect 372396 269940 372402 269952
rect 401870 269940 401876 269952
rect 372396 269912 401876 269940
rect 372396 269900 372402 269912
rect 401870 269900 401876 269912
rect 401928 269900 401934 269952
rect 402946 269940 402974 270048
rect 403066 270036 403072 270088
rect 403124 270076 403130 270088
rect 444374 270076 444380 270088
rect 403124 270048 444380 270076
rect 403124 270036 403130 270048
rect 444374 270036 444380 270048
rect 444432 270036 444438 270088
rect 447778 270036 447784 270088
rect 447836 270076 447842 270088
rect 449894 270076 449900 270088
rect 447836 270048 449900 270076
rect 447836 270036 447842 270048
rect 449894 270036 449900 270048
rect 449952 270036 449958 270088
rect 457714 270036 457720 270088
rect 457772 270076 457778 270088
rect 482278 270076 482284 270088
rect 457772 270048 482284 270076
rect 457772 270036 457778 270048
rect 482278 270036 482284 270048
rect 482336 270036 482342 270088
rect 482646 270036 482652 270088
rect 482704 270076 482710 270088
rect 538674 270076 538680 270088
rect 482704 270048 538680 270076
rect 482704 270036 482710 270048
rect 538674 270036 538680 270048
rect 538732 270036 538738 270088
rect 633618 270076 633624 270088
rect 543016 270048 633624 270076
rect 404262 269940 404268 269952
rect 402946 269912 404268 269940
rect 404262 269900 404268 269912
rect 404320 269900 404326 269952
rect 417142 269900 417148 269952
rect 417200 269940 417206 269952
rect 465074 269940 465080 269952
rect 417200 269912 465080 269940
rect 417200 269900 417206 269912
rect 465074 269900 465080 269912
rect 465132 269900 465138 269952
rect 465994 269900 466000 269952
rect 466052 269940 466058 269952
rect 531314 269940 531320 269952
rect 466052 269912 531320 269940
rect 466052 269900 466058 269912
rect 531314 269900 531320 269912
rect 531372 269900 531378 269952
rect 531682 269900 531688 269952
rect 531740 269940 531746 269952
rect 537846 269940 537852 269952
rect 531740 269912 537852 269940
rect 531740 269900 531746 269912
rect 537846 269900 537852 269912
rect 537904 269900 537910 269952
rect 538030 269900 538036 269952
rect 538088 269940 538094 269952
rect 543016 269940 543044 270048
rect 633618 270036 633624 270048
rect 633676 270036 633682 270088
rect 538088 269912 543044 269940
rect 538088 269900 538094 269912
rect 543182 269900 543188 269952
rect 543240 269940 543246 269952
rect 548702 269940 548708 269952
rect 543240 269912 548708 269940
rect 543240 269900 543246 269912
rect 548702 269900 548708 269912
rect 548760 269900 548766 269952
rect 548886 269900 548892 269952
rect 548944 269940 548950 269952
rect 641898 269940 641904 269952
rect 548944 269912 641904 269940
rect 548944 269900 548950 269912
rect 641898 269900 641904 269912
rect 641956 269900 641962 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 139946 269764 139952 269816
rect 140004 269804 140010 269816
rect 181162 269804 181168 269816
rect 140004 269776 181168 269804
rect 140004 269764 140010 269776
rect 181162 269764 181168 269776
rect 181220 269764 181226 269816
rect 182082 269764 182088 269816
rect 182140 269804 182146 269816
rect 186958 269804 186964 269816
rect 182140 269776 186964 269804
rect 182140 269764 182146 269776
rect 186958 269764 186964 269776
rect 187016 269764 187022 269816
rect 187326 269764 187332 269816
rect 187384 269804 187390 269816
rect 191926 269804 191932 269816
rect 187384 269776 191932 269804
rect 187384 269764 187390 269776
rect 191926 269764 191932 269776
rect 191984 269764 191990 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 84102 269628 84108 269680
rect 84160 269668 84166 269680
rect 119798 269668 119804 269680
rect 84160 269640 119804 269668
rect 84160 269628 84166 269640
rect 119798 269628 119804 269640
rect 119856 269628 119862 269680
rect 173710 269668 173716 269680
rect 122806 269640 173716 269668
rect 119062 269492 119068 269544
rect 119120 269532 119126 269544
rect 122806 269532 122834 269640
rect 173710 269628 173716 269640
rect 173768 269628 173774 269680
rect 184750 269628 184756 269680
rect 184808 269668 184814 269680
rect 213822 269668 213828 269680
rect 184808 269640 213828 269668
rect 184808 269628 184814 269640
rect 213822 269628 213828 269640
rect 213880 269628 213886 269680
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 251450 269764 251456 269816
rect 251508 269804 251514 269816
rect 267274 269804 267280 269816
rect 251508 269776 267280 269804
rect 251508 269764 251514 269776
rect 267274 269764 267280 269776
rect 267332 269764 267338 269816
rect 269206 269764 269212 269816
rect 269264 269804 269270 269816
rect 279694 269804 279700 269816
rect 269264 269776 279700 269804
rect 269264 269764 269270 269776
rect 279694 269764 279700 269776
rect 279752 269764 279758 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318794 269804 318800 269816
rect 314528 269776 318800 269804
rect 314528 269764 314534 269776
rect 318794 269764 318800 269776
rect 318852 269764 318858 269816
rect 321922 269764 321928 269816
rect 321980 269804 321986 269816
rect 328454 269804 328460 269816
rect 321980 269776 328460 269804
rect 321980 269764 321986 269776
rect 328454 269764 328460 269776
rect 328512 269764 328518 269816
rect 329374 269764 329380 269816
rect 329432 269804 329438 269816
rect 339494 269804 339500 269816
rect 329432 269776 339500 269804
rect 329432 269764 329438 269776
rect 339494 269764 339500 269776
rect 339552 269764 339558 269816
rect 341794 269764 341800 269816
rect 341852 269804 341858 269816
rect 357434 269804 357440 269816
rect 341852 269776 357440 269804
rect 341852 269764 341858 269776
rect 357434 269764 357440 269776
rect 357492 269764 357498 269816
rect 364978 269764 364984 269816
rect 365036 269804 365042 269816
rect 390554 269804 390560 269816
rect 365036 269776 390560 269804
rect 365036 269764 365042 269776
rect 390554 269764 390560 269776
rect 390612 269764 390618 269816
rect 392302 269764 392308 269816
rect 392360 269804 392366 269816
rect 429378 269804 429384 269816
rect 392360 269776 429384 269804
rect 392360 269764 392366 269776
rect 429378 269764 429384 269776
rect 429436 269764 429442 269816
rect 434438 269764 434444 269816
rect 434496 269804 434502 269816
rect 469214 269804 469220 269816
rect 434496 269776 469220 269804
rect 434496 269764 434502 269776
rect 469214 269764 469220 269776
rect 469272 269764 469278 269816
rect 470962 269764 470968 269816
rect 471020 269804 471026 269816
rect 471020 269776 475608 269804
rect 471020 269764 471026 269776
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 250898 269628 250904 269680
rect 250956 269668 250962 269680
rect 258166 269668 258172 269680
rect 250956 269640 258172 269668
rect 250956 269628 250962 269640
rect 258166 269628 258172 269640
rect 258224 269628 258230 269680
rect 351638 269628 351644 269680
rect 351696 269668 351702 269680
rect 364334 269668 364340 269680
rect 351696 269640 364340 269668
rect 351696 269628 351702 269640
rect 364334 269628 364340 269640
rect 364392 269628 364398 269680
rect 384022 269628 384028 269680
rect 384080 269668 384086 269680
rect 388070 269668 388076 269680
rect 384080 269640 388076 269668
rect 384080 269628 384086 269640
rect 388070 269628 388076 269640
rect 388128 269628 388134 269680
rect 394694 269628 394700 269680
rect 394752 269668 394758 269680
rect 416774 269668 416780 269680
rect 394752 269640 416780 269668
rect 394752 269628 394758 269640
rect 416774 269628 416780 269640
rect 416832 269628 416838 269680
rect 424594 269628 424600 269680
rect 424652 269668 424658 269680
rect 475378 269668 475384 269680
rect 424652 269640 475384 269668
rect 424652 269628 424658 269640
rect 475378 269628 475384 269640
rect 475436 269628 475442 269680
rect 475580 269668 475608 269776
rect 476022 269764 476028 269816
rect 476080 269804 476086 269816
rect 482646 269804 482652 269816
rect 476080 269776 482652 269804
rect 476080 269764 476086 269776
rect 482646 269764 482652 269776
rect 482704 269764 482710 269816
rect 541434 269804 541440 269816
rect 482848 269776 541440 269804
rect 482848 269668 482876 269776
rect 541434 269764 541440 269776
rect 541492 269764 541498 269816
rect 542998 269764 543004 269816
rect 543056 269804 543062 269816
rect 644474 269804 644480 269816
rect 543056 269776 644480 269804
rect 543056 269764 543062 269776
rect 644474 269764 644480 269776
rect 644532 269764 644538 269816
rect 475580 269640 482876 269668
rect 485038 269628 485044 269680
rect 485096 269668 485102 269680
rect 485096 269640 548564 269668
rect 485096 269628 485102 269640
rect 119120 269504 122834 269532
rect 119120 269492 119126 269504
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 187326 269532 187332 269544
rect 183520 269504 187332 269532
rect 183520 269492 183526 269504
rect 187326 269492 187332 269504
rect 187384 269492 187390 269544
rect 208302 269492 208308 269544
rect 208360 269532 208366 269544
rect 230750 269532 230756 269544
rect 208360 269504 230756 269532
rect 208360 269492 208366 269504
rect 230750 269492 230756 269504
rect 230808 269492 230814 269544
rect 390462 269492 390468 269544
rect 390520 269532 390526 269544
rect 390520 269504 393314 269532
rect 390520 269492 390526 269504
rect 118602 269356 118608 269408
rect 118660 269396 118666 269408
rect 166902 269396 166908 269408
rect 118660 269368 166908 269396
rect 118660 269356 118666 269368
rect 166902 269356 166908 269368
rect 166960 269356 166966 269408
rect 335630 269356 335636 269408
rect 335688 269396 335694 269408
rect 343818 269396 343824 269408
rect 335688 269368 343824 269396
rect 335688 269356 335694 269368
rect 343818 269356 343824 269368
rect 343876 269356 343882 269408
rect 393286 269396 393314 269504
rect 401594 269492 401600 269544
rect 401652 269532 401658 269544
rect 426618 269532 426624 269544
rect 401652 269504 426624 269532
rect 401652 269492 401658 269504
rect 426618 269492 426624 269504
rect 426676 269492 426682 269544
rect 427354 269492 427360 269544
rect 427412 269532 427418 269544
rect 475746 269532 475752 269544
rect 427412 269504 475752 269532
rect 427412 269492 427418 269504
rect 475746 269492 475752 269504
rect 475804 269492 475810 269544
rect 489868 269532 489874 269544
rect 475948 269504 489874 269532
rect 402422 269396 402428 269408
rect 393286 269368 402428 269396
rect 402422 269356 402428 269368
rect 402480 269356 402486 269408
rect 419626 269356 419632 269408
rect 419684 269396 419690 269408
rect 468294 269396 468300 269408
rect 419684 269368 468300 269396
rect 419684 269356 419690 269368
rect 468294 269356 468300 269368
rect 468352 269356 468358 269408
rect 469214 269356 469220 269408
rect 469272 269396 469278 269408
rect 475948 269396 475976 269504
rect 489868 269492 489874 269504
rect 489926 269492 489932 269544
rect 490006 269492 490012 269544
rect 490064 269532 490070 269544
rect 494514 269532 494520 269544
rect 490064 269504 494520 269532
rect 490064 269492 490070 269504
rect 494514 269492 494520 269504
rect 494572 269492 494578 269544
rect 494698 269492 494704 269544
rect 494756 269532 494762 269544
rect 504910 269532 504916 269544
rect 494756 269504 504916 269532
rect 494756 269492 494762 269504
rect 504910 269492 504916 269504
rect 504968 269492 504974 269544
rect 505048 269492 505054 269544
rect 505106 269532 505112 269544
rect 505106 269504 545620 269532
rect 505106 269492 505112 269504
rect 545592 269464 545620 269504
rect 545850 269492 545856 269544
rect 545908 269532 545914 269544
rect 546494 269532 546500 269544
rect 545908 269504 546500 269532
rect 545908 269492 545914 269504
rect 546494 269492 546500 269504
rect 546552 269492 546558 269544
rect 548536 269532 548564 269640
rect 548702 269628 548708 269680
rect 548760 269668 548766 269680
rect 564434 269668 564440 269680
rect 548760 269640 564440 269668
rect 548760 269628 548766 269640
rect 564434 269628 564440 269640
rect 564492 269628 564498 269680
rect 553394 269532 553400 269544
rect 548536 269504 553400 269532
rect 553394 269492 553400 269504
rect 553452 269492 553458 269544
rect 558914 269492 558920 269544
rect 558972 269532 558978 269544
rect 572714 269532 572720 269544
rect 558972 269504 572720 269532
rect 558972 269492 558978 269504
rect 572714 269492 572720 269504
rect 572772 269492 572778 269544
rect 545592 269436 545712 269464
rect 479058 269396 479064 269408
rect 469272 269368 475976 269396
rect 476086 269368 479064 269396
rect 469272 269356 469278 269368
rect 136818 269220 136824 269272
rect 136876 269260 136882 269272
rect 182174 269260 182180 269272
rect 136876 269232 182180 269260
rect 136876 269220 136882 269232
rect 182174 269220 182180 269232
rect 182232 269220 182238 269272
rect 264882 269220 264888 269272
rect 264940 269260 264946 269272
rect 269114 269260 269120 269272
rect 264940 269232 269120 269260
rect 264940 269220 264946 269232
rect 269114 269220 269120 269232
rect 269172 269220 269178 269272
rect 295334 269220 295340 269272
rect 295392 269260 295398 269272
rect 297910 269260 297916 269272
rect 295392 269232 297916 269260
rect 295392 269220 295398 269232
rect 297910 269220 297916 269232
rect 297968 269220 297974 269272
rect 420914 269220 420920 269272
rect 420972 269260 420978 269272
rect 448514 269260 448520 269272
rect 420972 269232 448520 269260
rect 420972 269220 420978 269232
rect 448514 269220 448520 269232
rect 448572 269220 448578 269272
rect 450722 269220 450728 269272
rect 450780 269260 450786 269272
rect 471974 269260 471980 269272
rect 450780 269232 471980 269260
rect 450780 269220 450786 269232
rect 471974 269220 471980 269232
rect 472032 269220 472038 269272
rect 474274 269220 474280 269272
rect 474332 269260 474338 269272
rect 476086 269260 476114 269368
rect 479058 269356 479064 269368
rect 479116 269356 479122 269408
rect 479242 269356 479248 269408
rect 479300 269396 479306 269408
rect 480162 269396 480168 269408
rect 479300 269368 480168 269396
rect 479300 269356 479306 269368
rect 480162 269356 480168 269368
rect 480220 269356 480226 269408
rect 480346 269356 480352 269408
rect 480404 269396 480410 269408
rect 480404 269368 538444 269396
rect 480404 269356 480410 269368
rect 474332 269232 476114 269260
rect 474332 269220 474338 269232
rect 476758 269220 476764 269272
rect 476816 269260 476822 269272
rect 538214 269260 538220 269272
rect 476816 269232 538220 269260
rect 476816 269220 476822 269232
rect 538214 269220 538220 269232
rect 538272 269220 538278 269272
rect 538416 269192 538444 269368
rect 538582 269356 538588 269408
rect 538640 269396 538646 269408
rect 543366 269396 543372 269408
rect 538640 269368 543372 269396
rect 538640 269356 538646 269368
rect 543366 269356 543372 269368
rect 543424 269356 543430 269408
rect 543550 269356 543556 269408
rect 543608 269396 543614 269408
rect 545298 269396 545304 269408
rect 543608 269368 545304 269396
rect 543608 269356 543614 269368
rect 545298 269356 545304 269368
rect 545356 269356 545362 269408
rect 541618 269220 541624 269272
rect 541676 269260 541682 269272
rect 545482 269260 545488 269272
rect 541676 269232 545488 269260
rect 541676 269220 541682 269232
rect 545482 269220 545488 269232
rect 545540 269220 545546 269272
rect 541434 269192 541440 269204
rect 538416 269164 541440 269192
rect 541434 269152 541440 269164
rect 541492 269152 541498 269204
rect 545684 269192 545712 269436
rect 545850 269356 545856 269408
rect 545908 269396 545914 269408
rect 548886 269396 548892 269408
rect 545908 269368 548892 269396
rect 545908 269356 545914 269368
rect 548886 269356 548892 269368
rect 548944 269356 548950 269408
rect 549254 269356 549260 269408
rect 549312 269396 549318 269408
rect 568574 269396 568580 269408
rect 549312 269368 568580 269396
rect 549312 269356 549318 269368
rect 568574 269356 568580 269368
rect 568632 269356 568638 269408
rect 557534 269260 557540 269272
rect 557506 269220 557540 269260
rect 557592 269220 557598 269272
rect 557506 269192 557534 269220
rect 545684 269164 557534 269192
rect 282730 269084 282736 269136
rect 282788 269124 282794 269136
rect 288802 269124 288808 269136
rect 282788 269096 288808 269124
rect 282788 269084 282794 269096
rect 288802 269084 288808 269096
rect 288860 269084 288866 269136
rect 294046 269084 294052 269136
rect 294104 269124 294110 269136
rect 297082 269124 297088 269136
rect 294104 269096 297088 269124
rect 294104 269084 294110 269096
rect 297082 269084 297088 269096
rect 297140 269084 297146 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 502610 269084 502616 269136
rect 502668 269124 502674 269136
rect 505002 269124 505008 269136
rect 502668 269096 505008 269124
rect 502668 269084 502674 269096
rect 505002 269084 505008 269096
rect 505060 269084 505066 269136
rect 108942 269016 108948 269068
rect 109000 269056 109006 269068
rect 166258 269056 166264 269068
rect 109000 269028 166264 269056
rect 109000 269016 109006 269028
rect 166258 269016 166264 269028
rect 166316 269016 166322 269068
rect 185578 269016 185584 269068
rect 185636 269056 185642 269068
rect 196894 269056 196900 269068
rect 185636 269028 196900 269056
rect 185636 269016 185642 269028
rect 196894 269016 196900 269028
rect 196952 269016 196958 269068
rect 422294 269056 422300 269068
rect 412606 269028 422300 269056
rect 86862 268880 86868 268932
rect 86920 268920 86926 268932
rect 144730 268920 144736 268932
rect 86920 268892 144736 268920
rect 86920 268880 86926 268892
rect 144730 268880 144736 268892
rect 144788 268880 144794 268932
rect 179322 268880 179328 268932
rect 179380 268920 179386 268932
rect 215938 268920 215944 268932
rect 179380 268892 215944 268920
rect 179380 268880 179386 268892
rect 215938 268880 215944 268892
rect 215996 268880 216002 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 400582 268920 400588 268932
rect 382424 268892 400588 268920
rect 382424 268880 382430 268892
rect 400582 268880 400588 268892
rect 400640 268880 400646 268932
rect 102502 268744 102508 268796
rect 102560 268784 102566 268796
rect 162946 268784 162952 268796
rect 102560 268756 162952 268784
rect 102560 268744 102566 268756
rect 162946 268744 162952 268756
rect 163004 268744 163010 268796
rect 163130 268744 163136 268796
rect 163188 268784 163194 268796
rect 203518 268784 203524 268796
rect 163188 268756 203524 268784
rect 163188 268744 163194 268756
rect 203518 268744 203524 268756
rect 203576 268744 203582 268796
rect 203978 268744 203984 268796
rect 204036 268784 204042 268796
rect 227714 268784 227720 268796
rect 204036 268756 227720 268784
rect 204036 268744 204042 268756
rect 227714 268744 227720 268756
rect 227772 268744 227778 268796
rect 227898 268744 227904 268796
rect 227956 268784 227962 268796
rect 250714 268784 250720 268796
rect 227956 268756 250720 268784
rect 227956 268744 227962 268756
rect 250714 268744 250720 268756
rect 250772 268744 250778 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 412606 268784 412634 269028
rect 422294 269016 422300 269028
rect 422352 269016 422358 269068
rect 443914 269016 443920 269068
rect 443972 269056 443978 269068
rect 502334 269056 502340 269068
rect 443972 269028 502340 269056
rect 443972 269016 443978 269028
rect 502334 269016 502340 269028
rect 502392 269016 502398 269068
rect 506106 269016 506112 269068
rect 506164 269056 506170 269068
rect 591022 269056 591028 269068
rect 506164 269028 591028 269056
rect 506164 269016 506170 269028
rect 591022 269016 591028 269028
rect 591080 269016 591086 269068
rect 418982 268880 418988 268932
rect 419040 268920 419046 268932
rect 440234 268920 440240 268932
rect 419040 268892 440240 268920
rect 419040 268880 419046 268892
rect 440234 268880 440240 268892
rect 440292 268880 440298 268932
rect 441154 268880 441160 268932
rect 441212 268920 441218 268932
rect 499574 268920 499580 268932
rect 441212 268892 499580 268920
rect 441212 268880 441218 268892
rect 499574 268880 499580 268892
rect 499632 268880 499638 268932
rect 503254 268880 503260 268932
rect 503312 268920 503318 268932
rect 587894 268920 587900 268932
rect 503312 268892 587900 268920
rect 503312 268880 503318 268892
rect 587894 268880 587900 268892
rect 587952 268880 587958 268932
rect 387392 268756 412634 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268796
rect 422352 268784 422358 268796
rect 436094 268784 436100 268796
rect 422352 268756 436100 268784
rect 422352 268744 422358 268756
rect 436094 268744 436100 268756
rect 436152 268744 436158 268796
rect 446122 268744 446128 268796
rect 446180 268784 446186 268796
rect 505186 268784 505192 268796
rect 446180 268756 505192 268784
rect 446180 268744 446186 268756
rect 505186 268744 505192 268756
rect 505244 268744 505250 268796
rect 508222 268744 508228 268796
rect 508280 268784 508286 268796
rect 514018 268784 514024 268796
rect 508280 268756 514024 268784
rect 508280 268744 508286 268756
rect 514018 268744 514024 268756
rect 514076 268744 514082 268796
rect 598842 268784 598848 268796
rect 514772 268756 598848 268784
rect 99282 268608 99288 268660
rect 99340 268648 99346 268660
rect 160462 268648 160468 268660
rect 99340 268620 160468 268648
rect 99340 268608 99346 268620
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 162762 268608 162768 268660
rect 162820 268648 162826 268660
rect 205174 268648 205180 268660
rect 162820 268620 205180 268648
rect 162820 268608 162826 268620
rect 205174 268608 205180 268620
rect 205232 268608 205238 268660
rect 219526 268608 219532 268660
rect 219584 268648 219590 268660
rect 244918 268648 244924 268660
rect 219584 268620 244924 268648
rect 219584 268608 219590 268620
rect 244918 268608 244924 268620
rect 244976 268608 244982 268660
rect 363046 268608 363052 268660
rect 363104 268648 363110 268660
rect 386414 268648 386420 268660
rect 363104 268620 386420 268648
rect 363104 268608 363110 268620
rect 386414 268608 386420 268620
rect 386472 268608 386478 268660
rect 397638 268608 397644 268660
rect 397696 268648 397702 268660
rect 433334 268648 433340 268660
rect 397696 268620 433340 268648
rect 397696 268608 397702 268620
rect 433334 268608 433340 268620
rect 433392 268608 433398 268660
rect 448606 268608 448612 268660
rect 448664 268648 448670 268660
rect 509326 268648 509332 268660
rect 448664 268620 509332 268648
rect 448664 268608 448670 268620
rect 509326 268608 509332 268620
rect 509384 268608 509390 268660
rect 510706 268608 510712 268660
rect 510764 268648 510770 268660
rect 514772 268648 514800 268756
rect 598842 268744 598848 268756
rect 598900 268744 598906 268796
rect 510764 268620 514800 268648
rect 510764 268608 510770 268620
rect 514938 268608 514944 268660
rect 514996 268648 515002 268660
rect 517514 268648 517520 268660
rect 514996 268620 517520 268648
rect 514996 268608 515002 268620
rect 517514 268608 517520 268620
rect 517572 268608 517578 268660
rect 518434 268608 518440 268660
rect 518492 268648 518498 268660
rect 608686 268648 608692 268660
rect 518492 268620 608692 268648
rect 518492 268608 518498 268620
rect 608686 268608 608692 268620
rect 608744 268608 608750 268660
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 155862 268472 155868 268524
rect 155920 268512 155926 268524
rect 200206 268512 200212 268524
rect 155920 268484 200212 268512
rect 155920 268472 155926 268484
rect 200206 268472 200212 268484
rect 200264 268472 200270 268524
rect 202966 268472 202972 268524
rect 203024 268512 203030 268524
rect 233326 268512 233332 268524
rect 203024 268484 233332 268512
rect 203024 268472 203030 268484
rect 233326 268472 233332 268484
rect 233384 268472 233390 268524
rect 245562 268472 245568 268524
rect 245620 268512 245626 268524
rect 263134 268512 263140 268524
rect 245620 268484 263140 268512
rect 245620 268472 245626 268484
rect 263134 268472 263140 268484
rect 263192 268472 263198 268524
rect 263502 268472 263508 268524
rect 263560 268512 263566 268524
rect 275554 268512 275560 268524
rect 263560 268484 275560 268512
rect 263560 268472 263566 268484
rect 275554 268472 275560 268484
rect 275612 268472 275618 268524
rect 328546 268472 328552 268524
rect 328604 268512 328610 268524
rect 334342 268512 334348 268524
rect 328604 268484 334348 268512
rect 328604 268472 328610 268484
rect 334342 268472 334348 268484
rect 334400 268472 334406 268524
rect 345934 268472 345940 268524
rect 345992 268512 345998 268524
rect 360286 268512 360292 268524
rect 345992 268484 360292 268512
rect 345992 268472 345998 268484
rect 360286 268472 360292 268484
rect 360344 268472 360350 268524
rect 360746 268472 360752 268524
rect 360804 268512 360810 268524
rect 369854 268512 369860 268524
rect 360804 268484 369860 268512
rect 360804 268472 360810 268484
rect 369854 268472 369860 268484
rect 369912 268472 369918 268524
rect 370314 268472 370320 268524
rect 370372 268512 370378 268524
rect 397454 268512 397460 268524
rect 370372 268484 397460 268512
rect 370372 268472 370378 268484
rect 397454 268472 397460 268484
rect 397512 268472 397518 268524
rect 400582 268472 400588 268524
rect 400640 268512 400646 268524
rect 441614 268512 441620 268524
rect 400640 268484 441620 268512
rect 400640 268472 400646 268484
rect 441614 268472 441620 268484
rect 441672 268472 441678 268524
rect 456058 268472 456064 268524
rect 456116 268512 456122 268524
rect 456116 268484 512592 268512
rect 456116 268472 456122 268484
rect 66254 268336 66260 268388
rect 66312 268376 66318 268388
rect 137278 268376 137284 268388
rect 66312 268348 137284 268376
rect 66312 268336 66318 268348
rect 137278 268336 137284 268348
rect 137336 268336 137342 268388
rect 147582 268336 147588 268388
rect 147640 268376 147646 268388
rect 193582 268376 193588 268388
rect 147640 268348 193588 268376
rect 147640 268336 147646 268348
rect 193582 268336 193588 268348
rect 193640 268336 193646 268388
rect 197262 268336 197268 268388
rect 197320 268376 197326 268388
rect 229186 268376 229192 268388
rect 197320 268348 229192 268376
rect 197320 268336 197326 268348
rect 229186 268336 229192 268348
rect 229244 268336 229250 268388
rect 233694 268336 233700 268388
rect 233752 268376 233758 268388
rect 254854 268376 254860 268388
rect 233752 268348 254860 268376
rect 233752 268336 233758 268348
rect 254854 268336 254860 268348
rect 254912 268336 254918 268388
rect 255222 268336 255228 268388
rect 255280 268376 255286 268388
rect 269758 268376 269764 268388
rect 255280 268348 269764 268376
rect 255280 268336 255286 268348
rect 269758 268336 269764 268348
rect 269816 268336 269822 268388
rect 335170 268336 335176 268388
rect 335228 268376 335234 268388
rect 347774 268376 347780 268388
rect 335228 268348 347780 268376
rect 335228 268336 335234 268348
rect 347774 268336 347780 268348
rect 347832 268336 347838 268388
rect 350074 268336 350080 268388
rect 350132 268376 350138 268388
rect 367094 268376 367100 268388
rect 350132 268348 367100 268376
rect 350132 268336 350138 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 374914 268336 374920 268388
rect 374972 268376 374978 268388
rect 404446 268376 404452 268388
rect 374972 268348 404452 268376
rect 374972 268336 374978 268348
rect 404446 268336 404452 268348
rect 404504 268336 404510 268388
rect 407206 268336 407212 268388
rect 407264 268376 407270 268388
rect 451458 268376 451464 268388
rect 407264 268348 451464 268376
rect 407264 268336 407270 268348
rect 451458 268336 451464 268348
rect 451516 268336 451522 268388
rect 466822 268336 466828 268388
rect 466880 268376 466886 268388
rect 512362 268376 512368 268388
rect 466880 268348 512368 268376
rect 466880 268336 466886 268348
rect 512362 268336 512368 268348
rect 512420 268336 512426 268388
rect 512564 268376 512592 268484
rect 512730 268472 512736 268524
rect 512788 268512 512794 268524
rect 523678 268512 523684 268524
rect 512788 268484 523684 268512
rect 512788 268472 512794 268484
rect 523678 268472 523684 268484
rect 523736 268472 523742 268524
rect 525334 268472 525340 268524
rect 525392 268512 525398 268524
rect 527174 268512 527180 268524
rect 525392 268484 527180 268512
rect 525392 268472 525398 268484
rect 527174 268472 527180 268484
rect 527232 268472 527238 268524
rect 527358 268472 527364 268524
rect 527416 268512 527422 268524
rect 527416 268484 528784 268512
rect 527416 268472 527422 268484
rect 513834 268376 513840 268388
rect 512564 268348 513840 268376
rect 513834 268336 513840 268348
rect 513892 268336 513898 268388
rect 514018 268336 514024 268388
rect 514076 268376 514082 268388
rect 528756 268376 528784 268484
rect 528922 268472 528928 268524
rect 528980 268512 528986 268524
rect 619726 268512 619732 268524
rect 528980 268484 619732 268512
rect 528980 268472 528986 268484
rect 619726 268472 619732 268484
rect 619784 268472 619790 268524
rect 543688 268376 543694 268388
rect 514076 268348 528692 268376
rect 528756 268348 543694 268376
rect 514076 268336 514082 268348
rect 122742 268200 122748 268252
rect 122800 268240 122806 268252
rect 176194 268240 176200 268252
rect 122800 268212 176200 268240
rect 122800 268200 122806 268212
rect 176194 268200 176200 268212
rect 176252 268200 176258 268252
rect 326062 268200 326068 268252
rect 326120 268240 326126 268252
rect 331398 268240 331404 268252
rect 326120 268212 331404 268240
rect 326120 268200 326126 268212
rect 331398 268200 331404 268212
rect 331456 268200 331462 268252
rect 420454 268200 420460 268252
rect 420512 268240 420518 268252
rect 469398 268240 469404 268252
rect 420512 268212 469404 268240
rect 420512 268200 420518 268212
rect 469398 268200 469404 268212
rect 469456 268200 469462 268252
rect 470134 268200 470140 268252
rect 470192 268240 470198 268252
rect 523494 268240 523500 268252
rect 470192 268212 523500 268240
rect 470192 268200 470198 268212
rect 523494 268200 523500 268212
rect 523552 268200 523558 268252
rect 523678 268200 523684 268252
rect 523736 268240 523742 268252
rect 528508 268240 528514 268252
rect 523736 268212 528514 268240
rect 523736 268200 523742 268212
rect 528508 268200 528514 268212
rect 528566 268200 528572 268252
rect 528664 268240 528692 268348
rect 543688 268336 543694 268348
rect 543746 268336 543752 268388
rect 543826 268336 543832 268388
rect 543884 268376 543890 268388
rect 543884 268348 548656 268376
rect 543884 268336 543890 268348
rect 548426 268240 548432 268252
rect 528664 268212 548432 268240
rect 548426 268200 548432 268212
rect 548484 268200 548490 268252
rect 548628 268240 548656 268348
rect 548794 268336 548800 268388
rect 548852 268376 548858 268388
rect 594794 268376 594800 268388
rect 548852 268348 594800 268376
rect 548852 268336 548858 268348
rect 594794 268336 594800 268348
rect 594852 268336 594858 268388
rect 638954 268240 638960 268252
rect 548628 268212 638960 268240
rect 638954 268200 638960 268212
rect 639012 268200 639018 268252
rect 133782 268064 133788 268116
rect 133840 268104 133846 268116
rect 183646 268104 183652 268116
rect 133840 268076 183652 268104
rect 133840 268064 133846 268076
rect 183646 268064 183652 268076
rect 183704 268064 183710 268116
rect 436186 268064 436192 268116
rect 436244 268104 436250 268116
rect 488534 268104 488540 268116
rect 436244 268076 488540 268104
rect 436244 268064 436250 268076
rect 488534 268064 488540 268076
rect 488592 268064 488598 268116
rect 489886 268076 494744 268104
rect 125502 267928 125508 267980
rect 125560 267968 125566 267980
rect 147582 267968 147588 267980
rect 125560 267940 147588 267968
rect 125560 267928 125566 267940
rect 147582 267928 147588 267940
rect 147640 267928 147646 267980
rect 442810 267928 442816 267980
rect 442868 267968 442874 267980
rect 460842 267968 460848 267980
rect 442868 267940 460848 267968
rect 442868 267928 442874 267940
rect 460842 267928 460848 267940
rect 460900 267928 460906 267980
rect 431954 267792 431960 267844
rect 432012 267832 432018 267844
rect 447134 267832 447140 267844
rect 432012 267804 447140 267832
rect 432012 267792 432018 267804
rect 447134 267792 447140 267804
rect 447192 267792 447198 267844
rect 489178 267792 489184 267844
rect 489236 267832 489242 267844
rect 489886 267832 489914 268076
rect 494054 267900 494060 267912
rect 489236 267804 489914 267832
rect 492646 267872 494060 267900
rect 489236 267792 489242 267804
rect 88978 267656 88984 267708
rect 89036 267696 89042 267708
rect 144546 267696 144552 267708
rect 89036 267668 144552 267696
rect 89036 267656 89042 267668
rect 144546 267656 144552 267668
rect 144604 267656 144610 267708
rect 144914 267656 144920 267708
rect 144972 267696 144978 267708
rect 150526 267696 150532 267708
rect 144972 267668 150532 267696
rect 144972 267656 144978 267668
rect 150526 267656 150532 267668
rect 150584 267656 150590 267708
rect 171778 267656 171784 267708
rect 171836 267696 171842 267708
rect 199378 267696 199384 267708
rect 171836 267668 199384 267696
rect 171836 267656 171842 267668
rect 199378 267656 199384 267668
rect 199436 267656 199442 267708
rect 207658 267656 207664 267708
rect 207716 267696 207722 267708
rect 213454 267696 213460 267708
rect 207716 267668 213460 267696
rect 207716 267656 207722 267668
rect 213454 267656 213460 267668
rect 213512 267656 213518 267708
rect 216122 267656 216128 267708
rect 216180 267696 216186 267708
rect 223390 267696 223396 267708
rect 216180 267668 223396 267696
rect 216180 267656 216186 267668
rect 223390 267656 223396 267668
rect 223448 267656 223454 267708
rect 370774 267656 370780 267708
rect 370832 267696 370838 267708
rect 381354 267696 381360 267708
rect 370832 267668 381360 267696
rect 370832 267656 370838 267668
rect 381354 267656 381360 267668
rect 381412 267656 381418 267708
rect 393130 267656 393136 267708
rect 393188 267696 393194 267708
rect 402054 267696 402060 267708
rect 393188 267668 402060 267696
rect 393188 267656 393194 267668
rect 402054 267656 402060 267668
rect 402112 267656 402118 267708
rect 405550 267656 405556 267708
rect 405608 267696 405614 267708
rect 420914 267696 420920 267708
rect 405608 267668 420920 267696
rect 405608 267656 405614 267668
rect 420914 267656 420920 267668
rect 420972 267656 420978 267708
rect 440326 267656 440332 267708
rect 440384 267696 440390 267708
rect 492646 267696 492674 267872
rect 494054 267860 494060 267872
rect 494112 267860 494118 267912
rect 494716 267832 494744 268076
rect 500770 268064 500776 268116
rect 500828 268104 500834 268116
rect 583846 268104 583852 268116
rect 500828 268076 583852 268104
rect 500828 268064 500834 268076
rect 583846 268064 583852 268076
rect 583904 268064 583910 268116
rect 496446 267928 496452 267980
rect 496504 267968 496510 267980
rect 498194 267968 498200 267980
rect 496504 267940 498200 267968
rect 496504 267928 496510 267940
rect 498194 267928 498200 267940
rect 498252 267928 498258 267980
rect 499114 267928 499120 267980
rect 499172 267968 499178 267980
rect 582374 267968 582380 267980
rect 499172 267940 582380 267968
rect 499172 267928 499178 267940
rect 582374 267928 582380 267940
rect 582432 267928 582438 267980
rect 567654 267832 567660 267844
rect 494716 267804 567660 267832
rect 567654 267792 567660 267804
rect 567712 267792 567718 267844
rect 440384 267668 492674 267696
rect 440384 267656 440390 267668
rect 493318 267656 493324 267708
rect 493376 267696 493382 267708
rect 495618 267696 495624 267708
rect 493376 267668 495624 267696
rect 493376 267656 493382 267668
rect 495618 267656 495624 267668
rect 495676 267656 495682 267708
rect 495802 267656 495808 267708
rect 495860 267696 495866 267708
rect 496630 267696 496636 267708
rect 495860 267668 496636 267696
rect 495860 267656 495866 267668
rect 496630 267656 496636 267668
rect 496688 267656 496694 267708
rect 497458 267656 497464 267708
rect 497516 267696 497522 267708
rect 543688 267696 543694 267708
rect 497516 267668 543694 267696
rect 497516 267656 497522 267668
rect 543688 267656 543694 267668
rect 543746 267656 543752 267708
rect 543826 267656 543832 267708
rect 543884 267696 543890 267708
rect 571978 267696 571984 267708
rect 543884 267668 571984 267696
rect 543884 267656 543890 267668
rect 571978 267656 571984 267668
rect 572036 267656 572042 267708
rect 581270 267656 581276 267708
rect 581328 267696 581334 267708
rect 585778 267696 585784 267708
rect 581328 267668 585784 267696
rect 581328 267656 581334 267668
rect 585778 267656 585784 267668
rect 585836 267656 585842 267708
rect 95878 267520 95884 267572
rect 95936 267560 95942 267572
rect 154666 267560 154672 267572
rect 95936 267532 154672 267560
rect 95936 267520 95942 267532
rect 154666 267520 154672 267532
rect 154724 267520 154730 267572
rect 162118 267520 162124 267572
rect 162176 267560 162182 267572
rect 169570 267560 169576 267572
rect 162176 267532 169576 267560
rect 162176 267520 162182 267532
rect 169570 267520 169576 267532
rect 169628 267520 169634 267572
rect 187142 267520 187148 267572
rect 187200 267560 187206 267572
rect 221734 267560 221740 267572
rect 187200 267532 221740 267560
rect 187200 267520 187206 267532
rect 221734 267520 221740 267532
rect 221792 267520 221798 267572
rect 365806 267520 365812 267572
rect 365864 267560 365870 267572
rect 377582 267560 377588 267572
rect 365864 267532 377588 267560
rect 365864 267520 365870 267532
rect 377582 267520 377588 267532
rect 377640 267520 377646 267572
rect 383194 267520 383200 267572
rect 383252 267560 383258 267572
rect 394694 267560 394700 267572
rect 383252 267532 394700 267560
rect 383252 267520 383258 267532
rect 394694 267520 394700 267532
rect 394752 267520 394758 267572
rect 399754 267520 399760 267572
rect 399812 267560 399818 267572
rect 418982 267560 418988 267572
rect 399812 267532 418988 267560
rect 399812 267520 399818 267532
rect 418982 267520 418988 267532
rect 419040 267520 419046 267572
rect 430390 267520 430396 267572
rect 430448 267560 430454 267572
rect 457438 267560 457444 267572
rect 430448 267532 457444 267560
rect 430448 267520 430454 267532
rect 457438 267520 457444 267532
rect 457496 267520 457502 267572
rect 459186 267520 459192 267572
rect 459244 267560 459250 267572
rect 464338 267560 464344 267572
rect 459244 267532 464344 267560
rect 459244 267520 459250 267532
rect 464338 267520 464344 267532
rect 464396 267520 464402 267572
rect 465166 267520 465172 267572
rect 465224 267560 465230 267572
rect 531498 267560 531504 267572
rect 465224 267532 531504 267560
rect 465224 267520 465230 267532
rect 531498 267520 531504 267532
rect 531556 267520 531562 267572
rect 531866 267520 531872 267572
rect 531924 267560 531930 267572
rect 538168 267560 538174 267572
rect 531924 267532 538174 267560
rect 531924 267520 531930 267532
rect 538168 267520 538174 267532
rect 538226 267520 538232 267572
rect 538306 267520 538312 267572
rect 538364 267560 538370 267572
rect 621658 267560 621664 267572
rect 538364 267532 621664 267560
rect 538364 267520 538370 267532
rect 621658 267520 621664 267532
rect 621716 267520 621722 267572
rect 107562 267384 107568 267436
rect 107620 267424 107626 267436
rect 167086 267424 167092 267436
rect 107620 267396 167092 267424
rect 107620 267384 107626 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 167730 267384 167736 267436
rect 167788 267424 167794 267436
rect 204346 267424 204352 267436
rect 167788 267396 204352 267424
rect 167788 267384 167794 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 211798 267384 211804 267436
rect 211856 267424 211862 267436
rect 222562 267424 222568 267436
rect 211856 267396 222568 267424
rect 211856 267384 211862 267396
rect 222562 267384 222568 267396
rect 222620 267384 222626 267436
rect 224218 267384 224224 267436
rect 224276 267424 224282 267436
rect 231670 267424 231676 267436
rect 224276 267396 231676 267424
rect 224276 267384 224282 267396
rect 231670 267384 231676 267396
rect 231728 267384 231734 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 246574 267424 246580 267436
rect 233936 267396 246580 267424
rect 233936 267384 233942 267396
rect 246574 267384 246580 267396
rect 246632 267384 246638 267436
rect 313642 267384 313648 267436
rect 313700 267424 313706 267436
rect 317782 267424 317788 267436
rect 313700 267396 317788 267424
rect 313700 267384 313706 267396
rect 317782 267384 317788 267396
rect 317840 267384 317846 267436
rect 334342 267384 334348 267436
rect 334400 267424 334406 267436
rect 342898 267424 342904 267436
rect 334400 267396 342904 267424
rect 334400 267384 334406 267396
rect 342898 267384 342904 267396
rect 342956 267384 342962 267436
rect 350902 267384 350908 267436
rect 350960 267424 350966 267436
rect 360746 267424 360752 267436
rect 350960 267396 360752 267424
rect 350960 267384 350966 267396
rect 360746 267384 360752 267396
rect 360804 267384 360810 267436
rect 363322 267384 363328 267436
rect 363380 267424 363386 267436
rect 370498 267424 370504 267436
rect 363380 267396 370504 267424
rect 363380 267384 363386 267396
rect 370498 267384 370504 267396
rect 370556 267384 370562 267436
rect 373258 267384 373264 267436
rect 373316 267424 373322 267436
rect 390462 267424 390468 267436
rect 373316 267396 390468 267424
rect 373316 267384 373322 267396
rect 390462 267384 390468 267396
rect 390520 267384 390526 267436
rect 390646 267384 390652 267436
rect 390704 267424 390710 267436
rect 401594 267424 401600 267436
rect 390704 267396 401600 267424
rect 390704 267384 390710 267396
rect 401594 267384 401600 267396
rect 401652 267384 401658 267436
rect 409598 267384 409604 267436
rect 409656 267424 409662 267436
rect 435358 267424 435364 267436
rect 409656 267396 435364 267424
rect 409656 267384 409662 267396
rect 435358 267384 435364 267396
rect 435416 267384 435422 267436
rect 445938 267384 445944 267436
rect 445996 267424 446002 267436
rect 450722 267424 450728 267436
rect 445996 267396 450728 267424
rect 445996 267384 446002 267396
rect 450722 267384 450728 267396
rect 450780 267384 450786 267436
rect 450906 267384 450912 267436
rect 450964 267424 450970 267436
rect 496446 267424 496452 267436
rect 450964 267396 496452 267424
rect 450964 267384 450970 267396
rect 496446 267384 496452 267396
rect 496504 267384 496510 267436
rect 496814 267384 496820 267436
rect 496872 267424 496878 267436
rect 507854 267424 507860 267436
rect 496872 267396 507860 267424
rect 496872 267384 496878 267396
rect 507854 267384 507860 267396
rect 507912 267384 507918 267436
rect 508038 267384 508044 267436
rect 508096 267424 508102 267436
rect 570598 267424 570604 267436
rect 508096 267396 570604 267424
rect 508096 267384 508102 267396
rect 570598 267384 570604 267396
rect 570656 267384 570662 267436
rect 571978 267384 571984 267436
rect 572036 267424 572042 267436
rect 602338 267424 602344 267436
rect 572036 267396 602344 267424
rect 572036 267384 572042 267396
rect 602338 267384 602344 267396
rect 602396 267384 602402 267436
rect 100662 267248 100668 267300
rect 100720 267288 100726 267300
rect 162118 267288 162124 267300
rect 100720 267260 162124 267288
rect 100720 267248 100726 267260
rect 162118 267248 162124 267260
rect 162176 267248 162182 267300
rect 166902 267248 166908 267300
rect 166960 267288 166966 267300
rect 174538 267288 174544 267300
rect 166960 267260 174544 267288
rect 166960 267248 166966 267260
rect 174538 267248 174544 267260
rect 174596 267248 174602 267300
rect 175090 267248 175096 267300
rect 175148 267288 175154 267300
rect 214282 267288 214288 267300
rect 175148 267260 214288 267288
rect 175148 267248 175154 267260
rect 214282 267248 214288 267260
rect 214340 267248 214346 267300
rect 220078 267248 220084 267300
rect 220136 267288 220142 267300
rect 239122 267288 239128 267300
rect 220136 267260 239128 267288
rect 220136 267248 220142 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 253658 267248 253664 267300
rect 253716 267288 253722 267300
rect 265618 267288 265624 267300
rect 253716 267260 265624 267288
rect 253716 267248 253722 267260
rect 265618 267248 265624 267260
rect 265676 267248 265682 267300
rect 312814 267248 312820 267300
rect 312872 267288 312878 267300
rect 316034 267288 316040 267300
rect 312872 267260 316040 267288
rect 312872 267248 312878 267260
rect 316034 267248 316040 267260
rect 316092 267248 316098 267300
rect 343450 267248 343456 267300
rect 343508 267288 343514 267300
rect 353938 267288 353944 267300
rect 343508 267260 353944 267288
rect 343508 267248 343514 267260
rect 353938 267248 353944 267260
rect 353996 267248 354002 267300
rect 368198 267248 368204 267300
rect 368256 267288 368262 267300
rect 385494 267288 385500 267300
rect 368256 267260 385500 267288
rect 368256 267248 368262 267260
rect 385494 267248 385500 267260
rect 385552 267248 385558 267300
rect 397086 267248 397092 267300
rect 397144 267288 397150 267300
rect 422294 267288 422300 267300
rect 397144 267260 422300 267288
rect 397144 267248 397150 267260
rect 422294 267248 422300 267260
rect 422352 267248 422358 267300
rect 427906 267248 427912 267300
rect 427964 267288 427970 267300
rect 427964 267260 446444 267288
rect 427964 267248 427970 267260
rect 73798 267112 73804 267164
rect 73856 267152 73862 267164
rect 141418 267152 141424 267164
rect 73856 267124 141424 267152
rect 73856 267112 73862 267124
rect 141418 267112 141424 267124
rect 141476 267112 141482 267164
rect 144546 267112 144552 267164
rect 144604 267152 144610 267164
rect 147398 267152 147404 267164
rect 144604 267124 147404 267152
rect 144604 267112 144610 267124
rect 147398 267112 147404 267124
rect 147456 267112 147462 267164
rect 147582 267112 147588 267164
rect 147640 267152 147646 267164
rect 149054 267152 149060 267164
rect 147640 267124 149060 267152
rect 147640 267112 147646 267124
rect 149054 267112 149060 267124
rect 149112 267112 149118 267164
rect 149882 267112 149888 267164
rect 149940 267152 149946 267164
rect 194410 267152 194416 267164
rect 149940 267124 194416 267152
rect 149940 267112 149946 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 199654 267112 199660 267164
rect 199712 267152 199718 267164
rect 218422 267152 218428 267164
rect 199712 267124 218428 267152
rect 199712 267112 199718 267124
rect 218422 267112 218428 267124
rect 218480 267112 218486 267164
rect 221458 267112 221464 267164
rect 221516 267152 221522 267164
rect 241606 267152 241612 267164
rect 221516 267124 241612 267152
rect 221516 267112 221522 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 335998 267112 336004 267164
rect 336056 267152 336062 267164
rect 347038 267152 347044 267164
rect 336056 267124 347044 267152
rect 336056 267112 336062 267124
rect 347038 267112 347044 267124
rect 347096 267112 347102 267164
rect 355870 267112 355876 267164
rect 355928 267152 355934 267164
rect 369118 267152 369124 267164
rect 355928 267124 369124 267152
rect 355928 267112 355934 267124
rect 369118 267112 369124 267124
rect 369176 267112 369182 267164
rect 375742 267112 375748 267164
rect 375800 267152 375806 267164
rect 393958 267152 393964 267164
rect 375800 267124 393964 267152
rect 375800 267112 375806 267124
rect 393958 267112 393964 267124
rect 394016 267112 394022 267164
rect 404722 267112 404728 267164
rect 404780 267152 404786 267164
rect 431954 267152 431960 267164
rect 404780 267124 431960 267152
rect 404780 267112 404786 267124
rect 431954 267112 431960 267124
rect 432012 267112 432018 267164
rect 432322 267112 432328 267164
rect 432380 267152 432386 267164
rect 440878 267152 440884 267164
rect 432380 267124 440884 267152
rect 432380 267112 432386 267124
rect 440878 267112 440884 267124
rect 440936 267112 440942 267164
rect 71038 266976 71044 267028
rect 71096 267016 71102 267028
rect 138106 267016 138112 267028
rect 71096 266988 138112 267016
rect 71096 266976 71102 266988
rect 138106 266976 138112 266988
rect 138164 266976 138170 267028
rect 141602 266976 141608 267028
rect 141660 267016 141666 267028
rect 184014 267016 184020 267028
rect 141660 266988 184020 267016
rect 141660 266976 141666 266988
rect 184014 266976 184020 266988
rect 184072 266976 184078 267028
rect 184198 266976 184204 267028
rect 184256 267016 184262 267028
rect 184256 266988 190454 267016
rect 184256 266976 184262 266988
rect 132402 266840 132408 266892
rect 132460 266880 132466 266892
rect 184474 266880 184480 266892
rect 132460 266852 184480 266880
rect 132460 266840 132466 266852
rect 184474 266840 184480 266852
rect 184532 266840 184538 266892
rect 190426 266880 190454 266988
rect 193858 266976 193864 267028
rect 193916 267016 193922 267028
rect 201862 267016 201868 267028
rect 193916 266988 201868 267016
rect 193916 266976 193922 266988
rect 201862 266976 201868 266988
rect 201920 266976 201926 267028
rect 227714 266976 227720 267028
rect 227772 267016 227778 267028
rect 234154 267016 234160 267028
rect 227772 266988 234160 267016
rect 227772 266976 227778 266988
rect 234154 266976 234160 266988
rect 234212 266976 234218 267028
rect 237282 266976 237288 267028
rect 237340 267016 237346 267028
rect 254026 267016 254032 267028
rect 237340 266988 254032 267016
rect 237340 266976 237346 266988
rect 254026 266976 254032 266988
rect 254084 266976 254090 267028
rect 271414 267016 271420 267028
rect 258046 266988 271420 267016
rect 258046 266892 258074 266988
rect 271414 266976 271420 266988
rect 271472 266976 271478 267028
rect 276658 266976 276664 267028
rect 276716 267016 276722 267028
rect 278038 267016 278044 267028
rect 276716 266988 278044 267016
rect 276716 266976 276722 266988
rect 278038 266976 278044 266988
rect 278096 266976 278102 267028
rect 286962 266976 286968 267028
rect 287020 267016 287026 267028
rect 291286 267016 291292 267028
rect 287020 266988 291292 267016
rect 287020 266976 287026 266988
rect 291286 266976 291292 266988
rect 291344 266976 291350 267028
rect 324406 266976 324412 267028
rect 324464 267016 324470 267028
rect 332502 267016 332508 267028
rect 324464 266988 332508 267016
rect 324464 266976 324470 266988
rect 332502 266976 332508 266988
rect 332560 266976 332566 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 355318 267016 355324 267028
rect 353444 266988 355324 267016
rect 353444 266976 353450 266988
rect 355318 266976 355324 266988
rect 355376 266976 355382 267028
rect 378226 266976 378232 267028
rect 378284 267016 378290 267028
rect 409138 267016 409144 267028
rect 378284 266988 409144 267016
rect 378284 266976 378290 266988
rect 409138 266976 409144 266988
rect 409196 266976 409202 267028
rect 421282 266976 421288 267028
rect 421340 267016 421346 267028
rect 422110 267016 422116 267028
rect 421340 266988 422116 267016
rect 421340 266976 421346 266988
rect 422110 266976 422116 266988
rect 422168 266976 422174 267028
rect 422294 266976 422300 267028
rect 422352 267016 422358 267028
rect 445938 267016 445944 267028
rect 422352 266988 445944 267016
rect 422352 266976 422358 266988
rect 445938 266976 445944 266988
rect 445996 266976 446002 267028
rect 446416 267016 446444 267260
rect 449434 267248 449440 267300
rect 449492 267288 449498 267300
rect 453298 267288 453304 267300
rect 449492 267260 453304 267288
rect 449492 267248 449498 267260
rect 453298 267248 453304 267260
rect 453356 267248 453362 267300
rect 455230 267248 455236 267300
rect 455288 267288 455294 267300
rect 511718 267288 511724 267300
rect 455288 267260 511724 267288
rect 455288 267248 455294 267260
rect 511718 267248 511724 267260
rect 511776 267248 511782 267300
rect 519170 267248 519176 267300
rect 519228 267288 519234 267300
rect 528508 267288 528514 267300
rect 519228 267260 528514 267288
rect 519228 267248 519234 267260
rect 528508 267248 528514 267260
rect 528566 267248 528572 267300
rect 528646 267248 528652 267300
rect 528704 267288 528710 267300
rect 613378 267288 613384 267300
rect 528704 267260 613384 267288
rect 528704 267248 528710 267260
rect 613378 267248 613384 267260
rect 613436 267248 613442 267300
rect 512196 267192 518894 267220
rect 450262 267112 450268 267164
rect 450320 267152 450326 267164
rect 507118 267152 507124 267164
rect 450320 267124 507124 267152
rect 450320 267112 450326 267124
rect 507118 267112 507124 267124
rect 507176 267112 507182 267164
rect 507394 267112 507400 267164
rect 507452 267152 507458 267164
rect 512196 267152 512224 267192
rect 507452 267124 512224 267152
rect 507452 267112 507458 267124
rect 512362 267044 512368 267096
rect 512420 267084 512426 267096
rect 514662 267084 514668 267096
rect 512420 267056 514668 267084
rect 512420 267044 512426 267056
rect 514662 267044 514668 267056
rect 514720 267044 514726 267096
rect 514846 267044 514852 267096
rect 514904 267084 514910 267096
rect 516318 267084 516324 267096
rect 514904 267056 516324 267084
rect 514904 267044 514910 267056
rect 516318 267044 516324 267056
rect 516376 267044 516382 267096
rect 516502 267044 516508 267096
rect 516560 267084 516566 267096
rect 517330 267084 517336 267096
rect 516560 267056 517336 267084
rect 516560 267044 516566 267056
rect 517330 267044 517336 267056
rect 517388 267044 517394 267096
rect 517514 267044 517520 267096
rect 517572 267084 517578 267096
rect 518710 267084 518716 267096
rect 517572 267056 518716 267084
rect 517572 267044 517578 267056
rect 518710 267044 518716 267056
rect 518768 267044 518774 267096
rect 451734 267016 451740 267028
rect 446416 266988 451740 267016
rect 451734 266976 451740 266988
rect 451792 266976 451798 267028
rect 454402 266976 454408 267028
rect 454460 267016 454466 267028
rect 459554 267016 459560 267028
rect 454460 266988 459560 267016
rect 454460 266976 454466 266988
rect 459554 266976 459560 266988
rect 459612 266976 459618 267028
rect 460198 266976 460204 267028
rect 460256 267016 460262 267028
rect 487246 267016 487252 267028
rect 460256 266988 487252 267016
rect 460256 266976 460262 266988
rect 487246 266976 487252 266988
rect 487304 266976 487310 267028
rect 487430 266976 487436 267028
rect 487488 267016 487494 267028
rect 487488 266988 489914 267016
rect 487488 266976 487494 266988
rect 209314 266880 209320 266892
rect 190426 266852 209320 266880
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 209498 266840 209504 266892
rect 209556 266880 209562 266892
rect 210970 266880 210976 266892
rect 209556 266852 210976 266880
rect 209556 266840 209562 266852
rect 210970 266840 210976 266852
rect 211028 266840 211034 266892
rect 257982 266840 257988 266892
rect 258040 266852 258074 266892
rect 258040 266840 258046 266852
rect 271138 266840 271144 266892
rect 271196 266880 271202 266892
rect 280522 266880 280528 266892
rect 271196 266852 280528 266880
rect 271196 266840 271202 266852
rect 280522 266840 280528 266852
rect 280580 266840 280586 266892
rect 316126 266840 316132 266892
rect 316184 266880 316190 266892
rect 320174 266880 320180 266892
rect 316184 266852 320180 266880
rect 316184 266840 316190 266852
rect 320174 266840 320180 266852
rect 320232 266840 320238 266892
rect 331858 266840 331864 266892
rect 331916 266880 331922 266892
rect 335630 266880 335636 266892
rect 331916 266852 335636 266880
rect 331916 266840 331922 266852
rect 335630 266840 335636 266852
rect 335688 266840 335694 266892
rect 342622 266840 342628 266892
rect 342680 266880 342686 266892
rect 356514 266880 356520 266892
rect 342680 266852 356520 266880
rect 342680 266840 342686 266852
rect 356514 266840 356520 266852
rect 356572 266840 356578 266892
rect 359182 266840 359188 266892
rect 359240 266880 359246 266892
rect 373074 266880 373080 266892
rect 359240 266852 373080 266880
rect 359240 266840 359246 266852
rect 373074 266840 373080 266852
rect 373132 266840 373138 266892
rect 388162 266840 388168 266892
rect 388220 266880 388226 266892
rect 396258 266880 396264 266892
rect 388220 266852 396264 266880
rect 388220 266840 388226 266852
rect 396258 266840 396264 266852
rect 396316 266840 396322 266892
rect 402238 266840 402244 266892
rect 402296 266880 402302 266892
rect 404998 266880 405004 266892
rect 402296 266852 405004 266880
rect 402296 266840 402302 266852
rect 404998 266840 405004 266852
rect 405056 266840 405062 266892
rect 412174 266840 412180 266892
rect 412232 266880 412238 266892
rect 428458 266880 428464 266892
rect 412232 266852 428464 266880
rect 412232 266840 412238 266852
rect 428458 266840 428464 266852
rect 428516 266840 428522 266892
rect 435358 266840 435364 266892
rect 435416 266880 435422 266892
rect 439682 266880 439688 266892
rect 435416 266852 439688 266880
rect 435416 266840 435422 266852
rect 439682 266840 439688 266852
rect 439740 266840 439746 266892
rect 441798 266840 441804 266892
rect 441856 266880 441862 266892
rect 447594 266880 447600 266892
rect 441856 266852 447600 266880
rect 441856 266840 441862 266852
rect 447594 266840 447600 266852
rect 447652 266840 447658 266892
rect 452746 266840 452752 266892
rect 452804 266880 452810 266892
rect 455874 266880 455880 266892
rect 452804 266852 455880 266880
rect 452804 266840 452810 266852
rect 455874 266840 455880 266852
rect 455932 266840 455938 266892
rect 461026 266840 461032 266892
rect 461084 266880 461090 266892
rect 470134 266880 470140 266892
rect 461084 266852 470140 266880
rect 461084 266840 461090 266852
rect 470134 266840 470140 266852
rect 470192 266840 470198 266892
rect 471790 266840 471796 266892
rect 471848 266880 471854 266892
rect 475562 266880 475568 266892
rect 471848 266852 475568 266880
rect 471848 266840 471854 266852
rect 475562 266840 475568 266852
rect 475620 266840 475626 266892
rect 477586 266840 477592 266892
rect 477644 266880 477650 266892
rect 489362 266880 489368 266892
rect 477644 266852 489368 266880
rect 477644 266840 477650 266852
rect 489362 266840 489368 266852
rect 489420 266840 489426 266892
rect 489886 266880 489914 266988
rect 492490 266976 492496 267028
rect 492548 267016 492554 267028
rect 500218 267016 500224 267028
rect 492548 266988 500224 267016
rect 492548 266976 492554 266988
rect 500218 266976 500224 266988
rect 500276 266976 500282 267028
rect 502426 266976 502432 267028
rect 502484 267016 502490 267028
rect 504910 267016 504916 267028
rect 502484 266988 504916 267016
rect 502484 266976 502490 266988
rect 504910 266976 504916 266988
rect 504968 266976 504974 267028
rect 509234 267016 509240 267028
rect 505066 266988 509240 267016
rect 495434 266880 495440 266892
rect 489886 266852 495440 266880
rect 495434 266840 495440 266852
rect 495492 266840 495498 266892
rect 495618 266840 495624 266892
rect 495676 266880 495682 266892
rect 505066 266880 505094 266988
rect 509234 266976 509240 266988
rect 509292 266976 509298 267028
rect 518710 266948 518716 266960
rect 509436 266920 518716 266948
rect 495676 266852 505094 266880
rect 495676 266840 495682 266852
rect 506566 266840 506572 266892
rect 506624 266880 506630 266892
rect 507670 266880 507676 266892
rect 506624 266852 507676 266880
rect 506624 266840 506630 266852
rect 507670 266840 507676 266852
rect 507728 266840 507734 266892
rect 507854 266840 507860 266892
rect 507912 266880 507918 266892
rect 509436 266880 509464 266920
rect 518710 266908 518716 266920
rect 518768 266908 518774 266960
rect 507912 266852 509464 266880
rect 518866 266880 518894 267192
rect 518986 267112 518992 267164
rect 519044 267152 519050 267164
rect 581270 267152 581276 267164
rect 519044 267124 581276 267152
rect 519044 267112 519050 267124
rect 581270 267112 581276 267124
rect 581328 267112 581334 267164
rect 581638 267112 581644 267164
rect 581696 267152 581702 267164
rect 622394 267152 622400 267164
rect 581696 267124 622400 267152
rect 581696 267112 581702 267124
rect 622394 267112 622400 267124
rect 622452 267112 622458 267164
rect 518986 266976 518992 267028
rect 519044 267016 519050 267028
rect 520182 267016 520188 267028
rect 519044 266988 520188 267016
rect 519044 266976 519050 266988
rect 520182 266976 520188 266988
rect 520240 266976 520246 267028
rect 523126 266976 523132 267028
rect 523184 267016 523190 267028
rect 524322 267016 524328 267028
rect 523184 266988 524328 267016
rect 523184 266976 523190 266988
rect 524322 266976 524328 266988
rect 524380 266976 524386 267028
rect 524782 266976 524788 267028
rect 524840 267016 524846 267028
rect 525518 267016 525524 267028
rect 524840 266988 525524 267016
rect 524840 266976 524846 266988
rect 525518 266976 525524 266988
rect 525576 266976 525582 267028
rect 527266 266976 527272 267028
rect 527324 267016 527330 267028
rect 528462 267016 528468 267028
rect 527324 266988 528468 267016
rect 527324 266976 527330 266988
rect 528462 266976 528468 266988
rect 528520 266976 528526 267028
rect 528738 266976 528744 267028
rect 528796 267016 528802 267028
rect 540422 267016 540428 267028
rect 528796 266988 540428 267016
rect 528796 266976 528802 266988
rect 540422 266976 540428 266988
rect 540480 266976 540486 267028
rect 540882 266976 540888 267028
rect 540940 267016 540946 267028
rect 629294 267016 629300 267028
rect 540940 266988 629300 267016
rect 540940 266976 540946 266988
rect 629294 266976 629300 266988
rect 629352 266976 629358 267028
rect 518866 266852 572024 266880
rect 507912 266840 507918 266852
rect 120718 266704 120724 266756
rect 120776 266744 120782 266756
rect 156414 266744 156420 266756
rect 120776 266716 156420 266744
rect 120776 266704 120782 266716
rect 156414 266704 156420 266716
rect 156472 266704 156478 266756
rect 156598 266704 156604 266756
rect 156656 266744 156662 266756
rect 159634 266744 159640 266756
rect 156656 266716 159640 266744
rect 156656 266704 156662 266716
rect 159634 266704 159640 266716
rect 159692 266704 159698 266756
rect 169018 266704 169024 266756
rect 169076 266744 169082 266756
rect 172054 266744 172060 266756
rect 169076 266716 172060 266744
rect 169076 266704 169082 266716
rect 172054 266704 172060 266716
rect 172112 266704 172118 266756
rect 184014 266704 184020 266756
rect 184072 266744 184078 266756
rect 189442 266744 189448 266756
rect 184072 266716 189448 266744
rect 184072 266704 184078 266716
rect 189442 266704 189448 266716
rect 189500 266704 189506 266756
rect 206278 266704 206284 266756
rect 206336 266744 206342 266756
rect 228358 266744 228364 266756
rect 206336 266716 228364 266744
rect 206336 266704 206342 266716
rect 228358 266704 228364 266716
rect 228416 266704 228422 266756
rect 240686 266704 240692 266756
rect 240744 266744 240750 266756
rect 245746 266744 245752 266756
rect 240744 266716 245752 266744
rect 240744 266704 240750 266716
rect 245746 266704 245752 266716
rect 245804 266704 245810 266756
rect 249058 266704 249064 266756
rect 249116 266744 249122 266756
rect 251542 266744 251548 266756
rect 249116 266716 251548 266744
rect 249116 266704 249122 266716
rect 251542 266704 251548 266716
rect 251600 266704 251606 266756
rect 265066 266704 265072 266756
rect 265124 266744 265130 266756
rect 268930 266744 268936 266756
rect 265124 266716 268936 266744
rect 265124 266704 265130 266716
rect 268930 266704 268936 266716
rect 268988 266704 268994 266756
rect 320266 266704 320272 266756
rect 320324 266744 320330 266756
rect 327074 266744 327080 266756
rect 320324 266716 327080 266744
rect 320324 266704 320330 266716
rect 327074 266704 327080 266716
rect 327132 266704 327138 266756
rect 355042 266704 355048 266756
rect 355100 266744 355106 266756
rect 359918 266744 359924 266756
rect 355100 266716 359924 266744
rect 355100 266704 355106 266716
rect 359918 266704 359924 266716
rect 359976 266704 359982 266756
rect 398098 266704 398104 266756
rect 398156 266744 398162 266756
rect 411898 266744 411904 266756
rect 398156 266716 411904 266744
rect 398156 266704 398162 266716
rect 411898 266704 411904 266716
rect 411956 266704 411962 266756
rect 413002 266704 413008 266756
rect 413060 266744 413066 266756
rect 428274 266744 428280 266756
rect 413060 266716 428280 266744
rect 413060 266704 413066 266716
rect 428274 266704 428280 266716
rect 428332 266704 428338 266756
rect 428734 266704 428740 266756
rect 428792 266744 428798 266756
rect 465718 266744 465724 266756
rect 428792 266716 465724 266744
rect 428792 266704 428798 266716
rect 465718 266704 465724 266716
rect 465776 266704 465782 266756
rect 476574 266744 476580 266756
rect 466426 266716 476580 266744
rect 138658 266568 138664 266620
rect 138716 266608 138722 266620
rect 138716 266580 145328 266608
rect 138716 266568 138722 266580
rect 119798 266432 119804 266484
rect 119856 266472 119862 266484
rect 144914 266472 144920 266484
rect 119856 266444 144920 266472
rect 119856 266432 119862 266444
rect 144914 266432 144920 266444
rect 144972 266432 144978 266484
rect 145300 266404 145328 266580
rect 149054 266568 149060 266620
rect 149112 266608 149118 266620
rect 179506 266608 179512 266620
rect 149112 266580 179512 266608
rect 149112 266568 149118 266580
rect 179506 266568 179512 266580
rect 179564 266568 179570 266620
rect 213822 266568 213828 266620
rect 213880 266608 213886 266620
rect 220078 266608 220084 266620
rect 213880 266580 220084 266608
rect 213880 266568 213886 266580
rect 220078 266568 220084 266580
rect 220136 266568 220142 266620
rect 245102 266568 245108 266620
rect 245160 266608 245166 266620
rect 249058 266608 249064 266620
rect 245160 266580 249064 266608
rect 245160 266568 245166 266580
rect 249058 266568 249064 266580
rect 249116 266568 249122 266620
rect 358354 266568 358360 266620
rect 358412 266608 358418 266620
rect 362218 266608 362224 266620
rect 358412 266580 362224 266608
rect 358412 266568 358418 266580
rect 362218 266568 362224 266580
rect 362276 266568 362282 266620
rect 422938 266568 422944 266620
rect 422996 266608 423002 266620
rect 441798 266608 441804 266620
rect 422996 266580 441804 266608
rect 422996 266568 423002 266580
rect 441798 266568 441804 266580
rect 441856 266568 441862 266620
rect 441982 266568 441988 266620
rect 442040 266608 442046 266620
rect 443638 266608 443644 266620
rect 442040 266580 443644 266608
rect 442040 266568 442046 266580
rect 443638 266568 443644 266580
rect 443696 266568 443702 266620
rect 444466 266568 444472 266620
rect 444524 266608 444530 266620
rect 445662 266608 445668 266620
rect 444524 266580 445668 266608
rect 444524 266568 444530 266580
rect 445662 266568 445668 266580
rect 445720 266568 445726 266620
rect 445846 266568 445852 266620
rect 445904 266608 445910 266620
rect 450906 266608 450912 266620
rect 445904 266580 450912 266608
rect 445904 266568 445910 266580
rect 450906 266568 450912 266580
rect 450964 266568 450970 266620
rect 451918 266568 451924 266620
rect 451976 266608 451982 266620
rect 454678 266608 454684 266620
rect 451976 266580 454684 266608
rect 451976 266568 451982 266580
rect 454678 266568 454684 266580
rect 454736 266568 454742 266620
rect 456886 266568 456892 266620
rect 456944 266608 456950 266620
rect 458082 266608 458088 266620
rect 456944 266580 458088 266608
rect 456944 266568 456950 266580
rect 458082 266568 458088 266580
rect 458140 266568 458146 266620
rect 458542 266568 458548 266620
rect 458600 266608 458606 266620
rect 459370 266608 459376 266620
rect 458600 266580 459376 266608
rect 458600 266568 458606 266580
rect 459370 266568 459376 266580
rect 459428 266568 459434 266620
rect 459554 266568 459560 266620
rect 459612 266608 459618 266620
rect 461578 266608 461584 266620
rect 459612 266580 461584 266608
rect 459612 266568 459618 266580
rect 461578 266568 461584 266580
rect 461636 266568 461642 266620
rect 145558 266500 145564 266552
rect 145616 266540 145622 266552
rect 148870 266540 148876 266552
rect 145616 266512 148876 266540
rect 145616 266500 145622 266512
rect 148870 266500 148876 266512
rect 148928 266500 148934 266552
rect 269114 266500 269120 266552
rect 269172 266540 269178 266552
rect 276382 266540 276388 266552
rect 269172 266512 276388 266540
rect 269172 266500 269178 266512
rect 276382 266500 276388 266512
rect 276440 266500 276446 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 330202 266500 330208 266552
rect 330260 266540 330266 266552
rect 334802 266540 334808 266552
rect 330260 266512 334808 266540
rect 330260 266500 330266 266512
rect 334802 266500 334808 266512
rect 334860 266500 334866 266552
rect 346762 266500 346768 266552
rect 346820 266540 346826 266552
rect 351638 266540 351644 266552
rect 346820 266512 351644 266540
rect 346820 266500 346826 266512
rect 351638 266500 351644 266512
rect 351696 266500 351702 266552
rect 380526 266500 380532 266552
rect 380584 266540 380590 266552
rect 382918 266540 382924 266552
rect 380584 266512 382924 266540
rect 380584 266500 380590 266512
rect 382918 266500 382924 266512
rect 382976 266500 382982 266552
rect 394786 266500 394792 266552
rect 394844 266540 394850 266552
rect 397638 266540 397644 266552
rect 394844 266512 397644 266540
rect 394844 266500 394850 266512
rect 397638 266500 397644 266512
rect 397696 266500 397702 266552
rect 151078 266432 151084 266484
rect 151136 266472 151142 266484
rect 172882 266472 172888 266484
rect 151136 266444 172888 266472
rect 151136 266432 151142 266444
rect 172882 266432 172888 266444
rect 172940 266432 172946 266484
rect 361666 266432 361672 266484
rect 361724 266472 361730 266484
rect 362770 266472 362776 266484
rect 361724 266444 362776 266472
rect 361724 266432 361730 266444
rect 362770 266432 362776 266444
rect 362828 266432 362834 266484
rect 439682 266432 439688 266484
rect 439740 266472 439746 266484
rect 466426 266472 466454 266716
rect 476574 266704 476580 266716
rect 476632 266704 476638 266756
rect 481726 266704 481732 266756
rect 481784 266744 481790 266756
rect 484854 266744 484860 266756
rect 481784 266716 484860 266744
rect 481784 266704 481790 266716
rect 484854 266704 484860 266716
rect 484912 266704 484918 266756
rect 485038 266704 485044 266756
rect 485096 266744 485102 266756
rect 496814 266744 496820 266756
rect 485096 266716 496820 266744
rect 485096 266704 485102 266716
rect 496814 266704 496820 266716
rect 496872 266704 496878 266756
rect 496998 266704 497004 266756
rect 497056 266744 497062 266756
rect 549254 266744 549260 266756
rect 497056 266716 549260 266744
rect 497056 266704 497062 266716
rect 549254 266704 549260 266716
rect 549312 266704 549318 266756
rect 571996 266744 572024 266852
rect 572162 266840 572168 266892
rect 572220 266880 572226 266892
rect 581638 266880 581644 266892
rect 572220 266852 581644 266880
rect 572220 266840 572226 266852
rect 581638 266840 581644 266852
rect 581696 266840 581702 266892
rect 578878 266744 578884 266756
rect 557506 266716 567194 266744
rect 571996 266716 578884 266744
rect 470134 266568 470140 266620
rect 470192 266608 470198 266620
rect 528738 266608 528744 266620
rect 470192 266580 528744 266608
rect 470192 266568 470198 266580
rect 528738 266568 528744 266580
rect 528796 266568 528802 266620
rect 528922 266568 528928 266620
rect 528980 266608 528986 266620
rect 529842 266608 529848 266620
rect 528980 266580 529848 266608
rect 528980 266568 528986 266580
rect 529842 266568 529848 266580
rect 529900 266568 529906 266620
rect 532234 266568 532240 266620
rect 532292 266608 532298 266620
rect 540238 266608 540244 266620
rect 532292 266580 540244 266608
rect 532292 266568 532298 266580
rect 540238 266568 540244 266580
rect 540296 266568 540302 266620
rect 540422 266568 540428 266620
rect 540480 266608 540486 266620
rect 557506 266608 557534 266716
rect 540480 266580 557534 266608
rect 567166 266608 567194 266716
rect 578878 266704 578884 266716
rect 578936 266704 578942 266756
rect 572162 266608 572168 266620
rect 567166 266580 572168 266608
rect 540480 266568 540486 266580
rect 572162 266568 572168 266580
rect 572220 266568 572226 266620
rect 439740 266444 466454 266472
rect 439740 266432 439746 266444
rect 469306 266432 469312 266484
rect 469364 266472 469370 266484
rect 474734 266472 474740 266484
rect 469364 266444 474740 266472
rect 469364 266432 469370 266444
rect 474734 266432 474740 266444
rect 474792 266432 474798 266484
rect 475930 266432 475936 266484
rect 475988 266472 475994 266484
rect 485038 266472 485044 266484
rect 475988 266444 485044 266472
rect 475988 266432 475994 266444
rect 485038 266432 485044 266444
rect 485096 266432 485102 266484
rect 487246 266432 487252 266484
rect 487304 266472 487310 266484
rect 493318 266472 493324 266484
rect 487304 266444 493324 266472
rect 487304 266432 487310 266444
rect 493318 266432 493324 266444
rect 493376 266432 493382 266484
rect 500218 266432 500224 266484
rect 500276 266472 500282 266484
rect 558914 266472 558920 266484
rect 500276 266444 558920 266472
rect 500276 266432 500282 266444
rect 558914 266432 558920 266444
rect 558972 266432 558978 266484
rect 147214 266404 147220 266416
rect 145300 266376 147220 266404
rect 147214 266364 147220 266376
rect 147272 266364 147278 266416
rect 148318 266364 148324 266416
rect 148376 266404 148382 266416
rect 149698 266404 149704 266416
rect 148376 266376 149704 266404
rect 148376 266364 148382 266376
rect 149698 266364 149704 266376
rect 149756 266364 149762 266416
rect 182174 266364 182180 266416
rect 182232 266404 182238 266416
rect 186130 266404 186136 266416
rect 182232 266376 186136 266404
rect 182232 266364 182238 266376
rect 186130 266364 186136 266376
rect 186188 266364 186194 266416
rect 202138 266364 202144 266416
rect 202196 266404 202202 266416
rect 206830 266404 206836 266416
rect 202196 266376 206836 266404
rect 202196 266364 202202 266376
rect 206830 266364 206836 266376
rect 206888 266364 206894 266416
rect 210418 266364 210424 266416
rect 210476 266404 210482 266416
rect 211798 266404 211804 266416
rect 210476 266376 211804 266404
rect 210476 266364 210482 266376
rect 211798 266364 211804 266376
rect 211856 266364 211862 266416
rect 222838 266364 222844 266416
rect 222896 266404 222902 266416
rect 224218 266404 224224 266416
rect 222896 266376 224224 266404
rect 222896 266364 222902 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 230750 266364 230756 266416
rect 230808 266404 230814 266416
rect 236638 266404 236644 266416
rect 230808 266376 236644 266404
rect 230808 266364 230814 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 242250 266364 242256 266416
rect 242308 266404 242314 266416
rect 243262 266404 243268 266416
rect 242308 266376 243268 266404
rect 242308 266364 242314 266376
rect 243262 266364 243268 266376
rect 243320 266364 243326 266416
rect 252002 266364 252008 266416
rect 252060 266404 252066 266416
rect 257338 266404 257344 266416
rect 252060 266376 257344 266404
rect 252060 266364 252066 266376
rect 257338 266364 257344 266376
rect 257396 266364 257402 266416
rect 268378 266364 268384 266416
rect 268436 266404 268442 266416
rect 273070 266404 273076 266416
rect 268436 266376 273076 266404
rect 268436 266364 268442 266376
rect 273070 266364 273076 266376
rect 273128 266364 273134 266416
rect 278590 266364 278596 266416
rect 278648 266404 278654 266416
rect 286318 266404 286324 266416
rect 278648 266376 286324 266404
rect 278648 266364 278654 266376
rect 286318 266364 286324 266376
rect 286376 266364 286382 266416
rect 290458 266364 290464 266416
rect 290516 266404 290522 266416
rect 292942 266404 292948 266416
rect 290516 266376 292948 266404
rect 290516 266364 290522 266376
rect 292942 266364 292948 266376
rect 293000 266364 293006 266416
rect 293862 266364 293868 266416
rect 293920 266404 293926 266416
rect 296254 266404 296260 266416
rect 293920 266376 296260 266404
rect 293920 266364 293926 266376
rect 296254 266364 296260 266376
rect 296312 266364 296318 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 312354 266364 312360 266416
rect 312412 266404 312418 266416
rect 314654 266404 314660 266416
rect 312412 266376 314660 266404
rect 312412 266364 312418 266376
rect 314654 266364 314660 266376
rect 314712 266364 314718 266416
rect 317782 266364 317788 266416
rect 317840 266404 317846 266416
rect 323118 266404 323124 266416
rect 317840 266376 323124 266404
rect 317840 266364 317846 266376
rect 323118 266364 323124 266376
rect 323176 266364 323182 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333606 266404 333612 266416
rect 332744 266376 333612 266404
rect 332744 266364 332750 266376
rect 333606 266364 333612 266376
rect 333664 266364 333670 266416
rect 340966 266364 340972 266416
rect 341024 266404 341030 266416
rect 342162 266404 342168 266416
rect 341024 266376 342168 266404
rect 341024 266364 341030 266376
rect 342162 266364 342168 266376
rect 342220 266364 342226 266416
rect 345106 266364 345112 266416
rect 345164 266404 345170 266416
rect 346118 266404 346124 266416
rect 345164 266376 346124 266404
rect 345164 266364 345170 266376
rect 346118 266364 346124 266376
rect 346176 266364 346182 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350258 266404 350264 266416
rect 349304 266376 350264 266404
rect 349304 266364 349310 266376
rect 350258 266364 350264 266376
rect 350316 266364 350322 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 358630 266404 358636 266416
rect 357584 266376 358636 266404
rect 357584 266364 357590 266376
rect 358630 266364 358636 266376
rect 358688 266364 358694 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368382 266404 368388 266416
rect 367520 266376 368388 266404
rect 367520 266364 367526 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375098 266404 375104 266416
rect 374144 266376 375104 266404
rect 374144 266364 374150 266376
rect 375098 266364 375104 266376
rect 375156 266364 375162 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 380710 266404 380716 266416
rect 379940 266376 380716 266404
rect 379940 266364 379946 266376
rect 380710 266364 380716 266376
rect 380768 266364 380774 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412450 266404 412456 266416
rect 411404 266376 412456 266404
rect 411404 266364 411410 266376
rect 412450 266364 412456 266376
rect 412508 266364 412514 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 423766 266364 423772 266416
rect 423824 266404 423830 266416
rect 424962 266404 424968 266416
rect 423824 266376 424968 266404
rect 423824 266364 423830 266376
rect 424962 266364 424968 266376
rect 425020 266364 425026 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 433702 266364 433708 266416
rect 433760 266404 433766 266416
rect 434622 266404 434628 266416
rect 433760 266376 434628 266404
rect 433760 266364 433766 266376
rect 434622 266364 434628 266376
rect 434680 266364 434686 266416
rect 437842 266364 437848 266416
rect 437900 266404 437906 266416
rect 439498 266404 439504 266416
rect 437900 266376 439504 266404
rect 437900 266364 437906 266376
rect 439498 266364 439504 266376
rect 439556 266364 439562 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 487062 266404 487068 266416
rect 485924 266376 487068 266404
rect 485924 266364 485930 266376
rect 487062 266364 487068 266376
rect 487120 266364 487126 266416
rect 496998 266404 497004 266416
rect 493520 266376 497004 266404
rect 490282 266296 490288 266348
rect 490340 266336 490346 266348
rect 493520 266336 493548 266376
rect 496998 266364 497004 266376
rect 497056 266364 497062 266416
rect 497200 266376 500080 266404
rect 490340 266308 493548 266336
rect 490340 266296 490346 266308
rect 495434 266228 495440 266280
rect 495492 266268 495498 266280
rect 497200 266268 497228 266376
rect 500052 266336 500080 266376
rect 502610 266336 502616 266348
rect 500052 266308 502616 266336
rect 502610 266296 502616 266308
rect 502668 266296 502674 266348
rect 495492 266240 497228 266268
rect 495492 266228 495498 266240
rect 498562 266160 498568 266212
rect 498620 266200 498626 266212
rect 500954 266200 500960 266212
rect 498620 266172 500960 266200
rect 498620 266160 498626 266172
rect 500954 266160 500960 266172
rect 501012 266160 501018 266212
rect 475102 266024 475108 266076
rect 475160 266064 475166 266076
rect 547874 266064 547880 266076
rect 475160 266036 547880 266064
rect 475160 266024 475166 266036
rect 547874 266024 547880 266036
rect 547932 266024 547938 266076
rect 485038 265888 485044 265940
rect 485096 265928 485102 265940
rect 561674 265928 561680 265940
rect 485096 265900 561680 265928
rect 485096 265888 485102 265900
rect 561674 265888 561680 265900
rect 561732 265888 561738 265940
rect 494974 265752 494980 265804
rect 495032 265792 495038 265804
rect 575842 265792 575848 265804
rect 495032 265764 575848 265792
rect 495032 265752 495038 265764
rect 575842 265752 575848 265764
rect 575900 265752 575906 265804
rect 187694 265616 187700 265668
rect 187752 265656 187758 265668
rect 188246 265656 188252 265668
rect 187752 265628 188252 265656
rect 187752 265616 187758 265628
rect 188246 265616 188252 265628
rect 188304 265616 188310 265668
rect 247218 265616 247224 265668
rect 247276 265656 247282 265668
rect 247862 265656 247868 265668
rect 247276 265628 247868 265656
rect 247276 265616 247282 265628
rect 247862 265616 247868 265628
rect 247920 265616 247926 265668
rect 255498 265616 255504 265668
rect 255556 265656 255562 265668
rect 256142 265656 256148 265668
rect 255556 265628 256148 265656
rect 255556 265616 255562 265628
rect 256142 265616 256148 265628
rect 256200 265616 256206 265668
rect 259546 265616 259552 265668
rect 259604 265656 259610 265668
rect 260374 265656 260380 265668
rect 259604 265628 260380 265656
rect 259604 265616 259610 265628
rect 260374 265616 260380 265628
rect 260432 265616 260438 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 480070 265616 480076 265668
rect 480128 265656 480134 265668
rect 554774 265656 554780 265668
rect 480128 265628 554780 265656
rect 480128 265616 480134 265628
rect 554774 265616 554780 265628
rect 554832 265616 554838 265668
rect 558178 265616 558184 265668
rect 558236 265656 558242 265668
rect 647234 265656 647240 265668
rect 558236 265628 647240 265656
rect 558236 265616 558242 265628
rect 647234 265616 647240 265628
rect 647292 265616 647298 265668
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 565078 259468 565084 259480
rect 554372 259440 565084 259468
rect 554372 259428 554378 259440
rect 565078 259428 565084 259440
rect 565136 259428 565142 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 560938 256748 560944 256760
rect 554004 256720 560944 256748
rect 554004 256708 554010 256720
rect 560938 256708 560944 256720
rect 560996 256708 561002 256760
rect 553486 255552 553492 255604
rect 553544 255592 553550 255604
rect 555418 255592 555424 255604
rect 553544 255564 555424 255592
rect 553544 255552 553550 255564
rect 555418 255552 555424 255564
rect 555476 255552 555482 255604
rect 39022 252968 39028 253020
rect 39080 253008 39086 253020
rect 41506 253008 41512 253020
rect 39080 252980 41512 253008
rect 39080 252968 39086 252980
rect 41506 252968 41512 252980
rect 41564 252968 41570 253020
rect 35802 252832 35808 252884
rect 35860 252872 35866 252884
rect 40678 252872 40684 252884
rect 35860 252844 40684 252872
rect 35860 252832 35866 252844
rect 40678 252832 40684 252844
rect 40736 252832 40742 252884
rect 35618 252696 35624 252748
rect 35676 252736 35682 252748
rect 39022 252736 39028 252748
rect 35676 252708 39028 252736
rect 35676 252696 35682 252708
rect 39022 252696 39028 252708
rect 39080 252696 39086 252748
rect 39224 252640 40080 252668
rect 35434 252560 35440 252612
rect 35492 252600 35498 252612
rect 39224 252600 39252 252640
rect 35492 252572 39252 252600
rect 35492 252560 35498 252572
rect 40052 252532 40080 252640
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 563698 252600 563704 252612
rect 554464 252572 563704 252600
rect 554464 252560 554470 252572
rect 563698 252560 563704 252572
rect 563756 252560 563762 252612
rect 41690 252532 41696 252544
rect 40052 252504 41696 252532
rect 41690 252492 41696 252504
rect 41748 252492 41754 252544
rect 676030 252356 676036 252408
rect 676088 252396 676094 252408
rect 678422 252396 678428 252408
rect 676088 252368 678428 252396
rect 676088 252356 676094 252368
rect 678422 252356 678428 252368
rect 678480 252356 678486 252408
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 36538 251240 36544 251252
rect 35860 251212 36544 251240
rect 35860 251200 35866 251212
rect 36538 251200 36544 251212
rect 36596 251200 36602 251252
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 553854 246304 553860 246356
rect 553912 246344 553918 246356
rect 632698 246344 632704 246356
rect 553912 246316 632704 246344
rect 553912 246304 553918 246316
rect 632698 246304 632704 246316
rect 632756 246304 632762 246356
rect 554406 245624 554412 245676
rect 554464 245664 554470 245676
rect 598198 245664 598204 245676
rect 554464 245636 598204 245664
rect 554464 245624 554470 245636
rect 598198 245624 598204 245636
rect 598256 245624 598262 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 623038 244304 623044 244316
rect 554556 244276 623044 244304
rect 554556 244264 554562 244276
rect 623038 244264 623044 244276
rect 623096 244264 623102 244316
rect 36538 242836 36544 242888
rect 36596 242876 36602 242888
rect 41690 242876 41696 242888
rect 36596 242848 41696 242876
rect 36596 242836 36602 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 587158 242156 587164 242208
rect 587216 242196 587222 242208
rect 648614 242196 648620 242208
rect 587216 242168 648620 242196
rect 587216 242156 587222 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553946 241476 553952 241528
rect 554004 241516 554010 241528
rect 631318 241516 631324 241528
rect 554004 241488 631324 241516
rect 554004 241476 554010 241488
rect 631318 241476 631324 241488
rect 631376 241476 631382 241528
rect 553854 240116 553860 240168
rect 553912 240156 553918 240168
rect 577498 240156 577504 240168
rect 553912 240128 577504 240156
rect 553912 240116 553918 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 587158 238728 587164 238740
rect 554372 238700 587164 238728
rect 554372 238688 554378 238700
rect 587158 238688 587164 238700
rect 587216 238688 587222 238740
rect 671890 237804 671896 237856
rect 671948 237844 671954 237856
rect 672756 237844 672784 238102
rect 671948 237816 672784 237844
rect 671948 237804 671954 237816
rect 672258 237600 672264 237652
rect 672316 237640 672322 237652
rect 672874 237640 672902 237898
rect 672316 237612 672902 237640
rect 672316 237600 672322 237612
rect 668762 237192 668768 237244
rect 668820 237232 668826 237244
rect 672966 237232 672994 237694
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 668820 237204 672994 237232
rect 668820 237192 668826 237204
rect 671522 236988 671528 237040
rect 671580 237028 671586 237040
rect 673196 237028 673224 237286
rect 673304 237108 673356 237114
rect 673304 237050 673356 237056
rect 671580 237000 673224 237028
rect 671580 236988 671586 237000
rect 672902 236852 672908 236904
rect 672960 236892 672966 236904
rect 673270 236892 673276 236904
rect 672960 236864 673276 236892
rect 672960 236852 672966 236864
rect 673270 236852 673276 236864
rect 673328 236852 673334 236904
rect 673426 236564 673454 236878
rect 673528 236700 673580 236706
rect 673528 236642 673580 236648
rect 673426 236524 673460 236564
rect 673454 236512 673460 236524
rect 673512 236512 673518 236564
rect 672534 236172 672540 236224
rect 672592 236212 672598 236224
rect 673656 236212 673684 236470
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 672592 236184 673684 236212
rect 672592 236172 672598 236184
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 671706 236036 671712 236088
rect 671764 236076 671770 236088
rect 671764 236048 673900 236076
rect 671764 236036 671770 236048
rect 673730 235900 673736 235952
rect 673788 235940 673794 235952
rect 673788 235912 673992 235940
rect 673788 235900 673794 235912
rect 672902 235696 672908 235748
rect 672960 235736 672966 235748
rect 672960 235708 674114 235736
rect 672960 235696 672966 235708
rect 669774 235492 669780 235544
rect 669832 235532 669838 235544
rect 669832 235504 674222 235532
rect 669832 235492 669838 235504
rect 668118 235288 668124 235340
rect 668176 235328 668182 235340
rect 668176 235300 674338 235328
rect 668176 235288 668182 235300
rect 598198 235220 598204 235272
rect 598256 235260 598262 235272
rect 633618 235260 633624 235272
rect 598256 235232 633624 235260
rect 598256 235220 598262 235232
rect 633618 235220 633624 235232
rect 633676 235220 633682 235272
rect 674306 234948 674312 235000
rect 674364 234988 674370 235000
rect 674438 234988 674466 235110
rect 674364 234960 674466 234988
rect 674364 234948 674370 234960
rect 672810 234812 672816 234864
rect 672868 234852 672874 234864
rect 674548 234852 674576 234906
rect 672868 234824 674576 234852
rect 672868 234812 672874 234824
rect 674576 234688 674682 234716
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 671338 234540 671344 234592
rect 671396 234580 671402 234592
rect 671396 234552 672074 234580
rect 671396 234540 671402 234552
rect 668394 234404 668400 234456
rect 668452 234444 668458 234456
rect 671890 234444 671896 234456
rect 668452 234416 671896 234444
rect 668452 234404 668458 234416
rect 671890 234404 671896 234416
rect 671948 234404 671954 234456
rect 672046 234376 672074 234552
rect 674576 234376 674604 234688
rect 675846 234540 675852 234592
rect 675904 234580 675910 234592
rect 678238 234580 678244 234592
rect 675904 234552 678244 234580
rect 675904 234540 675910 234552
rect 678238 234540 678244 234552
rect 678296 234540 678302 234592
rect 674748 234524 674800 234530
rect 674748 234466 674800 234472
rect 672046 234348 674604 234376
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 667934 234064 667940 234116
rect 667992 234104 667998 234116
rect 667992 234076 675004 234104
rect 667992 234064 667998 234076
rect 675236 233912 675288 233918
rect 670786 233860 670792 233912
rect 670844 233900 670850 233912
rect 670844 233872 675122 233900
rect 670844 233860 670850 233872
rect 675236 233854 675288 233860
rect 675846 233792 675852 233844
rect 675904 233832 675910 233844
rect 677778 233832 677784 233844
rect 675904 233804 677784 233832
rect 675904 233792 675910 233804
rect 677778 233792 677784 233804
rect 677836 233792 677842 233844
rect 675846 233520 675852 233572
rect 675904 233560 675910 233572
rect 683482 233560 683488 233572
rect 675904 233532 683488 233560
rect 675904 233520 675910 233532
rect 683482 233520 683488 233532
rect 683540 233520 683546 233572
rect 670602 233452 670608 233504
rect 670660 233492 670666 233504
rect 670660 233464 675372 233492
rect 670660 233452 670666 233464
rect 669590 233316 669596 233368
rect 669648 233356 669654 233368
rect 671338 233356 671344 233368
rect 669648 233328 671344 233356
rect 669648 233316 669654 233328
rect 671338 233316 671344 233328
rect 671396 233316 671402 233368
rect 676030 233248 676036 233300
rect 676088 233288 676094 233300
rect 678422 233288 678428 233300
rect 676088 233260 678428 233288
rect 676088 233248 676094 233260
rect 678422 233248 678428 233260
rect 678480 233248 678486 233300
rect 671338 233180 671344 233232
rect 671396 233220 671402 233232
rect 673086 233220 673092 233232
rect 671396 233192 673092 233220
rect 671396 233180 671402 233192
rect 673086 233180 673092 233192
rect 673144 233180 673150 233232
rect 671154 233044 671160 233096
rect 671212 233084 671218 233096
rect 674834 233084 674840 233096
rect 671212 233056 674840 233084
rect 671212 233044 671218 233056
rect 674834 233044 674840 233056
rect 674892 233044 674898 233096
rect 652018 232500 652024 232552
rect 652076 232540 652082 232552
rect 675478 232540 675484 232552
rect 652076 232512 675484 232540
rect 652076 232500 652082 232512
rect 675478 232500 675484 232512
rect 675536 232500 675542 232552
rect 662322 232364 662328 232416
rect 662380 232404 662386 232416
rect 662380 232376 663794 232404
rect 662380 232364 662386 232376
rect 663766 232336 663794 232376
rect 675846 232364 675852 232416
rect 675904 232404 675910 232416
rect 679250 232404 679256 232416
rect 675904 232376 679256 232404
rect 675904 232364 675910 232376
rect 679250 232364 679256 232376
rect 679308 232364 679314 232416
rect 672258 232336 672264 232348
rect 663766 232308 672264 232336
rect 672258 232296 672264 232308
rect 672316 232296 672322 232348
rect 665082 232160 665088 232212
rect 665140 232200 665146 232212
rect 665140 232172 675556 232200
rect 665140 232160 665146 232172
rect 672258 231956 672264 232008
rect 672316 231996 672322 232008
rect 672316 231968 675372 231996
rect 672316 231956 672322 231968
rect 675180 231804 675232 231810
rect 675180 231746 675232 231752
rect 675070 231600 675122 231606
rect 668210 231548 668216 231600
rect 668268 231588 668274 231600
rect 669406 231588 669412 231600
rect 668268 231560 669412 231588
rect 668268 231548 668274 231560
rect 669406 231548 669412 231560
rect 669464 231548 669470 231600
rect 675070 231542 675122 231548
rect 673454 231480 673460 231532
rect 673512 231520 673518 231532
rect 674742 231520 674748 231532
rect 673512 231492 674748 231520
rect 673512 231480 673518 231492
rect 674742 231480 674748 231492
rect 674800 231480 674806 231532
rect 674956 231328 675008 231334
rect 674956 231270 675008 231276
rect 674840 231260 674892 231266
rect 675846 231208 675852 231260
rect 675904 231248 675910 231260
rect 677594 231248 677600 231260
rect 675904 231220 677600 231248
rect 675904 231208 675910 231220
rect 677594 231208 677600 231220
rect 677652 231208 677658 231260
rect 674840 231202 674892 231208
rect 674732 230988 674784 230994
rect 674732 230930 674784 230936
rect 673270 230800 673276 230852
rect 673328 230840 673334 230852
rect 673328 230812 674636 230840
rect 673328 230800 673334 230812
rect 158254 230704 158260 230716
rect 157306 230676 158260 230704
rect 144638 230528 144644 230580
rect 144696 230568 144702 230580
rect 150526 230568 150532 230580
rect 144696 230540 150532 230568
rect 144696 230528 144702 230540
rect 150526 230528 150532 230540
rect 150584 230528 150590 230580
rect 152182 230528 152188 230580
rect 152240 230568 152246 230580
rect 157306 230568 157334 230676
rect 158254 230664 158260 230676
rect 158312 230664 158318 230716
rect 668946 230664 668952 230716
rect 669004 230704 669010 230716
rect 673454 230704 673460 230716
rect 669004 230676 673460 230704
rect 669004 230664 669010 230676
rect 673454 230664 673460 230676
rect 673512 230664 673518 230716
rect 674390 230636 674396 230648
rect 674300 230608 674396 230636
rect 152240 230540 157334 230568
rect 157536 230540 158760 230568
rect 152240 230528 152246 230540
rect 90358 230392 90364 230444
rect 90416 230432 90422 230444
rect 157536 230432 157564 230540
rect 90416 230404 157564 230432
rect 158732 230432 158760 230540
rect 166074 230528 166080 230580
rect 166132 230568 166138 230580
rect 168190 230568 168196 230580
rect 166132 230540 168196 230568
rect 166132 230528 166138 230540
rect 168190 230528 168196 230540
rect 168248 230528 168254 230580
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 161106 230432 161112 230444
rect 158732 230404 161112 230432
rect 90416 230392 90422 230404
rect 161106 230392 161112 230404
rect 161164 230392 161170 230444
rect 161290 230392 161296 230444
rect 161348 230432 161354 230444
rect 215202 230432 215208 230444
rect 161348 230404 215208 230432
rect 161348 230392 161354 230404
rect 215202 230392 215208 230404
rect 215260 230392 215266 230444
rect 223390 230392 223396 230444
rect 223448 230432 223454 230444
rect 271874 230432 271880 230444
rect 223448 230404 271880 230432
rect 223448 230392 223454 230404
rect 271874 230392 271880 230404
rect 271932 230392 271938 230444
rect 274174 230392 274180 230444
rect 274232 230432 274238 230444
rect 307938 230432 307944 230444
rect 274232 230404 307944 230432
rect 274232 230392 274238 230404
rect 307938 230392 307944 230404
rect 307996 230392 308002 230444
rect 312538 230392 312544 230444
rect 312596 230432 312602 230444
rect 315666 230432 315672 230444
rect 312596 230404 315672 230432
rect 312596 230392 312602 230404
rect 315666 230392 315672 230404
rect 315724 230392 315730 230444
rect 377398 230392 377404 230444
rect 377456 230432 377462 230444
rect 378778 230432 378784 230444
rect 377456 230404 378784 230432
rect 377456 230392 377462 230404
rect 378778 230392 378784 230404
rect 378836 230392 378842 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443546 230432 443552 230444
rect 441948 230404 443552 230432
rect 441948 230392 441954 230404
rect 443546 230392 443552 230404
rect 443604 230392 443610 230444
rect 468294 230392 468300 230444
rect 468352 230432 468358 230444
rect 469030 230432 469036 230444
rect 468352 230404 469036 230432
rect 468352 230392 468358 230404
rect 469030 230392 469036 230404
rect 469088 230392 469094 230444
rect 526898 230392 526904 230444
rect 526956 230432 526962 230444
rect 537478 230432 537484 230444
rect 526956 230404 537484 230432
rect 526956 230392 526962 230404
rect 537478 230392 537484 230404
rect 537536 230392 537542 230444
rect 674300 230432 674328 230608
rect 674390 230596 674396 230608
rect 674448 230596 674454 230648
rect 674518 230580 674570 230586
rect 674518 230522 674570 230528
rect 674208 230404 674328 230432
rect 674396 230444 674448 230450
rect 404262 230324 404268 230376
rect 404320 230364 404326 230376
rect 412266 230364 412272 230376
rect 404320 230336 412272 230364
rect 404320 230324 404326 230336
rect 412266 230324 412272 230336
rect 412324 230324 412330 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444834 230364 444840 230376
rect 443880 230336 444840 230364
rect 443880 230324 443886 230336
rect 444834 230324 444840 230336
rect 444892 230324 444898 230376
rect 446398 230324 446404 230376
rect 446456 230364 446462 230376
rect 449158 230364 449164 230376
rect 446456 230336 449164 230364
rect 446456 230324 446462 230336
rect 449158 230324 449164 230336
rect 449216 230324 449222 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 476666 230324 476672 230376
rect 476724 230364 476730 230376
rect 479702 230364 479708 230376
rect 476724 230336 479708 230364
rect 476724 230324 476730 230336
rect 479702 230324 479708 230336
rect 479760 230324 479766 230376
rect 480530 230324 480536 230376
rect 480588 230364 480594 230376
rect 481542 230364 481548 230376
rect 480588 230336 481548 230364
rect 480588 230324 480594 230336
rect 481542 230324 481548 230336
rect 481600 230324 481606 230376
rect 483106 230324 483112 230376
rect 483164 230364 483170 230376
rect 484302 230364 484308 230376
rect 483164 230336 484308 230364
rect 483164 230324 483170 230336
rect 484302 230324 484308 230336
rect 484360 230324 484366 230376
rect 490190 230324 490196 230376
rect 490248 230364 490254 230376
rect 491202 230364 491208 230376
rect 490248 230336 491208 230364
rect 490248 230324 490254 230336
rect 491202 230324 491208 230336
rect 491260 230324 491266 230376
rect 492766 230324 492772 230376
rect 492824 230364 492830 230376
rect 493778 230364 493784 230376
rect 492824 230336 493784 230364
rect 492824 230324 492830 230336
rect 493778 230324 493784 230336
rect 493836 230324 493842 230376
rect 494698 230324 494704 230376
rect 494756 230364 494762 230376
rect 496354 230364 496360 230376
rect 494756 230336 496360 230364
rect 494756 230324 494762 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 499850 230324 499856 230376
rect 499908 230364 499914 230376
rect 501322 230364 501328 230376
rect 499908 230336 501328 230364
rect 499908 230324 499914 230336
rect 501322 230324 501328 230336
rect 501380 230324 501386 230376
rect 505002 230324 505008 230376
rect 505060 230364 505066 230376
rect 505738 230364 505744 230376
rect 505060 230336 505744 230364
rect 505060 230324 505066 230336
rect 505738 230324 505744 230336
rect 505796 230324 505802 230376
rect 516594 230324 516600 230376
rect 516652 230364 516658 230376
rect 517422 230364 517428 230376
rect 516652 230336 517428 230364
rect 516652 230324 516658 230336
rect 517422 230324 517428 230336
rect 517480 230324 517486 230376
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521562 230364 521568 230376
rect 520516 230336 521568 230364
rect 520516 230324 520522 230336
rect 521562 230324 521568 230336
rect 521620 230324 521626 230376
rect 669038 230324 669044 230376
rect 669096 230364 669102 230376
rect 673638 230364 673644 230376
rect 669096 230336 673644 230364
rect 669096 230324 669102 230336
rect 673638 230324 673644 230336
rect 673696 230324 673702 230376
rect 118418 230256 118424 230308
rect 118476 230296 118482 230308
rect 189442 230296 189448 230308
rect 118476 230268 189448 230296
rect 118476 230256 118482 230268
rect 189442 230256 189448 230268
rect 189500 230256 189506 230308
rect 190914 230256 190920 230308
rect 190972 230296 190978 230308
rect 190972 230268 195974 230296
rect 190972 230256 190978 230268
rect 111058 230120 111064 230172
rect 111116 230160 111122 230172
rect 184290 230160 184296 230172
rect 111116 230132 184296 230160
rect 111116 230120 111122 230132
rect 184290 230120 184296 230132
rect 184348 230120 184354 230172
rect 191282 230160 191288 230172
rect 186286 230132 191288 230160
rect 88242 229984 88248 230036
rect 88300 230024 88306 230036
rect 166258 230024 166264 230036
rect 88300 229996 166264 230024
rect 88300 229984 88306 229996
rect 166258 229984 166264 229996
rect 166316 229984 166322 230036
rect 166626 229984 166632 230036
rect 166684 230024 166690 230036
rect 181714 230024 181720 230036
rect 166684 229996 181720 230024
rect 166684 229984 166690 229996
rect 181714 229984 181720 229996
rect 181772 229984 181778 230036
rect 184198 229984 184204 230036
rect 184256 230024 184262 230036
rect 186286 230024 186314 230132
rect 191282 230120 191288 230132
rect 191340 230120 191346 230172
rect 195946 230160 195974 230268
rect 196986 230256 196992 230308
rect 197044 230296 197050 230308
rect 197044 230268 204944 230296
rect 197044 230256 197050 230268
rect 202322 230160 202328 230172
rect 195946 230132 202328 230160
rect 202322 230120 202328 230132
rect 202380 230120 202386 230172
rect 204916 230160 204944 230268
rect 205358 230256 205364 230308
rect 205416 230296 205422 230308
rect 256418 230296 256424 230308
rect 205416 230268 256424 230296
rect 205416 230256 205422 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 261386 230256 261392 230308
rect 261444 230296 261450 230308
rect 297634 230296 297640 230308
rect 261444 230268 297640 230296
rect 261444 230256 261450 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 302878 230256 302884 230308
rect 302936 230296 302942 230308
rect 305362 230296 305368 230308
rect 302936 230268 305368 230296
rect 302936 230256 302942 230268
rect 305362 230256 305368 230268
rect 305420 230256 305426 230308
rect 307846 230256 307852 230308
rect 307904 230296 307910 230308
rect 323394 230296 323400 230308
rect 307904 230268 323400 230296
rect 307904 230256 307910 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 497918 230256 497924 230308
rect 497976 230296 497982 230308
rect 497976 230268 499712 230296
rect 497976 230256 497982 230268
rect 408862 230188 408868 230240
rect 408920 230228 408926 230240
rect 410978 230228 410984 230240
rect 408920 230200 410984 230228
rect 408920 230188 408926 230200
rect 410978 230188 410984 230200
rect 411036 230188 411042 230240
rect 447042 230188 447048 230240
rect 447100 230228 447106 230240
rect 449894 230228 449900 230240
rect 447100 230200 449900 230228
rect 447100 230188 447106 230200
rect 449894 230188 449900 230200
rect 449952 230188 449958 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 454126 230188 454132 230240
rect 454184 230228 454190 230240
rect 455230 230228 455236 230240
rect 454184 230200 455236 230228
rect 454184 230188 454190 230200
rect 455230 230188 455236 230200
rect 455288 230188 455294 230240
rect 470870 230188 470876 230240
rect 470928 230228 470934 230240
rect 471882 230228 471888 230240
rect 470928 230200 471888 230228
rect 470928 230188 470934 230200
rect 471882 230188 471888 230200
rect 471940 230188 471946 230240
rect 475378 230188 475384 230240
rect 475436 230228 475442 230240
rect 479058 230228 479064 230240
rect 475436 230200 479064 230228
rect 475436 230188 475442 230200
rect 479058 230188 479064 230200
rect 479116 230188 479122 230240
rect 499684 230228 499712 230268
rect 532694 230256 532700 230308
rect 532752 230296 532758 230308
rect 547138 230296 547144 230308
rect 532752 230268 547144 230296
rect 532752 230256 532758 230268
rect 547138 230256 547144 230268
rect 547196 230256 547202 230308
rect 504358 230228 504364 230240
rect 499684 230200 504364 230228
rect 504358 230188 504364 230200
rect 504416 230188 504422 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 516778 230228 516784 230240
rect 511500 230200 516784 230228
rect 511500 230188 511506 230200
rect 516778 230188 516784 230200
rect 516836 230188 516842 230240
rect 521102 230188 521108 230240
rect 521160 230228 521166 230240
rect 530302 230228 530308 230240
rect 521160 230200 530308 230228
rect 521160 230188 521166 230200
rect 530302 230188 530308 230200
rect 530360 230188 530366 230240
rect 674208 230228 674236 230404
rect 674396 230386 674448 230392
rect 674208 230200 674314 230228
rect 251266 230160 251272 230172
rect 204916 230132 251272 230160
rect 251266 230120 251272 230132
rect 251324 230120 251330 230172
rect 276842 230120 276848 230172
rect 276900 230160 276906 230172
rect 313090 230160 313096 230172
rect 276900 230132 313096 230160
rect 276900 230120 276906 230132
rect 313090 230120 313096 230132
rect 313148 230120 313154 230172
rect 315298 230120 315304 230172
rect 315356 230160 315362 230172
rect 340138 230160 340144 230172
rect 315356 230132 340144 230160
rect 315356 230120 315362 230132
rect 340138 230120 340144 230132
rect 340196 230120 340202 230172
rect 488258 230120 488264 230172
rect 488316 230160 488322 230172
rect 488316 230132 499574 230160
rect 488316 230120 488322 230132
rect 499546 230104 499574 230132
rect 533522 230120 533528 230172
rect 533580 230160 533586 230172
rect 543918 230160 543924 230172
rect 533580 230132 543924 230160
rect 533580 230120 533586 230132
rect 543918 230120 543924 230132
rect 543976 230120 543982 230172
rect 555418 230120 555424 230172
rect 555476 230160 555482 230172
rect 571334 230160 571340 230172
rect 555476 230132 571340 230160
rect 555476 230120 555482 230132
rect 571334 230120 571340 230132
rect 571392 230120 571398 230172
rect 345658 230052 345664 230104
rect 345716 230092 345722 230104
rect 353018 230092 353024 230104
rect 345716 230064 353024 230092
rect 345716 230052 345722 230064
rect 353018 230052 353024 230064
rect 353076 230052 353082 230104
rect 444466 230052 444472 230104
rect 444524 230092 444530 230104
rect 447594 230092 447600 230104
rect 444524 230064 447600 230092
rect 444524 230052 444530 230064
rect 447594 230052 447600 230064
rect 447652 230052 447658 230104
rect 499546 230064 499580 230104
rect 499574 230052 499580 230064
rect 499632 230052 499638 230104
rect 673592 230052 673598 230104
rect 673650 230092 673656 230104
rect 673650 230064 674198 230092
rect 673650 230052 673656 230064
rect 184256 229996 186314 230024
rect 184256 229984 184262 229996
rect 190270 229984 190276 230036
rect 190328 230024 190334 230036
rect 246114 230024 246120 230036
rect 190328 229996 246120 230024
rect 190328 229984 190334 229996
rect 246114 229984 246120 229996
rect 246172 229984 246178 230036
rect 251726 229984 251732 230036
rect 251784 230024 251790 230036
rect 292482 230024 292488 230036
rect 251784 229996 292488 230024
rect 251784 229984 251790 229996
rect 292482 229984 292488 229996
rect 292540 229984 292546 230036
rect 296990 229984 296996 230036
rect 297048 230024 297054 230036
rect 302510 230024 302516 230036
rect 297048 229996 302516 230024
rect 297048 229984 297054 229996
rect 302510 229984 302516 229996
rect 302568 229984 302574 230036
rect 305638 229984 305644 230036
rect 305696 230024 305702 230036
rect 334986 230024 334992 230036
rect 305696 229996 334992 230024
rect 305696 229984 305702 229996
rect 334986 229984 334992 229996
rect 335044 229984 335050 230036
rect 380434 229984 380440 230036
rect 380492 230024 380498 230036
rect 389082 230024 389088 230036
rect 380492 229996 389088 230024
rect 380492 229984 380498 229996
rect 389082 229984 389088 229996
rect 389140 229984 389146 230036
rect 410886 229984 410892 230036
rect 410944 230024 410950 230036
rect 417418 230024 417424 230036
rect 410944 229996 417424 230024
rect 410944 229984 410950 229996
rect 417418 229984 417424 229996
rect 417476 229984 417482 230036
rect 467006 229984 467012 230036
rect 467064 230024 467070 230036
rect 473998 230024 474004 230036
rect 467064 229996 474004 230024
rect 467064 229984 467070 229996
rect 473998 229984 474004 229996
rect 474056 229984 474062 230036
rect 484762 229984 484768 230036
rect 484820 230024 484826 230036
rect 484820 229996 490696 230024
rect 484820 229984 484826 229996
rect 74442 229848 74448 229900
rect 74500 229888 74506 229900
rect 155954 229888 155960 229900
rect 74500 229860 155960 229888
rect 74500 229848 74506 229860
rect 155954 229848 155960 229860
rect 156012 229848 156018 229900
rect 156598 229848 156604 229900
rect 156656 229888 156662 229900
rect 176562 229888 176568 229900
rect 156656 229860 176568 229888
rect 156656 229848 156662 229860
rect 176562 229848 176568 229860
rect 176620 229848 176626 229900
rect 177574 229848 177580 229900
rect 177632 229888 177638 229900
rect 177632 229860 191144 229888
rect 177632 229848 177638 229860
rect 67542 229712 67548 229764
rect 67600 229752 67606 229764
rect 144638 229752 144644 229764
rect 67600 229724 144644 229752
rect 67600 229712 67606 229724
rect 144638 229712 144644 229724
rect 144696 229712 144702 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 144880 229724 147168 229752
rect 144880 229712 144886 229724
rect 140038 229576 140044 229628
rect 140096 229616 140102 229628
rect 146938 229616 146944 229628
rect 140096 229588 146944 229616
rect 140096 229576 140102 229588
rect 146938 229576 146944 229588
rect 146996 229576 147002 229628
rect 147140 229616 147168 229724
rect 148778 229712 148784 229764
rect 148836 229752 148842 229764
rect 151906 229752 151912 229764
rect 148836 229724 151912 229752
rect 148836 229712 148842 229724
rect 151906 229712 151912 229724
rect 151964 229712 151970 229764
rect 152366 229712 152372 229764
rect 152424 229752 152430 229764
rect 190914 229752 190920 229764
rect 152424 229724 190920 229752
rect 152424 229712 152430 229724
rect 190914 229712 190920 229724
rect 190972 229712 190978 229764
rect 191116 229752 191144 229860
rect 191282 229848 191288 229900
rect 191340 229888 191346 229900
rect 240962 229888 240968 229900
rect 191340 229860 240968 229888
rect 191340 229848 191346 229860
rect 240962 229848 240968 229860
rect 241020 229848 241026 229900
rect 245654 229848 245660 229900
rect 245712 229888 245718 229900
rect 287330 229888 287336 229900
rect 245712 229860 287336 229888
rect 245712 229848 245718 229860
rect 287330 229848 287336 229860
rect 287388 229848 287394 229900
rect 300118 229848 300124 229900
rect 300176 229888 300182 229900
rect 329834 229888 329840 229900
rect 300176 229860 329840 229888
rect 300176 229848 300182 229860
rect 329834 229848 329840 229860
rect 329892 229848 329898 229900
rect 334250 229848 334256 229900
rect 334308 229888 334314 229900
rect 345290 229888 345296 229900
rect 334308 229860 345296 229888
rect 334308 229848 334314 229860
rect 345290 229848 345296 229860
rect 345348 229848 345354 229900
rect 352558 229848 352564 229900
rect 352616 229888 352622 229900
rect 358170 229888 358176 229900
rect 352616 229860 358176 229888
rect 352616 229848 352622 229860
rect 358170 229848 358176 229860
rect 358228 229848 358234 229900
rect 364150 229848 364156 229900
rect 364208 229888 364214 229900
rect 381354 229888 381360 229900
rect 364208 229860 381360 229888
rect 364208 229848 364214 229860
rect 381354 229848 381360 229860
rect 381412 229848 381418 229900
rect 384298 229848 384304 229900
rect 384356 229888 384362 229900
rect 394234 229888 394240 229900
rect 384356 229860 394240 229888
rect 384356 229848 384362 229860
rect 394234 229848 394240 229860
rect 394292 229848 394298 229900
rect 469582 229848 469588 229900
rect 469640 229888 469646 229900
rect 476850 229888 476856 229900
rect 469640 229860 476856 229888
rect 469640 229848 469646 229860
rect 476850 229848 476856 229860
rect 476908 229848 476914 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 489914 229888 489920 229900
rect 481876 229860 489920 229888
rect 481876 229848 481882 229860
rect 489914 229848 489920 229860
rect 489972 229848 489978 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 235810 229752 235816 229764
rect 191116 229724 235816 229752
rect 235810 229712 235816 229724
rect 235868 229712 235874 229764
rect 236914 229712 236920 229764
rect 236972 229752 236978 229764
rect 282178 229752 282184 229764
rect 236972 229724 282184 229752
rect 236972 229712 236978 229724
rect 282178 229712 282184 229724
rect 282236 229712 282242 229764
rect 285306 229712 285312 229764
rect 285364 229752 285370 229764
rect 318242 229752 318248 229764
rect 285364 229724 318248 229752
rect 285364 229712 285370 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 324038 229712 324044 229764
rect 324096 229752 324102 229764
rect 350442 229752 350448 229764
rect 324096 229724 350448 229752
rect 324096 229712 324102 229724
rect 350442 229712 350448 229724
rect 350500 229712 350506 229764
rect 371050 229752 371056 229764
rect 354646 229724 371056 229752
rect 210050 229616 210056 229628
rect 147140 229588 210056 229616
rect 210050 229576 210056 229588
rect 210108 229576 210114 229628
rect 210234 229576 210240 229628
rect 210292 229616 210298 229628
rect 261570 229616 261576 229628
rect 210292 229588 261576 229616
rect 210292 229576 210298 229588
rect 261570 229576 261576 229588
rect 261628 229576 261634 229628
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 354646 229616 354674 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 386506 229752 386512 229764
rect 373966 229724 386512 229752
rect 350592 229588 354674 229616
rect 350592 229576 350598 229588
rect 370958 229576 370964 229628
rect 371016 229616 371022 229628
rect 373966 229616 373994 229724
rect 386506 229712 386512 229724
rect 386564 229712 386570 229764
rect 386966 229712 386972 229764
rect 387024 229752 387030 229764
rect 396810 229752 396816 229764
rect 387024 229724 396816 229752
rect 387024 229712 387030 229724
rect 396810 229712 396816 229724
rect 396868 229712 396874 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 412450 229712 412456 229764
rect 412508 229752 412514 229764
rect 419350 229752 419356 229764
rect 412508 229724 419356 229752
rect 412508 229712 412514 229724
rect 419350 229712 419356 229724
rect 419408 229712 419414 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 468846 229712 468852 229764
rect 468904 229752 468910 229764
rect 475378 229752 475384 229764
rect 468904 229724 475384 229752
rect 468904 229712 468910 229724
rect 475378 229712 475384 229724
rect 475436 229712 475442 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 487154 229752 487160 229764
rect 479300 229724 487160 229752
rect 479300 229712 479306 229724
rect 487154 229712 487160 229724
rect 487212 229712 487218 229764
rect 371016 229588 373994 229616
rect 371016 229576 371022 229588
rect 477954 229576 477960 229628
rect 478012 229616 478018 229628
rect 478506 229616 478512 229628
rect 478012 229588 478512 229616
rect 478012 229576 478018 229588
rect 478506 229576 478512 229588
rect 478564 229576 478570 229628
rect 490668 229616 490696 229996
rect 490834 229984 490840 230036
rect 490892 230024 490898 230036
rect 493962 230024 493968 230036
rect 490892 229996 493968 230024
rect 490892 229984 490898 229996
rect 493962 229984 493968 229996
rect 494020 229984 494026 230036
rect 505922 229984 505928 230036
rect 505980 230024 505986 230036
rect 515766 230024 515772 230036
rect 505980 229996 515772 230024
rect 505980 229984 505986 229996
rect 515766 229984 515772 229996
rect 515824 229984 515830 230036
rect 517238 229984 517244 230036
rect 517296 230024 517302 230036
rect 522298 230024 522304 230036
rect 517296 229996 522304 230024
rect 517296 229984 517302 229996
rect 522298 229984 522304 229996
rect 522356 229984 522362 230036
rect 523034 229984 523040 230036
rect 523092 230024 523098 230036
rect 534810 230024 534816 230036
rect 523092 229996 534816 230024
rect 523092 229984 523098 229996
rect 534810 229984 534816 229996
rect 534868 229984 534874 230036
rect 538490 229984 538496 230036
rect 538548 230024 538554 230036
rect 559558 230024 559564 230036
rect 538548 229996 559564 230024
rect 538548 229984 538554 229996
rect 559558 229984 559564 229996
rect 559616 229984 559622 230036
rect 673730 229916 673736 229968
rect 673788 229916 673794 229968
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 510614 229888 510620 229900
rect 496044 229860 510620 229888
rect 496044 229848 496050 229860
rect 510614 229848 510620 229860
rect 510672 229848 510678 229900
rect 513374 229848 513380 229900
rect 513432 229888 513438 229900
rect 525058 229888 525064 229900
rect 513432 229860 525064 229888
rect 513432 229848 513438 229860
rect 525058 229848 525064 229860
rect 525116 229848 525122 229900
rect 528830 229848 528836 229900
rect 528888 229888 528894 229900
rect 533522 229888 533528 229900
rect 528888 229860 533528 229888
rect 528888 229848 528894 229860
rect 533522 229848 533528 229860
rect 533580 229848 533586 229900
rect 534626 229848 534632 229900
rect 534684 229888 534690 229900
rect 555234 229888 555240 229900
rect 534684 229860 555240 229888
rect 534684 229848 534690 229860
rect 555234 229848 555240 229860
rect 555292 229848 555298 229900
rect 673748 229820 673776 229916
rect 675846 229848 675852 229900
rect 675904 229888 675910 229900
rect 677226 229888 677232 229900
rect 675904 229860 677232 229888
rect 675904 229848 675910 229860
rect 677226 229848 677232 229860
rect 677284 229848 677290 229900
rect 673748 229792 674084 229820
rect 494330 229712 494336 229764
rect 494388 229752 494394 229764
rect 509878 229752 509884 229764
rect 494388 229724 509884 229752
rect 494388 229712 494394 229724
rect 509878 229712 509884 229724
rect 509936 229712 509942 229764
rect 525242 229712 525248 229764
rect 525300 229752 525306 229764
rect 528922 229752 528928 229764
rect 525300 229724 528928 229752
rect 525300 229712 525306 229724
rect 528922 229712 528928 229724
rect 528980 229712 528986 229764
rect 536558 229712 536564 229764
rect 536616 229752 536622 229764
rect 562318 229752 562324 229764
rect 536616 229724 562324 229752
rect 536616 229712 536622 229724
rect 562318 229712 562324 229724
rect 562376 229712 562382 229764
rect 669406 229712 669412 229764
rect 669464 229752 669470 229764
rect 670510 229752 670516 229764
rect 669464 229724 670516 229752
rect 669464 229712 669470 229724
rect 670510 229712 670516 229724
rect 670568 229712 670574 229764
rect 670712 229656 673974 229684
rect 497458 229616 497464 229628
rect 490668 229588 497464 229616
rect 497458 229576 497464 229588
rect 497516 229576 497522 229628
rect 503714 229576 503720 229628
rect 503772 229616 503778 229628
rect 508498 229616 508504 229628
rect 503772 229588 508504 229616
rect 503772 229576 503778 229588
rect 508498 229576 508504 229588
rect 508556 229576 508562 229628
rect 515306 229576 515312 229628
rect 515364 229616 515370 229628
rect 526070 229616 526076 229628
rect 515364 229588 526076 229616
rect 515364 229576 515370 229588
rect 526070 229576 526076 229588
rect 526128 229576 526134 229628
rect 530762 229576 530768 229628
rect 530820 229616 530826 229628
rect 540238 229616 540244 229628
rect 530820 229588 540244 229616
rect 530820 229576 530826 229588
rect 540238 229576 540244 229588
rect 540296 229576 540302 229628
rect 666830 229576 666836 229628
rect 666888 229616 666894 229628
rect 670712 229616 670740 229656
rect 666888 229588 670740 229616
rect 666888 229576 666894 229588
rect 131114 229440 131120 229492
rect 131172 229480 131178 229492
rect 197170 229480 197176 229492
rect 131172 229452 197176 229480
rect 131172 229440 131178 229452
rect 197170 229440 197176 229452
rect 197228 229440 197234 229492
rect 203886 229440 203892 229492
rect 203944 229480 203950 229492
rect 205358 229480 205364 229492
rect 203944 229452 205364 229480
rect 203944 229440 203950 229452
rect 205358 229440 205364 229452
rect 205416 229440 205422 229492
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 277026 229480 277032 229492
rect 231176 229452 277032 229480
rect 231176 229440 231182 229452
rect 277026 229440 277032 229452
rect 277084 229440 277090 229492
rect 509510 229440 509516 229492
rect 509568 229480 509574 229492
rect 518158 229480 518164 229492
rect 509568 229452 518164 229480
rect 509568 229440 509574 229452
rect 518158 229440 518164 229452
rect 518216 229440 518222 229492
rect 519170 229440 519176 229492
rect 519228 229480 519234 229492
rect 527818 229480 527824 229492
rect 519228 229452 527824 229480
rect 519228 229440 519234 229452
rect 527818 229440 527824 229452
rect 527876 229440 527882 229492
rect 673408 229440 673414 229492
rect 673466 229480 673472 229492
rect 673466 229452 673854 229480
rect 673466 229440 673472 229452
rect 436094 229372 436100 229424
rect 436152 229412 436158 229424
rect 436738 229412 436744 229424
rect 436152 229384 436744 229412
rect 436152 229372 436158 229384
rect 436738 229372 436744 229384
rect 436796 229372 436802 229424
rect 448974 229372 448980 229424
rect 449032 229412 449038 229424
rect 451366 229412 451372 229424
rect 449032 229384 451372 229412
rect 449032 229372 449038 229384
rect 451366 229372 451372 229384
rect 451424 229372 451430 229424
rect 122926 229304 122932 229356
rect 122984 229344 122990 229356
rect 179138 229344 179144 229356
rect 122984 229316 179144 229344
rect 122984 229304 122990 229316
rect 179138 229304 179144 229316
rect 179196 229304 179202 229356
rect 182082 229304 182088 229356
rect 182140 229344 182146 229356
rect 230658 229344 230664 229356
rect 182140 229316 230664 229344
rect 182140 229304 182146 229316
rect 230658 229304 230664 229316
rect 230716 229304 230722 229356
rect 453482 229304 453488 229356
rect 453540 229344 453546 229356
rect 455782 229344 455788 229356
rect 453540 229316 455788 229344
rect 453540 229304 453546 229316
rect 455782 229304 455788 229316
rect 455840 229304 455846 229356
rect 673736 229288 673788 229294
rect 358078 229236 358084 229288
rect 358136 229276 358142 229288
rect 360746 229276 360752 229288
rect 358136 229248 360752 229276
rect 358136 229236 358142 229248
rect 360746 229236 360752 229248
rect 360804 229236 360810 229288
rect 360930 229236 360936 229288
rect 360988 229276 360994 229288
rect 363322 229276 363328 229288
rect 360988 229248 363328 229276
rect 360988 229236 360994 229248
rect 363322 229236 363328 229248
rect 363380 229236 363386 229288
rect 419442 229236 419448 229288
rect 419500 229276 419506 229288
rect 424502 229276 424508 229288
rect 419500 229248 424508 229276
rect 419500 229236 419506 229248
rect 424502 229236 424508 229248
rect 424560 229236 424566 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451826 229276 451832 229288
rect 450320 229248 451832 229276
rect 450320 229236 450326 229248
rect 451826 229236 451832 229248
rect 451884 229236 451890 229288
rect 479886 229236 479892 229288
rect 479944 229276 479950 229288
rect 482278 229276 482284 229288
rect 479944 229248 482284 229276
rect 479944 229236 479950 229248
rect 482278 229236 482284 229248
rect 482336 229236 482342 229288
rect 501782 229236 501788 229288
rect 501840 229276 501846 229288
rect 507118 229276 507124 229288
rect 501840 229248 507124 229276
rect 501840 229236 501846 229248
rect 507118 229236 507124 229248
rect 507176 229236 507182 229288
rect 673736 229230 673788 229236
rect 92474 229168 92480 229220
rect 92532 229208 92538 229220
rect 146294 229208 146300 229220
rect 92532 229180 146300 229208
rect 92532 229168 92538 229180
rect 146294 229168 146300 229180
rect 146352 229168 146358 229220
rect 146938 229168 146944 229220
rect 146996 229208 147002 229220
rect 153378 229208 153384 229220
rect 146996 229180 153384 229208
rect 146996 229168 147002 229180
rect 153378 229168 153384 229180
rect 153436 229168 153442 229220
rect 153838 229168 153844 229220
rect 153896 229208 153902 229220
rect 163682 229208 163688 229220
rect 153896 229180 163688 229208
rect 153896 229168 153902 229180
rect 163682 229168 163688 229180
rect 163740 229168 163746 229220
rect 163866 229168 163872 229220
rect 163924 229208 163930 229220
rect 166626 229208 166632 229220
rect 163924 229180 166632 229208
rect 163924 229168 163930 229180
rect 166626 229168 166632 229180
rect 166684 229168 166690 229220
rect 167638 229168 167644 229220
rect 167696 229208 167702 229220
rect 220354 229208 220360 229220
rect 167696 229180 220360 229208
rect 167696 229168 167702 229180
rect 220354 229168 220360 229180
rect 220412 229168 220418 229220
rect 476022 229168 476028 229220
rect 476080 229208 476086 229220
rect 478690 229208 478696 229220
rect 476080 229180 478696 229208
rect 476080 229168 476086 229180
rect 478690 229168 478696 229180
rect 478748 229168 478754 229220
rect 378962 229100 378968 229152
rect 379020 229140 379026 229152
rect 383930 229140 383936 229152
rect 379020 229112 383936 229140
rect 379020 229100 379026 229112
rect 383930 229100 383936 229112
rect 383988 229100 383994 229152
rect 419994 229140 420000 229152
rect 418126 229112 420000 229140
rect 102042 229032 102048 229084
rect 102100 229072 102106 229084
rect 175274 229072 175280 229084
rect 102100 229044 175280 229072
rect 102100 229032 102106 229044
rect 175274 229032 175280 229044
rect 175332 229032 175338 229084
rect 175642 229032 175648 229084
rect 175700 229072 175706 229084
rect 175700 229044 181576 229072
rect 175700 229032 175706 229044
rect 97902 228896 97908 228948
rect 97960 228936 97966 228948
rect 97960 228908 108344 228936
rect 97960 228896 97966 228908
rect 108114 228800 108120 228812
rect 84166 228772 108120 228800
rect 82078 228624 82084 228676
rect 82136 228664 82142 228676
rect 84166 228664 84194 228772
rect 108114 228760 108120 228772
rect 108172 228760 108178 228812
rect 108316 228800 108344 228908
rect 108482 228896 108488 228948
rect 108540 228936 108546 228948
rect 170950 228936 170956 228948
rect 108540 228908 170956 228936
rect 108540 228896 108546 228908
rect 170950 228896 170956 228908
rect 171008 228896 171014 228948
rect 173894 228936 173900 228948
rect 171336 228908 173900 228936
rect 171336 228800 171364 228908
rect 173894 228896 173900 228908
rect 173952 228896 173958 228948
rect 174078 228896 174084 228948
rect 174136 228936 174142 228948
rect 174136 228908 181484 228936
rect 174136 228896 174142 228908
rect 108316 228772 171364 228800
rect 171594 228760 171600 228812
rect 171652 228800 171658 228812
rect 181254 228800 181260 228812
rect 171652 228772 181260 228800
rect 171652 228760 171658 228772
rect 181254 228760 181260 228772
rect 181312 228760 181318 228812
rect 82136 228636 84194 228664
rect 82136 228624 82142 228636
rect 96522 228624 96528 228676
rect 96580 228664 96586 228676
rect 172054 228664 172060 228676
rect 96580 228636 172060 228664
rect 96580 228624 96586 228636
rect 172054 228624 172060 228636
rect 172112 228624 172118 228676
rect 172238 228624 172244 228676
rect 172296 228664 172302 228676
rect 179782 228664 179788 228676
rect 172296 228636 179788 228664
rect 172296 228624 172302 228636
rect 179782 228624 179788 228636
rect 179840 228624 179846 228676
rect 181456 228664 181484 228908
rect 181548 228800 181576 229044
rect 181714 229032 181720 229084
rect 181772 229072 181778 229084
rect 190546 229072 190552 229084
rect 181772 229044 190552 229072
rect 181772 229032 181778 229044
rect 190546 229032 190552 229044
rect 190604 229032 190610 229084
rect 191374 229032 191380 229084
rect 191432 229072 191438 229084
rect 194594 229072 194600 229084
rect 191432 229044 194600 229072
rect 191432 229032 191438 229044
rect 194594 229032 194600 229044
rect 194652 229032 194658 229084
rect 195698 229032 195704 229084
rect 195756 229072 195762 229084
rect 250622 229072 250628 229084
rect 195756 229044 250628 229072
rect 195756 229032 195762 229044
rect 250622 229032 250628 229044
rect 250680 229032 250686 229084
rect 259270 229032 259276 229084
rect 259328 229072 259334 229084
rect 298278 229072 298284 229084
rect 259328 229044 298284 229072
rect 259328 229032 259334 229044
rect 298278 229032 298284 229044
rect 298336 229032 298342 229084
rect 413738 229032 413744 229084
rect 413796 229072 413802 229084
rect 418126 229072 418154 229112
rect 419994 229100 420000 229112
rect 420052 229100 420058 229152
rect 420178 229100 420184 229152
rect 420236 229140 420242 229152
rect 421926 229140 421932 229152
rect 420236 229112 421932 229140
rect 420236 229100 420242 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 424318 229100 424324 229152
rect 424376 229140 424382 229152
rect 427722 229140 427728 229152
rect 424376 229112 427728 229140
rect 424376 229100 424382 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 413796 229044 418154 229072
rect 413796 229032 413802 229044
rect 519814 229032 519820 229084
rect 519872 229072 519878 229084
rect 543182 229072 543188 229084
rect 519872 229044 543188 229072
rect 519872 229032 519878 229044
rect 543182 229032 543188 229044
rect 543240 229032 543246 229084
rect 673382 229032 673388 229084
rect 673440 229072 673446 229084
rect 673440 229044 673624 229072
rect 673440 229032 673446 229044
rect 675846 229032 675852 229084
rect 675904 229072 675910 229084
rect 676214 229072 676220 229084
rect 675904 229044 676220 229072
rect 675904 229032 675910 229044
rect 676214 229032 676220 229044
rect 676272 229032 676278 229084
rect 181898 228896 181904 228948
rect 181956 228936 181962 228948
rect 181956 228908 191144 228936
rect 181956 228896 181962 228908
rect 190914 228800 190920 228812
rect 181548 228772 190920 228800
rect 190914 228760 190920 228772
rect 190972 228760 190978 228812
rect 191116 228800 191144 228908
rect 192202 228896 192208 228948
rect 192260 228936 192266 228948
rect 241606 228936 241612 228948
rect 192260 228908 241612 228936
rect 192260 228896 192266 228908
rect 241606 228896 241612 228908
rect 241664 228896 241670 228948
rect 251082 228896 251088 228948
rect 251140 228936 251146 228948
rect 291194 228936 291200 228948
rect 251140 228908 291200 228936
rect 251140 228896 251146 228908
rect 291194 228896 291200 228908
rect 291252 228896 291258 228948
rect 319806 228896 319812 228948
rect 319864 228936 319870 228948
rect 345934 228936 345940 228948
rect 319864 228908 345940 228936
rect 319864 228896 319870 228908
rect 345934 228896 345940 228908
rect 345992 228896 345998 228948
rect 349982 228896 349988 228948
rect 350040 228936 350046 228948
rect 369118 228936 369124 228948
rect 350040 228908 369124 228936
rect 350040 228896 350046 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 517882 228896 517888 228948
rect 517940 228936 517946 228948
rect 540054 228936 540060 228948
rect 517940 228908 540060 228936
rect 517940 228896 517946 228908
rect 540054 228896 540060 228908
rect 540112 228896 540118 228948
rect 212626 228800 212632 228812
rect 191116 228772 212632 228800
rect 212626 228760 212632 228772
rect 212684 228760 212690 228812
rect 219158 228760 219164 228812
rect 219216 228800 219222 228812
rect 224034 228800 224040 228812
rect 219216 228772 224040 228800
rect 219216 228760 219222 228772
rect 224034 228760 224040 228772
rect 224092 228760 224098 228812
rect 231302 228800 231308 228812
rect 224236 228772 231308 228800
rect 224236 228664 224264 228772
rect 231302 228760 231308 228772
rect 231360 228760 231366 228812
rect 246206 228760 246212 228812
rect 246264 228800 246270 228812
rect 253842 228800 253848 228812
rect 246264 228772 253848 228800
rect 246264 228760 246270 228772
rect 253842 228760 253848 228772
rect 253900 228760 253906 228812
rect 255038 228760 255044 228812
rect 255096 228800 255102 228812
rect 295702 228800 295708 228812
rect 255096 228772 295708 228800
rect 255096 228760 255102 228772
rect 295702 228760 295708 228772
rect 295760 228760 295766 228812
rect 318058 228760 318064 228812
rect 318116 228800 318122 228812
rect 344646 228800 344652 228812
rect 318116 228772 344652 228800
rect 318116 228760 318122 228772
rect 344646 228760 344652 228772
rect 344704 228760 344710 228812
rect 346118 228760 346124 228812
rect 346176 228800 346182 228812
rect 366174 228800 366180 228812
rect 346176 228772 366180 228800
rect 346176 228760 346182 228772
rect 366174 228760 366180 228772
rect 366232 228760 366238 228812
rect 373810 228760 373816 228812
rect 373868 228800 373874 228812
rect 387242 228800 387248 228812
rect 373868 228772 387248 228800
rect 373868 228760 373874 228772
rect 387242 228760 387248 228772
rect 387300 228760 387306 228812
rect 401318 228760 401324 228812
rect 401376 228800 401382 228812
rect 408402 228800 408408 228812
rect 401376 228772 408408 228800
rect 401376 228760 401382 228772
rect 408402 228760 408408 228772
rect 408460 228760 408466 228812
rect 487154 228760 487160 228812
rect 487212 228800 487218 228812
rect 489914 228800 489920 228812
rect 487212 228772 489920 228800
rect 487212 228760 487218 228772
rect 489914 228760 489920 228772
rect 489972 228760 489978 228812
rect 493962 228760 493968 228812
rect 494020 228800 494026 228812
rect 505922 228800 505928 228812
rect 494020 228772 505928 228800
rect 494020 228760 494026 228772
rect 505922 228760 505928 228772
rect 505980 228760 505986 228812
rect 507118 228760 507124 228812
rect 507176 228800 507182 228812
rect 519722 228800 519728 228812
rect 507176 228772 519728 228800
rect 507176 228760 507182 228772
rect 519722 228760 519728 228772
rect 519780 228760 519786 228812
rect 526254 228760 526260 228812
rect 526312 228800 526318 228812
rect 551186 228800 551192 228812
rect 526312 228772 551192 228800
rect 526312 228760 526318 228772
rect 551186 228760 551192 228772
rect 551244 228760 551250 228812
rect 673506 228744 673558 228750
rect 673506 228686 673558 228692
rect 237190 228664 237196 228676
rect 181456 228636 224264 228664
rect 224328 228636 237196 228664
rect 62758 228488 62764 228540
rect 62816 228528 62822 228540
rect 140774 228528 140780 228540
rect 62816 228500 140780 228528
rect 62816 228488 62822 228500
rect 140774 228488 140780 228500
rect 140832 228488 140838 228540
rect 140958 228488 140964 228540
rect 141016 228528 141022 228540
rect 156414 228528 156420 228540
rect 141016 228500 156420 228528
rect 141016 228488 141022 228500
rect 156414 228488 156420 228500
rect 156472 228488 156478 228540
rect 204714 228528 204720 228540
rect 156800 228500 204720 228528
rect 65978 228352 65984 228404
rect 66036 228392 66042 228404
rect 150158 228392 150164 228404
rect 66036 228364 150164 228392
rect 66036 228352 66042 228364
rect 150158 228352 150164 228364
rect 150216 228352 150222 228404
rect 150342 228352 150348 228404
rect 150400 228392 150406 228404
rect 156800 228392 156828 228500
rect 204714 228488 204720 228500
rect 204772 228488 204778 228540
rect 204898 228488 204904 228540
rect 204956 228528 204962 228540
rect 204956 228500 212396 228528
rect 204956 228488 204962 228500
rect 150400 228364 156828 228392
rect 150400 228352 150406 228364
rect 156966 228352 156972 228404
rect 157024 228392 157030 228404
rect 157426 228392 157432 228404
rect 157024 228364 157432 228392
rect 157024 228352 157030 228364
rect 157426 228352 157432 228364
rect 157484 228352 157490 228404
rect 157794 228352 157800 228404
rect 157852 228392 157858 228404
rect 212166 228392 212172 228404
rect 157852 228364 212172 228392
rect 157852 228352 157858 228364
rect 212166 228352 212172 228364
rect 212224 228352 212230 228404
rect 212368 228392 212396 228500
rect 212626 228488 212632 228540
rect 212684 228528 212690 228540
rect 224328 228528 224356 228636
rect 237190 228624 237196 228636
rect 237248 228624 237254 228676
rect 239398 228624 239404 228676
rect 239456 228664 239462 228676
rect 284110 228664 284116 228676
rect 239456 228636 284116 228664
rect 239456 228624 239462 228636
rect 284110 228624 284116 228636
rect 284168 228624 284174 228676
rect 292390 228624 292396 228676
rect 292448 228664 292454 228676
rect 326614 228664 326620 228676
rect 292448 228636 326620 228664
rect 292448 228624 292454 228636
rect 326614 228624 326620 228636
rect 326672 228624 326678 228676
rect 333238 228624 333244 228676
rect 333296 228664 333302 228676
rect 355594 228664 355600 228676
rect 333296 228636 355600 228664
rect 333296 228624 333302 228636
rect 355594 228624 355600 228636
rect 355652 228624 355658 228676
rect 369762 228664 369768 228676
rect 359016 228636 369768 228664
rect 267366 228528 267372 228540
rect 212684 228500 224356 228528
rect 224420 228500 267372 228528
rect 212684 228488 212690 228500
rect 222746 228392 222752 228404
rect 212368 228364 222752 228392
rect 222746 228352 222752 228364
rect 222804 228352 222810 228404
rect 224034 228352 224040 228404
rect 224092 228392 224098 228404
rect 224420 228392 224448 228500
rect 267366 228488 267372 228500
rect 267424 228488 267430 228540
rect 267550 228488 267556 228540
rect 267608 228528 267614 228540
rect 307294 228528 307300 228540
rect 267608 228500 307300 228528
rect 267608 228488 267614 228500
rect 307294 228488 307300 228500
rect 307352 228488 307358 228540
rect 307662 228488 307668 228540
rect 307720 228528 307726 228540
rect 335630 228528 335636 228540
rect 307720 228500 335636 228528
rect 307720 228488 307726 228500
rect 335630 228488 335636 228500
rect 335688 228488 335694 228540
rect 336642 228488 336648 228540
rect 336700 228528 336706 228540
rect 358814 228528 358820 228540
rect 336700 228500 358820 228528
rect 336700 228488 336706 228500
rect 358814 228488 358820 228500
rect 358872 228488 358878 228540
rect 224092 228364 224448 228392
rect 224092 228352 224098 228364
rect 225690 228352 225696 228404
rect 225748 228392 225754 228404
rect 273806 228392 273812 228404
rect 225748 228364 273812 228392
rect 225748 228352 225754 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 283926 228352 283932 228404
rect 283984 228392 283990 228404
rect 320174 228392 320180 228404
rect 283984 228364 320180 228392
rect 283984 228352 283990 228364
rect 320174 228352 320180 228364
rect 320232 228352 320238 228404
rect 326798 228352 326804 228404
rect 326856 228392 326862 228404
rect 351086 228392 351092 228404
rect 326856 228364 351092 228392
rect 326856 228352 326862 228364
rect 351086 228352 351092 228364
rect 351144 228352 351150 228404
rect 355318 228352 355324 228404
rect 355376 228392 355382 228404
rect 359016 228392 359044 228636
rect 369762 228624 369768 228636
rect 369820 228624 369826 228676
rect 376478 228624 376484 228676
rect 376536 228664 376542 228676
rect 389726 228664 389732 228676
rect 376536 228636 389732 228664
rect 376536 228624 376542 228636
rect 389726 228624 389732 228636
rect 389784 228624 389790 228676
rect 390278 228624 390284 228676
rect 390336 228664 390342 228676
rect 400030 228664 400036 228676
rect 390336 228636 400036 228664
rect 390336 228624 390342 228636
rect 400030 228624 400036 228636
rect 400088 228624 400094 228676
rect 411070 228624 411076 228676
rect 411128 228664 411134 228676
rect 416130 228664 416136 228676
rect 411128 228636 416136 228664
rect 411128 228624 411134 228636
rect 416130 228624 416136 228636
rect 416188 228624 416194 228676
rect 479702 228624 479708 228676
rect 479760 228664 479766 228676
rect 487430 228664 487436 228676
rect 479760 228636 487436 228664
rect 479760 228624 479766 228636
rect 487430 228624 487436 228636
rect 487488 228624 487494 228676
rect 495342 228624 495348 228676
rect 495400 228664 495406 228676
rect 511442 228664 511448 228676
rect 495400 228636 511448 228664
rect 495400 228624 495406 228636
rect 511442 228624 511448 228636
rect 511500 228624 511506 228676
rect 528186 228624 528192 228676
rect 528244 228664 528250 228676
rect 553670 228664 553676 228676
rect 528244 228636 553676 228664
rect 528244 228624 528250 228636
rect 553670 228624 553676 228636
rect 553728 228624 553734 228676
rect 672718 228556 672724 228608
rect 672776 228596 672782 228608
rect 672902 228596 672908 228608
rect 672776 228568 672908 228596
rect 672776 228556 672782 228568
rect 672902 228556 672908 228568
rect 672960 228556 672966 228608
rect 673388 228540 673440 228546
rect 366910 228488 366916 228540
rect 366968 228528 366974 228540
rect 381998 228528 382004 228540
rect 366968 228500 382004 228528
rect 366968 228488 366974 228500
rect 381998 228488 382004 228500
rect 382056 228488 382062 228540
rect 392854 228528 392860 228540
rect 383626 228500 392860 228528
rect 355376 228364 359044 228392
rect 355376 228352 355382 228364
rect 362862 228352 362868 228404
rect 362920 228392 362926 228404
rect 379422 228392 379428 228404
rect 362920 228364 379428 228392
rect 362920 228352 362926 228364
rect 379422 228352 379428 228364
rect 379480 228352 379486 228404
rect 381906 228352 381912 228404
rect 381964 228392 381970 228404
rect 383626 228392 383654 228500
rect 392854 228488 392860 228500
rect 392912 228488 392918 228540
rect 393038 228488 393044 228540
rect 393096 228528 393102 228540
rect 393096 228500 397960 228528
rect 393096 228488 393102 228500
rect 381964 228364 383654 228392
rect 381964 228352 381970 228364
rect 391842 228352 391848 228404
rect 391900 228392 391906 228404
rect 397932 228392 397960 228500
rect 400030 228488 400036 228540
rect 400088 228528 400094 228540
rect 407758 228528 407764 228540
rect 400088 228500 407764 228528
rect 400088 228488 400094 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 482462 228488 482468 228540
rect 482520 228528 482526 228540
rect 494698 228528 494704 228540
rect 482520 228500 494704 228528
rect 482520 228488 482526 228500
rect 494698 228488 494704 228500
rect 494756 228488 494762 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 520918 228528 520924 228540
rect 502484 228500 520924 228528
rect 502484 228488 502490 228500
rect 520918 228488 520924 228500
rect 520976 228488 520982 228540
rect 531406 228488 531412 228540
rect 531464 228528 531470 228540
rect 558178 228528 558184 228540
rect 531464 228500 558184 228528
rect 531464 228488 531470 228500
rect 558178 228488 558184 228500
rect 558236 228488 558242 228540
rect 673388 228482 673440 228488
rect 672258 228420 672264 228472
rect 672316 228460 672322 228472
rect 672316 228432 673302 228460
rect 672316 228420 672322 228432
rect 402606 228392 402612 228404
rect 391900 228364 393314 228392
rect 397932 228364 402612 228392
rect 391900 228352 391906 228364
rect 108114 228216 108120 228268
rect 108172 228256 108178 228268
rect 140958 228256 140964 228268
rect 108172 228228 140964 228256
rect 108172 228216 108178 228228
rect 140958 228216 140964 228228
rect 141016 228216 141022 228268
rect 141142 228216 141148 228268
rect 141200 228256 141206 228268
rect 190914 228256 190920 228268
rect 141200 228228 190920 228256
rect 141200 228216 141206 228228
rect 190914 228216 190920 228228
rect 190972 228216 190978 228268
rect 204898 228256 204904 228268
rect 191116 228228 204904 228256
rect 106182 228080 106188 228132
rect 106240 228120 106246 228132
rect 108482 228120 108488 228132
rect 106240 228092 108488 228120
rect 106240 228080 106246 228092
rect 108482 228080 108488 228092
rect 108540 228080 108546 228132
rect 113082 228080 113088 228132
rect 113140 228120 113146 228132
rect 181070 228120 181076 228132
rect 113140 228092 181076 228120
rect 113140 228080 113146 228092
rect 181070 228080 181076 228092
rect 181128 228080 181134 228132
rect 181254 228080 181260 228132
rect 181312 228120 181318 228132
rect 191116 228120 191144 228228
rect 204898 228216 204904 228228
rect 204956 228216 204962 228268
rect 252554 228256 252560 228268
rect 205100 228228 252560 228256
rect 201034 228120 201040 228132
rect 181312 228092 191144 228120
rect 195946 228092 201040 228120
rect 181312 228080 181318 228092
rect 122742 227944 122748 227996
rect 122800 227984 122806 227996
rect 181714 227984 181720 227996
rect 122800 227956 181720 227984
rect 122800 227944 122806 227956
rect 181714 227944 181720 227956
rect 181772 227944 181778 227996
rect 181898 227944 181904 227996
rect 181956 227984 181962 227996
rect 184934 227984 184940 227996
rect 181956 227956 184940 227984
rect 181956 227944 181962 227956
rect 184934 227944 184940 227956
rect 184992 227944 184998 227996
rect 190914 227944 190920 227996
rect 190972 227984 190978 227996
rect 195946 227984 195974 228092
rect 201034 228080 201040 228092
rect 201092 228080 201098 228132
rect 201402 228080 201408 228132
rect 201460 228120 201466 228132
rect 205100 228120 205128 228228
rect 252554 228216 252560 228228
rect 252612 228216 252618 228268
rect 277118 228216 277124 228268
rect 277176 228256 277182 228268
rect 311802 228256 311808 228268
rect 277176 228228 311808 228256
rect 277176 228216 277182 228228
rect 311802 228216 311808 228228
rect 311860 228216 311866 228268
rect 393286 228256 393314 228364
rect 402606 228352 402612 228364
rect 402664 228352 402670 228404
rect 409598 228352 409604 228404
rect 409656 228392 409662 228404
rect 415486 228392 415492 228404
rect 409656 228364 415492 228392
rect 409656 228352 409662 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 486970 228352 486976 228404
rect 487028 228392 487034 228404
rect 501690 228392 501696 228404
rect 487028 228364 501696 228392
rect 487028 228352 487034 228364
rect 501690 228352 501696 228364
rect 501748 228352 501754 228404
rect 506290 228352 506296 228404
rect 506348 228392 506354 228404
rect 526530 228392 526536 228404
rect 506348 228364 526536 228392
rect 506348 228352 506354 228364
rect 526530 228352 526536 228364
rect 526588 228352 526594 228404
rect 537846 228352 537852 228404
rect 537904 228392 537910 228404
rect 566182 228392 566188 228404
rect 537904 228364 566188 228392
rect 537904 228352 537910 228364
rect 566182 228352 566188 228364
rect 566240 228352 566246 228404
rect 403894 228256 403900 228268
rect 393286 228228 403900 228256
rect 403894 228216 403900 228228
rect 403952 228216 403958 228268
rect 478690 228216 478696 228268
rect 478748 228256 478754 228268
rect 487062 228256 487068 228268
rect 478748 228228 487068 228256
rect 478748 228216 478754 228228
rect 487062 228216 487068 228228
rect 487120 228216 487126 228268
rect 512086 228216 512092 228268
rect 512144 228256 512150 228268
rect 533522 228256 533528 228268
rect 512144 228228 533528 228256
rect 512144 228216 512150 228228
rect 533522 228216 533528 228228
rect 533580 228216 533586 228268
rect 671338 228216 671344 228268
rect 671396 228256 671402 228268
rect 671396 228228 673190 228256
rect 671396 228216 671402 228228
rect 201460 228092 205128 228120
rect 201460 228080 201466 228092
rect 205450 228080 205456 228132
rect 205508 228120 205514 228132
rect 257062 228120 257068 228132
rect 205508 228092 257068 228120
rect 205508 228080 205514 228092
rect 257062 228080 257068 228092
rect 257120 228080 257126 228132
rect 288066 228080 288072 228132
rect 288124 228120 288130 228132
rect 321462 228120 321468 228132
rect 288124 228092 321468 228120
rect 288124 228080 288130 228092
rect 321462 228080 321468 228092
rect 321520 228080 321526 228132
rect 671890 228012 671896 228064
rect 671948 228052 671954 228064
rect 671948 228024 673072 228052
rect 671948 228012 671954 228024
rect 190972 227956 195974 227984
rect 190972 227944 190978 227956
rect 197998 227944 198004 227996
rect 198056 227984 198062 227996
rect 204530 227984 204536 227996
rect 198056 227956 204536 227984
rect 198056 227944 198062 227956
rect 204530 227944 204536 227956
rect 204588 227944 204594 227996
rect 212166 227944 212172 227996
rect 212224 227984 212230 227996
rect 218422 227984 218428 227996
rect 212224 227956 218428 227984
rect 212224 227944 212230 227956
rect 218422 227944 218428 227956
rect 218480 227944 218486 227996
rect 222746 227944 222752 227996
rect 222804 227984 222810 227996
rect 226150 227984 226156 227996
rect 222804 227956 226156 227984
rect 222804 227944 222810 227956
rect 226150 227944 226156 227956
rect 226208 227944 226214 227996
rect 272518 227984 272524 227996
rect 229066 227956 272524 227984
rect 133782 227808 133788 227860
rect 133840 227848 133846 227860
rect 200390 227848 200396 227860
rect 133840 227820 200396 227848
rect 133840 227808 133846 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 204714 227808 204720 227860
rect 204772 227848 204778 227860
rect 210694 227848 210700 227860
rect 204772 227820 210700 227848
rect 204772 227808 204778 227820
rect 210694 227808 210700 227820
rect 210752 227808 210758 227860
rect 226150 227808 226156 227860
rect 226208 227848 226214 227860
rect 229066 227848 229094 227956
rect 272518 227944 272524 227956
rect 272576 227944 272582 227996
rect 369118 227876 369124 227928
rect 369176 227916 369182 227928
rect 375558 227916 375564 227928
rect 369176 227888 375564 227916
rect 369176 227876 369182 227888
rect 375558 227876 375564 227888
rect 375616 227876 375622 227928
rect 407758 227876 407764 227928
rect 407816 227916 407822 227928
rect 411622 227916 411628 227928
rect 407816 227888 411628 227916
rect 407816 227876 407822 227888
rect 411622 227876 411628 227888
rect 411680 227876 411686 227928
rect 471514 227876 471520 227928
rect 471572 227916 471578 227928
rect 479242 227916 479248 227928
rect 471572 227888 479248 227916
rect 471572 227876 471578 227888
rect 479242 227876 479248 227888
rect 479300 227876 479306 227928
rect 226208 227820 229094 227848
rect 226208 227808 226214 227820
rect 672954 227792 673006 227798
rect 242526 227740 242532 227792
rect 242584 227780 242590 227792
rect 245654 227780 245660 227792
rect 242584 227752 245660 227780
rect 242584 227740 242590 227752
rect 245654 227740 245660 227752
rect 245712 227740 245718 227792
rect 255958 227740 255964 227792
rect 256016 227780 256022 227792
rect 258994 227780 259000 227792
rect 256016 227752 259000 227780
rect 256016 227740 256022 227752
rect 258994 227740 259000 227752
rect 259052 227740 259058 227792
rect 366266 227740 366272 227792
rect 366324 227780 366330 227792
rect 372982 227780 372988 227792
rect 366324 227752 372988 227780
rect 366324 227740 366330 227752
rect 372982 227740 372988 227752
rect 373040 227740 373046 227792
rect 393958 227740 393964 227792
rect 394016 227780 394022 227792
rect 395522 227780 395528 227792
rect 394016 227752 395528 227780
rect 394016 227740 394022 227752
rect 395522 227740 395528 227752
rect 395580 227740 395586 227792
rect 396718 227740 396724 227792
rect 396776 227780 396782 227792
rect 397454 227780 397460 227792
rect 396776 227752 397460 227780
rect 396776 227740 396782 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 402238 227740 402244 227792
rect 402296 227780 402302 227792
rect 403250 227780 403256 227792
rect 402296 227752 403256 227780
rect 402296 227740 402302 227752
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 404078 227740 404084 227792
rect 404136 227780 404142 227792
rect 408862 227780 408868 227792
rect 404136 227752 408868 227780
rect 404136 227740 404142 227752
rect 408862 227740 408868 227752
rect 408920 227740 408926 227792
rect 409138 227740 409144 227792
rect 409196 227780 409202 227792
rect 410334 227780 410340 227792
rect 409196 227752 410340 227780
rect 409196 227740 409202 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416590 227740 416596 227792
rect 416648 227780 416654 227792
rect 420638 227780 420644 227792
rect 416648 227752 420644 227780
rect 416648 227740 416654 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 475010 227740 475016 227792
rect 475068 227780 475074 227792
rect 482830 227780 482836 227792
rect 475068 227752 482836 227780
rect 475068 227740 475074 227752
rect 482830 227740 482836 227752
rect 482888 227740 482894 227792
rect 510614 227740 510620 227792
rect 510672 227780 510678 227792
rect 513006 227780 513012 227792
rect 510672 227752 513012 227780
rect 510672 227740 510678 227752
rect 513006 227740 513012 227752
rect 513064 227740 513070 227792
rect 663702 227740 663708 227792
rect 663760 227780 663766 227792
rect 665266 227780 665272 227792
rect 663760 227752 665272 227780
rect 663760 227740 663766 227752
rect 665266 227740 665272 227752
rect 665324 227740 665330 227792
rect 672954 227734 673006 227740
rect 109862 227672 109868 227724
rect 109920 227712 109926 227724
rect 182358 227712 182364 227724
rect 109920 227684 182364 227712
rect 109920 227672 109926 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 184566 227672 184572 227724
rect 184624 227712 184630 227724
rect 187510 227712 187516 227724
rect 184624 227684 187516 227712
rect 184624 227672 184630 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 191742 227672 191748 227724
rect 191800 227712 191806 227724
rect 191800 227684 238754 227712
rect 191800 227672 191806 227684
rect 238726 227644 238754 227684
rect 270310 227672 270316 227724
rect 270368 227712 270374 227724
rect 306650 227712 306656 227724
rect 270368 227684 306656 227712
rect 270368 227672 270374 227684
rect 306650 227672 306656 227684
rect 306708 227672 306714 227724
rect 321370 227672 321376 227724
rect 321428 227712 321434 227724
rect 346578 227712 346584 227724
rect 321428 227684 346584 227712
rect 321428 227672 321434 227684
rect 346578 227672 346584 227684
rect 346636 227672 346642 227724
rect 528922 227672 528928 227724
rect 528980 227712 528986 227724
rect 549898 227712 549904 227724
rect 528980 227684 549904 227712
rect 528980 227672 528986 227684
rect 549898 227672 549904 227684
rect 549956 227672 549962 227724
rect 248046 227644 248052 227656
rect 238726 227616 248052 227644
rect 248046 227604 248052 227616
rect 248104 227604 248110 227656
rect 670510 227604 670516 227656
rect 670568 227644 670574 227656
rect 670568 227616 672842 227644
rect 670568 227604 670574 227616
rect 100662 227536 100668 227588
rect 100720 227576 100726 227588
rect 174630 227576 174636 227588
rect 100720 227548 174636 227576
rect 100720 227536 100726 227548
rect 174630 227536 174636 227548
rect 174688 227536 174694 227588
rect 179322 227536 179328 227588
rect 179380 227576 179386 227588
rect 236454 227576 236460 227588
rect 179380 227548 236460 227576
rect 179380 227536 179386 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 252278 227536 252284 227588
rect 252336 227576 252342 227588
rect 293126 227576 293132 227588
rect 252336 227548 293132 227576
rect 252336 227536 252342 227548
rect 293126 227536 293132 227548
rect 293184 227536 293190 227588
rect 299198 227536 299204 227588
rect 299256 227576 299262 227588
rect 328546 227576 328552 227588
rect 299256 227548 328552 227576
rect 299256 227536 299262 227548
rect 328546 227536 328552 227548
rect 328604 227536 328610 227588
rect 359458 227536 359464 227588
rect 359516 227576 359522 227588
rect 374914 227576 374920 227588
rect 359516 227548 374920 227576
rect 359516 227536 359522 227548
rect 374914 227536 374920 227548
rect 374972 227536 374978 227588
rect 465902 227536 465908 227588
rect 465960 227576 465966 227588
rect 469858 227576 469864 227588
rect 465960 227548 469864 227576
rect 465960 227536 465966 227548
rect 469858 227536 469864 227548
rect 469916 227536 469922 227588
rect 518526 227536 518532 227588
rect 518584 227576 518590 227588
rect 541618 227576 541624 227588
rect 518584 227548 541624 227576
rect 518584 227536 518590 227548
rect 541618 227536 541624 227548
rect 541676 227536 541682 227588
rect 560938 227536 560944 227588
rect 560996 227576 561002 227588
rect 567654 227576 567660 227588
rect 560996 227548 567660 227576
rect 560996 227536 561002 227548
rect 567654 227536 567660 227548
rect 567712 227536 567718 227588
rect 89622 227400 89628 227452
rect 89680 227440 89686 227452
rect 159634 227440 159640 227452
rect 89680 227412 159640 227440
rect 89680 227400 89686 227412
rect 159634 227400 159640 227412
rect 159692 227400 159698 227452
rect 160002 227400 160008 227452
rect 160060 227440 160066 227452
rect 166902 227440 166908 227452
rect 160060 227412 166908 227440
rect 160060 227400 160066 227412
rect 166902 227400 166908 227412
rect 166960 227400 166966 227452
rect 171106 227412 173756 227440
rect 86678 227264 86684 227316
rect 86736 227304 86742 227316
rect 164326 227304 164332 227316
rect 86736 227276 164332 227304
rect 86736 227264 86742 227276
rect 164326 227264 164332 227276
rect 164384 227264 164390 227316
rect 165338 227264 165344 227316
rect 165396 227304 165402 227316
rect 171106 227304 171134 227412
rect 165396 227276 171134 227304
rect 173728 227304 173756 227412
rect 174998 227400 175004 227452
rect 175056 227440 175062 227452
rect 231946 227440 231952 227452
rect 175056 227412 231952 227440
rect 175056 227400 175062 227412
rect 231946 227400 231952 227412
rect 232004 227400 232010 227452
rect 248138 227400 248144 227452
rect 248196 227440 248202 227452
rect 291838 227440 291844 227452
rect 248196 227412 291844 227440
rect 248196 227400 248202 227412
rect 291838 227400 291844 227412
rect 291896 227400 291902 227452
rect 293678 227400 293684 227452
rect 293736 227440 293742 227452
rect 325326 227440 325332 227452
rect 293736 227412 325332 227440
rect 293736 227400 293742 227412
rect 325326 227400 325332 227412
rect 325384 227400 325390 227452
rect 340598 227400 340604 227452
rect 340656 227440 340662 227452
rect 361390 227440 361396 227452
rect 340656 227412 361396 227440
rect 340656 227400 340662 227412
rect 361390 227400 361396 227412
rect 361448 227400 361454 227452
rect 377214 227440 377220 227452
rect 362052 227412 377220 227440
rect 227438 227304 227444 227316
rect 173728 227276 227444 227304
rect 165396 227264 165402 227276
rect 227438 227264 227444 227276
rect 227496 227264 227502 227316
rect 233234 227304 233240 227316
rect 228928 227276 233240 227304
rect 75822 227128 75828 227180
rect 75880 227168 75886 227180
rect 151722 227168 151728 227180
rect 75880 227140 151728 227168
rect 75880 227128 75886 227140
rect 151722 227128 151728 227140
rect 151780 227128 151786 227180
rect 152274 227128 152280 227180
rect 152332 227168 152338 227180
rect 156506 227168 156512 227180
rect 152332 227140 156512 227168
rect 152332 227128 152338 227140
rect 156506 227128 156512 227140
rect 156564 227128 156570 227180
rect 168834 227168 168840 227180
rect 156800 227140 168840 227168
rect 57698 226992 57704 227044
rect 57756 227032 57762 227044
rect 135254 227032 135260 227044
rect 57756 227004 135260 227032
rect 57756 226992 57762 227004
rect 135254 226992 135260 227004
rect 135312 226992 135318 227044
rect 135438 226992 135444 227044
rect 135496 227032 135502 227044
rect 156800 227032 156828 227140
rect 168834 227128 168840 227140
rect 168892 227128 168898 227180
rect 169478 227128 169484 227180
rect 169536 227168 169542 227180
rect 228726 227168 228732 227180
rect 169536 227140 228732 227168
rect 169536 227128 169542 227140
rect 228726 227128 228732 227140
rect 228784 227128 228790 227180
rect 135496 227004 156828 227032
rect 135496 226992 135502 227004
rect 156966 226992 156972 227044
rect 157024 227032 157030 227044
rect 213270 227032 213276 227044
rect 157024 227004 213276 227032
rect 157024 226992 157030 227004
rect 213270 226992 213276 227004
rect 213328 226992 213334 227044
rect 226978 226992 226984 227044
rect 227036 227032 227042 227044
rect 228928 227032 228956 227276
rect 233234 227264 233240 227276
rect 233292 227264 233298 227316
rect 234522 227264 234528 227316
rect 234580 227304 234586 227316
rect 278314 227304 278320 227316
rect 234580 227276 278320 227304
rect 234580 227264 234586 227276
rect 278314 227264 278320 227276
rect 278372 227264 278378 227316
rect 280798 227264 280804 227316
rect 280856 227304 280862 227316
rect 312078 227304 312084 227316
rect 280856 227276 312084 227304
rect 280856 227264 280862 227276
rect 312078 227264 312084 227276
rect 312136 227264 312142 227316
rect 326338 227264 326344 227316
rect 326396 227304 326402 227316
rect 352374 227304 352380 227316
rect 326396 227276 352380 227304
rect 326396 227264 326402 227276
rect 352374 227264 352380 227276
rect 352432 227264 352438 227316
rect 361298 227264 361304 227316
rect 361356 227304 361362 227316
rect 362052 227304 362080 227412
rect 377214 227400 377220 227412
rect 377272 227400 377278 227452
rect 383286 227440 383292 227452
rect 378612 227412 383292 227440
rect 361356 227276 362080 227304
rect 361356 227264 361362 227276
rect 362218 227264 362224 227316
rect 362276 227304 362282 227316
rect 372338 227304 372344 227316
rect 362276 227276 372344 227304
rect 362276 227264 362282 227276
rect 372338 227264 372344 227276
rect 372396 227264 372402 227316
rect 373258 227264 373264 227316
rect 373316 227304 373322 227316
rect 378612 227304 378640 227412
rect 383286 227400 383292 227412
rect 383344 227400 383350 227452
rect 515950 227400 515956 227452
rect 516008 227440 516014 227452
rect 538490 227440 538496 227452
rect 516008 227412 538496 227440
rect 516008 227400 516014 227412
rect 538490 227400 538496 227412
rect 538548 227400 538554 227452
rect 672724 227384 672776 227390
rect 672258 227332 672264 227384
rect 672316 227372 672322 227384
rect 672316 227344 672488 227372
rect 672316 227332 672322 227344
rect 373316 227276 378640 227304
rect 373316 227264 373322 227276
rect 382826 227264 382832 227316
rect 382884 227304 382890 227316
rect 391658 227304 391664 227316
rect 382884 227276 391664 227304
rect 382884 227264 382890 227276
rect 391658 227264 391664 227276
rect 391716 227264 391722 227316
rect 395982 227264 395988 227316
rect 396040 227304 396046 227316
rect 406470 227304 406476 227316
rect 396040 227276 406476 227304
rect 396040 227264 396046 227276
rect 406470 227264 406476 227276
rect 406528 227264 406534 227316
rect 485038 227264 485044 227316
rect 485096 227304 485102 227316
rect 498838 227304 498844 227316
rect 485096 227276 498844 227304
rect 485096 227264 485102 227276
rect 498838 227264 498844 227276
rect 498896 227264 498902 227316
rect 501322 227264 501328 227316
rect 501380 227304 501386 227316
rect 517790 227304 517796 227316
rect 501380 227276 517796 227304
rect 501380 227264 501386 227276
rect 517790 227264 517796 227276
rect 517848 227264 517854 227316
rect 521746 227264 521752 227316
rect 521804 227304 521810 227316
rect 545758 227304 545764 227316
rect 521804 227276 545764 227304
rect 521804 227264 521810 227276
rect 545758 227264 545764 227276
rect 545816 227264 545822 227316
rect 672460 227236 672488 227344
rect 672724 227326 672776 227332
rect 672460 227208 672630 227236
rect 235718 227128 235724 227180
rect 235776 227168 235782 227180
rect 280246 227168 280252 227180
rect 235776 227140 280252 227168
rect 235776 227128 235782 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 296162 227128 296168 227180
rect 296220 227168 296226 227180
rect 329190 227168 329196 227180
rect 296220 227140 329196 227168
rect 296220 227128 296226 227140
rect 329190 227128 329196 227140
rect 329248 227128 329254 227180
rect 329742 227128 329748 227180
rect 329800 227168 329806 227180
rect 353662 227168 353668 227180
rect 329800 227140 353668 227168
rect 329800 227128 329806 227140
rect 353662 227128 353668 227140
rect 353720 227128 353726 227180
rect 354582 227128 354588 227180
rect 354640 227168 354646 227180
rect 373626 227168 373632 227180
rect 354640 227140 373632 227168
rect 354640 227128 354646 227140
rect 373626 227128 373632 227140
rect 373684 227128 373690 227180
rect 382090 227128 382096 227180
rect 382148 227168 382154 227180
rect 396166 227168 396172 227180
rect 382148 227140 396172 227168
rect 382148 227128 382154 227140
rect 396166 227128 396172 227140
rect 396224 227128 396230 227180
rect 498562 227128 498568 227180
rect 498620 227168 498626 227180
rect 516042 227168 516048 227180
rect 498620 227140 516048 227168
rect 498620 227128 498626 227140
rect 516042 227128 516048 227140
rect 516100 227128 516106 227180
rect 533982 227128 533988 227180
rect 534040 227168 534046 227180
rect 561490 227168 561496 227180
rect 534040 227140 561496 227168
rect 534040 227128 534046 227140
rect 561490 227128 561496 227140
rect 561548 227128 561554 227180
rect 227036 227004 228956 227032
rect 227036 226992 227042 227004
rect 229048 226992 229054 227044
rect 229106 227032 229112 227044
rect 271230 227032 271236 227044
rect 229106 227004 271236 227032
rect 229106 226992 229112 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 336274 227032 336280 227044
rect 316006 227004 336280 227032
rect 106918 226856 106924 226908
rect 106976 226896 106982 226908
rect 125778 226896 125784 226908
rect 106976 226868 125784 226896
rect 106976 226856 106982 226868
rect 125778 226856 125784 226868
rect 125836 226856 125842 226908
rect 190454 226896 190460 226908
rect 125980 226868 190460 226896
rect 121362 226720 121368 226772
rect 121420 226760 121426 226772
rect 125980 226760 126008 226868
rect 190454 226856 190460 226868
rect 190512 226856 190518 226908
rect 200022 226856 200028 226908
rect 200080 226896 200086 226908
rect 252002 226896 252008 226908
rect 200080 226868 252008 226896
rect 200080 226856 200086 226868
rect 252002 226856 252008 226868
rect 252060 226856 252066 226908
rect 272518 226856 272524 226908
rect 272576 226896 272582 226908
rect 284754 226896 284760 226908
rect 272576 226868 284760 226896
rect 272576 226856 272582 226868
rect 284754 226856 284760 226868
rect 284812 226856 284818 226908
rect 308582 226856 308588 226908
rect 308640 226896 308646 226908
rect 316006 226896 316034 227004
rect 336274 226992 336280 227004
rect 336332 226992 336338 227044
rect 336458 226992 336464 227044
rect 336516 227032 336522 227044
rect 360102 227032 360108 227044
rect 336516 227004 360108 227032
rect 336516 226992 336522 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 369762 226992 369768 227044
rect 369820 227032 369826 227044
rect 385862 227032 385868 227044
rect 369820 227004 385868 227032
rect 369820 226992 369826 227004
rect 385862 226992 385868 227004
rect 385920 226992 385926 227044
rect 386322 226992 386328 227044
rect 386380 227032 386386 227044
rect 398742 227032 398748 227044
rect 386380 227004 398748 227032
rect 386380 226992 386386 227004
rect 398742 226992 398748 227004
rect 398800 226992 398806 227044
rect 472158 226992 472164 227044
rect 472216 227032 472222 227044
rect 480806 227032 480812 227044
rect 472216 227004 480812 227032
rect 472216 226992 472222 227004
rect 480806 226992 480812 227004
rect 480864 226992 480870 227044
rect 481174 226992 481180 227044
rect 481232 227032 481238 227044
rect 493962 227032 493968 227044
rect 481232 227004 493968 227032
rect 481232 226992 481238 227004
rect 493962 226992 493968 227004
rect 494020 226992 494026 227044
rect 497274 226992 497280 227044
rect 497332 227032 497338 227044
rect 513834 227032 513840 227044
rect 497332 227004 513840 227032
rect 497332 226992 497338 227004
rect 513834 226992 513840 227004
rect 513892 226992 513898 227044
rect 514018 226992 514024 227044
rect 514076 227032 514082 227044
rect 536098 227032 536104 227044
rect 514076 227004 536104 227032
rect 514076 226992 514082 227004
rect 536098 226992 536104 227004
rect 536156 226992 536162 227044
rect 537202 226992 537208 227044
rect 537260 227032 537266 227044
rect 565354 227032 565360 227044
rect 537260 227004 565360 227032
rect 537260 226992 537266 227004
rect 565354 226992 565360 227004
rect 565412 226992 565418 227044
rect 670510 226992 670516 227044
rect 670568 227032 670574 227044
rect 670568 227004 672520 227032
rect 670568 226992 670574 227004
rect 308640 226868 316034 226896
rect 308640 226856 308646 226868
rect 355502 226856 355508 226908
rect 355560 226896 355566 226908
rect 362218 226896 362224 226908
rect 355560 226868 362224 226896
rect 355560 226856 355566 226868
rect 362218 226856 362224 226868
rect 362276 226856 362282 226908
rect 398742 226856 398748 226908
rect 398800 226896 398806 226908
rect 408678 226896 408684 226908
rect 398800 226868 408684 226896
rect 398800 226856 398806 226868
rect 408678 226856 408684 226868
rect 408736 226856 408742 226908
rect 671890 226788 671896 226840
rect 671948 226828 671954 226840
rect 671948 226800 672406 226828
rect 671948 226788 671954 226800
rect 190086 226760 190092 226772
rect 121420 226732 126008 226760
rect 126072 226732 190092 226760
rect 121420 226720 121426 226732
rect 119798 226584 119804 226636
rect 119856 226624 119862 226636
rect 126072 226624 126100 226732
rect 190086 226720 190092 226732
rect 190144 226720 190150 226772
rect 195882 226720 195888 226772
rect 195940 226760 195946 226772
rect 199286 226760 199292 226772
rect 195940 226732 199292 226760
rect 195940 226720 195946 226732
rect 199286 226720 199292 226732
rect 199344 226720 199350 226772
rect 212350 226720 212356 226772
rect 212408 226760 212414 226772
rect 262214 226760 262220 226772
rect 212408 226732 262220 226760
rect 212408 226720 212414 226732
rect 262214 226720 262220 226732
rect 262272 226720 262278 226772
rect 135438 226624 135444 226636
rect 119856 226596 126100 226624
rect 126164 226596 135444 226624
rect 119856 226584 119862 226596
rect 125778 226448 125784 226500
rect 125836 226488 125842 226500
rect 126164 226488 126192 226596
rect 135438 226584 135444 226596
rect 135496 226584 135502 226636
rect 135622 226584 135628 226636
rect 135680 226624 135686 226636
rect 135680 226596 137416 226624
rect 135680 226584 135686 226596
rect 125836 226460 126192 226488
rect 125836 226448 125842 226460
rect 129642 226448 129648 226500
rect 129700 226488 129706 226500
rect 137186 226488 137192 226500
rect 129700 226460 137192 226488
rect 129700 226448 129706 226460
rect 137186 226448 137192 226460
rect 137244 226448 137250 226500
rect 137388 226488 137416 226596
rect 137554 226584 137560 226636
rect 137612 226624 137618 226636
rect 197354 226624 197360 226636
rect 137612 226596 197360 226624
rect 137612 226584 137618 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 222010 226584 222016 226636
rect 222068 226624 222074 226636
rect 269942 226624 269948 226636
rect 222068 226596 269948 226624
rect 222068 226584 222074 226596
rect 269942 226584 269948 226596
rect 270000 226584 270006 226636
rect 672046 226596 672290 226624
rect 672046 226556 672074 226596
rect 671908 226528 672074 226556
rect 142108 226488 142114 226500
rect 137388 226460 142114 226488
rect 142108 226448 142114 226460
rect 142166 226448 142172 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 205174 226488 205180 226500
rect 142304 226460 205180 226488
rect 142304 226448 142310 226460
rect 205174 226448 205180 226460
rect 205232 226448 205238 226500
rect 213178 226448 213184 226500
rect 213236 226488 213242 226500
rect 217778 226488 217784 226500
rect 213236 226460 217784 226488
rect 213236 226448 213242 226460
rect 217778 226448 217784 226460
rect 217836 226448 217842 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 229002 226488 229008 226500
rect 221884 226460 229008 226488
rect 221884 226448 221890 226460
rect 229002 226448 229008 226460
rect 229060 226448 229066 226500
rect 232498 226448 232504 226500
rect 232556 226488 232562 226500
rect 266722 226488 266728 226500
rect 232556 226460 266728 226488
rect 232556 226448 232562 226460
rect 266722 226448 266728 226460
rect 266780 226448 266786 226500
rect 291838 226380 291844 226432
rect 291896 226420 291902 226432
rect 295058 226420 295064 226432
rect 291896 226392 295064 226420
rect 291896 226380 291902 226392
rect 295058 226380 295064 226392
rect 295116 226380 295122 226432
rect 671908 226364 671936 226528
rect 672156 226500 672208 226506
rect 672156 226442 672208 226448
rect 154408 226324 154620 226352
rect 83458 226244 83464 226296
rect 83516 226284 83522 226296
rect 154206 226284 154212 226296
rect 83516 226256 154212 226284
rect 83516 226244 83522 226256
rect 154206 226244 154212 226256
rect 154264 226244 154270 226296
rect 69658 226108 69664 226160
rect 69716 226148 69722 226160
rect 143534 226148 143540 226160
rect 69716 226120 143540 226148
rect 69716 226108 69722 226120
rect 143534 226108 143540 226120
rect 143592 226108 143598 226160
rect 146938 226108 146944 226160
rect 146996 226148 147002 226160
rect 154408 226148 154436 226324
rect 154592 226284 154620 226324
rect 166948 226312 166954 226364
rect 167006 226352 167012 226364
rect 220998 226352 221004 226364
rect 167006 226324 221004 226352
rect 167006 226312 167012 226324
rect 220998 226312 221004 226324
rect 221056 226312 221062 226364
rect 490098 226312 490104 226364
rect 490156 226352 490162 226364
rect 494882 226352 494888 226364
rect 490156 226324 494888 226352
rect 490156 226312 490162 226324
rect 494882 226312 494888 226324
rect 494940 226312 494946 226364
rect 671890 226312 671896 226364
rect 671948 226312 671954 226364
rect 672034 226296 672086 226302
rect 161934 226284 161940 226296
rect 154592 226256 161940 226284
rect 161934 226244 161940 226256
rect 161992 226244 161998 226296
rect 162302 226244 162308 226296
rect 162360 226284 162366 226296
rect 166810 226284 166816 226296
rect 162360 226256 166816 226284
rect 162360 226244 162366 226256
rect 166810 226244 166816 226256
rect 166868 226244 166874 226296
rect 222470 226244 222476 226296
rect 222528 226284 222534 226296
rect 225506 226284 225512 226296
rect 222528 226256 225512 226284
rect 222528 226244 222534 226256
rect 225506 226244 225512 226256
rect 225564 226244 225570 226296
rect 228910 226244 228916 226296
rect 228968 226284 228974 226296
rect 275094 226284 275100 226296
rect 228968 226256 275100 226284
rect 228968 226244 228974 226256
rect 275094 226244 275100 226256
rect 275152 226244 275158 226296
rect 278406 226244 278412 226296
rect 278464 226284 278470 226296
rect 315022 226284 315028 226296
rect 278464 226256 315028 226284
rect 278464 226244 278470 226256
rect 315022 226244 315028 226256
rect 315080 226244 315086 226296
rect 317322 226244 317328 226296
rect 317380 226284 317386 226296
rect 334250 226284 334256 226296
rect 317380 226256 334256 226284
rect 317380 226244 317386 226256
rect 334250 226244 334256 226256
rect 334308 226244 334314 226296
rect 672034 226238 672086 226244
rect 146996 226120 154436 226148
rect 146996 226108 147002 226120
rect 154758 226108 154764 226160
rect 154816 226148 154822 226160
rect 157426 226148 157432 226160
rect 154816 226120 157432 226148
rect 154816 226108 154822 226120
rect 157426 226108 157432 226120
rect 157484 226108 157490 226160
rect 157610 226108 157616 226160
rect 157668 226148 157674 226160
rect 215846 226148 215852 226160
rect 157668 226120 215852 226148
rect 157668 226108 157674 226120
rect 215846 226108 215852 226120
rect 215904 226108 215910 226160
rect 216490 226108 216496 226160
rect 216548 226148 216554 226160
rect 264790 226148 264796 226160
rect 216548 226120 264796 226148
rect 216548 226108 216554 226120
rect 264790 226108 264796 226120
rect 264848 226108 264854 226160
rect 266262 226108 266268 226160
rect 266320 226148 266326 226160
rect 303430 226148 303436 226160
rect 266320 226120 303436 226148
rect 266320 226108 266326 226120
rect 303430 226108 303436 226120
rect 303488 226108 303494 226160
rect 325602 226108 325608 226160
rect 325660 226148 325666 226160
rect 349154 226148 349160 226160
rect 325660 226120 349160 226148
rect 325660 226108 325666 226120
rect 349154 226108 349160 226120
rect 349212 226108 349218 226160
rect 514662 226108 514668 226160
rect 514720 226148 514726 226160
rect 535454 226148 535460 226160
rect 514720 226120 535460 226148
rect 514720 226108 514726 226120
rect 535454 226108 535460 226120
rect 535512 226108 535518 226160
rect 667842 226040 667848 226092
rect 667900 226080 667906 226092
rect 667900 226052 671968 226080
rect 667900 226040 667906 226052
rect 93762 225972 93768 226024
rect 93820 226012 93826 226024
rect 161566 226012 161572 226024
rect 93820 225984 161572 226012
rect 93820 225972 93826 225984
rect 161566 225972 161572 225984
rect 161624 225972 161630 226024
rect 161934 225972 161940 226024
rect 161992 226012 161998 226024
rect 171042 226012 171048 226024
rect 161992 225984 171048 226012
rect 161992 225972 161998 225984
rect 171042 225972 171048 225984
rect 171100 225972 171106 226024
rect 171226 225972 171232 226024
rect 171284 226012 171290 226024
rect 186406 226012 186412 226024
rect 171284 225984 186412 226012
rect 171284 225972 171290 225984
rect 186406 225972 186412 225984
rect 186464 225972 186470 226024
rect 186590 225972 186596 226024
rect 186648 226012 186654 226024
rect 224218 226012 224224 226024
rect 186648 225984 224224 226012
rect 186648 225972 186654 225984
rect 224218 225972 224224 225984
rect 224276 225972 224282 226024
rect 233878 226012 233884 226024
rect 229066 225984 233884 226012
rect 94958 225836 94964 225888
rect 95016 225876 95022 225888
rect 166810 225876 166816 225888
rect 95016 225848 166816 225876
rect 95016 225836 95022 225848
rect 166810 225836 166816 225848
rect 166868 225836 166874 225888
rect 166948 225836 166954 225888
rect 167006 225876 167012 225888
rect 167006 225848 176148 225876
rect 167006 225836 167012 225848
rect 64782 225700 64788 225752
rect 64840 225740 64846 225752
rect 92474 225740 92480 225752
rect 64840 225712 92480 225740
rect 64840 225700 64846 225712
rect 92474 225700 92480 225712
rect 92532 225700 92538 225752
rect 108298 225700 108304 225752
rect 108356 225740 108362 225752
rect 171042 225740 171048 225752
rect 108356 225712 171048 225740
rect 108356 225700 108362 225712
rect 171042 225700 171048 225712
rect 171100 225700 171106 225752
rect 171226 225700 171232 225752
rect 171284 225740 171290 225752
rect 175918 225740 175924 225752
rect 171284 225712 175924 225740
rect 171284 225700 171290 225712
rect 175918 225700 175924 225712
rect 175976 225700 175982 225752
rect 176120 225740 176148 225848
rect 176286 225836 176292 225888
rect 176344 225876 176350 225888
rect 176608 225876 176614 225888
rect 176344 225848 176614 225876
rect 176344 225836 176350 225848
rect 176608 225836 176614 225848
rect 176666 225836 176672 225888
rect 176746 225836 176752 225888
rect 176804 225876 176810 225888
rect 181070 225876 181076 225888
rect 176804 225848 181076 225876
rect 176804 225836 176810 225848
rect 181070 225836 181076 225848
rect 181128 225836 181134 225888
rect 181622 225876 181628 225888
rect 181272 225848 181628 225876
rect 181272 225740 181300 225848
rect 181622 225836 181628 225848
rect 181680 225836 181686 225888
rect 183278 225836 183284 225888
rect 183336 225876 183342 225888
rect 186130 225876 186136 225888
rect 183336 225848 186136 225876
rect 183336 225836 183342 225848
rect 186130 225836 186136 225848
rect 186188 225836 186194 225888
rect 186268 225836 186274 225888
rect 186326 225876 186332 225888
rect 229066 225876 229094 225984
rect 233878 225972 233884 225984
rect 233936 225972 233942 226024
rect 243538 225972 243544 226024
rect 243596 226012 243602 226024
rect 248690 226012 248696 226024
rect 243596 225984 248696 226012
rect 243596 225972 243602 225984
rect 248690 225972 248696 225984
rect 248748 225972 248754 226024
rect 267550 225972 267556 226024
rect 267608 226012 267614 226024
rect 304074 226012 304080 226024
rect 267608 225984 304080 226012
rect 267608 225972 267614 225984
rect 304074 225972 304080 225984
rect 304132 225972 304138 226024
rect 313090 225972 313096 226024
rect 313148 226012 313154 226024
rect 340782 226012 340788 226024
rect 313148 225984 340788 226012
rect 313148 225972 313154 225984
rect 340782 225972 340788 225984
rect 340840 225972 340846 226024
rect 347866 226012 347872 226024
rect 344986 225984 347872 226012
rect 239030 225876 239036 225888
rect 186326 225848 229094 225876
rect 232700 225848 239036 225876
rect 186326 225836 186332 225848
rect 176120 225712 181300 225740
rect 181438 225700 181444 225752
rect 181496 225740 181502 225752
rect 184566 225740 184572 225752
rect 181496 225712 184572 225740
rect 181496 225700 181502 225712
rect 184566 225700 184572 225712
rect 184624 225700 184630 225752
rect 187050 225700 187056 225752
rect 187108 225740 187114 225752
rect 232700 225740 232728 225848
rect 239030 225836 239036 225848
rect 239088 225836 239094 225888
rect 249702 225836 249708 225888
rect 249760 225876 249766 225888
rect 290550 225876 290556 225888
rect 249760 225848 290556 225876
rect 249760 225836 249766 225848
rect 290550 225836 290556 225848
rect 290608 225836 290614 225888
rect 295242 225836 295248 225888
rect 295300 225876 295306 225888
rect 325970 225876 325976 225888
rect 295300 225848 325976 225876
rect 295300 225836 295306 225848
rect 325970 225836 325976 225848
rect 326028 225836 326034 225888
rect 340138 225836 340144 225888
rect 340196 225876 340202 225888
rect 344986 225876 345014 225984
rect 347866 225972 347872 225984
rect 347924 225972 347930 226024
rect 349062 225972 349068 226024
rect 349120 226012 349126 226024
rect 367186 226012 367192 226024
rect 349120 225984 367192 226012
rect 349120 225972 349126 225984
rect 367186 225972 367192 225984
rect 367244 225972 367250 226024
rect 501138 225972 501144 226024
rect 501196 226012 501202 226024
rect 501196 225984 503300 226012
rect 501196 225972 501202 225984
rect 340196 225848 345014 225876
rect 340196 225836 340202 225848
rect 347038 225836 347044 225888
rect 347096 225876 347102 225888
rect 365898 225876 365904 225888
rect 347096 225848 365904 225876
rect 347096 225836 347102 225848
rect 365898 225836 365904 225848
rect 365956 225836 365962 225888
rect 367738 225836 367744 225888
rect 367796 225876 367802 225888
rect 379606 225876 379612 225888
rect 367796 225848 379612 225876
rect 367796 225836 367802 225848
rect 379606 225836 379612 225848
rect 379664 225836 379670 225888
rect 488902 225836 488908 225888
rect 488960 225876 488966 225888
rect 502978 225876 502984 225888
rect 488960 225848 502984 225876
rect 488960 225836 488966 225848
rect 502978 225836 502984 225848
rect 503036 225836 503042 225888
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462590 225808 462596 225820
rect 458692 225780 462596 225808
rect 458692 225768 458698 225780
rect 462590 225768 462596 225780
rect 462648 225768 462654 225820
rect 242894 225740 242900 225752
rect 187108 225712 232728 225740
rect 232792 225712 242900 225740
rect 187108 225700 187114 225712
rect 61378 225564 61384 225616
rect 61436 225604 61442 225616
rect 136818 225604 136824 225616
rect 61436 225576 136824 225604
rect 61436 225564 61442 225576
rect 136818 225564 136824 225576
rect 136876 225564 136882 225616
rect 137002 225564 137008 225616
rect 137060 225604 137066 225616
rect 146938 225604 146944 225616
rect 137060 225576 146944 225604
rect 137060 225564 137066 225576
rect 146938 225564 146944 225576
rect 146996 225564 147002 225616
rect 147398 225564 147404 225616
rect 147456 225604 147462 225616
rect 204070 225604 204076 225616
rect 147456 225576 186268 225604
rect 147456 225564 147462 225576
rect 186240 225536 186268 225576
rect 186332 225576 204076 225604
rect 186332 225536 186360 225576
rect 204070 225564 204076 225576
rect 204128 225564 204134 225616
rect 204898 225564 204904 225616
rect 204956 225604 204962 225616
rect 222470 225604 222476 225616
rect 204956 225576 222476 225604
rect 204956 225564 204962 225576
rect 222470 225564 222476 225576
rect 222528 225564 222534 225616
rect 224218 225564 224224 225616
rect 224276 225604 224282 225616
rect 232792 225604 232820 225712
rect 242894 225700 242900 225712
rect 242952 225700 242958 225752
rect 257798 225700 257804 225752
rect 257856 225740 257862 225752
rect 299566 225740 299572 225752
rect 257856 225712 299572 225740
rect 257856 225700 257862 225712
rect 299566 225700 299572 225712
rect 299624 225700 299630 225752
rect 304902 225700 304908 225752
rect 304960 225740 304966 225752
rect 333698 225740 333704 225752
rect 304960 225712 333704 225740
rect 304960 225700 304966 225712
rect 333698 225700 333704 225712
rect 333756 225700 333762 225752
rect 335078 225700 335084 225752
rect 335136 225740 335142 225752
rect 356882 225740 356888 225752
rect 335136 225712 356888 225740
rect 335136 225700 335142 225712
rect 356882 225700 356888 225712
rect 356940 225700 356946 225752
rect 379330 225700 379336 225752
rect 379388 225740 379394 225752
rect 393590 225740 393596 225752
rect 379388 225712 393596 225740
rect 379388 225700 379394 225712
rect 393590 225700 393596 225712
rect 393648 225700 393654 225752
rect 394602 225700 394608 225752
rect 394660 225740 394666 225752
rect 404538 225740 404544 225752
rect 394660 225712 404544 225740
rect 394660 225700 394666 225712
rect 404538 225700 404544 225712
rect 404596 225700 404602 225752
rect 487614 225700 487620 225752
rect 487672 225740 487678 225752
rect 501506 225740 501512 225752
rect 487672 225712 501512 225740
rect 487672 225700 487678 225712
rect 501506 225700 501512 225712
rect 501564 225700 501570 225752
rect 503272 225740 503300 225984
rect 524322 225972 524328 226024
rect 524380 226012 524386 226024
rect 547874 226012 547880 226024
rect 524380 225984 547880 226012
rect 524380 225972 524386 225984
rect 547874 225972 547880 225984
rect 547932 225972 547938 226024
rect 508866 225836 508872 225888
rect 508924 225876 508930 225888
rect 528922 225876 528928 225888
rect 508924 225848 528928 225876
rect 508924 225836 508930 225848
rect 528922 225836 528928 225848
rect 528980 225836 528986 225888
rect 530118 225836 530124 225888
rect 530176 225876 530182 225888
rect 556154 225876 556160 225888
rect 530176 225848 556160 225876
rect 530176 225836 530182 225848
rect 556154 225836 556160 225848
rect 556212 225836 556218 225888
rect 671820 225752 671872 225758
rect 519354 225740 519360 225752
rect 503272 225712 519360 225740
rect 519354 225700 519360 225712
rect 519412 225700 519418 225752
rect 527542 225700 527548 225752
rect 527600 225740 527606 225752
rect 553302 225740 553308 225752
rect 527600 225712 553308 225740
rect 527600 225700 527606 225712
rect 553302 225700 553308 225712
rect 553360 225700 553366 225752
rect 556798 225700 556804 225752
rect 556856 225740 556862 225752
rect 570690 225740 570696 225752
rect 556856 225712 570696 225740
rect 556856 225700 556862 225712
rect 570690 225700 570696 225712
rect 570748 225700 570754 225752
rect 671820 225694 671872 225700
rect 671338 225632 671344 225684
rect 671396 225672 671402 225684
rect 671396 225644 671738 225672
rect 671396 225632 671402 225644
rect 224276 225576 232820 225604
rect 224276 225564 224282 225576
rect 234338 225564 234344 225616
rect 234396 225604 234402 225616
rect 281534 225604 281540 225616
rect 234396 225576 281540 225604
rect 234396 225564 234402 225576
rect 281534 225564 281540 225576
rect 281592 225564 281598 225616
rect 285490 225564 285496 225616
rect 285548 225604 285554 225616
rect 318886 225604 318892 225616
rect 285548 225576 318892 225604
rect 285548 225564 285554 225576
rect 318886 225564 318892 225576
rect 318944 225564 318950 225616
rect 322658 225564 322664 225616
rect 322716 225604 322722 225616
rect 349798 225604 349804 225616
rect 322716 225576 349804 225604
rect 322716 225564 322722 225576
rect 349798 225564 349804 225576
rect 349856 225564 349862 225616
rect 351178 225564 351184 225616
rect 351236 225604 351242 225616
rect 370406 225604 370412 225616
rect 351236 225576 370412 225604
rect 351236 225564 351242 225576
rect 370406 225564 370412 225576
rect 370464 225564 370470 225616
rect 372338 225564 372344 225616
rect 372396 225604 372402 225616
rect 388070 225604 388076 225616
rect 372396 225576 388076 225604
rect 372396 225564 372402 225576
rect 388070 225564 388076 225576
rect 388128 225564 388134 225616
rect 388438 225564 388444 225616
rect 388496 225604 388502 225616
rect 399386 225604 399392 225616
rect 388496 225576 399392 225604
rect 388496 225564 388502 225576
rect 399386 225564 399392 225576
rect 399444 225564 399450 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476666 225604 476672 225616
rect 467708 225576 476672 225604
rect 467708 225564 467714 225576
rect 476666 225564 476672 225576
rect 476724 225564 476730 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488534 225604 488540 225616
rect 477368 225576 488540 225604
rect 477368 225564 477374 225576
rect 488534 225564 488540 225576
rect 488592 225564 488598 225616
rect 494146 225564 494152 225616
rect 494204 225604 494210 225616
rect 509694 225604 509700 225616
rect 494204 225576 509700 225604
rect 494204 225564 494210 225576
rect 509694 225564 509700 225576
rect 509752 225564 509758 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530578 225604 530584 225616
rect 510212 225576 530584 225604
rect 510212 225564 510218 225576
rect 530578 225564 530584 225576
rect 530636 225564 530642 225616
rect 535914 225564 535920 225616
rect 535972 225604 535978 225616
rect 564710 225604 564716 225616
rect 535972 225576 564716 225604
rect 535972 225564 535978 225576
rect 564710 225564 564716 225576
rect 564768 225564 564774 225616
rect 186240 225508 186360 225536
rect 103238 225428 103244 225480
rect 103296 225468 103302 225480
rect 108298 225468 108304 225480
rect 103296 225440 108304 225468
rect 103296 225428 103302 225440
rect 108298 225428 108304 225440
rect 108356 225428 108362 225480
rect 127434 225468 127440 225480
rect 113146 225440 127440 225468
rect 105722 225292 105728 225344
rect 105780 225332 105786 225344
rect 113146 225332 113174 225440
rect 127434 225428 127440 225440
rect 127492 225428 127498 225480
rect 181438 225468 181444 225480
rect 127636 225440 181444 225468
rect 105780 225304 113174 225332
rect 105780 225292 105786 225304
rect 117222 225292 117228 225344
rect 117280 225332 117286 225344
rect 127636 225332 127664 225440
rect 181438 225428 181444 225440
rect 181496 225428 181502 225480
rect 181622 225428 181628 225480
rect 181680 225468 181686 225480
rect 185578 225468 185584 225480
rect 181680 225440 185584 225468
rect 181680 225428 181686 225440
rect 185578 225428 185584 225440
rect 185636 225428 185642 225480
rect 187694 225428 187700 225480
rect 187752 225468 187758 225480
rect 190546 225468 190552 225480
rect 187752 225440 190552 225468
rect 187752 225428 187758 225440
rect 190546 225428 190552 225440
rect 190604 225428 190610 225480
rect 190730 225428 190736 225480
rect 190788 225468 190794 225480
rect 242250 225468 242256 225480
rect 190788 225440 242256 225468
rect 190788 225428 190794 225440
rect 242250 225428 242256 225440
rect 242308 225428 242314 225480
rect 667014 225428 667020 225480
rect 667072 225468 667078 225480
rect 667072 225440 671622 225468
rect 667072 225428 667078 225440
rect 137002 225332 137008 225344
rect 117280 225304 127664 225332
rect 127728 225304 137008 225332
rect 117280 225292 117286 225304
rect 127434 225156 127440 225208
rect 127492 225196 127498 225208
rect 127728 225196 127756 225304
rect 137002 225292 137008 225304
rect 137060 225292 137066 225344
rect 142108 225332 142114 225344
rect 137204 225304 142114 225332
rect 127492 225168 127756 225196
rect 127492 225156 127498 225168
rect 128078 225156 128084 225208
rect 128136 225196 128142 225208
rect 137204 225196 137232 225304
rect 142108 225292 142114 225304
rect 142166 225292 142172 225344
rect 142246 225292 142252 225344
rect 142304 225332 142310 225344
rect 202966 225332 202972 225344
rect 142304 225304 202972 225332
rect 142304 225292 142310 225304
rect 202966 225292 202972 225304
rect 203024 225292 203030 225344
rect 204070 225292 204076 225344
rect 204128 225332 204134 225344
rect 207750 225332 207756 225344
rect 204128 225304 207756 225332
rect 204128 225292 204134 225304
rect 207750 225292 207756 225304
rect 207808 225292 207814 225344
rect 208118 225292 208124 225344
rect 208176 225332 208182 225344
rect 260926 225332 260932 225344
rect 208176 225304 260932 225332
rect 208176 225292 208182 225304
rect 260926 225292 260932 225304
rect 260984 225292 260990 225344
rect 463142 225224 463148 225276
rect 463200 225264 463206 225276
rect 467098 225264 467104 225276
rect 463200 225236 467104 225264
rect 463200 225224 463206 225236
rect 467098 225224 467104 225236
rect 467156 225224 467162 225276
rect 670510 225224 670516 225276
rect 670568 225264 670574 225276
rect 670568 225236 671508 225264
rect 670568 225224 670574 225236
rect 187694 225196 187700 225208
rect 128136 225168 137232 225196
rect 137296 225168 187700 225196
rect 128136 225156 128142 225168
rect 126882 225020 126888 225072
rect 126940 225060 126946 225072
rect 137296 225060 137324 225168
rect 187694 225156 187700 225168
rect 187752 225156 187758 225208
rect 188062 225156 188068 225208
rect 188120 225196 188126 225208
rect 195882 225196 195888 225208
rect 188120 225168 195888 225196
rect 188120 225156 188126 225168
rect 195882 225156 195888 225168
rect 195940 225156 195946 225208
rect 199378 225156 199384 225208
rect 199436 225196 199442 225208
rect 204898 225196 204904 225208
rect 199436 225168 204904 225196
rect 199436 225156 199442 225168
rect 204898 225156 204904 225168
rect 204956 225156 204962 225208
rect 205082 225156 205088 225208
rect 205140 225196 205146 225208
rect 254486 225196 254492 225208
rect 205140 225168 254492 225196
rect 205140 225156 205146 225168
rect 254486 225156 254492 225168
rect 254544 225156 254550 225208
rect 126940 225032 137324 225060
rect 126940 225020 126946 225032
rect 137462 225020 137468 225072
rect 137520 225060 137526 225072
rect 141510 225060 141516 225072
rect 137520 225032 141516 225060
rect 137520 225020 137526 225032
rect 141510 225020 141516 225032
rect 141568 225020 141574 225072
rect 141878 225020 141884 225072
rect 141936 225060 141942 225072
rect 141936 225032 142292 225060
rect 141936 225020 141942 225032
rect 116854 224884 116860 224936
rect 116912 224924 116918 224936
rect 122926 224924 122932 224936
rect 116912 224896 122932 224924
rect 116912 224884 116918 224896
rect 122926 224884 122932 224896
rect 122984 224884 122990 224936
rect 126514 224884 126520 224936
rect 126572 224924 126578 224936
rect 142062 224924 142068 224936
rect 126572 224896 142068 224924
rect 126572 224884 126578 224896
rect 142062 224884 142068 224896
rect 142120 224884 142126 224936
rect 142264 224924 142292 225032
rect 142430 225020 142436 225072
rect 142488 225060 142494 225072
rect 162302 225060 162308 225072
rect 142488 225032 162308 225060
rect 142488 225020 142494 225032
rect 162302 225020 162308 225032
rect 162360 225020 162366 225072
rect 162762 225020 162768 225072
rect 162820 225060 162826 225072
rect 166534 225060 166540 225072
rect 162820 225032 166540 225060
rect 162820 225020 162826 225032
rect 166534 225020 166540 225032
rect 166592 225020 166598 225072
rect 166718 225020 166724 225072
rect 166776 225060 166782 225072
rect 169018 225060 169024 225072
rect 166776 225032 169024 225060
rect 166776 225020 166782 225032
rect 169018 225020 169024 225032
rect 169076 225020 169082 225072
rect 169202 225020 169208 225072
rect 169260 225060 169266 225072
rect 170858 225060 170864 225072
rect 169260 225032 170864 225060
rect 169260 225020 169266 225032
rect 170858 225020 170864 225032
rect 170916 225020 170922 225072
rect 171042 225020 171048 225072
rect 171100 225060 171106 225072
rect 223574 225060 223580 225072
rect 171100 225032 223580 225060
rect 171100 225020 171106 225032
rect 223574 225020 223580 225032
rect 223632 225020 223638 225072
rect 224678 225020 224684 225072
rect 224736 225060 224742 225072
rect 270586 225060 270592 225072
rect 224736 225032 270592 225060
rect 224736 225020 224742 225032
rect 270586 225020 270592 225032
rect 270644 225020 270650 225072
rect 671246 225020 671252 225072
rect 671304 225060 671310 225072
rect 671304 225032 671398 225060
rect 671304 225020 671310 225032
rect 275646 224952 275652 225004
rect 275704 224992 275710 225004
rect 276842 224992 276848 225004
rect 275704 224964 276848 224992
rect 275704 224952 275710 224964
rect 276842 224952 276848 224964
rect 276900 224952 276906 225004
rect 282822 224952 282828 225004
rect 282880 224992 282886 225004
rect 285306 224992 285312 225004
rect 282880 224964 285312 224992
rect 282880 224952 282886 224964
rect 285306 224952 285312 224964
rect 285364 224952 285370 225004
rect 209406 224924 209412 224936
rect 142264 224896 209412 224924
rect 209406 224884 209412 224896
rect 209464 224884 209470 224936
rect 209682 224884 209688 224936
rect 209740 224924 209746 224936
rect 259638 224924 259644 224936
rect 209740 224896 259644 224924
rect 209740 224884 209746 224896
rect 259638 224884 259644 224896
rect 259696 224884 259702 224936
rect 264238 224884 264244 224936
rect 264296 224924 264302 224936
rect 269298 224924 269304 224936
rect 264296 224896 269304 224924
rect 264296 224884 264302 224896
rect 269298 224884 269304 224896
rect 269356 224884 269362 224936
rect 288250 224884 288256 224936
rect 288308 224924 288314 224936
rect 322382 224924 322388 224936
rect 288308 224896 322388 224924
rect 288308 224884 288314 224896
rect 322382 224884 322388 224896
rect 322440 224884 322446 224936
rect 407022 224884 407028 224936
rect 407080 224924 407086 224936
rect 414842 224924 414848 224936
rect 407080 224896 414848 224924
rect 407080 224884 407086 224896
rect 414842 224884 414848 224896
rect 414900 224884 414906 224936
rect 426434 224884 426440 224936
rect 426492 224924 426498 224936
rect 426986 224924 426992 224936
rect 426492 224896 426992 224924
rect 426492 224884 426498 224896
rect 426986 224884 426992 224896
rect 427044 224884 427050 224936
rect 118602 224748 118608 224800
rect 118660 224788 118666 224800
rect 181254 224788 181260 224800
rect 118660 224760 181260 224788
rect 118660 224748 118666 224760
rect 181254 224748 181260 224760
rect 181312 224748 181318 224800
rect 187050 224788 187056 224800
rect 181502 224760 187056 224788
rect 115658 224612 115664 224664
rect 115716 224652 115722 224664
rect 181502 224652 181530 224760
rect 187050 224748 187056 224760
rect 187108 224748 187114 224800
rect 187510 224748 187516 224800
rect 187568 224788 187574 224800
rect 190730 224788 190736 224800
rect 187568 224760 190736 224788
rect 187568 224748 187574 224760
rect 190730 224748 190736 224760
rect 190788 224748 190794 224800
rect 194318 224748 194324 224800
rect 194376 224788 194382 224800
rect 247402 224788 247408 224800
rect 194376 224760 247408 224788
rect 194376 224748 194382 224760
rect 247402 224748 247408 224760
rect 247460 224748 247466 224800
rect 282638 224748 282644 224800
rect 282696 224788 282702 224800
rect 316310 224788 316316 224800
rect 282696 224760 316316 224788
rect 282696 224748 282702 224760
rect 316310 224748 316316 224760
rect 316368 224748 316374 224800
rect 515766 224748 515772 224800
rect 515824 224788 515830 224800
rect 525242 224788 525248 224800
rect 515824 224760 525248 224788
rect 515824 224748 515830 224760
rect 525242 224748 525248 224760
rect 525300 224748 525306 224800
rect 526070 224748 526076 224800
rect 526128 224788 526134 224800
rect 537110 224788 537116 224800
rect 526128 224760 537116 224788
rect 526128 224748 526134 224760
rect 537110 224748 537116 224760
rect 537168 224748 537174 224800
rect 671252 224732 671304 224738
rect 460566 224680 460572 224732
rect 460624 224720 460630 224732
rect 462958 224720 462964 224732
rect 460624 224692 462964 224720
rect 460624 224680 460630 224692
rect 462958 224680 462964 224692
rect 463016 224680 463022 224732
rect 671252 224674 671304 224680
rect 115716 224624 181530 224652
rect 115716 224612 115722 224624
rect 181806 224612 181812 224664
rect 181864 224652 181870 224664
rect 191374 224652 191380 224664
rect 181864 224624 191380 224652
rect 181864 224612 181870 224624
rect 191374 224612 191380 224624
rect 191432 224612 191438 224664
rect 192478 224612 192484 224664
rect 192536 224652 192542 224664
rect 194502 224652 194508 224664
rect 192536 224624 194508 224652
rect 192536 224612 192542 224624
rect 194502 224612 194508 224624
rect 194560 224612 194566 224664
rect 195698 224612 195704 224664
rect 195756 224652 195762 224664
rect 248874 224652 248880 224664
rect 195756 224624 248880 224652
rect 195756 224612 195762 224624
rect 248874 224612 248880 224624
rect 248932 224612 248938 224664
rect 249058 224612 249064 224664
rect 249116 224652 249122 224664
rect 263870 224652 263876 224664
rect 249116 224624 263876 224652
rect 249116 224612 249122 224624
rect 263870 224612 263876 224624
rect 263928 224612 263934 224664
rect 271322 224612 271328 224664
rect 271380 224652 271386 224664
rect 309870 224652 309876 224664
rect 271380 224624 309876 224652
rect 271380 224612 271386 224624
rect 309870 224612 309876 224624
rect 309928 224612 309934 224664
rect 315850 224612 315856 224664
rect 315908 224652 315914 224664
rect 341426 224652 341432 224664
rect 315908 224624 341432 224652
rect 315908 224612 315914 224624
rect 341426 224612 341432 224624
rect 341484 224612 341490 224664
rect 344922 224612 344928 224664
rect 344980 224652 344986 224664
rect 364610 224652 364616 224664
rect 344980 224624 364616 224652
rect 344980 224612 344986 224624
rect 364610 224612 364616 224624
rect 364668 224612 364674 224664
rect 486602 224612 486608 224664
rect 486660 224652 486666 224664
rect 500402 224652 500408 224664
rect 486660 224624 500408 224652
rect 486660 224612 486666 224624
rect 500402 224612 500408 224624
rect 500460 224612 500466 224664
rect 508222 224612 508228 224664
rect 508280 224652 508286 224664
rect 528002 224652 528008 224664
rect 508280 224624 528008 224652
rect 508280 224612 508286 224624
rect 528002 224612 528008 224624
rect 528060 224612 528066 224664
rect 670510 224612 670516 224664
rect 670568 224652 670574 224664
rect 670568 224624 671186 224652
rect 670568 224612 670574 224624
rect 60642 224476 60648 224528
rect 60700 224516 60706 224528
rect 103606 224516 103612 224528
rect 60700 224488 103612 224516
rect 60700 224476 60706 224488
rect 103606 224476 103612 224488
rect 103664 224476 103670 224528
rect 108942 224476 108948 224528
rect 109000 224516 109006 224528
rect 183646 224516 183652 224528
rect 109000 224488 183652 224516
rect 109000 224476 109006 224488
rect 183646 224476 183652 224488
rect 183704 224476 183710 224528
rect 184014 224476 184020 224528
rect 184072 224516 184078 224528
rect 233694 224516 233700 224528
rect 184072 224488 233700 224516
rect 184072 224476 184078 224488
rect 233694 224476 233700 224488
rect 233752 224476 233758 224528
rect 233878 224476 233884 224528
rect 233936 224516 233942 224528
rect 246758 224516 246764 224528
rect 233936 224488 246764 224516
rect 233936 224476 233942 224488
rect 246758 224476 246764 224488
rect 246816 224476 246822 224528
rect 247678 224476 247684 224528
rect 247736 224516 247742 224528
rect 289262 224516 289268 224528
rect 247736 224488 289268 224516
rect 247736 224476 247742 224488
rect 289262 224476 289268 224488
rect 289320 224476 289326 224528
rect 319990 224476 319996 224528
rect 320048 224516 320054 224528
rect 347222 224516 347228 224528
rect 320048 224488 347228 224516
rect 320048 224476 320054 224488
rect 347222 224476 347228 224488
rect 347280 224476 347286 224528
rect 491478 224476 491484 224528
rect 491536 224516 491542 224528
rect 506474 224516 506480 224528
rect 491536 224488 506480 224516
rect 491536 224476 491542 224488
rect 506474 224476 506480 224488
rect 506532 224476 506538 224528
rect 510798 224476 510804 224528
rect 510856 224516 510862 224528
rect 531774 224516 531780 224528
rect 510856 224488 531780 224516
rect 510856 224476 510862 224488
rect 531774 224476 531780 224488
rect 531832 224476 531838 224528
rect 532050 224476 532056 224528
rect 532108 224516 532114 224528
rect 558914 224516 558920 224528
rect 532108 224488 558920 224516
rect 532108 224476 532114 224488
rect 558914 224476 558920 224488
rect 558972 224476 558978 224528
rect 670602 224408 670608 224460
rect 670660 224448 670666 224460
rect 670660 224420 671048 224448
rect 670660 224408 670666 224420
rect 82538 224340 82544 224392
rect 82596 224380 82602 224392
rect 126514 224380 126520 224392
rect 82596 224352 126520 224380
rect 82596 224340 82602 224352
rect 126514 224340 126520 224352
rect 126572 224340 126578 224392
rect 126698 224340 126704 224392
rect 126756 224380 126762 224392
rect 131114 224380 131120 224392
rect 126756 224352 131120 224380
rect 126756 224340 126762 224352
rect 131114 224340 131120 224352
rect 131172 224340 131178 224392
rect 131298 224340 131304 224392
rect 131356 224380 131362 224392
rect 193950 224380 193956 224392
rect 131356 224352 193956 224380
rect 131356 224340 131362 224352
rect 193950 224340 193956 224352
rect 194008 224340 194014 224392
rect 194134 224340 194140 224392
rect 194192 224380 194198 224392
rect 204898 224380 204904 224392
rect 194192 224352 204904 224380
rect 194192 224340 194198 224352
rect 204898 224340 204904 224352
rect 204956 224340 204962 224392
rect 205082 224340 205088 224392
rect 205140 224380 205146 224392
rect 255774 224380 255780 224392
rect 205140 224352 255780 224380
rect 205140 224340 205146 224352
rect 255774 224340 255780 224352
rect 255832 224340 255838 224392
rect 262122 224340 262128 224392
rect 262180 224380 262186 224392
rect 300854 224380 300860 224392
rect 262180 224352 300860 224380
rect 262180 224340 262186 224352
rect 300854 224340 300860 224352
rect 300912 224340 300918 224392
rect 303430 224340 303436 224392
rect 303488 224380 303494 224392
rect 333054 224380 333060 224392
rect 303488 224352 333060 224380
rect 303488 224340 303494 224352
rect 333054 224340 333060 224352
rect 333112 224340 333118 224392
rect 333882 224340 333888 224392
rect 333940 224380 333946 224392
rect 356238 224380 356244 224392
rect 333940 224352 356244 224380
rect 333940 224340 333946 224352
rect 356238 224340 356244 224352
rect 356296 224340 356302 224392
rect 357342 224340 357348 224392
rect 357400 224380 357406 224392
rect 374270 224380 374276 224392
rect 357400 224352 374276 224380
rect 357400 224340 357406 224352
rect 374270 224340 374276 224352
rect 374328 224340 374334 224392
rect 375282 224340 375288 224392
rect 375340 224380 375346 224392
rect 387794 224380 387800 224392
rect 375340 224352 387800 224380
rect 375340 224340 375346 224352
rect 387794 224340 387800 224352
rect 387852 224340 387858 224392
rect 456150 224340 456156 224392
rect 456208 224380 456214 224392
rect 459646 224380 459652 224392
rect 456208 224352 459652 224380
rect 456208 224340 456214 224352
rect 459646 224340 459652 224352
rect 459704 224340 459710 224392
rect 479058 224340 479064 224392
rect 479116 224380 479122 224392
rect 485774 224380 485780 224392
rect 479116 224352 485780 224380
rect 479116 224340 479122 224352
rect 485774 224340 485780 224352
rect 485832 224340 485838 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516410 224380 516416 224392
rect 499264 224352 516416 224380
rect 499264 224340 499270 224352
rect 516410 224340 516416 224352
rect 516468 224340 516474 224392
rect 525610 224340 525616 224392
rect 525668 224380 525674 224392
rect 550634 224380 550640 224392
rect 525668 224352 550640 224380
rect 525668 224340 525674 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 59262 224204 59268 224256
rect 59320 224244 59326 224256
rect 141602 224244 141608 224256
rect 59320 224216 141608 224244
rect 59320 224204 59326 224216
rect 141602 224204 141608 224216
rect 141660 224204 141666 224256
rect 142062 224204 142068 224256
rect 142120 224244 142126 224256
rect 157288 224244 157294 224256
rect 142120 224216 157294 224244
rect 142120 224204 142126 224216
rect 157288 224204 157294 224216
rect 157346 224204 157352 224256
rect 157426 224204 157432 224256
rect 157484 224244 157490 224256
rect 170950 224244 170956 224256
rect 157484 224216 170956 224244
rect 157484 224204 157490 224216
rect 170950 224204 170956 224216
rect 171008 224204 171014 224256
rect 171088 224204 171094 224256
rect 171146 224244 171152 224256
rect 186866 224244 186872 224256
rect 171146 224216 186872 224244
rect 171146 224204 171152 224216
rect 186866 224204 186872 224216
rect 186924 224204 186930 224256
rect 187050 224204 187056 224256
rect 187108 224244 187114 224256
rect 188798 224244 188804 224256
rect 187108 224216 188804 224244
rect 187108 224204 187114 224216
rect 188798 224204 188804 224216
rect 188856 224204 188862 224256
rect 188982 224204 188988 224256
rect 189040 224244 189046 224256
rect 243814 224244 243820 224256
rect 189040 224216 243820 224244
rect 189040 224204 189046 224216
rect 243814 224204 243820 224216
rect 243872 224204 243878 224256
rect 246942 224204 246948 224256
rect 247000 224244 247006 224256
rect 288618 224244 288624 224256
rect 247000 224216 288624 224244
rect 247000 224204 247006 224216
rect 288618 224204 288624 224216
rect 288676 224204 288682 224256
rect 289538 224204 289544 224256
rect 289596 224244 289602 224256
rect 307846 224244 307852 224256
rect 289596 224216 307852 224244
rect 289596 224204 289602 224216
rect 307846 224204 307852 224216
rect 307904 224204 307910 224256
rect 308950 224204 308956 224256
rect 309008 224244 309014 224256
rect 339494 224244 339500 224256
rect 309008 224216 339500 224244
rect 309008 224204 309014 224216
rect 339494 224204 339500 224216
rect 339552 224204 339558 224256
rect 341886 224204 341892 224256
rect 341944 224244 341950 224256
rect 364794 224244 364800 224256
rect 341944 224216 364800 224244
rect 341944 224204 341950 224216
rect 364794 224204 364800 224216
rect 364852 224204 364858 224256
rect 364978 224204 364984 224256
rect 365036 224244 365042 224256
rect 378134 224244 378140 224256
rect 365036 224216 378140 224244
rect 365036 224204 365042 224216
rect 378134 224204 378140 224216
rect 378192 224204 378198 224256
rect 388898 224204 388904 224256
rect 388956 224244 388962 224256
rect 400950 224244 400956 224256
rect 388956 224216 400956 224244
rect 388956 224204 388962 224216
rect 400950 224204 400956 224216
rect 401008 224204 401014 224256
rect 416406 224204 416412 224256
rect 416464 224244 416470 224256
rect 422202 224244 422208 224256
rect 416464 224216 422208 224244
rect 416464 224204 416470 224216
rect 422202 224204 422208 224216
rect 422260 224204 422266 224256
rect 451366 224204 451372 224256
rect 451424 224244 451430 224256
rect 452010 224244 452016 224256
rect 451424 224216 452016 224244
rect 451424 224204 451430 224216
rect 452010 224204 452016 224216
rect 452068 224204 452074 224256
rect 462406 224204 462412 224256
rect 462464 224244 462470 224256
rect 469674 224244 469680 224256
rect 462464 224216 469680 224244
rect 462464 224204 462470 224216
rect 469674 224204 469680 224216
rect 469732 224204 469738 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 479518 224244 479524 224256
rect 470284 224216 479524 224244
rect 470284 224204 470290 224216
rect 479518 224204 479524 224216
rect 479576 224204 479582 224256
rect 483750 224204 483756 224256
rect 483808 224244 483814 224256
rect 497274 224244 497280 224256
rect 483808 224216 497280 224244
rect 483808 224204 483814 224216
rect 497274 224204 497280 224216
rect 497332 224204 497338 224256
rect 513190 224204 513196 224256
rect 513248 224244 513254 224256
rect 534442 224244 534448 224256
rect 513248 224216 534448 224244
rect 513248 224204 513254 224216
rect 534442 224204 534448 224216
rect 534500 224204 534506 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 563974 224244 563980 224256
rect 535328 224216 563980 224244
rect 535328 224204 535334 224216
rect 563974 224204 563980 224216
rect 564032 224204 564038 224256
rect 423582 224136 423588 224188
rect 423640 224176 423646 224188
rect 424318 224176 424324 224188
rect 423640 224148 424324 224176
rect 423640 224136 423646 224148
rect 424318 224136 424324 224148
rect 424376 224136 424382 224188
rect 667014 224136 667020 224188
rect 667072 224176 667078 224188
rect 667072 224148 670956 224176
rect 667072 224136 667078 224148
rect 104802 224068 104808 224120
rect 104860 224108 104866 224120
rect 116854 224108 116860 224120
rect 104860 224080 116860 224108
rect 104860 224068 104866 224080
rect 116854 224068 116860 224080
rect 116912 224068 116918 224120
rect 117038 224068 117044 224120
rect 117096 224108 117102 224120
rect 118418 224108 118424 224120
rect 117096 224080 118424 224108
rect 117096 224068 117102 224080
rect 118418 224068 118424 224080
rect 118476 224068 118482 224120
rect 122282 224068 122288 224120
rect 122340 224108 122346 224120
rect 131298 224108 131304 224120
rect 122340 224080 131304 224108
rect 122340 224068 122346 224080
rect 131298 224068 131304 224080
rect 131356 224068 131362 224120
rect 131482 224068 131488 224120
rect 131540 224108 131546 224120
rect 192478 224108 192484 224120
rect 131540 224080 192484 224108
rect 131540 224068 131546 224080
rect 192478 224068 192484 224080
rect 192536 224068 192542 224120
rect 192662 224068 192668 224120
rect 192720 224108 192726 224120
rect 194134 224108 194140 224120
rect 192720 224080 194140 224108
rect 192720 224068 192726 224080
rect 194134 224068 194140 224080
rect 194192 224068 194198 224120
rect 194502 224068 194508 224120
rect 194560 224108 194566 224120
rect 196526 224108 196532 224120
rect 194560 224080 196532 224108
rect 194560 224068 194566 224080
rect 196526 224068 196532 224080
rect 196584 224068 196590 224120
rect 201218 224068 201224 224120
rect 201276 224108 201282 224120
rect 204714 224108 204720 224120
rect 201276 224080 204720 224108
rect 201276 224068 201282 224080
rect 204714 224068 204720 224080
rect 204772 224068 204778 224120
rect 204898 224068 204904 224120
rect 204956 224108 204962 224120
rect 233878 224108 233884 224120
rect 204956 224080 233884 224108
rect 204956 224068 204962 224080
rect 233878 224068 233884 224080
rect 233936 224068 233942 224120
rect 278958 224108 278964 224120
rect 234080 224080 278964 224108
rect 76466 223932 76472 223984
rect 76524 223972 76530 223984
rect 141418 223972 141424 223984
rect 76524 223944 141424 223972
rect 76524 223932 76530 223944
rect 141418 223932 141424 223944
rect 141476 223932 141482 223984
rect 141602 223932 141608 223984
rect 141660 223972 141666 223984
rect 145190 223972 145196 223984
rect 141660 223944 145196 223972
rect 141660 223932 141666 223944
rect 145190 223932 145196 223944
rect 145248 223932 145254 223984
rect 145374 223932 145380 223984
rect 145432 223972 145438 223984
rect 147214 223972 147220 223984
rect 145432 223944 147220 223972
rect 145432 223932 145438 223944
rect 147214 223932 147220 223944
rect 147272 223932 147278 223984
rect 147674 223932 147680 223984
rect 147732 223972 147738 223984
rect 154574 223972 154580 223984
rect 147732 223944 154580 223972
rect 147732 223932 147738 223944
rect 154574 223932 154580 223944
rect 154632 223932 154638 223984
rect 156874 223932 156880 223984
rect 156932 223972 156938 223984
rect 217042 223972 217048 223984
rect 156932 223944 217048 223972
rect 156932 223932 156938 223944
rect 217042 223932 217048 223944
rect 217100 223932 217106 223984
rect 217226 223932 217232 223984
rect 217284 223972 217290 223984
rect 228082 223972 228088 223984
rect 217284 223944 228088 223972
rect 217284 223932 217290 223944
rect 228082 223932 228088 223944
rect 228140 223932 228146 223984
rect 231578 223932 231584 223984
rect 231636 223972 231642 223984
rect 234080 223972 234108 224080
rect 278958 224068 278964 224080
rect 279016 224068 279022 224120
rect 286962 224068 286968 224120
rect 287020 224108 287026 224120
rect 319530 224108 319536 224120
rect 287020 224080 319536 224108
rect 287020 224068 287026 224080
rect 319530 224068 319536 224080
rect 319588 224068 319594 224120
rect 231636 223944 234108 223972
rect 231636 223932 231642 223944
rect 238662 223932 238668 223984
rect 238720 223972 238726 223984
rect 282454 223972 282460 223984
rect 238720 223944 282460 223972
rect 238720 223932 238726 223944
rect 282454 223932 282460 223944
rect 282512 223932 282518 223984
rect 125134 223796 125140 223848
rect 125192 223836 125198 223848
rect 131482 223836 131488 223848
rect 125192 223808 131488 223836
rect 125192 223796 125198 223808
rect 131482 223796 131488 223808
rect 131540 223796 131546 223848
rect 134978 223796 134984 223848
rect 135036 223836 135042 223848
rect 204254 223836 204260 223848
rect 135036 223808 204260 223836
rect 135036 223796 135042 223808
rect 204254 223796 204260 223808
rect 204312 223796 204318 223848
rect 205266 223796 205272 223848
rect 205324 223836 205330 223848
rect 212810 223836 212816 223848
rect 205324 223808 212816 223836
rect 205324 223796 205330 223808
rect 212810 223796 212816 223808
rect 212868 223796 212874 223848
rect 215938 223796 215944 223848
rect 215996 223836 216002 223848
rect 222930 223836 222936 223848
rect 215996 223808 222936 223836
rect 215996 223796 216002 223808
rect 222930 223796 222936 223808
rect 222988 223796 222994 223848
rect 233694 223796 233700 223848
rect 233752 223836 233758 223848
rect 239674 223836 239680 223848
rect 233752 223808 239680 223836
rect 233752 223796 233758 223808
rect 239674 223796 239680 223808
rect 239732 223796 239738 223848
rect 242710 223796 242716 223848
rect 242768 223836 242774 223848
rect 285030 223836 285036 223848
rect 242768 223808 285036 223836
rect 242768 223796 242774 223808
rect 285030 223796 285036 223808
rect 285088 223796 285094 223848
rect 132218 223660 132224 223712
rect 132276 223700 132282 223712
rect 201678 223700 201684 223712
rect 132276 223672 201684 223700
rect 132276 223660 132282 223672
rect 201678 223660 201684 223672
rect 201736 223660 201742 223712
rect 297652 223672 300348 223700
rect 88058 223524 88064 223576
rect 88116 223564 88122 223576
rect 164970 223564 164976 223576
rect 88116 223536 164976 223564
rect 88116 223524 88122 223536
rect 164970 223524 164976 223536
rect 165028 223524 165034 223576
rect 166258 223524 166264 223576
rect 166316 223564 166322 223576
rect 168098 223564 168104 223576
rect 166316 223536 168104 223564
rect 166316 223524 166322 223536
rect 168098 223524 168104 223536
rect 168156 223524 168162 223576
rect 168282 223524 168288 223576
rect 168340 223564 168346 223576
rect 226794 223564 226800 223576
rect 168340 223536 226800 223564
rect 168340 223524 168346 223536
rect 226794 223524 226800 223536
rect 226852 223524 226858 223576
rect 268838 223524 268844 223576
rect 268896 223564 268902 223576
rect 297652 223564 297680 223672
rect 268896 223536 297680 223564
rect 268896 223524 268902 223536
rect 297818 223524 297824 223576
rect 297876 223564 297882 223576
rect 300118 223564 300124 223576
rect 297876 223536 300124 223564
rect 297876 223524 297882 223536
rect 300118 223524 300124 223536
rect 300176 223524 300182 223576
rect 300320 223564 300348 223672
rect 563698 223592 563704 223644
rect 563756 223632 563762 223644
rect 571242 223632 571248 223644
rect 563756 223604 571248 223632
rect 563756 223592 563762 223604
rect 571242 223592 571248 223604
rect 571300 223592 571306 223644
rect 306006 223564 306012 223576
rect 300320 223536 306012 223564
rect 306006 223524 306012 223536
rect 306064 223524 306070 223576
rect 329006 223524 329012 223576
rect 329064 223564 329070 223576
rect 342714 223564 342720 223576
rect 329064 223536 342720 223564
rect 329064 223524 329070 223536
rect 342714 223524 342720 223536
rect 342772 223524 342778 223576
rect 457990 223524 457996 223576
rect 458048 223564 458054 223576
rect 460198 223564 460204 223576
rect 458048 223536 460204 223564
rect 458048 223524 458054 223536
rect 460198 223524 460204 223536
rect 460256 223524 460262 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475746 223564 475752 223576
rect 473504 223536 475752 223564
rect 473504 223524 473510 223536
rect 475746 223524 475752 223536
rect 475804 223524 475810 223576
rect 499574 223524 499580 223576
rect 499632 223564 499638 223576
rect 503162 223564 503168 223576
rect 499632 223536 503168 223564
rect 499632 223524 499638 223536
rect 503162 223524 503168 223536
rect 503220 223524 503226 223576
rect 81342 223388 81348 223440
rect 81400 223428 81406 223440
rect 157242 223428 157248 223440
rect 81400 223400 157248 223428
rect 81400 223388 81406 223400
rect 157242 223388 157248 223400
rect 157300 223388 157306 223440
rect 157426 223388 157432 223440
rect 157484 223428 157490 223440
rect 159818 223428 159824 223440
rect 157484 223400 159824 223428
rect 157484 223388 157490 223400
rect 159818 223388 159824 223400
rect 159876 223388 159882 223440
rect 161106 223388 161112 223440
rect 161164 223428 161170 223440
rect 162302 223428 162308 223440
rect 161164 223400 162308 223428
rect 161164 223388 161170 223400
rect 162302 223388 162308 223400
rect 162360 223388 162366 223440
rect 164142 223388 164148 223440
rect 164200 223428 164206 223440
rect 224034 223428 224040 223440
rect 164200 223400 224040 223428
rect 164200 223388 164206 223400
rect 224034 223388 224040 223400
rect 224092 223388 224098 223440
rect 260558 223388 260564 223440
rect 260616 223428 260622 223440
rect 298922 223428 298928 223440
rect 260616 223400 298928 223428
rect 260616 223388 260622 223400
rect 298922 223388 298928 223400
rect 298980 223388 298986 223440
rect 301958 223388 301964 223440
rect 302016 223428 302022 223440
rect 331122 223428 331128 223440
rect 302016 223400 331128 223428
rect 302016 223388 302022 223400
rect 331122 223388 331128 223400
rect 331180 223388 331186 223440
rect 516778 223388 516784 223440
rect 516836 223428 516842 223440
rect 532142 223428 532148 223440
rect 516836 223400 532148 223428
rect 516836 223388 516842 223400
rect 532142 223388 532148 223400
rect 532200 223388 532206 223440
rect 543918 223388 543924 223440
rect 543976 223428 543982 223440
rect 554866 223428 554872 223440
rect 543976 223400 554872 223428
rect 543976 223388 543982 223400
rect 554866 223388 554872 223400
rect 554924 223388 554930 223440
rect 96706 223252 96712 223304
rect 96764 223292 96770 223304
rect 117958 223292 117964 223304
rect 96764 223264 117964 223292
rect 96764 223252 96770 223264
rect 117958 223252 117964 223264
rect 118016 223252 118022 223304
rect 118142 223252 118148 223304
rect 118200 223292 118206 223304
rect 166258 223292 166264 223304
rect 118200 223264 166264 223292
rect 118200 223252 118206 223264
rect 166258 223252 166264 223264
rect 166316 223252 166322 223304
rect 168098 223252 168104 223304
rect 168156 223292 168162 223304
rect 185762 223292 185768 223304
rect 168156 223264 185768 223292
rect 168156 223252 168162 223264
rect 185762 223252 185768 223264
rect 185820 223252 185826 223304
rect 186038 223252 186044 223304
rect 186096 223292 186102 223304
rect 192202 223292 192208 223304
rect 186096 223264 192208 223292
rect 186096 223252 186102 223264
rect 192202 223252 192208 223264
rect 192260 223252 192266 223304
rect 192478 223252 192484 223304
rect 192536 223292 192542 223304
rect 196066 223292 196072 223304
rect 192536 223264 196072 223292
rect 192536 223252 192542 223264
rect 196066 223252 196072 223264
rect 196124 223252 196130 223304
rect 204070 223252 204076 223304
rect 204128 223292 204134 223304
rect 254854 223292 254860 223304
rect 204128 223264 254860 223292
rect 204128 223252 204134 223264
rect 254854 223252 254860 223264
rect 254912 223252 254918 223304
rect 264698 223252 264704 223304
rect 264756 223292 264762 223304
rect 304718 223292 304724 223304
rect 264756 223264 304724 223292
rect 264756 223252 264762 223264
rect 304718 223252 304724 223264
rect 304776 223252 304782 223304
rect 306098 223252 306104 223304
rect 306156 223292 306162 223304
rect 336918 223292 336924 223304
rect 306156 223264 336924 223292
rect 306156 223252 306162 223264
rect 336918 223252 336924 223264
rect 336976 223252 336982 223304
rect 343358 223252 343364 223304
rect 343416 223292 343422 223304
rect 363966 223292 363972 223304
rect 343416 223264 363972 223292
rect 343416 223252 343422 223264
rect 363966 223252 363972 223264
rect 364024 223252 364030 223304
rect 506934 223252 506940 223304
rect 506992 223292 506998 223304
rect 526346 223292 526352 223304
rect 506992 223264 526352 223292
rect 506992 223252 506998 223264
rect 526346 223252 526352 223264
rect 526404 223252 526410 223304
rect 530302 223252 530308 223304
rect 530360 223292 530366 223304
rect 544930 223292 544936 223304
rect 530360 223264 544936 223292
rect 530360 223252 530366 223264
rect 544930 223252 544936 223264
rect 544988 223252 544994 223304
rect 78398 223116 78404 223168
rect 78456 223156 78462 223168
rect 152274 223156 152280 223168
rect 78456 223128 152280 223156
rect 78456 223116 78462 223128
rect 152274 223116 152280 223128
rect 152332 223116 152338 223168
rect 152458 223116 152464 223168
rect 152516 223156 152522 223168
rect 166258 223156 166264 223168
rect 152516 223128 166264 223156
rect 152516 223116 152522 223128
rect 166258 223116 166264 223128
rect 166316 223116 166322 223168
rect 166442 223116 166448 223168
rect 166500 223156 166506 223168
rect 222286 223156 222292 223168
rect 166500 223128 222292 223156
rect 166500 223116 166506 223128
rect 222286 223116 222292 223128
rect 222344 223116 222350 223168
rect 224218 223116 224224 223168
rect 224276 223156 224282 223168
rect 238386 223156 238392 223168
rect 224276 223128 238392 223156
rect 224276 223116 224282 223128
rect 238386 223116 238392 223128
rect 238444 223116 238450 223168
rect 245562 223116 245568 223168
rect 245620 223156 245626 223168
rect 287606 223156 287612 223168
rect 245620 223128 287612 223156
rect 245620 223116 245626 223128
rect 287606 223116 287612 223128
rect 287664 223116 287670 223168
rect 291102 223116 291108 223168
rect 291160 223156 291166 223168
rect 323670 223156 323676 223168
rect 291160 223128 323676 223156
rect 291160 223116 291166 223128
rect 323670 223116 323676 223128
rect 323728 223116 323734 223168
rect 330478 223116 330484 223168
rect 330536 223156 330542 223168
rect 354950 223156 354956 223168
rect 330536 223128 354956 223156
rect 330536 223116 330542 223128
rect 354950 223116 354956 223128
rect 355008 223116 355014 223168
rect 357158 223116 357164 223168
rect 357216 223156 357222 223168
rect 376202 223156 376208 223168
rect 357216 223128 376208 223156
rect 357216 223116 357222 223128
rect 376202 223116 376208 223128
rect 376260 223116 376266 223168
rect 522666 223116 522672 223168
rect 522724 223156 522730 223168
rect 546770 223156 546776 223168
rect 522724 223128 546776 223156
rect 522724 223116 522730 223128
rect 546770 223116 546776 223128
rect 546828 223116 546834 223168
rect 92382 222980 92388 223032
rect 92440 223020 92446 223032
rect 96706 223020 96712 223032
rect 92440 222992 96712 223020
rect 92440 222980 92446 222992
rect 96706 222980 96712 222992
rect 96764 222980 96770 223032
rect 98638 222980 98644 223032
rect 98696 223020 98702 223032
rect 166074 223020 166080 223032
rect 98696 222992 166080 223020
rect 98696 222980 98702 222992
rect 166074 222980 166080 222992
rect 166132 222980 166138 223032
rect 166810 222980 166816 223032
rect 166868 223020 166874 223032
rect 181622 223020 181628 223032
rect 166868 222992 181628 223020
rect 166868 222980 166874 222992
rect 181622 222980 181628 222992
rect 181680 222980 181686 223032
rect 181806 222980 181812 223032
rect 181864 223020 181870 223032
rect 234798 223020 234804 223032
rect 181864 222992 234804 223020
rect 181864 222980 181870 222992
rect 234798 222980 234804 222992
rect 234856 222980 234862 223032
rect 235258 222980 235264 223032
rect 235316 223020 235322 223032
rect 243262 223020 243268 223032
rect 235316 222992 243268 223020
rect 235316 222980 235322 222992
rect 243262 222980 243268 222992
rect 243320 222980 243326 223032
rect 250898 222980 250904 223032
rect 250956 223020 250962 223032
rect 294414 223020 294420 223032
rect 250956 222992 294420 223020
rect 250956 222980 250962 222992
rect 294414 222980 294420 222992
rect 294472 222980 294478 223032
rect 300302 222980 300308 223032
rect 300360 223020 300366 223032
rect 331306 223020 331312 223032
rect 300360 222992 331312 223020
rect 300360 222980 300366 222992
rect 331306 222980 331312 222992
rect 331364 222980 331370 223032
rect 337930 222980 337936 223032
rect 337988 223020 337994 223032
rect 359182 223020 359188 223032
rect 337988 222992 359188 223020
rect 337988 222980 337994 222992
rect 359182 222980 359188 222992
rect 359240 222980 359246 223032
rect 370498 222980 370504 223032
rect 370556 223020 370562 223032
rect 384574 223020 384580 223032
rect 370556 222992 384580 223020
rect 370556 222980 370562 222992
rect 384574 222980 384580 222992
rect 384632 222980 384638 223032
rect 387702 222980 387708 223032
rect 387760 223020 387766 223032
rect 398098 223020 398104 223032
rect 387760 222992 398104 223020
rect 387760 222980 387766 222992
rect 398098 222980 398104 222992
rect 398156 222980 398162 223032
rect 478322 222980 478328 223032
rect 478380 223020 478386 223032
rect 485038 223020 485044 223032
rect 478380 222992 485044 223020
rect 478380 222980 478386 222992
rect 485038 222980 485044 222992
rect 485096 222980 485102 223032
rect 485590 222980 485596 223032
rect 485648 223020 485654 223032
rect 498194 223020 498200 223032
rect 485648 222992 498200 223020
rect 485648 222980 485654 222992
rect 498194 222980 498200 222992
rect 498252 222980 498258 223032
rect 503346 222980 503352 223032
rect 503404 223020 503410 223032
rect 521930 223020 521936 223032
rect 503404 222992 521936 223020
rect 503404 222980 503410 222992
rect 521930 222980 521936 222992
rect 521988 222980 521994 223032
rect 523678 222980 523684 223032
rect 523736 223020 523742 223032
rect 548150 223020 548156 223032
rect 523736 222992 548156 223020
rect 523736 222980 523742 222992
rect 548150 222980 548156 222992
rect 548208 222980 548214 223032
rect 570322 222980 570328 223032
rect 570380 223020 570386 223032
rect 575382 223020 575388 223032
rect 570380 222992 575388 223020
rect 570380 222980 570386 222992
rect 575382 222980 575388 222992
rect 575440 222980 575446 223032
rect 56502 222844 56508 222896
rect 56560 222884 56566 222896
rect 137094 222884 137100 222896
rect 56560 222856 137100 222884
rect 56560 222844 56566 222856
rect 137094 222844 137100 222856
rect 137152 222844 137158 222896
rect 137278 222844 137284 222896
rect 137336 222884 137342 222896
rect 152458 222884 152464 222896
rect 137336 222856 152464 222884
rect 137336 222844 137342 222856
rect 152458 222844 152464 222856
rect 152516 222844 152522 222896
rect 154482 222844 154488 222896
rect 154540 222884 154546 222896
rect 212166 222884 212172 222896
rect 154540 222856 166396 222884
rect 154540 222844 154546 222856
rect 166368 222816 166396 222856
rect 166736 222856 212172 222884
rect 166736 222816 166764 222856
rect 212166 222844 212172 222856
rect 212224 222844 212230 222896
rect 221642 222884 221648 222896
rect 212368 222856 221648 222884
rect 166368 222788 166764 222816
rect 85482 222708 85488 222760
rect 85540 222748 85546 222760
rect 162118 222748 162124 222760
rect 85540 222720 162124 222748
rect 85540 222708 85546 222720
rect 162118 222708 162124 222720
rect 162176 222708 162182 222760
rect 162302 222708 162308 222760
rect 162360 222748 162366 222760
rect 162360 222720 166304 222748
rect 162360 222708 162366 222720
rect 166276 222680 166304 222720
rect 168098 222708 168104 222760
rect 168156 222748 168162 222760
rect 168156 222720 181484 222748
rect 168156 222708 168162 222720
rect 166810 222680 166816 222692
rect 166276 222652 166816 222680
rect 166810 222640 166816 222652
rect 166868 222640 166874 222692
rect 89162 222572 89168 222624
rect 89220 222612 89226 222624
rect 98638 222612 98644 222624
rect 89220 222584 98644 222612
rect 89220 222572 89226 222584
rect 98638 222572 98644 222584
rect 98696 222572 98702 222624
rect 99098 222572 99104 222624
rect 99156 222612 99162 222624
rect 166074 222612 166080 222624
rect 99156 222584 166080 222612
rect 99156 222572 99162 222584
rect 166074 222572 166080 222584
rect 166132 222572 166138 222624
rect 166994 222572 167000 222624
rect 167052 222612 167058 222624
rect 174814 222612 174820 222624
rect 167052 222584 174820 222612
rect 167052 222572 167058 222584
rect 174814 222572 174820 222584
rect 174872 222572 174878 222624
rect 174998 222572 175004 222624
rect 175056 222612 175062 222624
rect 181254 222612 181260 222624
rect 175056 222584 181260 222612
rect 175056 222572 175062 222584
rect 181254 222572 181260 222584
rect 181312 222572 181318 222624
rect 181456 222612 181484 222720
rect 181622 222708 181628 222760
rect 181680 222748 181686 222760
rect 181680 222720 195468 222748
rect 181680 222708 181686 222720
rect 195440 222680 195468 222720
rect 196066 222708 196072 222760
rect 196124 222748 196130 222760
rect 203702 222748 203708 222760
rect 196124 222720 203708 222748
rect 196124 222708 196130 222720
rect 203702 222708 203708 222720
rect 203760 222708 203766 222760
rect 212368 222748 212396 222856
rect 221642 222844 221648 222856
rect 221700 222844 221706 222896
rect 233142 222844 233148 222896
rect 233200 222884 233206 222896
rect 277670 222884 277676 222896
rect 233200 222856 277676 222884
rect 233200 222844 233206 222856
rect 277670 222844 277676 222856
rect 277728 222844 277734 222896
rect 284110 222844 284116 222896
rect 284168 222884 284174 222896
rect 316678 222884 316684 222896
rect 284168 222856 316684 222884
rect 284168 222844 284174 222856
rect 316678 222844 316684 222856
rect 316736 222844 316742 222896
rect 316862 222844 316868 222896
rect 316920 222884 316926 222896
rect 343174 222884 343180 222896
rect 316920 222856 343180 222884
rect 316920 222844 316926 222856
rect 343174 222844 343180 222856
rect 343232 222844 343238 222896
rect 347498 222844 347504 222896
rect 347556 222884 347562 222896
rect 368474 222884 368480 222896
rect 347556 222856 368480 222884
rect 347556 222844 347562 222856
rect 368474 222844 368480 222856
rect 368532 222844 368538 222896
rect 375098 222844 375104 222896
rect 375156 222884 375162 222896
rect 391014 222884 391020 222896
rect 375156 222856 391020 222884
rect 375156 222844 375162 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 397178 222844 397184 222896
rect 397236 222884 397242 222896
rect 407206 222884 407212 222896
rect 397236 222856 407212 222884
rect 397236 222844 397242 222856
rect 407206 222844 407212 222856
rect 407264 222844 407270 222896
rect 408402 222844 408408 222896
rect 408460 222884 408466 222896
rect 416774 222884 416780 222896
rect 408460 222856 416780 222884
rect 408460 222844 408466 222856
rect 416774 222844 416780 222856
rect 416832 222844 416838 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 466730 222884 466736 222896
rect 459980 222856 466736 222884
rect 459980 222844 459986 222856
rect 466730 222844 466736 222856
rect 466788 222844 466794 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473446 222884 473452 222896
rect 467524 222856 473452 222884
rect 467524 222844 467530 222856
rect 473446 222844 473452 222856
rect 473504 222844 473510 222896
rect 474734 222844 474740 222896
rect 474792 222884 474798 222896
rect 484854 222884 484860 222896
rect 474792 222856 484860 222884
rect 474792 222844 474798 222856
rect 484854 222844 484860 222856
rect 484912 222844 484918 222896
rect 489546 222844 489552 222896
rect 489604 222884 489610 222896
rect 503990 222884 503996 222896
rect 489604 222856 503996 222884
rect 489604 222844 489610 222856
rect 503990 222844 503996 222856
rect 504048 222844 504054 222896
rect 504634 222844 504640 222896
rect 504692 222884 504698 222896
rect 523770 222884 523776 222896
rect 504692 222856 523776 222884
rect 504692 222844 504698 222856
rect 523770 222844 523776 222856
rect 523828 222844 523834 222896
rect 533706 222844 533712 222896
rect 533764 222884 533770 222896
rect 560662 222884 560668 222896
rect 533764 222856 560668 222884
rect 533764 222844 533770 222856
rect 560662 222844 560668 222856
rect 560720 222884 560726 222896
rect 562962 222884 562968 222896
rect 560720 222856 562968 222884
rect 560720 222844 560726 222856
rect 562962 222844 562968 222856
rect 563020 222844 563026 222896
rect 571426 222844 571432 222896
rect 571484 222884 571490 222896
rect 571886 222884 571892 222896
rect 571484 222856 571892 222884
rect 571484 222844 571490 222856
rect 571886 222844 571892 222856
rect 571944 222844 571950 222896
rect 204916 222720 212396 222748
rect 195440 222652 195560 222680
rect 192018 222612 192024 222624
rect 181456 222584 192024 222612
rect 192018 222572 192024 222584
rect 192076 222572 192082 222624
rect 195532 222612 195560 222652
rect 204916 222612 204944 222720
rect 213822 222708 213828 222760
rect 213880 222748 213886 222760
rect 262858 222748 262864 222760
rect 213880 222720 262864 222748
rect 213880 222708 213886 222720
rect 262858 222708 262864 222720
rect 262916 222708 262922 222760
rect 263502 222708 263508 222760
rect 263560 222748 263566 222760
rect 296990 222748 296996 222760
rect 263560 222720 296996 222748
rect 263560 222708 263566 222720
rect 296990 222708 296996 222720
rect 297048 222708 297054 222760
rect 563974 222640 563980 222692
rect 564032 222680 564038 222692
rect 574646 222680 574652 222692
rect 564032 222652 574652 222680
rect 564032 222640 564038 222652
rect 574646 222640 574652 222652
rect 574704 222640 574710 222692
rect 195532 222584 204944 222612
rect 205082 222572 205088 222624
rect 205140 222612 205146 222624
rect 208762 222612 208768 222624
rect 205140 222584 208768 222612
rect 205140 222572 205146 222584
rect 208762 222572 208768 222584
rect 208820 222572 208826 222624
rect 209498 222572 209504 222624
rect 209556 222612 209562 222624
rect 210234 222612 210240 222624
rect 209556 222584 210240 222612
rect 209556 222572 209562 222584
rect 210234 222572 210240 222584
rect 210292 222572 210298 222624
rect 210878 222572 210884 222624
rect 210936 222612 210942 222624
rect 260282 222612 260288 222624
rect 210936 222584 260288 222612
rect 210936 222572 210942 222584
rect 260282 222572 260288 222584
rect 260340 222572 260346 222624
rect 572254 222544 572260 222556
rect 563026 222516 572260 222544
rect 117958 222436 117964 222488
rect 118016 222476 118022 222488
rect 137278 222476 137284 222488
rect 118016 222448 137284 222476
rect 118016 222436 118022 222448
rect 137278 222436 137284 222448
rect 137336 222436 137342 222488
rect 137462 222436 137468 222488
rect 137520 222476 137526 222488
rect 151354 222476 151360 222488
rect 137520 222448 151360 222476
rect 137520 222436 137526 222448
rect 151354 222436 151360 222448
rect 151412 222436 151418 222488
rect 152274 222436 152280 222488
rect 152332 222476 152338 222488
rect 157058 222476 157064 222488
rect 152332 222448 157064 222476
rect 152332 222436 152338 222448
rect 157058 222436 157064 222448
rect 157116 222436 157122 222488
rect 157242 222436 157248 222488
rect 157300 222476 157306 222488
rect 219710 222476 219716 222488
rect 157300 222448 219716 222476
rect 157300 222436 157306 222448
rect 219710 222436 219716 222448
rect 219768 222436 219774 222488
rect 220078 222436 220084 222488
rect 220136 222476 220142 222488
rect 268654 222476 268660 222488
rect 220136 222448 268660 222476
rect 220136 222436 220142 222448
rect 268654 222436 268660 222448
rect 268712 222436 268718 222488
rect 555234 222368 555240 222420
rect 555292 222408 555298 222420
rect 562134 222408 562140 222420
rect 555292 222380 562140 222408
rect 555292 222368 555298 222380
rect 562134 222368 562140 222380
rect 562192 222408 562198 222420
rect 563026 222408 563054 222516
rect 572254 222504 572260 222516
rect 572312 222504 572318 222556
rect 562192 222380 563054 222408
rect 562192 222368 562198 222380
rect 565078 222368 565084 222420
rect 565136 222408 565142 222420
rect 568666 222408 568672 222420
rect 565136 222380 568672 222408
rect 565136 222368 565142 222380
rect 568666 222368 568672 222380
rect 568724 222368 568730 222420
rect 570138 222368 570144 222420
rect 570196 222408 570202 222420
rect 574462 222408 574468 222420
rect 570196 222380 574468 222408
rect 570196 222368 570202 222380
rect 574462 222368 574468 222380
rect 574520 222368 574526 222420
rect 112898 222300 112904 222352
rect 112956 222340 112962 222352
rect 118142 222340 118148 222352
rect 112956 222312 118148 222340
rect 112956 222300 112962 222312
rect 118142 222300 118148 222312
rect 118200 222300 118206 222352
rect 133598 222300 133604 222352
rect 133656 222340 133662 222352
rect 136910 222340 136916 222352
rect 133656 222312 136916 222340
rect 133656 222300 133662 222312
rect 136910 222300 136916 222312
rect 136968 222300 136974 222352
rect 137094 222300 137100 222352
rect 137152 222340 137158 222352
rect 142614 222340 142620 222352
rect 137152 222312 142620 222340
rect 137152 222300 137158 222312
rect 142614 222300 142620 222312
rect 142672 222300 142678 222352
rect 145006 222300 145012 222352
rect 145064 222340 145070 222352
rect 145064 222312 200114 222340
rect 145064 222300 145070 222312
rect 143442 222232 143448 222284
rect 143500 222272 143506 222284
rect 144822 222272 144828 222284
rect 143500 222244 144828 222272
rect 143500 222232 143506 222244
rect 144822 222232 144828 222244
rect 144880 222232 144886 222284
rect 200086 222272 200114 222312
rect 203702 222300 203708 222352
rect 203760 222340 203766 222352
rect 207474 222340 207480 222352
rect 203760 222312 207480 222340
rect 203760 222300 203766 222312
rect 207474 222300 207480 222312
rect 207532 222300 207538 222352
rect 212166 222300 212172 222352
rect 212224 222340 212230 222352
rect 216214 222340 216220 222352
rect 212224 222312 216220 222340
rect 212224 222300 212230 222312
rect 216214 222300 216220 222312
rect 216272 222300 216278 222352
rect 220722 222300 220728 222352
rect 220780 222340 220786 222352
rect 268010 222340 268016 222352
rect 220780 222312 268016 222340
rect 220780 222300 220786 222312
rect 268010 222300 268016 222312
rect 268068 222300 268074 222352
rect 203518 222272 203524 222284
rect 200086 222244 203524 222272
rect 203518 222232 203524 222244
rect 203576 222232 203582 222284
rect 593966 222272 593972 222284
rect 528526 222244 593972 222272
rect 171134 222204 171140 222216
rect 171106 222164 171140 222204
rect 171192 222164 171198 222216
rect 482830 222164 482836 222216
rect 482888 222204 482894 222216
rect 528526 222204 528554 222244
rect 593966 222232 593972 222244
rect 594024 222232 594030 222284
rect 596634 222232 596640 222284
rect 596692 222272 596698 222284
rect 596692 222244 597048 222272
rect 596692 222232 596698 222244
rect 482888 222176 528554 222204
rect 482888 222164 482894 222176
rect 117958 222136 117964 222148
rect 103486 222108 117964 222136
rect 95694 221960 95700 222012
rect 95752 222000 95758 222012
rect 103486 222000 103514 222108
rect 117958 222096 117964 222108
rect 118016 222096 118022 222148
rect 118142 222096 118148 222148
rect 118200 222136 118206 222148
rect 171106 222136 171134 222164
rect 118200 222108 171134 222136
rect 118200 222096 118206 222108
rect 171318 222096 171324 222148
rect 171376 222136 171382 222148
rect 177390 222136 177396 222148
rect 171376 222108 177396 222136
rect 171376 222096 171382 222108
rect 177390 222096 177396 222108
rect 177448 222096 177454 222148
rect 177574 222096 177580 222148
rect 177632 222136 177638 222148
rect 179966 222136 179972 222148
rect 177632 222108 179972 222136
rect 177632 222096 177638 222108
rect 179966 222096 179972 222108
rect 180024 222096 180030 222148
rect 180150 222096 180156 222148
rect 180208 222136 180214 222148
rect 180208 222108 181668 222136
rect 180208 222096 180214 222108
rect 95752 221972 103514 222000
rect 95752 221960 95758 221972
rect 104618 221960 104624 222012
rect 104676 222000 104682 222012
rect 171042 222000 171048 222012
rect 104676 221972 171048 222000
rect 104676 221960 104682 221972
rect 171042 221960 171048 221972
rect 171100 221960 171106 222012
rect 172974 222000 172980 222012
rect 171244 221972 172980 222000
rect 71682 221824 71688 221876
rect 71740 221864 71746 221876
rect 142798 221864 142804 221876
rect 71740 221836 142804 221864
rect 71740 221824 71746 221836
rect 142798 221824 142804 221836
rect 142856 221824 142862 221876
rect 143166 221824 143172 221876
rect 143224 221864 143230 221876
rect 171244 221864 171272 221972
rect 172974 221960 172980 221972
rect 173032 221960 173038 222012
rect 176286 221960 176292 222012
rect 176344 222000 176350 222012
rect 181438 222000 181444 222012
rect 176344 221972 181444 222000
rect 176344 221960 176350 221972
rect 181438 221960 181444 221972
rect 181496 221960 181502 222012
rect 181640 222000 181668 222108
rect 181806 222096 181812 222148
rect 181864 222136 181870 222148
rect 240134 222136 240140 222148
rect 181864 222108 240140 222136
rect 181864 222096 181870 222108
rect 240134 222096 240140 222108
rect 240192 222096 240198 222148
rect 256326 222096 256332 222148
rect 256384 222136 256390 222148
rect 261202 222136 261208 222148
rect 256384 222108 261208 222136
rect 256384 222096 256390 222108
rect 261202 222096 261208 222108
rect 261260 222096 261266 222148
rect 261386 222096 261392 222148
rect 261444 222136 261450 222148
rect 301682 222136 301688 222148
rect 261444 222108 301688 222136
rect 261444 222096 261450 222108
rect 301682 222096 301688 222108
rect 301740 222096 301746 222148
rect 331674 222096 331680 222148
rect 331732 222136 331738 222148
rect 353938 222136 353944 222148
rect 331732 222108 353944 222136
rect 331732 222096 331738 222108
rect 353938 222096 353944 222108
rect 353996 222096 354002 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468478 222136 468484 222148
rect 462188 222108 468484 222136
rect 462188 222096 462194 222108
rect 468478 222096 468484 222108
rect 468536 222096 468542 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477586 222136 477592 222148
rect 471940 222108 477592 222136
rect 471940 222096 471946 222108
rect 477586 222096 477592 222108
rect 477644 222096 477650 222148
rect 547138 222096 547144 222148
rect 547196 222136 547202 222148
rect 557994 222136 558000 222148
rect 547196 222108 558000 222136
rect 547196 222096 547202 222108
rect 557994 222096 558000 222108
rect 558052 222096 558058 222148
rect 558178 222096 558184 222148
rect 558236 222136 558242 222148
rect 562870 222136 562876 222148
rect 558236 222108 562876 222136
rect 558236 222096 558242 222108
rect 562870 222096 562876 222108
rect 562928 222096 562934 222148
rect 564894 222136 564900 222148
rect 563164 222108 564900 222136
rect 237374 222000 237380 222012
rect 181640 221972 237380 222000
rect 237374 221960 237380 221972
rect 237432 221960 237438 222012
rect 243906 221960 243912 222012
rect 243964 222000 243970 222012
rect 285674 222000 285680 222012
rect 243964 221972 285680 222000
rect 243964 221960 243970 221972
rect 285674 221960 285680 221972
rect 285732 221960 285738 222012
rect 310146 221960 310152 222012
rect 310204 222000 310210 222012
rect 338114 222000 338120 222012
rect 310204 221972 338120 222000
rect 310204 221960 310210 221972
rect 338114 221960 338120 221972
rect 338172 221960 338178 222012
rect 517606 221960 517612 222012
rect 517664 222000 517670 222012
rect 518526 222000 518532 222012
rect 517664 221972 518532 222000
rect 517664 221960 517670 221972
rect 518526 221960 518532 221972
rect 518584 222000 518590 222012
rect 562686 222000 562692 222012
rect 518584 221972 562692 222000
rect 518584 221960 518590 221972
rect 562686 221960 562692 221972
rect 562744 221960 562750 222012
rect 424962 221892 424968 221944
rect 425020 221932 425026 221944
rect 429194 221932 429200 221944
rect 425020 221904 429200 221932
rect 425020 221892 425026 221904
rect 429194 221892 429200 221904
rect 429252 221892 429258 221944
rect 563164 221932 563192 222108
rect 564894 222096 564900 222108
rect 564952 222096 564958 222148
rect 565354 222096 565360 222148
rect 565412 222136 565418 222148
rect 596818 222136 596824 222148
rect 565412 222108 596824 222136
rect 565412 222096 565418 222108
rect 596818 222096 596824 222108
rect 596876 222096 596882 222148
rect 597020 222136 597048 222244
rect 600406 222136 600412 222148
rect 597020 222108 600412 222136
rect 600406 222096 600412 222108
rect 600464 222096 600470 222148
rect 563514 221960 563520 222012
rect 563572 222000 563578 222012
rect 591942 222000 591948 222012
rect 563572 221972 591948 222000
rect 563572 221960 563578 221972
rect 591942 221960 591948 221972
rect 592000 221960 592006 222012
rect 592126 221960 592132 222012
rect 592184 222000 592190 222012
rect 599118 222000 599124 222012
rect 592184 221972 599124 222000
rect 592184 221960 592190 221972
rect 599118 221960 599124 221972
rect 599176 221960 599182 222012
rect 599302 221960 599308 222012
rect 599360 222000 599366 222012
rect 600590 222000 600596 222012
rect 599360 221972 600596 222000
rect 599360 221960 599366 221972
rect 600590 221960 600596 221972
rect 600648 221960 600654 222012
rect 562888 221904 563192 221932
rect 143224 221836 171272 221864
rect 143224 221824 143230 221836
rect 171410 221824 171416 221876
rect 171468 221864 171474 221876
rect 229646 221864 229652 221876
rect 171468 221836 229652 221864
rect 171468 221824 171474 221836
rect 229646 221824 229652 221836
rect 229704 221824 229710 221876
rect 237282 221824 237288 221876
rect 237340 221864 237346 221876
rect 280430 221864 280436 221876
rect 237340 221836 280436 221864
rect 237340 221824 237346 221836
rect 280430 221824 280436 221836
rect 280488 221824 280494 221876
rect 285674 221824 285680 221876
rect 285732 221864 285738 221876
rect 286318 221864 286324 221876
rect 285732 221836 286324 221864
rect 285732 221824 285738 221836
rect 286318 221824 286324 221836
rect 286376 221824 286382 221876
rect 304718 221824 304724 221876
rect 304776 221864 304782 221876
rect 334066 221864 334072 221876
rect 304776 221836 334072 221864
rect 304776 221824 304782 221836
rect 334066 221824 334072 221836
rect 334124 221824 334130 221876
rect 505738 221824 505744 221876
rect 505796 221864 505802 221876
rect 523954 221864 523960 221876
rect 505796 221836 523960 221864
rect 505796 221824 505802 221836
rect 523954 221824 523960 221836
rect 524012 221824 524018 221876
rect 529842 221824 529848 221876
rect 529900 221864 529906 221876
rect 555694 221864 555700 221876
rect 529900 221836 555700 221864
rect 529900 221824 529906 221836
rect 555694 221824 555700 221836
rect 555752 221824 555758 221876
rect 559558 221824 559564 221876
rect 559616 221864 559622 221876
rect 562888 221864 562916 221904
rect 559616 221836 562916 221864
rect 559616 221824 559622 221836
rect 563330 221824 563336 221876
rect 563388 221864 563394 221876
rect 609974 221864 609980 221876
rect 563388 221836 609980 221864
rect 563388 221824 563394 221836
rect 609974 221824 609980 221836
rect 610032 221824 610038 221876
rect 68370 221688 68376 221740
rect 68428 221728 68434 221740
rect 147490 221728 147496 221740
rect 68428 221700 147496 221728
rect 68428 221688 68434 221700
rect 147490 221688 147496 221700
rect 147548 221688 147554 221740
rect 154546 221700 157334 221728
rect 61746 221552 61752 221604
rect 61804 221592 61810 221604
rect 137278 221592 137284 221604
rect 61804 221564 137284 221592
rect 61804 221552 61810 221564
rect 137278 221552 137284 221564
rect 137336 221552 137342 221604
rect 137462 221552 137468 221604
rect 137520 221592 137526 221604
rect 137520 221564 142660 221592
rect 137520 221552 137526 221564
rect 64598 221416 64604 221468
rect 64656 221456 64662 221468
rect 138566 221456 138572 221468
rect 64656 221428 138572 221456
rect 64656 221416 64662 221428
rect 138566 221416 138572 221428
rect 138624 221416 138630 221468
rect 138750 221416 138756 221468
rect 138808 221456 138814 221468
rect 142430 221456 142436 221468
rect 138808 221428 142436 221456
rect 138808 221416 138814 221428
rect 142430 221416 142436 221428
rect 142488 221416 142494 221468
rect 142632 221456 142660 221564
rect 142798 221552 142804 221604
rect 142856 221592 142862 221604
rect 147306 221592 147312 221604
rect 142856 221564 147312 221592
rect 142856 221552 142862 221564
rect 147306 221552 147312 221564
rect 147364 221552 147370 221604
rect 154546 221592 154574 221700
rect 147784 221564 154574 221592
rect 157306 221592 157334 221700
rect 161750 221688 161756 221740
rect 161808 221728 161814 221740
rect 224402 221728 224408 221740
rect 161808 221700 224408 221728
rect 161808 221688 161814 221700
rect 224402 221688 224408 221700
rect 224460 221688 224466 221740
rect 230382 221688 230388 221740
rect 230440 221728 230446 221740
rect 275186 221728 275192 221740
rect 230440 221700 275192 221728
rect 230440 221688 230446 221700
rect 275186 221688 275192 221700
rect 275244 221688 275250 221740
rect 275370 221688 275376 221740
rect 275428 221728 275434 221740
rect 310882 221728 310888 221740
rect 275428 221700 310888 221728
rect 275428 221688 275434 221700
rect 310882 221688 310888 221700
rect 310940 221688 310946 221740
rect 311526 221688 311532 221740
rect 311584 221728 311590 221740
rect 338390 221728 338396 221740
rect 311584 221700 338396 221728
rect 311584 221688 311590 221700
rect 338390 221688 338396 221700
rect 338448 221688 338454 221740
rect 341610 221728 341616 221740
rect 338592 221700 341616 221728
rect 204898 221592 204904 221604
rect 157306 221564 204904 221592
rect 143166 221456 143172 221468
rect 142632 221428 143172 221456
rect 143166 221416 143172 221428
rect 143224 221416 143230 221468
rect 145374 221416 145380 221468
rect 145432 221456 145438 221468
rect 147784 221456 147812 221564
rect 204898 221552 204904 221564
rect 204956 221552 204962 221604
rect 205082 221552 205088 221604
rect 205140 221592 205146 221604
rect 205140 221564 212304 221592
rect 205140 221552 205146 221564
rect 145432 221428 147812 221456
rect 145432 221416 145438 221428
rect 148778 221416 148784 221468
rect 148836 221456 148842 221468
rect 211982 221456 211988 221468
rect 148836 221428 211988 221456
rect 148836 221416 148842 221428
rect 211982 221416 211988 221428
rect 212040 221416 212046 221468
rect 212276 221456 212304 221564
rect 214926 221552 214932 221604
rect 214984 221592 214990 221604
rect 265710 221592 265716 221604
rect 214984 221564 265716 221592
rect 214984 221552 214990 221564
rect 265710 221552 265716 221564
rect 265768 221552 265774 221604
rect 267734 221552 267740 221604
rect 267792 221592 267798 221604
rect 273990 221592 273996 221604
rect 267792 221564 273996 221592
rect 267792 221552 267798 221564
rect 273990 221552 273996 221564
rect 274048 221552 274054 221604
rect 278222 221552 278228 221604
rect 278280 221592 278286 221604
rect 313274 221592 313280 221604
rect 278280 221564 313280 221592
rect 278280 221552 278286 221564
rect 313274 221552 313280 221564
rect 313332 221552 313338 221604
rect 314562 221552 314568 221604
rect 314620 221592 314626 221604
rect 338592 221592 338620 221700
rect 341610 221688 341616 221700
rect 341668 221688 341674 221740
rect 359826 221688 359832 221740
rect 359884 221728 359890 221740
rect 376846 221728 376852 221740
rect 359884 221700 376852 221728
rect 359884 221688 359890 221700
rect 376846 221688 376852 221700
rect 376904 221688 376910 221740
rect 496170 221688 496176 221740
rect 496228 221728 496234 221740
rect 513558 221728 513564 221740
rect 496228 221700 513564 221728
rect 496228 221688 496234 221700
rect 513558 221688 513564 221700
rect 513616 221688 513622 221740
rect 527818 221688 527824 221740
rect 527876 221728 527882 221740
rect 542446 221728 542452 221740
rect 527876 221700 542452 221728
rect 527876 221688 527882 221700
rect 542446 221688 542452 221700
rect 542504 221688 542510 221740
rect 553210 221688 553216 221740
rect 553268 221728 553274 221740
rect 608962 221728 608968 221740
rect 553268 221700 608968 221728
rect 553268 221688 553274 221700
rect 608962 221688 608968 221700
rect 609020 221688 609026 221740
rect 314620 221564 338620 221592
rect 314620 221552 314626 221564
rect 341610 221552 341616 221604
rect 341668 221592 341674 221604
rect 361574 221592 361580 221604
rect 341668 221564 361580 221592
rect 341668 221552 341674 221564
rect 361574 221552 361580 221564
rect 361632 221552 361638 221604
rect 378042 221552 378048 221604
rect 378100 221592 378106 221604
rect 390002 221592 390008 221604
rect 378100 221564 390008 221592
rect 378100 221552 378106 221564
rect 390002 221552 390008 221564
rect 390060 221552 390066 221604
rect 456702 221552 456708 221604
rect 456760 221592 456766 221604
rect 461762 221592 461768 221604
rect 456760 221564 461768 221592
rect 456760 221552 456766 221564
rect 461762 221552 461768 221564
rect 461820 221552 461826 221604
rect 484302 221552 484308 221604
rect 484360 221592 484366 221604
rect 495802 221592 495808 221604
rect 484360 221564 495808 221592
rect 484360 221552 484366 221564
rect 495802 221552 495808 221564
rect 495860 221552 495866 221604
rect 500034 221552 500040 221604
rect 500092 221592 500098 221604
rect 517606 221592 517612 221604
rect 500092 221564 517612 221592
rect 500092 221552 500098 221564
rect 517606 221552 517612 221564
rect 517664 221552 517670 221604
rect 518158 221552 518164 221604
rect 518216 221592 518222 221604
rect 530026 221592 530032 221604
rect 518216 221564 530032 221592
rect 518216 221552 518222 221564
rect 530026 221552 530032 221564
rect 530084 221552 530090 221604
rect 534810 221552 534816 221604
rect 534868 221592 534874 221604
rect 547414 221592 547420 221604
rect 534868 221564 547420 221592
rect 534868 221552 534874 221564
rect 547414 221552 547420 221564
rect 547472 221552 547478 221604
rect 552658 221552 552664 221604
rect 552716 221592 552722 221604
rect 553670 221592 553676 221604
rect 552716 221564 553676 221592
rect 552716 221552 552722 221564
rect 553670 221552 553676 221564
rect 553728 221552 553734 221604
rect 553854 221552 553860 221604
rect 553912 221592 553918 221604
rect 557074 221592 557080 221604
rect 553912 221564 557080 221592
rect 553912 221552 553918 221564
rect 557074 221552 557080 221564
rect 557132 221552 557138 221604
rect 557994 221552 558000 221604
rect 558052 221592 558058 221604
rect 559834 221592 559840 221604
rect 558052 221564 559840 221592
rect 558052 221552 558058 221564
rect 559834 221552 559840 221564
rect 559892 221592 559898 221604
rect 563146 221592 563152 221604
rect 559892 221564 563152 221592
rect 559892 221552 559898 221564
rect 563146 221552 563152 221564
rect 563204 221552 563210 221604
rect 563698 221552 563704 221604
rect 563756 221592 563762 221604
rect 608778 221592 608784 221604
rect 563756 221564 608784 221592
rect 563756 221552 563762 221564
rect 608778 221552 608784 221564
rect 608836 221552 608842 221604
rect 232130 221456 232136 221468
rect 212276 221428 232136 221456
rect 232130 221416 232136 221428
rect 232188 221416 232194 221468
rect 241238 221416 241244 221468
rect 241296 221456 241302 221468
rect 285674 221456 285680 221468
rect 241296 221428 285680 221456
rect 241296 221416 241302 221428
rect 285674 221416 285680 221428
rect 285732 221416 285738 221468
rect 286042 221416 286048 221468
rect 286100 221456 286106 221468
rect 289906 221456 289912 221468
rect 286100 221428 289912 221456
rect 286100 221416 286106 221428
rect 289906 221416 289912 221428
rect 289964 221416 289970 221468
rect 290274 221416 290280 221468
rect 290332 221456 290338 221468
rect 321738 221456 321744 221468
rect 290332 221428 321744 221456
rect 290332 221416 290338 221428
rect 321738 221416 321744 221428
rect 321796 221416 321802 221468
rect 339126 221416 339132 221468
rect 339184 221456 339190 221468
rect 362034 221456 362040 221468
rect 339184 221428 362040 221456
rect 339184 221416 339190 221428
rect 362034 221416 362040 221428
rect 362092 221416 362098 221468
rect 362310 221416 362316 221468
rect 362368 221456 362374 221468
rect 380250 221456 380256 221468
rect 362368 221428 380256 221456
rect 362368 221416 362374 221428
rect 380250 221416 380256 221428
rect 380308 221416 380314 221468
rect 391290 221416 391296 221468
rect 391348 221456 391354 221468
rect 400398 221456 400404 221468
rect 391348 221428 400404 221456
rect 391348 221416 391354 221428
rect 400398 221416 400404 221428
rect 400456 221416 400462 221468
rect 405366 221416 405372 221468
rect 405424 221456 405430 221468
rect 414198 221456 414204 221468
rect 405424 221428 414204 221456
rect 405424 221416 405430 221428
rect 414198 221416 414204 221428
rect 414256 221416 414262 221468
rect 452562 221416 452568 221468
rect 452620 221456 452626 221468
rect 456702 221456 456708 221468
rect 452620 221428 456708 221456
rect 452620 221416 452626 221428
rect 456702 221416 456708 221428
rect 456760 221416 456766 221468
rect 484026 221416 484032 221468
rect 484084 221456 484090 221468
rect 538674 221456 538680 221468
rect 484084 221428 538680 221456
rect 484084 221416 484090 221428
rect 538674 221416 538680 221428
rect 538732 221416 538738 221468
rect 540054 221416 540060 221468
rect 540112 221456 540118 221468
rect 540882 221456 540888 221468
rect 540112 221428 540888 221456
rect 540112 221416 540118 221428
rect 540882 221416 540888 221428
rect 540940 221456 540946 221468
rect 606018 221456 606024 221468
rect 540940 221428 606024 221456
rect 540940 221416 540946 221428
rect 606018 221416 606024 221428
rect 606076 221416 606082 221468
rect 114462 221280 114468 221332
rect 114520 221320 114526 221332
rect 178310 221320 178316 221332
rect 114520 221292 178316 221320
rect 114520 221280 114526 221292
rect 178310 221280 178316 221292
rect 178368 221280 178374 221332
rect 178494 221280 178500 221332
rect 178552 221320 178558 221332
rect 180150 221320 180156 221332
rect 178552 221292 180156 221320
rect 178552 221280 178558 221292
rect 180150 221280 180156 221292
rect 180208 221280 180214 221332
rect 181438 221280 181444 221332
rect 181496 221320 181502 221332
rect 195238 221320 195244 221332
rect 181496 221292 195244 221320
rect 181496 221280 181502 221292
rect 195238 221280 195244 221292
rect 195296 221280 195302 221332
rect 195422 221280 195428 221332
rect 195480 221320 195486 221332
rect 245102 221320 245108 221332
rect 195480 221292 245108 221320
rect 195480 221280 195486 221292
rect 245102 221280 245108 221292
rect 245160 221280 245166 221332
rect 273714 221280 273720 221332
rect 273772 221320 273778 221332
rect 309226 221320 309232 221332
rect 273772 221292 309232 221320
rect 273772 221280 273778 221292
rect 309226 221280 309232 221292
rect 309284 221280 309290 221332
rect 525058 221280 525064 221332
rect 525116 221320 525122 221332
rect 535086 221320 535092 221332
rect 525116 221292 535092 221320
rect 525116 221280 525122 221292
rect 535086 221280 535092 221292
rect 535144 221320 535150 221332
rect 543550 221320 543556 221332
rect 535144 221292 543556 221320
rect 535144 221280 535150 221292
rect 543550 221280 543556 221292
rect 543608 221280 543614 221332
rect 547874 221212 547880 221264
rect 547932 221252 547938 221264
rect 549070 221252 549076 221264
rect 547932 221224 549076 221252
rect 547932 221212 547938 221224
rect 549070 221212 549076 221224
rect 549128 221212 549134 221264
rect 550634 221212 550640 221264
rect 550692 221252 550698 221264
rect 607766 221252 607772 221264
rect 550692 221224 607772 221252
rect 550692 221212 550698 221224
rect 607766 221212 607772 221224
rect 607824 221212 607830 221264
rect 117958 221144 117964 221196
rect 118016 221184 118022 221196
rect 137094 221184 137100 221196
rect 118016 221156 137100 221184
rect 118016 221144 118022 221156
rect 137094 221144 137100 221156
rect 137152 221144 137158 221196
rect 137278 221144 137284 221196
rect 137336 221184 137342 221196
rect 143994 221184 144000 221196
rect 137336 221156 144000 221184
rect 137336 221144 137342 221156
rect 143994 221144 144000 221156
rect 144052 221144 144058 221196
rect 144178 221144 144184 221196
rect 144236 221184 144242 221196
rect 203242 221184 203248 221196
rect 144236 221156 203248 221184
rect 144236 221144 144242 221156
rect 203242 221144 203248 221156
rect 203300 221144 203306 221196
rect 205082 221184 205088 221196
rect 204732 221156 205088 221184
rect 108114 221008 108120 221060
rect 108172 221048 108178 221060
rect 118142 221048 118148 221060
rect 108172 221020 118148 221048
rect 108172 221008 108178 221020
rect 118142 221008 118148 221020
rect 118200 221008 118206 221060
rect 128814 221008 128820 221060
rect 128872 221048 128878 221060
rect 195054 221048 195060 221060
rect 128872 221020 195060 221048
rect 128872 221008 128878 221020
rect 195054 221008 195060 221020
rect 195112 221008 195118 221060
rect 195238 221008 195244 221060
rect 195296 221048 195302 221060
rect 204732 221048 204760 221156
rect 205082 221144 205088 221156
rect 205140 221144 205146 221196
rect 206002 221144 206008 221196
rect 206060 221184 206066 221196
rect 258074 221184 258080 221196
rect 206060 221156 258080 221184
rect 206060 221144 206066 221156
rect 258074 221144 258080 221156
rect 258132 221144 258138 221196
rect 530578 221076 530584 221128
rect 530636 221116 530642 221128
rect 603442 221116 603448 221128
rect 530636 221088 603448 221116
rect 530636 221076 530642 221088
rect 603442 221076 603448 221088
rect 603500 221076 603506 221128
rect 195296 221020 204760 221048
rect 195296 221008 195302 221020
rect 204898 221008 204904 221060
rect 204956 221048 204962 221060
rect 211614 221048 211620 221060
rect 204956 221020 211620 221048
rect 204956 221008 204962 221020
rect 211614 221008 211620 221020
rect 211672 221008 211678 221060
rect 211982 221008 211988 221060
rect 212040 221048 212046 221060
rect 214282 221048 214288 221060
rect 212040 221020 214288 221048
rect 212040 221008 212046 221020
rect 214282 221008 214288 221020
rect 214340 221008 214346 221060
rect 227346 221008 227352 221060
rect 227404 221048 227410 221060
rect 272702 221048 272708 221060
rect 227404 221020 272708 221048
rect 227404 221008 227410 221020
rect 272702 221008 272708 221020
rect 272760 221008 272766 221060
rect 415118 221008 415124 221060
rect 415176 221048 415182 221060
rect 420178 221048 420184 221060
rect 415176 221020 420184 221048
rect 415176 221008 415182 221020
rect 420178 221008 420184 221020
rect 420236 221008 420242 221060
rect 516042 220940 516048 220992
rect 516100 220980 516106 220992
rect 596634 220980 596640 220992
rect 516100 220952 596640 220980
rect 516100 220940 516106 220952
rect 596634 220940 596640 220952
rect 596692 220940 596698 220992
rect 107930 220872 107936 220924
rect 107988 220912 107994 220924
rect 107988 220884 108528 220912
rect 107988 220872 107994 220884
rect 97718 220736 97724 220788
rect 97776 220776 97782 220788
rect 108500 220776 108528 220884
rect 118050 220872 118056 220924
rect 118108 220912 118114 220924
rect 187878 220912 187884 220924
rect 118108 220884 187884 220912
rect 118108 220872 118114 220884
rect 187878 220872 187884 220884
rect 187936 220872 187942 220924
rect 188430 220872 188436 220924
rect 188488 220912 188494 220924
rect 195422 220912 195428 220924
rect 188488 220884 195428 220912
rect 188488 220872 188494 220884
rect 195422 220872 195428 220884
rect 195480 220872 195486 220924
rect 198918 220912 198924 220924
rect 195624 220884 198924 220912
rect 137278 220776 137284 220788
rect 97776 220748 108252 220776
rect 108500 220748 137284 220776
rect 97776 220736 97782 220748
rect 108224 220708 108252 220748
rect 137278 220736 137284 220748
rect 137336 220736 137342 220788
rect 137462 220736 137468 220788
rect 137520 220776 137526 220788
rect 194870 220776 194876 220788
rect 137520 220748 194876 220776
rect 137520 220736 137526 220748
rect 194870 220736 194876 220748
rect 194928 220736 194934 220788
rect 195054 220736 195060 220788
rect 195112 220776 195118 220788
rect 195624 220776 195652 220884
rect 198918 220872 198924 220884
rect 198976 220872 198982 220924
rect 203242 220872 203248 220924
rect 203300 220912 203306 220924
rect 206462 220912 206468 220924
rect 203300 220884 206468 220912
rect 203300 220872 203306 220884
rect 206462 220872 206468 220884
rect 206520 220872 206526 220924
rect 596818 220872 596824 220924
rect 596876 220912 596882 220924
rect 611630 220912 611636 220924
rect 596876 220884 611636 220912
rect 596876 220872 596882 220884
rect 611630 220872 611636 220884
rect 611688 220872 611694 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423766 220844 423772 220856
rect 420696 220816 423772 220844
rect 420696 220804 420702 220816
rect 423766 220804 423772 220816
rect 423824 220804 423830 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471698 220844 471704 220856
rect 466144 220816 471704 220844
rect 466144 220804 466150 220816
rect 471698 220804 471704 220816
rect 471756 220804 471762 220856
rect 513558 220804 513564 220856
rect 513616 220844 513622 220856
rect 592126 220844 592132 220856
rect 513616 220816 592132 220844
rect 513616 220804 513622 220816
rect 592126 220804 592132 220816
rect 592184 220804 592190 220856
rect 195112 220748 195652 220776
rect 195112 220736 195118 220748
rect 196066 220736 196072 220788
rect 196124 220776 196130 220788
rect 197814 220776 197820 220788
rect 196124 220748 197820 220776
rect 196124 220736 196130 220748
rect 197814 220736 197820 220748
rect 197872 220736 197878 220788
rect 198366 220736 198372 220788
rect 198424 220776 198430 220788
rect 252738 220776 252744 220788
rect 198424 220748 252744 220776
rect 198424 220736 198430 220748
rect 252738 220736 252744 220748
rect 252796 220736 252802 220788
rect 257154 220736 257160 220788
rect 257212 220776 257218 220788
rect 295886 220776 295892 220788
rect 257212 220748 295892 220776
rect 257212 220736 257218 220748
rect 295886 220736 295892 220748
rect 295944 220736 295950 220788
rect 306374 220736 306380 220788
rect 306432 220776 306438 220788
rect 320358 220776 320364 220788
rect 306432 220748 320364 220776
rect 306432 220736 306438 220748
rect 320358 220736 320364 220748
rect 320416 220736 320422 220788
rect 328822 220736 328828 220788
rect 328880 220776 328886 220788
rect 331950 220776 331956 220788
rect 328880 220748 331956 220776
rect 328880 220736 328886 220748
rect 331950 220736 331956 220748
rect 332008 220736 332014 220788
rect 414474 220736 414480 220788
rect 414532 220776 414538 220788
rect 418246 220776 418252 220788
rect 414532 220748 418252 220776
rect 414532 220736 414538 220748
rect 418246 220736 418252 220748
rect 418304 220736 418310 220788
rect 455230 220736 455236 220788
rect 455288 220776 455294 220788
rect 458542 220776 458548 220788
rect 455288 220748 458548 220776
rect 455288 220736 455294 220748
rect 458542 220736 458548 220748
rect 458600 220736 458606 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475102 220776 475108 220788
rect 474056 220748 475108 220776
rect 474056 220736 474062 220748
rect 475102 220736 475108 220748
rect 475160 220736 475166 220788
rect 475378 220736 475384 220788
rect 475436 220776 475442 220788
rect 476114 220776 476120 220788
rect 475436 220748 476120 220776
rect 475436 220736 475442 220748
rect 476114 220736 476120 220748
rect 476172 220736 476178 220788
rect 476850 220736 476856 220788
rect 476908 220776 476914 220788
rect 478414 220776 478420 220788
rect 476908 220748 478420 220776
rect 476908 220736 476914 220748
rect 478414 220736 478420 220748
rect 478472 220736 478478 220788
rect 592310 220736 592316 220788
rect 592368 220776 592374 220788
rect 601510 220776 601516 220788
rect 592368 220748 601516 220776
rect 592368 220736 592374 220748
rect 601510 220736 601516 220748
rect 601568 220736 601574 220788
rect 601694 220736 601700 220788
rect 601752 220776 601758 220788
rect 617518 220776 617524 220788
rect 601752 220748 617524 220776
rect 601752 220736 601758 220748
rect 617518 220736 617524 220748
rect 617576 220736 617582 220788
rect 108224 220680 108436 220708
rect 91554 220600 91560 220652
rect 91612 220640 91618 220652
rect 107930 220640 107936 220652
rect 91612 220612 107936 220640
rect 91612 220600 91618 220612
rect 107930 220600 107936 220612
rect 107988 220600 107994 220652
rect 108408 220640 108436 220680
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469306 220708 469312 220720
rect 465776 220680 469312 220708
rect 465776 220668 465782 220680
rect 469306 220668 469312 220680
rect 469364 220668 469370 220720
rect 172698 220640 172704 220652
rect 108408 220612 172704 220640
rect 172698 220600 172704 220612
rect 172756 220600 172762 220652
rect 177482 220600 177488 220652
rect 177540 220640 177546 220652
rect 182634 220640 182640 220652
rect 177540 220612 182640 220640
rect 177540 220600 177546 220612
rect 182634 220600 182640 220612
rect 182692 220600 182698 220652
rect 183462 220600 183468 220652
rect 183520 220640 183526 220652
rect 184198 220640 184204 220652
rect 183520 220612 184204 220640
rect 183520 220600 183526 220612
rect 184198 220600 184204 220612
rect 184256 220600 184262 220652
rect 184382 220600 184388 220652
rect 184440 220640 184446 220652
rect 234062 220640 234068 220652
rect 184440 220612 234068 220640
rect 184440 220600 184446 220612
rect 234062 220600 234068 220612
rect 234120 220600 234126 220652
rect 253842 220600 253848 220652
rect 253900 220640 253906 220652
rect 293402 220640 293408 220652
rect 253900 220612 293408 220640
rect 253900 220600 253906 220612
rect 293402 220600 293408 220612
rect 293460 220600 293466 220652
rect 296990 220600 296996 220652
rect 297048 220640 297054 220652
rect 310698 220640 310704 220652
rect 297048 220612 310704 220640
rect 297048 220600 297054 220612
rect 310698 220600 310704 220612
rect 310756 220600 310762 220652
rect 311710 220600 311716 220652
rect 311768 220640 311774 220652
rect 327258 220640 327264 220652
rect 311768 220612 327264 220640
rect 311768 220600 311774 220612
rect 327258 220600 327264 220612
rect 327316 220600 327322 220652
rect 508498 220600 508504 220652
rect 508556 220640 508562 220652
rect 522666 220640 522672 220652
rect 508556 220612 522672 220640
rect 508556 220600 508562 220612
rect 522666 220600 522672 220612
rect 522724 220600 522730 220652
rect 522850 220600 522856 220652
rect 522908 220640 522914 220652
rect 532878 220640 532884 220652
rect 522908 220612 532884 220640
rect 522908 220600 522914 220612
rect 532878 220600 532884 220612
rect 532936 220600 532942 220652
rect 533338 220600 533344 220652
rect 533396 220640 533402 220652
rect 618806 220640 618812 220652
rect 533396 220612 601556 220640
rect 533396 220600 533402 220612
rect 601528 220572 601556 220612
rect 601804 220612 618812 220640
rect 601804 220572 601832 220612
rect 618806 220600 618812 220612
rect 618864 220600 618870 220652
rect 601528 220544 601832 220572
rect 83274 220464 83280 220516
rect 83332 220504 83338 220516
rect 83332 220476 152504 220504
rect 83332 220464 83338 220476
rect 76650 220328 76656 220380
rect 76708 220368 76714 220380
rect 150618 220368 150624 220380
rect 76708 220340 150624 220368
rect 76708 220328 76714 220340
rect 150618 220328 150624 220340
rect 150676 220328 150682 220380
rect 152476 220368 152504 220476
rect 152642 220464 152648 220516
rect 152700 220504 152706 220516
rect 167178 220504 167184 220516
rect 152700 220476 167184 220504
rect 152700 220464 152706 220476
rect 167178 220464 167184 220476
rect 167236 220464 167242 220516
rect 171042 220464 171048 220516
rect 171100 220504 171106 220516
rect 229278 220504 229284 220516
rect 171100 220476 229284 220504
rect 171100 220464 171106 220476
rect 229278 220464 229284 220476
rect 229336 220464 229342 220516
rect 240594 220464 240600 220516
rect 240652 220504 240658 220516
rect 283006 220504 283012 220516
rect 240652 220476 283012 220504
rect 240652 220464 240658 220476
rect 283006 220464 283012 220476
rect 283064 220464 283070 220516
rect 296622 220464 296628 220516
rect 296680 220504 296686 220516
rect 327442 220504 327448 220516
rect 296680 220476 327448 220504
rect 296680 220464 296686 220476
rect 327442 220464 327448 220476
rect 327500 220464 327506 220516
rect 328178 220464 328184 220516
rect 328236 220504 328242 220516
rect 351362 220504 351368 220516
rect 328236 220476 351368 220504
rect 328236 220464 328242 220476
rect 351362 220464 351368 220476
rect 351420 220464 351426 220516
rect 371142 220464 371148 220516
rect 371200 220504 371206 220516
rect 385218 220504 385224 220516
rect 371200 220476 385224 220504
rect 371200 220464 371206 220476
rect 385218 220464 385224 220476
rect 385276 220464 385282 220516
rect 432230 220464 432236 220516
rect 432288 220504 432294 220516
rect 434806 220504 434812 220516
rect 432288 220476 434812 220504
rect 432288 220464 432294 220476
rect 434806 220464 434812 220476
rect 434864 220464 434870 220516
rect 496354 220464 496360 220516
rect 496412 220504 496418 220516
rect 496412 220476 507624 220504
rect 496412 220464 496418 220476
rect 157610 220368 157616 220380
rect 152476 220340 157616 220368
rect 157610 220328 157616 220340
rect 157668 220328 157674 220380
rect 157794 220328 157800 220380
rect 157852 220368 157858 220380
rect 218606 220368 218612 220380
rect 157852 220340 218612 220368
rect 157852 220328 157858 220340
rect 218606 220328 218612 220340
rect 218664 220328 218670 220380
rect 229186 220328 229192 220380
rect 229244 220368 229250 220380
rect 276106 220368 276112 220380
rect 229244 220340 276112 220368
rect 229244 220328 229250 220340
rect 276106 220328 276112 220340
rect 276164 220328 276170 220380
rect 281166 220328 281172 220380
rect 281224 220368 281230 220380
rect 317506 220368 317512 220380
rect 281224 220340 317512 220368
rect 281224 220328 281230 220340
rect 317506 220328 317512 220340
rect 317564 220328 317570 220380
rect 323394 220328 323400 220380
rect 323452 220368 323458 220380
rect 348142 220368 348148 220380
rect 323452 220340 348148 220368
rect 323452 220328 323458 220340
rect 348142 220328 348148 220340
rect 348200 220328 348206 220380
rect 353202 220328 353208 220380
rect 353260 220368 353266 220380
rect 371418 220368 371424 220380
rect 353260 220340 371424 220368
rect 353260 220328 353266 220340
rect 371418 220328 371424 220340
rect 371476 220328 371482 220380
rect 473262 220328 473268 220380
rect 473320 220368 473326 220380
rect 481726 220368 481732 220380
rect 473320 220340 481732 220368
rect 473320 220328 473326 220340
rect 481726 220328 481732 220340
rect 481784 220328 481790 220380
rect 482278 220328 482284 220380
rect 482336 220368 482342 220380
rect 491386 220368 491392 220380
rect 482336 220340 491392 220368
rect 482336 220328 482342 220340
rect 491386 220328 491392 220340
rect 491444 220328 491450 220380
rect 492582 220328 492588 220380
rect 492640 220368 492646 220380
rect 507394 220368 507400 220380
rect 492640 220340 507400 220368
rect 492640 220328 492646 220340
rect 507394 220328 507400 220340
rect 507452 220328 507458 220380
rect 66714 220192 66720 220244
rect 66772 220232 66778 220244
rect 147214 220232 147220 220244
rect 66772 220204 147220 220232
rect 66772 220192 66778 220204
rect 147214 220192 147220 220204
rect 147272 220192 147278 220244
rect 203242 220232 203248 220244
rect 147508 220204 203248 220232
rect 147508 220164 147536 220204
rect 203242 220192 203248 220204
rect 203300 220192 203306 220244
rect 211338 220232 211344 220244
rect 204916 220204 211344 220232
rect 147416 220136 147536 220164
rect 63402 220056 63408 220108
rect 63460 220096 63466 220108
rect 141050 220096 141056 220108
rect 63460 220068 141056 220096
rect 63460 220056 63466 220068
rect 141050 220056 141056 220068
rect 141108 220056 141114 220108
rect 141234 220056 141240 220108
rect 141292 220096 141298 220108
rect 147416 220096 147444 220136
rect 141292 220068 147444 220096
rect 141292 220056 141298 220068
rect 147628 220056 147634 220108
rect 147686 220096 147692 220108
rect 204916 220096 204944 220204
rect 211338 220192 211344 220204
rect 211396 220192 211402 220244
rect 211614 220192 211620 220244
rect 211672 220232 211678 220244
rect 263042 220232 263048 220244
rect 211672 220204 263048 220232
rect 211672 220192 211678 220204
rect 263042 220192 263048 220204
rect 263100 220192 263106 220244
rect 263318 220192 263324 220244
rect 263376 220232 263382 220244
rect 301038 220232 301044 220244
rect 263376 220204 301044 220232
rect 263376 220192 263382 220204
rect 301038 220192 301044 220204
rect 301096 220192 301102 220244
rect 318426 220192 318432 220244
rect 318484 220232 318490 220244
rect 343726 220232 343732 220244
rect 318484 220204 343732 220232
rect 318484 220192 318490 220204
rect 343726 220192 343732 220204
rect 343784 220192 343790 220244
rect 345842 220192 345848 220244
rect 345900 220232 345906 220244
rect 367370 220232 367376 220244
rect 345900 220204 367376 220232
rect 345900 220192 345906 220204
rect 367370 220192 367376 220204
rect 367428 220192 367434 220244
rect 368106 220192 368112 220244
rect 368164 220232 368170 220244
rect 382458 220232 382464 220244
rect 368164 220204 382464 220232
rect 368164 220192 368170 220204
rect 382458 220192 382464 220204
rect 382516 220192 382522 220244
rect 383010 220192 383016 220244
rect 383068 220232 383074 220244
rect 394786 220232 394792 220244
rect 383068 220204 394792 220232
rect 383068 220192 383074 220204
rect 394786 220192 394792 220204
rect 394844 220192 394850 220244
rect 397914 220192 397920 220244
rect 397972 220232 397978 220244
rect 405826 220232 405832 220244
rect 397972 220204 405832 220232
rect 397972 220192 397978 220204
rect 405826 220192 405832 220204
rect 405884 220192 405890 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465166 220232 465172 220244
rect 459520 220204 465172 220232
rect 459520 220192 459526 220204
rect 465166 220192 465172 220204
rect 465224 220192 465230 220244
rect 469030 220192 469036 220244
rect 469088 220232 469094 220244
rect 474274 220232 474280 220244
rect 469088 220204 474280 220232
rect 469088 220192 469094 220204
rect 474274 220192 474280 220204
rect 474332 220192 474338 220244
rect 478598 220192 478604 220244
rect 478656 220232 478662 220244
rect 489178 220232 489184 220244
rect 478656 220204 489184 220232
rect 478656 220192 478662 220204
rect 489178 220192 489184 220204
rect 489236 220192 489242 220244
rect 491202 220192 491208 220244
rect 491260 220232 491266 220244
rect 507596 220232 507624 220476
rect 515214 220464 515220 220516
rect 515272 220504 515278 220516
rect 601326 220504 601332 220516
rect 515272 220476 601332 220504
rect 515272 220464 515278 220476
rect 601326 220464 601332 220476
rect 601384 220464 601390 220516
rect 601970 220464 601976 220516
rect 602028 220504 602034 220516
rect 613286 220504 613292 220516
rect 602028 220476 613292 220504
rect 602028 220464 602034 220476
rect 613286 220464 613292 220476
rect 613344 220464 613350 220516
rect 507762 220328 507768 220380
rect 507820 220368 507826 220380
rect 527266 220368 527272 220380
rect 507820 220340 527272 220368
rect 507820 220328 507826 220340
rect 527266 220328 527272 220340
rect 527324 220328 527330 220380
rect 530026 220328 530032 220380
rect 530084 220368 530090 220380
rect 532694 220368 532700 220380
rect 530084 220340 532700 220368
rect 530084 220328 530090 220340
rect 532694 220328 532700 220340
rect 532752 220328 532758 220380
rect 532878 220328 532884 220380
rect 532936 220368 532942 220380
rect 534028 220368 534034 220380
rect 532936 220340 534034 220368
rect 532936 220328 532942 220340
rect 534028 220328 534034 220340
rect 534086 220328 534092 220380
rect 534166 220328 534172 220380
rect 534224 220368 534230 220380
rect 620462 220368 620468 220380
rect 534224 220340 620468 220368
rect 534224 220328 534230 220340
rect 620462 220328 620468 220340
rect 620520 220328 620526 220380
rect 510982 220232 510988 220244
rect 491260 220204 502380 220232
rect 507596 220204 510988 220232
rect 491260 220192 491266 220204
rect 244458 220096 244464 220108
rect 147686 220068 204944 220096
rect 205008 220068 244464 220096
rect 147686 220056 147692 220068
rect 111426 219920 111432 219972
rect 111484 219960 111490 219972
rect 177482 219960 177488 219972
rect 111484 219932 177488 219960
rect 111484 219920 111490 219932
rect 177482 219920 177488 219932
rect 177540 219920 177546 219972
rect 177666 219920 177672 219972
rect 177724 219960 177730 219972
rect 184382 219960 184388 219972
rect 177724 219932 184388 219960
rect 177724 219920 177730 219932
rect 184382 219920 184388 219932
rect 184440 219920 184446 219972
rect 190914 219920 190920 219972
rect 190972 219960 190978 219972
rect 205008 219960 205036 220068
rect 244458 220056 244464 220068
rect 244516 220056 244522 220108
rect 254670 220056 254676 220108
rect 254728 220096 254734 220108
rect 296806 220096 296812 220108
rect 254728 220068 296812 220096
rect 254728 220056 254734 220068
rect 296806 220056 296812 220068
rect 296864 220056 296870 220108
rect 300118 220056 300124 220108
rect 300176 220096 300182 220108
rect 330018 220096 330024 220108
rect 300176 220068 330024 220096
rect 300176 220056 300182 220068
rect 330018 220056 330024 220068
rect 330076 220056 330082 220108
rect 332502 220056 332508 220108
rect 332560 220096 332566 220108
rect 357526 220096 357532 220108
rect 332560 220068 357532 220096
rect 332560 220056 332566 220068
rect 357526 220056 357532 220068
rect 357584 220056 357590 220108
rect 360654 220056 360660 220108
rect 360712 220096 360718 220108
rect 377398 220096 377404 220108
rect 360712 220068 377404 220096
rect 360712 220056 360718 220068
rect 377398 220056 377404 220068
rect 377456 220056 377462 220108
rect 390462 220056 390468 220108
rect 390520 220096 390526 220108
rect 401686 220096 401692 220108
rect 390520 220068 401692 220096
rect 390520 220056 390526 220068
rect 401686 220056 401692 220068
rect 401744 220056 401750 220108
rect 421926 220056 421932 220108
rect 421984 220096 421990 220108
rect 426802 220096 426808 220108
rect 421984 220068 426808 220096
rect 421984 220056 421990 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 481542 220056 481548 220108
rect 481600 220096 481606 220108
rect 492766 220096 492772 220108
rect 481600 220068 492772 220096
rect 481600 220056 481606 220068
rect 492766 220056 492772 220068
rect 492824 220056 492830 220108
rect 502352 220096 502380 220204
rect 510982 220192 510988 220204
rect 511040 220232 511046 220244
rect 582742 220232 582748 220244
rect 511040 220204 582748 220232
rect 511040 220192 511046 220204
rect 582742 220192 582748 220204
rect 582800 220192 582806 220244
rect 582926 220192 582932 220244
rect 582984 220232 582990 220244
rect 591666 220232 591672 220244
rect 582984 220204 591672 220232
rect 582984 220192 582990 220204
rect 591666 220192 591672 220204
rect 591724 220192 591730 220244
rect 592494 220192 592500 220244
rect 592552 220232 592558 220244
rect 601510 220232 601516 220244
rect 592552 220204 601516 220232
rect 592552 220192 592558 220204
rect 601510 220192 601516 220204
rect 601568 220192 601574 220244
rect 601694 220192 601700 220244
rect 601752 220232 601758 220244
rect 612918 220232 612924 220244
rect 601752 220204 612924 220232
rect 601752 220192 601758 220204
rect 612918 220192 612924 220204
rect 612976 220192 612982 220244
rect 505186 220096 505192 220108
rect 502352 220068 505192 220096
rect 505186 220056 505192 220068
rect 505244 220056 505250 220108
rect 521562 220056 521568 220108
rect 521620 220096 521626 220108
rect 543366 220096 543372 220108
rect 521620 220068 543372 220096
rect 521620 220056 521626 220068
rect 543366 220056 543372 220068
rect 543424 220056 543430 220108
rect 548334 220096 548340 220108
rect 543660 220068 548340 220096
rect 543660 220028 543688 220068
rect 548334 220056 548340 220068
rect 548392 220056 548398 220108
rect 572622 220056 572628 220108
rect 572680 220096 572686 220108
rect 627086 220096 627092 220108
rect 572680 220068 627092 220096
rect 572680 220056 572686 220068
rect 627086 220056 627092 220068
rect 627144 220056 627150 220108
rect 647326 220056 647332 220108
rect 647384 220096 647390 220108
rect 652754 220096 652760 220108
rect 647384 220068 652760 220096
rect 647384 220056 647390 220068
rect 652754 220056 652760 220068
rect 652812 220056 652818 220108
rect 543568 220000 543688 220028
rect 249886 219960 249892 219972
rect 190972 219932 205036 219960
rect 205100 219932 249892 219960
rect 190972 219920 190978 219932
rect 124674 219784 124680 219836
rect 124732 219824 124738 219836
rect 193490 219824 193496 219836
rect 124732 219796 193496 219824
rect 124732 219784 124738 219796
rect 193490 219784 193496 219796
rect 193548 219784 193554 219836
rect 197262 219784 197268 219836
rect 197320 219824 197326 219836
rect 205100 219824 205128 219932
rect 249886 219920 249892 219932
rect 249944 219920 249950 219972
rect 280062 219920 280068 219972
rect 280120 219960 280126 219972
rect 313918 219960 313924 219972
rect 280120 219932 313924 219960
rect 280120 219920 280126 219932
rect 313918 219920 313924 219932
rect 313976 219920 313982 219972
rect 493778 219920 493784 219972
rect 493836 219960 493842 219972
rect 508222 219960 508228 219972
rect 493836 219932 508228 219960
rect 493836 219920 493842 219932
rect 508222 219920 508228 219932
rect 508280 219920 508286 219972
rect 522666 219920 522672 219972
rect 522724 219960 522730 219972
rect 533338 219960 533344 219972
rect 522724 219932 533344 219960
rect 522724 219920 522730 219932
rect 533338 219920 533344 219932
rect 533396 219920 533402 219972
rect 534074 219920 534080 219972
rect 534132 219960 534138 219972
rect 537294 219960 537300 219972
rect 534132 219932 537300 219960
rect 534132 219920 534138 219932
rect 537294 219920 537300 219932
rect 537352 219920 537358 219972
rect 537478 219852 537484 219904
rect 537536 219892 537542 219904
rect 543568 219892 543596 220000
rect 548518 219988 548524 220040
rect 548576 220028 548582 220040
rect 553854 220028 553860 220040
rect 548576 220000 553860 220028
rect 548576 219988 548582 220000
rect 553854 219988 553860 220000
rect 553912 219988 553918 220040
rect 554038 219988 554044 220040
rect 554096 220028 554102 220040
rect 562870 220028 562876 220040
rect 554096 220000 562876 220028
rect 554096 219988 554102 220000
rect 562870 219988 562876 220000
rect 562928 219988 562934 220040
rect 563238 219988 563244 220040
rect 563296 220028 563302 220040
rect 572070 220028 572076 220040
rect 563296 220000 572076 220028
rect 563296 219988 563302 220000
rect 572070 219988 572076 220000
rect 572128 219988 572134 220040
rect 592034 219920 592040 219972
rect 592092 219960 592098 219972
rect 592092 219932 598934 219960
rect 592092 219920 592098 219932
rect 537536 219864 543596 219892
rect 537536 219852 537542 219864
rect 543734 219852 543740 219904
rect 543792 219892 543798 219904
rect 572622 219892 572628 219904
rect 543792 219864 572628 219892
rect 543792 219852 543798 219864
rect 572622 219852 572628 219864
rect 572680 219852 572686 219904
rect 572806 219852 572812 219904
rect 572864 219892 572870 219904
rect 582190 219892 582196 219904
rect 572864 219864 582196 219892
rect 572864 219852 572870 219864
rect 582190 219852 582196 219864
rect 582248 219852 582254 219904
rect 582374 219852 582380 219904
rect 582432 219892 582438 219904
rect 591850 219892 591856 219904
rect 582432 219864 591856 219892
rect 582432 219852 582438 219864
rect 591850 219852 591856 219864
rect 591908 219852 591914 219904
rect 598906 219892 598934 219932
rect 621566 219892 621572 219904
rect 598906 219864 621572 219892
rect 621566 219852 621572 219864
rect 621624 219852 621630 219904
rect 197320 219796 205128 219824
rect 197320 219784 197326 219796
rect 207474 219784 207480 219836
rect 207532 219824 207538 219836
rect 257338 219824 257344 219836
rect 207532 219796 257344 219824
rect 207532 219784 207538 219796
rect 257338 219784 257344 219796
rect 257396 219784 257402 219836
rect 293862 219784 293868 219836
rect 293920 219824 293926 219836
rect 299934 219824 299940 219836
rect 293920 219796 299940 219824
rect 293920 219784 293926 219796
rect 299934 219784 299940 219796
rect 299992 219784 299998 219836
rect 504358 219784 504364 219836
rect 504416 219824 504422 219836
rect 515214 219824 515220 219836
rect 504416 219796 515220 219824
rect 504416 219784 504422 219796
rect 515214 219784 515220 219796
rect 515272 219784 515278 219836
rect 517422 219716 517428 219768
rect 517480 219756 517486 219768
rect 539042 219756 539048 219768
rect 517480 219728 539048 219756
rect 517480 219716 517486 219728
rect 539042 219716 539048 219728
rect 539100 219716 539106 219768
rect 540238 219716 540244 219768
rect 540296 219756 540302 219768
rect 548518 219756 548524 219768
rect 540296 219728 548524 219756
rect 540296 219716 540302 219728
rect 548518 219716 548524 219728
rect 548576 219716 548582 219768
rect 549898 219716 549904 219768
rect 549956 219756 549962 219768
rect 553210 219756 553216 219768
rect 549956 219728 553216 219756
rect 549956 219716 549962 219728
rect 553210 219716 553216 219728
rect 553268 219716 553274 219768
rect 553348 219716 553354 219768
rect 553406 219756 553412 219768
rect 570506 219756 570512 219768
rect 553406 219728 570512 219756
rect 553406 219716 553412 219728
rect 570506 219716 570512 219728
rect 570564 219716 570570 219768
rect 574830 219716 574836 219768
rect 574888 219756 574894 219768
rect 623774 219756 623780 219768
rect 574888 219728 623780 219756
rect 574888 219716 574894 219728
rect 623774 219716 623780 219728
rect 623832 219716 623838 219768
rect 137278 219648 137284 219700
rect 137336 219688 137342 219700
rect 152642 219688 152648 219700
rect 137336 219660 152648 219688
rect 137336 219648 137342 219660
rect 152642 219648 152648 219660
rect 152700 219648 152706 219700
rect 153102 219648 153108 219700
rect 153160 219688 153166 219700
rect 214098 219688 214104 219700
rect 153160 219660 214104 219688
rect 153160 219648 153166 219660
rect 214098 219648 214104 219660
rect 214156 219648 214162 219700
rect 217410 219648 217416 219700
rect 217468 219688 217474 219700
rect 265158 219688 265164 219700
rect 217468 219660 265164 219688
rect 217468 219648 217474 219660
rect 265158 219648 265164 219660
rect 265216 219648 265222 219700
rect 571076 219660 571840 219688
rect 273070 219580 273076 219632
rect 273128 219620 273134 219632
rect 279234 219620 279240 219632
rect 273128 219592 279240 219620
rect 273128 219580 273134 219592
rect 279234 219580 279240 219592
rect 279292 219580 279298 219632
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 471974 219620 471980 219632
rect 465040 219592 471980 219620
rect 465040 219580 465046 219592
rect 471974 219580 471980 219592
rect 472032 219580 472038 219632
rect 497274 219580 497280 219632
rect 497332 219620 497338 219632
rect 562870 219620 562876 219632
rect 497332 219592 562876 219620
rect 497332 219580 497338 219592
rect 562870 219580 562876 219592
rect 562928 219580 562934 219632
rect 563054 219580 563060 219632
rect 563112 219620 563118 219632
rect 571076 219620 571104 219660
rect 563112 219592 571104 219620
rect 571812 219620 571840 219660
rect 625430 219620 625436 219632
rect 571812 219592 625436 219620
rect 563112 219580 563118 219592
rect 625430 219580 625436 219592
rect 625488 219580 625494 219632
rect 131022 219512 131028 219564
rect 131080 219552 131086 219564
rect 137462 219552 137468 219564
rect 131080 219524 137468 219552
rect 131080 219512 131086 219524
rect 137462 219512 137468 219524
rect 137520 219512 137526 219564
rect 137922 219512 137928 219564
rect 137980 219552 137986 219564
rect 203058 219552 203064 219564
rect 137980 219524 203064 219552
rect 137980 219512 137986 219524
rect 203058 219512 203064 219524
rect 203116 219512 203122 219564
rect 203242 219512 203248 219564
rect 203300 219552 203306 219564
rect 205818 219552 205824 219564
rect 203300 219524 205824 219552
rect 203300 219512 203306 219524
rect 205818 219512 205824 219524
rect 205876 219512 205882 219564
rect 406194 219512 406200 219564
rect 406252 219552 406258 219564
rect 412726 219552 412732 219564
rect 406252 219524 412732 219552
rect 406252 219512 406258 219524
rect 412726 219512 412732 219524
rect 412784 219512 412790 219564
rect 432046 219552 432052 219564
rect 429212 219524 432052 219552
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 80790 219376 80796 219428
rect 80848 219416 80854 219428
rect 90358 219416 90364 219428
rect 80848 219388 90364 219416
rect 80848 219376 80854 219388
rect 90358 219376 90364 219388
rect 90416 219376 90422 219428
rect 90726 219376 90732 219428
rect 90784 219416 90790 219428
rect 106918 219416 106924 219428
rect 90784 219388 106924 219416
rect 90784 219376 90790 219388
rect 106918 219376 106924 219388
rect 106976 219376 106982 219428
rect 117866 219376 117872 219428
rect 117924 219416 117930 219428
rect 123478 219416 123484 219428
rect 117924 219388 123484 219416
rect 117924 219376 117930 219388
rect 123478 219376 123484 219388
rect 123536 219376 123542 219428
rect 132770 219376 132776 219428
rect 132828 219416 132834 219428
rect 140038 219416 140044 219428
rect 132828 219388 140044 219416
rect 132828 219376 132834 219388
rect 140038 219376 140044 219388
rect 140096 219376 140102 219428
rect 142798 219376 142804 219428
rect 142856 219416 142862 219428
rect 197998 219416 198004 219428
rect 142856 219388 198004 219416
rect 142856 219376 142862 219388
rect 197998 219376 198004 219388
rect 198056 219376 198062 219428
rect 199838 219376 199844 219428
rect 199896 219416 199902 219428
rect 204714 219416 204720 219428
rect 199896 219388 204720 219416
rect 199896 219376 199902 219388
rect 204714 219376 204720 219388
rect 204772 219376 204778 219428
rect 212994 219376 213000 219428
rect 213052 219416 213058 219428
rect 217226 219416 217232 219428
rect 213052 219388 217232 219416
rect 213052 219376 213058 219388
rect 217226 219376 217232 219388
rect 217284 219376 217290 219428
rect 217962 219376 217968 219428
rect 218020 219416 218026 219428
rect 220078 219416 220084 219428
rect 218020 219388 220084 219416
rect 218020 219376 218026 219388
rect 220078 219376 220084 219388
rect 220136 219376 220142 219428
rect 224034 219376 224040 219428
rect 224092 219416 224098 219428
rect 232498 219416 232504 219428
rect 224092 219388 232504 219416
rect 224092 219376 224098 219388
rect 232498 219376 232504 219388
rect 232556 219376 232562 219428
rect 232958 219376 232964 219428
rect 233016 219416 233022 219428
rect 233016 219388 243584 219416
rect 233016 219376 233022 219388
rect 93210 219240 93216 219292
rect 93268 219280 93274 219292
rect 93762 219280 93768 219292
rect 93268 219252 93768 219280
rect 93268 219240 93274 219252
rect 93762 219240 93768 219252
rect 93820 219240 93826 219292
rect 108298 219240 108304 219292
rect 108356 219280 108362 219292
rect 149974 219280 149980 219292
rect 108356 219252 149980 219280
rect 108356 219240 108362 219252
rect 149974 219240 149980 219252
rect 150032 219240 150038 219292
rect 150158 219240 150164 219292
rect 150216 219280 150222 219292
rect 161290 219280 161296 219292
rect 150216 219252 161296 219280
rect 150216 219240 150222 219252
rect 161290 219240 161296 219252
rect 161348 219240 161354 219292
rect 169018 219280 169024 219292
rect 162136 219252 169024 219280
rect 85298 219104 85304 219156
rect 85356 219144 85362 219156
rect 117866 219144 117872 219156
rect 85356 219116 117872 219144
rect 85356 219104 85362 219116
rect 117866 219104 117872 219116
rect 117924 219104 117930 219156
rect 123846 219104 123852 219156
rect 123904 219144 123910 219156
rect 127066 219144 127072 219156
rect 123904 219116 127072 219144
rect 123904 219104 123910 219116
rect 127066 219104 127072 219116
rect 127124 219104 127130 219156
rect 130470 219104 130476 219156
rect 130528 219144 130534 219156
rect 162136 219144 162164 219252
rect 169018 219240 169024 219252
rect 169076 219240 169082 219292
rect 169202 219240 169208 219292
rect 169260 219280 169266 219292
rect 169260 219252 181484 219280
rect 169260 219240 169266 219252
rect 130528 219116 162164 219144
rect 130528 219104 130534 219116
rect 162302 219104 162308 219156
rect 162360 219144 162366 219156
rect 180978 219144 180984 219156
rect 162360 219116 180984 219144
rect 162360 219104 162366 219116
rect 180978 219104 180984 219116
rect 181036 219104 181042 219156
rect 181456 219144 181484 219252
rect 182634 219240 182640 219292
rect 182692 219280 182698 219292
rect 183278 219280 183284 219292
rect 182692 219252 183284 219280
rect 182692 219240 182698 219252
rect 183278 219240 183284 219252
rect 183336 219240 183342 219292
rect 183646 219240 183652 219292
rect 183704 219280 183710 219292
rect 226978 219280 226984 219292
rect 183704 219252 226984 219280
rect 183704 219240 183710 219252
rect 226978 219240 226984 219252
rect 227036 219240 227042 219292
rect 238110 219240 238116 219292
rect 238168 219280 238174 219292
rect 239398 219280 239404 219292
rect 238168 219252 239404 219280
rect 238168 219240 238174 219252
rect 239398 219240 239404 219252
rect 239456 219240 239462 219292
rect 243556 219280 243584 219388
rect 246390 219376 246396 219428
rect 246448 219416 246454 219428
rect 286042 219416 286048 219428
rect 246448 219388 286048 219416
rect 246448 219376 246454 219388
rect 286042 219376 286048 219388
rect 286100 219376 286106 219428
rect 291654 219376 291660 219428
rect 291712 219416 291718 219428
rect 324682 219416 324688 219428
rect 291712 219388 324688 219416
rect 291712 219376 291718 219388
rect 324682 219376 324688 219388
rect 324740 219376 324746 219428
rect 345566 219416 345572 219428
rect 335326 219388 345572 219416
rect 273070 219280 273076 219292
rect 243556 219252 273076 219280
rect 273070 219240 273076 219252
rect 273128 219240 273134 219292
rect 325418 219240 325424 219292
rect 325476 219280 325482 219292
rect 326338 219280 326344 219292
rect 325476 219252 326344 219280
rect 325476 219240 325482 219252
rect 326338 219240 326344 219252
rect 326396 219240 326402 219292
rect 327534 219240 327540 219292
rect 327592 219280 327598 219292
rect 335326 219280 335354 219388
rect 345566 219376 345572 219388
rect 345624 219376 345630 219428
rect 352374 219376 352380 219428
rect 352432 219416 352438 219428
rect 352432 219388 358584 219416
rect 352432 219376 352438 219388
rect 327592 219252 335354 219280
rect 327592 219240 327598 219252
rect 344094 219240 344100 219292
rect 344152 219280 344158 219292
rect 347038 219280 347044 219292
rect 344152 219252 347044 219280
rect 344152 219240 344158 219252
rect 347038 219240 347044 219252
rect 347096 219240 347102 219292
rect 199378 219144 199384 219156
rect 181456 219116 199384 219144
rect 199378 219104 199384 219116
rect 199436 219104 199442 219156
rect 204714 219104 204720 219156
rect 204772 219144 204778 219156
rect 246206 219144 246212 219156
rect 204772 219116 246212 219144
rect 204772 219104 204778 219116
rect 246206 219104 246212 219116
rect 246264 219104 246270 219156
rect 262674 219104 262680 219156
rect 262732 219144 262738 219156
rect 291838 219144 291844 219156
rect 262732 219116 291844 219144
rect 262732 219104 262738 219116
rect 291838 219104 291844 219116
rect 291896 219104 291902 219156
rect 311710 219144 311716 219156
rect 296686 219116 311716 219144
rect 70854 218968 70860 219020
rect 70912 219008 70918 219020
rect 132770 219008 132776 219020
rect 70912 218980 132776 219008
rect 70912 218968 70918 218980
rect 132770 218968 132776 218980
rect 132828 218968 132834 219020
rect 132954 218968 132960 219020
rect 133012 219008 133018 219020
rect 133782 219008 133788 219020
rect 133012 218980 133788 219008
rect 133012 218968 133018 218980
rect 133782 218968 133788 218980
rect 133840 218968 133846 219020
rect 137094 218968 137100 219020
rect 137152 219008 137158 219020
rect 142798 219008 142804 219020
rect 137152 218980 142804 219008
rect 137152 218968 137158 218980
rect 142798 218968 142804 218980
rect 142856 218968 142862 219020
rect 143166 218968 143172 219020
rect 143224 219008 143230 219020
rect 143224 218980 152320 219008
rect 143224 218968 143230 218980
rect 62574 218832 62580 218884
rect 62632 218872 62638 218884
rect 76466 218872 76472 218884
rect 62632 218844 76472 218872
rect 62632 218832 62638 218844
rect 76466 218832 76472 218844
rect 76524 218832 76530 218884
rect 83918 218832 83924 218884
rect 83976 218872 83982 218884
rect 83976 218844 142936 218872
rect 83976 218832 83982 218844
rect 60090 218696 60096 218748
rect 60148 218736 60154 218748
rect 69658 218736 69664 218748
rect 60148 218708 69664 218736
rect 60148 218696 60154 218708
rect 69658 218696 69664 218708
rect 69716 218696 69722 218748
rect 77202 218696 77208 218748
rect 77260 218736 77266 218748
rect 142908 218736 142936 218844
rect 143626 218832 143632 218884
rect 143684 218872 143690 218884
rect 146202 218872 146208 218884
rect 143684 218844 146208 218872
rect 143684 218832 143690 218844
rect 146202 218832 146208 218844
rect 146260 218832 146266 218884
rect 152292 218872 152320 218980
rect 152458 218968 152464 219020
rect 152516 219008 152522 219020
rect 204898 219008 204904 219020
rect 152516 218980 204904 219008
rect 152516 218968 152522 218980
rect 204898 218968 204904 218980
rect 204956 218968 204962 219020
rect 206646 218968 206652 219020
rect 206704 219008 206710 219020
rect 255958 219008 255964 219020
rect 206704 218980 255964 219008
rect 206704 218968 206710 218980
rect 255958 218968 255964 218980
rect 256016 218968 256022 219020
rect 259086 218968 259092 219020
rect 259144 219008 259150 219020
rect 293862 219008 293868 219020
rect 259144 218980 293868 219008
rect 259144 218968 259150 218980
rect 293862 218968 293868 218980
rect 293920 218968 293926 219020
rect 294414 218968 294420 219020
rect 294472 219008 294478 219020
rect 296686 219008 296714 219116
rect 311710 219104 311716 219116
rect 311768 219104 311774 219156
rect 315666 219104 315672 219156
rect 315724 219144 315730 219156
rect 318058 219144 318064 219156
rect 315724 219116 318064 219144
rect 315724 219104 315730 219116
rect 318058 219104 318064 219116
rect 318116 219104 318122 219156
rect 320910 219104 320916 219156
rect 320968 219144 320974 219156
rect 340138 219144 340144 219156
rect 320968 219116 340144 219144
rect 320968 219104 320974 219116
rect 340138 219104 340144 219116
rect 340196 219104 340202 219156
rect 354398 219104 354404 219156
rect 354456 219144 354462 219156
rect 355502 219144 355508 219156
rect 354456 219116 355508 219144
rect 354456 219104 354462 219116
rect 355502 219104 355508 219116
rect 355560 219104 355566 219156
rect 358556 219144 358584 219388
rect 417786 219376 417792 219428
rect 417844 219416 417850 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 417844 219388 418200 219416
rect 417844 219376 417850 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 571168 219524 571748 219552
rect 437014 219484 437020 219496
rect 436480 219456 437020 219484
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 430206 219376 430212 219428
rect 430264 219416 430270 219428
rect 432690 219416 432696 219428
rect 430264 219388 432696 219416
rect 430264 219376 430270 219388
rect 432690 219376 432696 219388
rect 432748 219376 432754 219428
rect 435082 219376 435088 219428
rect 435140 219416 435146 219428
rect 436480 219416 436508 219456
rect 437014 219444 437020 219456
rect 437072 219444 437078 219496
rect 493962 219444 493968 219496
rect 494020 219484 494026 219496
rect 571168 219484 571196 219524
rect 494020 219456 497136 219484
rect 494020 219444 494026 219456
rect 435140 219388 436508 219416
rect 435140 219376 435146 219388
rect 497108 219348 497136 219456
rect 497798 219456 571196 219484
rect 571720 219484 571748 219524
rect 613102 219484 613108 219496
rect 571720 219456 613108 219484
rect 497798 219348 497826 219456
rect 613102 219444 613108 219456
rect 613160 219444 613166 219496
rect 613286 219444 613292 219496
rect 613344 219484 613350 219496
rect 628098 219484 628104 219496
rect 613344 219456 628104 219484
rect 613344 219444 613350 219456
rect 628098 219444 628104 219456
rect 628156 219444 628162 219496
rect 571260 219388 571656 219416
rect 497108 219320 497826 219348
rect 535454 219308 535460 219360
rect 535512 219348 535518 219360
rect 536374 219348 536380 219360
rect 535512 219320 536380 219348
rect 535512 219308 535518 219320
rect 536374 219308 536380 219320
rect 536432 219308 536438 219360
rect 537294 219308 537300 219360
rect 537352 219348 537358 219360
rect 539686 219348 539692 219360
rect 537352 219320 539692 219348
rect 537352 219308 537358 219320
rect 539686 219308 539692 219320
rect 539744 219308 539750 219360
rect 543366 219308 543372 219360
rect 543424 219348 543430 219360
rect 544286 219348 544292 219360
rect 543424 219320 544292 219348
rect 543424 219308 543430 219320
rect 544286 219308 544292 219320
rect 544344 219308 544350 219360
rect 562502 219348 562508 219360
rect 553780 219320 562508 219348
rect 358722 219240 358728 219292
rect 358780 219280 358786 219292
rect 364978 219280 364984 219292
rect 358780 219252 364984 219280
rect 358780 219240 358786 219252
rect 364978 219240 364984 219252
rect 365036 219240 365042 219292
rect 383562 219240 383568 219292
rect 383620 219280 383626 219292
rect 387058 219280 387064 219292
rect 383620 219252 387064 219280
rect 383620 219240 383626 219252
rect 387058 219240 387064 219252
rect 387116 219240 387122 219292
rect 475746 219240 475752 219292
rect 475804 219280 475810 219292
rect 482554 219280 482560 219292
rect 475804 219252 482560 219280
rect 475804 219240 475810 219252
rect 482554 219240 482560 219252
rect 482612 219240 482618 219292
rect 546310 219240 546316 219292
rect 546368 219280 546374 219292
rect 553486 219280 553492 219292
rect 546368 219252 553492 219280
rect 546368 219240 546374 219252
rect 553486 219240 553492 219252
rect 553544 219240 553550 219292
rect 513006 219172 513012 219224
rect 513064 219212 513070 219224
rect 519170 219212 519176 219224
rect 513064 219184 519176 219212
rect 513064 219172 513070 219184
rect 519170 219172 519176 219184
rect 519228 219172 519234 219224
rect 553780 219212 553808 219320
rect 562502 219308 562508 219320
rect 562560 219308 562566 219360
rect 562870 219308 562876 219360
rect 562928 219348 562934 219360
rect 563238 219348 563244 219360
rect 562928 219320 563244 219348
rect 562928 219308 562934 219320
rect 563238 219308 563244 219320
rect 563296 219308 563302 219360
rect 563422 219308 563428 219360
rect 563480 219348 563486 219360
rect 571260 219348 571288 219388
rect 563480 219320 571288 219348
rect 571628 219348 571656 219388
rect 573174 219348 573180 219360
rect 571628 219320 573180 219348
rect 563480 219308 563486 219320
rect 573174 219308 573180 219320
rect 573232 219308 573238 219360
rect 573450 219308 573456 219360
rect 573508 219348 573514 219360
rect 574830 219348 574836 219360
rect 573508 219320 574836 219348
rect 573508 219308 573514 219320
rect 574830 219308 574836 219320
rect 574888 219308 574894 219360
rect 582190 219308 582196 219360
rect 582248 219348 582254 219360
rect 582374 219348 582380 219360
rect 582248 219320 582380 219348
rect 582248 219308 582254 219320
rect 582374 219308 582380 219320
rect 582432 219308 582438 219360
rect 591850 219308 591856 219360
rect 591908 219348 591914 219360
rect 592310 219348 592316 219360
rect 591908 219320 592316 219348
rect 591908 219308 591914 219320
rect 592310 219308 592316 219320
rect 592368 219308 592374 219360
rect 553688 219184 553808 219212
rect 366266 219144 366272 219156
rect 358556 219116 366272 219144
rect 366266 219104 366272 219116
rect 366324 219104 366330 219156
rect 373074 219104 373080 219156
rect 373132 219144 373138 219156
rect 373810 219144 373816 219156
rect 373132 219116 373816 219144
rect 373132 219104 373138 219116
rect 373810 219104 373816 219116
rect 373868 219104 373874 219156
rect 407574 219104 407580 219156
rect 407632 219144 407638 219156
rect 411898 219144 411904 219156
rect 407632 219116 411904 219144
rect 407632 219104 407638 219116
rect 411898 219104 411904 219116
rect 411956 219104 411962 219156
rect 419258 219104 419264 219156
rect 419316 219144 419322 219156
rect 422662 219144 422668 219156
rect 419316 219116 422668 219144
rect 419316 219104 419322 219116
rect 422662 219104 422668 219116
rect 422720 219104 422726 219156
rect 507210 219104 507216 219156
rect 507268 219144 507274 219156
rect 509510 219144 509516 219156
rect 507268 219116 509516 219144
rect 507268 219104 507274 219116
rect 509510 219104 509516 219116
rect 509568 219104 509574 219156
rect 537110 219104 537116 219156
rect 537168 219144 537174 219156
rect 539226 219144 539232 219156
rect 537168 219116 539232 219144
rect 537168 219104 537174 219116
rect 539226 219104 539232 219116
rect 539284 219104 539290 219156
rect 543734 219104 543740 219156
rect 543792 219144 543798 219156
rect 553688 219144 553716 219184
rect 553946 219172 553952 219224
rect 554004 219212 554010 219224
rect 554004 219184 563468 219212
rect 554004 219172 554010 219184
rect 543792 219116 553716 219144
rect 543792 219104 543798 219116
rect 563440 219076 563468 219184
rect 563606 219172 563612 219224
rect 563664 219212 563670 219224
rect 570138 219212 570144 219224
rect 563664 219184 570144 219212
rect 563664 219172 563670 219184
rect 570138 219172 570144 219184
rect 570196 219172 570202 219224
rect 572346 219172 572352 219224
rect 572404 219212 572410 219224
rect 582926 219212 582932 219224
rect 572404 219184 582932 219212
rect 572404 219172 572410 219184
rect 582926 219172 582932 219184
rect 582984 219172 582990 219224
rect 591666 219172 591672 219224
rect 591724 219212 591730 219224
rect 592494 219212 592500 219224
rect 591724 219184 592500 219212
rect 591724 219172 591730 219184
rect 592494 219172 592500 219184
rect 592552 219172 592558 219224
rect 601510 219172 601516 219224
rect 601568 219212 601574 219224
rect 601694 219212 601700 219224
rect 601568 219184 601700 219212
rect 601568 219172 601574 219184
rect 601694 219172 601700 219184
rect 601752 219172 601758 219224
rect 571426 219144 571432 219156
rect 570340 219116 571432 219144
rect 570340 219076 570368 219116
rect 571426 219104 571432 219116
rect 571484 219104 571490 219156
rect 572346 219076 572352 219088
rect 563440 219048 570368 219076
rect 571628 219048 572352 219076
rect 294472 218980 296714 219008
rect 294472 218968 294478 218980
rect 300762 218968 300768 219020
rect 300820 219008 300826 219020
rect 328822 219008 328828 219020
rect 300820 218980 328828 219008
rect 300820 218968 300826 218980
rect 328822 218968 328828 218980
rect 328880 218968 328886 219020
rect 333698 218968 333704 219020
rect 333756 219008 333762 219020
rect 352558 219008 352564 219020
rect 333756 218980 352564 219008
rect 333756 218968 333762 218980
rect 352558 218968 352564 218980
rect 352616 218968 352622 219020
rect 355686 218968 355692 219020
rect 355744 219008 355750 219020
rect 369118 219008 369124 219020
rect 355744 218980 369124 219008
rect 355744 218968 355750 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 373718 218968 373724 219020
rect 373776 219008 373782 219020
rect 380158 219008 380164 219020
rect 373776 218980 380164 219008
rect 373776 218968 373782 218980
rect 380158 218968 380164 218980
rect 380216 218968 380222 219020
rect 384666 218968 384672 219020
rect 384724 219008 384730 219020
rect 393958 219008 393964 219020
rect 384724 218980 393964 219008
rect 384724 218968 384730 218980
rect 393958 218968 393964 218980
rect 394016 218968 394022 219020
rect 402054 218968 402060 219020
rect 402112 219008 402118 219020
rect 407758 219008 407764 219020
rect 402112 218980 407764 219008
rect 402112 218968 402118 218980
rect 407758 218968 407764 218980
rect 407816 218968 407822 219020
rect 460198 218968 460204 219020
rect 460256 219008 460262 219020
rect 461118 219008 461124 219020
rect 460256 218980 461124 219008
rect 460256 218968 460262 218980
rect 461118 218968 461124 218980
rect 461176 218968 461182 219020
rect 532142 218968 532148 219020
rect 532200 219008 532206 219020
rect 532602 219008 532608 219020
rect 532200 218980 532608 219008
rect 532200 218968 532206 218980
rect 532602 218968 532608 218980
rect 532660 219008 532666 219020
rect 538858 219008 538864 219020
rect 532660 218980 538864 219008
rect 532660 218968 532666 218980
rect 538858 218968 538864 218980
rect 538916 218968 538922 219020
rect 542446 218968 542452 219020
rect 542504 219008 542510 219020
rect 546586 219008 546592 219020
rect 542504 218980 546592 219008
rect 542504 218968 542510 218980
rect 546586 218968 546592 218980
rect 546644 218968 546650 219020
rect 546954 218968 546960 219020
rect 547012 219008 547018 219020
rect 552842 219008 552848 219020
rect 547012 218980 552848 219008
rect 547012 218968 547018 218980
rect 552842 218968 552848 218980
rect 552900 218968 552906 219020
rect 553486 218968 553492 219020
rect 553544 219008 553550 219020
rect 553544 218980 553992 219008
rect 553544 218968 553550 218980
rect 509510 218900 509516 218952
rect 509568 218940 509574 218952
rect 518710 218940 518716 218952
rect 509568 218912 518716 218940
rect 509568 218900 509574 218912
rect 518710 218900 518716 218912
rect 518768 218900 518774 218952
rect 531958 218940 531964 218952
rect 528526 218912 531964 218940
rect 162302 218872 162308 218884
rect 152292 218844 162308 218872
rect 162302 218832 162308 218844
rect 162360 218832 162366 218884
rect 162486 218832 162492 218884
rect 162544 218872 162550 218884
rect 215938 218872 215944 218884
rect 162544 218844 215944 218872
rect 162544 218832 162550 218844
rect 215938 218832 215944 218844
rect 215996 218832 216002 218884
rect 216306 218832 216312 218884
rect 216364 218872 216370 218884
rect 224034 218872 224040 218884
rect 216364 218844 224040 218872
rect 216364 218832 216370 218844
rect 224034 218832 224040 218844
rect 224092 218832 224098 218884
rect 225966 218832 225972 218884
rect 226024 218872 226030 218884
rect 226024 218844 264468 218872
rect 226024 218832 226030 218844
rect 149330 218736 149336 218748
rect 77260 218708 142844 218736
rect 142908 218708 149336 218736
rect 77260 218696 77266 218708
rect 93762 218560 93768 218612
rect 93820 218600 93826 218612
rect 140222 218600 140228 218612
rect 93820 218572 140228 218600
rect 93820 218560 93826 218572
rect 140222 218560 140228 218572
rect 140280 218560 140286 218612
rect 140406 218560 140412 218612
rect 140464 218600 140470 218612
rect 142614 218600 142620 218612
rect 140464 218572 142620 218600
rect 140464 218560 140470 218572
rect 142614 218560 142620 218572
rect 142672 218560 142678 218612
rect 142816 218600 142844 218708
rect 149330 218696 149336 218708
rect 149388 218696 149394 218748
rect 149514 218696 149520 218748
rect 149572 218736 149578 218748
rect 150342 218736 150348 218748
rect 149572 218708 150348 218736
rect 149572 218696 149578 218708
rect 150342 218696 150348 218708
rect 150400 218696 150406 218748
rect 156322 218736 156328 218748
rect 150544 218708 156328 218736
rect 148502 218600 148508 218612
rect 142816 218572 148508 218600
rect 148502 218560 148508 218572
rect 148560 218560 148566 218612
rect 149974 218560 149980 218612
rect 150032 218600 150038 218612
rect 150544 218600 150572 218708
rect 156322 218696 156328 218708
rect 156380 218696 156386 218748
rect 156966 218696 156972 218748
rect 157024 218736 157030 218748
rect 161934 218736 161940 218748
rect 157024 218708 161940 218736
rect 157024 218696 157030 218708
rect 161934 218696 161940 218708
rect 161992 218696 161998 218748
rect 213178 218736 213184 218748
rect 162136 218708 213184 218736
rect 150032 218572 150572 218600
rect 150032 218560 150038 218572
rect 151170 218560 151176 218612
rect 151228 218600 151234 218612
rect 153102 218600 153108 218612
rect 151228 218572 153108 218600
rect 151228 218560 151234 218572
rect 153102 218560 153108 218572
rect 153160 218560 153166 218612
rect 153654 218560 153660 218612
rect 153712 218600 153718 218612
rect 162136 218600 162164 218708
rect 213178 218696 213184 218708
rect 213236 218696 213242 218748
rect 219894 218696 219900 218748
rect 219952 218736 219958 218748
rect 264238 218736 264244 218748
rect 219952 218708 264244 218736
rect 219952 218696 219958 218708
rect 264238 218696 264244 218708
rect 264296 218696 264302 218748
rect 153712 218572 162164 218600
rect 153712 218560 153718 218572
rect 162302 218560 162308 218612
rect 162360 218600 162366 218612
rect 163958 218600 163964 218612
rect 162360 218572 163964 218600
rect 162360 218560 162366 218572
rect 163958 218560 163964 218572
rect 164016 218560 164022 218612
rect 165614 218560 165620 218612
rect 165672 218600 165678 218612
rect 166810 218600 166816 218612
rect 165672 218572 166816 218600
rect 165672 218560 165678 218572
rect 166810 218560 166816 218572
rect 166868 218560 166874 218612
rect 166994 218560 167000 218612
rect 167052 218600 167058 218612
rect 169202 218600 169208 218612
rect 167052 218572 169208 218600
rect 167052 218560 167058 218572
rect 169202 218560 169208 218572
rect 169260 218560 169266 218612
rect 170214 218560 170220 218612
rect 170272 218600 170278 218612
rect 180794 218600 180800 218612
rect 170272 218572 180800 218600
rect 170272 218560 170278 218572
rect 180794 218560 180800 218572
rect 180852 218560 180858 218612
rect 180978 218560 180984 218612
rect 181036 218600 181042 218612
rect 192478 218600 192484 218612
rect 181036 218572 192484 218600
rect 181036 218560 181042 218572
rect 192478 218560 192484 218572
rect 192536 218560 192542 218612
rect 193122 218560 193128 218612
rect 193180 218600 193186 218612
rect 243538 218600 243544 218612
rect 193180 218572 243544 218600
rect 193180 218560 193186 218572
rect 243538 218560 243544 218572
rect 243596 218560 243602 218612
rect 253014 218560 253020 218612
rect 253072 218600 253078 218612
rect 262674 218600 262680 218612
rect 253072 218572 262680 218600
rect 253072 218560 253078 218572
rect 262674 218560 262680 218572
rect 262732 218560 262738 218612
rect 264440 218600 264468 218844
rect 274542 218832 274548 218884
rect 274600 218872 274606 218884
rect 280798 218872 280804 218884
rect 274600 218844 280804 218872
rect 274600 218832 274606 218844
rect 280798 218832 280804 218844
rect 280856 218832 280862 218884
rect 280982 218832 280988 218884
rect 281040 218872 281046 218884
rect 312538 218872 312544 218884
rect 281040 218844 312544 218872
rect 281040 218832 281046 218844
rect 312538 218832 312544 218844
rect 312596 218832 312602 218884
rect 314286 218832 314292 218884
rect 314344 218872 314350 218884
rect 329006 218872 329012 218884
rect 314344 218844 329012 218872
rect 314344 218832 314350 218844
rect 329006 218832 329012 218844
rect 329064 218832 329070 218884
rect 337470 218832 337476 218884
rect 337528 218872 337534 218884
rect 358078 218872 358084 218884
rect 337528 218844 358084 218872
rect 337528 218832 337534 218844
rect 358078 218832 358084 218844
rect 358136 218832 358142 218884
rect 366726 218832 366732 218884
rect 366784 218872 366790 218884
rect 378686 218872 378692 218884
rect 366784 218844 378692 218872
rect 366784 218832 366790 218844
rect 378686 218832 378692 218844
rect 378744 218832 378750 218884
rect 386138 218832 386144 218884
rect 386196 218872 386202 218884
rect 396718 218872 396724 218884
rect 386196 218844 396724 218872
rect 386196 218832 386202 218844
rect 396718 218832 396724 218844
rect 396776 218832 396782 218884
rect 402698 218832 402704 218884
rect 402756 218872 402762 218884
rect 409138 218872 409144 218884
rect 402756 218844 409144 218872
rect 402756 218832 402762 218844
rect 409138 218832 409144 218844
rect 409196 218832 409202 218884
rect 411990 218832 411996 218884
rect 412048 218872 412054 218884
rect 412450 218872 412456 218884
rect 412048 218844 412456 218872
rect 412048 218832 412054 218844
rect 412450 218832 412456 218844
rect 412508 218832 412514 218884
rect 485038 218832 485044 218884
rect 485096 218872 485102 218884
rect 490650 218872 490656 218884
rect 485096 218844 490656 218872
rect 485096 218832 485102 218844
rect 490650 218832 490656 218844
rect 490708 218832 490714 218884
rect 266078 218696 266084 218748
rect 266136 218736 266142 218748
rect 302878 218736 302884 218748
rect 266136 218708 302884 218736
rect 266136 218696 266142 218708
rect 302878 218696 302884 218708
rect 302936 218696 302942 218748
rect 307478 218696 307484 218748
rect 307536 218736 307542 218748
rect 337102 218736 337108 218748
rect 307536 218708 337108 218736
rect 307536 218696 307542 218708
rect 337102 218696 337108 218708
rect 337160 218696 337166 218748
rect 340506 218696 340512 218748
rect 340564 218736 340570 218748
rect 360838 218736 360844 218748
rect 340564 218708 360844 218736
rect 340564 218696 340570 218708
rect 360838 218696 360844 218708
rect 360896 218696 360902 218748
rect 379146 218696 379152 218748
rect 379204 218736 379210 218748
rect 392118 218736 392124 218748
rect 379204 218708 392124 218736
rect 379204 218696 379210 218708
rect 392118 218696 392124 218708
rect 392176 218696 392182 218748
rect 395798 218696 395804 218748
rect 395856 218736 395862 218748
rect 404538 218736 404544 218748
rect 395856 218708 404544 218736
rect 395856 218696 395862 218708
rect 404538 218696 404544 218708
rect 404596 218696 404602 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 509234 218628 509240 218680
rect 509292 218668 509298 218680
rect 518848 218668 518854 218680
rect 509292 218640 518854 218668
rect 509292 218628 509298 218640
rect 518848 218628 518854 218640
rect 518906 218628 518912 218680
rect 527266 218628 527272 218680
rect 527324 218668 527330 218680
rect 528526 218668 528554 218912
rect 531958 218900 531964 218912
rect 532016 218900 532022 218952
rect 537846 218832 537852 218884
rect 537904 218872 537910 218884
rect 543918 218872 543924 218884
rect 537904 218844 543924 218872
rect 537904 218832 537910 218844
rect 543918 218832 543924 218844
rect 543976 218832 543982 218884
rect 544102 218832 544108 218884
rect 544160 218872 544166 218884
rect 553762 218872 553768 218884
rect 544160 218844 553768 218872
rect 544160 218832 544166 218844
rect 553762 218832 553768 218844
rect 553820 218832 553826 218884
rect 553964 218872 553992 218980
rect 554222 218968 554228 219020
rect 554280 219008 554286 219020
rect 554280 218980 563054 219008
rect 554280 218968 554286 218980
rect 563026 218940 563054 218980
rect 563026 218912 565814 218940
rect 562870 218872 562876 218884
rect 553964 218844 562876 218872
rect 562870 218832 562876 218844
rect 562928 218832 562934 218884
rect 565786 218872 565814 218912
rect 565786 218844 571288 218872
rect 528646 218764 528652 218816
rect 528704 218804 528710 218816
rect 534258 218804 534264 218816
rect 528704 218776 534264 218804
rect 528704 218764 528710 218776
rect 534258 218764 534264 218776
rect 534316 218764 534322 218816
rect 571260 218804 571288 218844
rect 571628 218804 571656 219048
rect 572346 219036 572352 219048
rect 572404 219036 572410 219088
rect 572990 219036 572996 219088
rect 573048 219076 573054 219088
rect 573048 219048 579614 219076
rect 573048 219036 573054 219048
rect 579586 219008 579614 219048
rect 579586 218980 582374 219008
rect 571794 218900 571800 218952
rect 571852 218940 571858 218952
rect 572530 218940 572536 218952
rect 571852 218912 572536 218940
rect 571852 218900 571858 218912
rect 572530 218900 572536 218912
rect 572588 218900 572594 218952
rect 573174 218900 573180 218952
rect 573232 218940 573238 218952
rect 575014 218940 575020 218952
rect 573232 218912 575020 218940
rect 573232 218900 573238 218912
rect 575014 218900 575020 218912
rect 575072 218900 575078 218952
rect 582346 218872 582374 218980
rect 605650 218872 605656 218884
rect 582346 218844 605656 218872
rect 605650 218832 605656 218844
rect 605708 218832 605714 218884
rect 571260 218776 571656 218804
rect 546954 218736 546960 218748
rect 527324 218640 528554 218668
rect 534460 218708 546960 218736
rect 527324 218628 527330 218640
rect 267734 218600 267740 218612
rect 264440 218572 267740 218600
rect 267734 218560 267740 218572
rect 267792 218560 267798 218612
rect 272886 218560 272892 218612
rect 272944 218600 272950 218612
rect 296990 218600 296996 218612
rect 272944 218572 296996 218600
rect 272944 218560 272950 218572
rect 296990 218560 296996 218572
rect 297048 218560 297054 218612
rect 351546 218560 351552 218612
rect 351604 218600 351610 218612
rect 355318 218600 355324 218612
rect 351604 218572 355324 218600
rect 351604 218560 351610 218572
rect 355318 218560 355324 218572
rect 355376 218560 355382 218612
rect 534460 218600 534488 218708
rect 546954 218696 546960 218708
rect 547012 218696 547018 218748
rect 547138 218696 547144 218748
rect 547196 218736 547202 218748
rect 552658 218736 552664 218748
rect 547196 218708 552664 218736
rect 547196 218696 547202 218708
rect 552658 218696 552664 218708
rect 552716 218696 552722 218748
rect 553256 218696 553262 218748
rect 553314 218736 553320 218748
rect 570322 218736 570328 218748
rect 553314 218708 570328 218736
rect 553314 218696 553320 218708
rect 570322 218696 570328 218708
rect 570380 218696 570386 218748
rect 575382 218696 575388 218748
rect 575440 218736 575446 218748
rect 597462 218736 597468 218748
rect 575440 218708 597468 218736
rect 575440 218696 575446 218708
rect 597462 218696 597468 218708
rect 597520 218696 597526 218748
rect 528664 218572 534488 218600
rect 469858 218492 469864 218544
rect 469916 218532 469922 218544
rect 470962 218532 470968 218544
rect 469916 218504 470968 218532
rect 469916 218492 469922 218504
rect 470962 218492 470968 218504
rect 471020 218492 471026 218544
rect 518710 218492 518716 218544
rect 518768 218532 518774 218544
rect 528664 218532 528692 218572
rect 538858 218560 538864 218612
rect 538916 218600 538922 218612
rect 538916 218572 571104 218600
rect 538916 218560 538922 218572
rect 518768 218504 528692 218532
rect 571076 218532 571104 218572
rect 571812 218572 572116 218600
rect 571812 218532 571840 218572
rect 571076 218504 571840 218532
rect 518768 218492 518774 218504
rect 100478 218424 100484 218476
rect 100536 218464 100542 218476
rect 108298 218464 108304 218476
rect 100536 218436 108304 218464
rect 100536 218424 100542 218436
rect 108298 218424 108304 218436
rect 108356 218424 108362 218476
rect 126330 218424 126336 218476
rect 126388 218464 126394 218476
rect 126882 218464 126888 218476
rect 126388 218436 126888 218464
rect 126388 218424 126394 218436
rect 126882 218424 126888 218436
rect 126940 218424 126946 218476
rect 127066 218424 127072 218476
rect 127124 218464 127130 218476
rect 174170 218464 174176 218476
rect 127124 218436 174176 218464
rect 127124 218424 127130 218436
rect 174170 218424 174176 218436
rect 174228 218424 174234 218476
rect 174354 218424 174360 218476
rect 174412 218464 174418 218476
rect 183646 218464 183652 218476
rect 174412 218436 183652 218464
rect 174412 218424 174418 218436
rect 183646 218424 183652 218436
rect 183704 218424 183710 218476
rect 186774 218424 186780 218476
rect 186832 218464 186838 218476
rect 235258 218464 235264 218476
rect 186832 218436 235264 218464
rect 186832 218424 186838 218436
rect 235258 218424 235264 218436
rect 235316 218424 235322 218476
rect 239766 218424 239772 218476
rect 239824 218464 239830 218476
rect 272518 218464 272524 218476
rect 239824 218436 272524 218464
rect 239824 218424 239830 218436
rect 272518 218424 272524 218436
rect 272576 218424 272582 218476
rect 279510 218424 279516 218476
rect 279568 218464 279574 218476
rect 280982 218464 280988 218476
rect 279568 218436 280988 218464
rect 279568 218424 279574 218436
rect 280982 218424 280988 218436
rect 281040 218424 281046 218476
rect 286134 218424 286140 218476
rect 286192 218464 286198 218476
rect 306374 218464 306380 218476
rect 286192 218436 306380 218464
rect 286192 218424 286198 218436
rect 306374 218424 306380 218436
rect 306432 218424 306438 218476
rect 380526 218424 380532 218476
rect 380584 218464 380590 218476
rect 384298 218464 384304 218476
rect 380584 218436 384304 218464
rect 380584 218424 380590 218436
rect 384298 218424 384304 218436
rect 384356 218424 384362 218476
rect 531958 218424 531964 218476
rect 532016 218464 532022 218476
rect 546310 218464 546316 218476
rect 532016 218436 533568 218464
rect 532016 218424 532022 218436
rect 450538 218356 450544 218408
rect 450596 218396 450602 218408
rect 453574 218396 453580 218408
rect 450596 218368 453580 218396
rect 450596 218356 450602 218368
rect 453574 218356 453580 218368
rect 453632 218356 453638 218408
rect 519078 218356 519084 218408
rect 519136 218396 519142 218408
rect 528554 218396 528560 218408
rect 519136 218368 528560 218396
rect 519136 218356 519142 218368
rect 528554 218356 528560 218368
rect 528612 218356 528618 218408
rect 75638 218288 75644 218340
rect 75696 218328 75702 218340
rect 83458 218328 83464 218340
rect 75696 218300 83464 218328
rect 75696 218288 75702 218300
rect 83458 218288 83464 218300
rect 83516 218288 83522 218340
rect 107286 218288 107292 218340
rect 107344 218328 107350 218340
rect 157978 218328 157984 218340
rect 107344 218300 157984 218328
rect 107344 218288 107350 218300
rect 157978 218288 157984 218300
rect 158036 218288 158042 218340
rect 161566 218328 161572 218340
rect 159652 218300 161572 218328
rect 56318 218152 56324 218204
rect 56376 218192 56382 218204
rect 62758 218192 62764 218204
rect 56376 218164 62764 218192
rect 56376 218152 56382 218164
rect 62758 218152 62764 218164
rect 62816 218152 62822 218204
rect 79778 218152 79784 218204
rect 79836 218192 79842 218204
rect 82078 218192 82084 218204
rect 79836 218164 82084 218192
rect 79836 218152 79842 218164
rect 82078 218152 82084 218164
rect 82136 218152 82142 218204
rect 113910 218152 113916 218204
rect 113968 218192 113974 218204
rect 159652 218192 159680 218300
rect 161566 218288 161572 218300
rect 161624 218288 161630 218340
rect 161934 218288 161940 218340
rect 161992 218328 161998 218340
rect 165154 218328 165160 218340
rect 161992 218300 165160 218328
rect 161992 218288 161998 218300
rect 165154 218288 165160 218300
rect 165212 218288 165218 218340
rect 212994 218328 213000 218340
rect 166828 218300 213000 218328
rect 166828 218204 166856 218300
rect 212994 218288 213000 218300
rect 213052 218288 213058 218340
rect 213270 218288 213276 218340
rect 213328 218328 213334 218340
rect 216674 218328 216680 218340
rect 213328 218300 216680 218328
rect 213328 218288 213334 218300
rect 216674 218288 216680 218300
rect 216732 218288 216738 218340
rect 224218 218328 224224 218340
rect 219406 218300 224224 218328
rect 113968 218164 159680 218192
rect 113968 218152 113974 218164
rect 159818 218152 159824 218204
rect 159876 218192 159882 218204
rect 162486 218192 162492 218204
rect 159876 218164 162492 218192
rect 159876 218152 159882 218164
rect 162486 218152 162492 218164
rect 162544 218152 162550 218204
rect 163590 218152 163596 218204
rect 163648 218192 163654 218204
rect 163648 218164 165936 218192
rect 163648 218152 163654 218164
rect 55950 218016 55956 218068
rect 56008 218056 56014 218068
rect 56502 218056 56508 218068
rect 56008 218028 56508 218056
rect 56008 218016 56014 218028
rect 56502 218016 56508 218028
rect 56560 218016 56566 218068
rect 58434 218016 58440 218068
rect 58492 218056 58498 218068
rect 61378 218056 61384 218068
rect 58492 218028 61384 218056
rect 58492 218016 58498 218028
rect 61378 218016 61384 218028
rect 61436 218016 61442 218068
rect 64230 218016 64236 218068
rect 64288 218056 64294 218068
rect 64782 218056 64788 218068
rect 64288 218028 64788 218056
rect 64288 218016 64294 218028
rect 64782 218016 64788 218028
rect 64840 218016 64846 218068
rect 72510 218016 72516 218068
rect 72568 218056 72574 218068
rect 73062 218056 73068 218068
rect 72568 218028 73068 218056
rect 72568 218016 72574 218028
rect 73062 218016 73068 218028
rect 73120 218016 73126 218068
rect 74994 218016 75000 218068
rect 75052 218056 75058 218068
rect 75822 218056 75828 218068
rect 75052 218028 75828 218056
rect 75052 218016 75058 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 79134 218016 79140 218068
rect 79192 218056 79198 218068
rect 79962 218056 79968 218068
rect 79192 218028 79968 218056
rect 79192 218016 79198 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 84930 218016 84936 218068
rect 84988 218056 84994 218068
rect 85482 218056 85488 218068
rect 84988 218028 85488 218056
rect 84988 218016 84994 218028
rect 85482 218016 85488 218028
rect 85540 218016 85546 218068
rect 87414 218016 87420 218068
rect 87472 218056 87478 218068
rect 88242 218056 88248 218068
rect 87472 218028 88248 218056
rect 87472 218016 87478 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 97350 218016 97356 218068
rect 97408 218056 97414 218068
rect 97902 218056 97908 218068
rect 97408 218028 97908 218056
rect 97408 218016 97414 218028
rect 97902 218016 97908 218028
rect 97960 218016 97966 218068
rect 99834 218016 99840 218068
rect 99892 218056 99898 218068
rect 100662 218056 100668 218068
rect 99892 218028 100668 218056
rect 99892 218016 99898 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 101490 218016 101496 218068
rect 101548 218056 101554 218068
rect 102042 218056 102048 218068
rect 101548 218028 102048 218056
rect 101548 218016 101554 218028
rect 102042 218016 102048 218028
rect 102100 218016 102106 218068
rect 103974 218016 103980 218068
rect 104032 218056 104038 218068
rect 104802 218056 104808 218068
rect 104032 218028 104808 218056
rect 104032 218016 104038 218028
rect 104802 218016 104808 218028
rect 104860 218016 104866 218068
rect 110322 218016 110328 218068
rect 110380 218056 110386 218068
rect 111058 218056 111064 218068
rect 110380 218028 111064 218056
rect 110380 218016 110386 218028
rect 111058 218016 111064 218028
rect 111116 218016 111122 218068
rect 112254 218016 112260 218068
rect 112312 218056 112318 218068
rect 112898 218056 112904 218068
rect 112312 218028 112904 218056
rect 112312 218016 112318 218028
rect 112898 218016 112904 218028
rect 112956 218016 112962 218068
rect 116394 218016 116400 218068
rect 116452 218056 116458 218068
rect 117222 218056 117228 218068
rect 116452 218028 117228 218056
rect 116452 218016 116458 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 120534 218016 120540 218068
rect 120592 218056 120598 218068
rect 120592 218028 159312 218056
rect 120592 218016 120598 218028
rect 159284 217920 159312 218028
rect 159450 218016 159456 218068
rect 159508 218056 159514 218068
rect 160002 218056 160008 218068
rect 159508 218028 160008 218056
rect 159508 218016 159514 218028
rect 160002 218016 160008 218028
rect 160060 218016 160066 218068
rect 165614 218056 165620 218068
rect 160204 218028 165620 218056
rect 160204 217920 160232 218028
rect 165614 218016 165620 218028
rect 165672 218016 165678 218068
rect 159284 217892 160232 217920
rect 165908 217920 165936 218164
rect 166810 218152 166816 218204
rect 166868 218152 166874 218204
rect 168098 218152 168104 218204
rect 168156 218192 168162 218204
rect 170858 218192 170864 218204
rect 168156 218164 170864 218192
rect 168156 218152 168162 218164
rect 170858 218152 170864 218164
rect 170916 218152 170922 218204
rect 171870 218152 171876 218204
rect 171928 218192 171934 218204
rect 171928 218164 175412 218192
rect 171928 218152 171934 218164
rect 166074 218084 166080 218136
rect 166132 218124 166138 218136
rect 166534 218124 166540 218136
rect 166132 218096 166540 218124
rect 166132 218084 166138 218096
rect 166534 218084 166540 218096
rect 166592 218084 166598 218136
rect 166994 218016 167000 218068
rect 167052 218016 167058 218068
rect 167730 218016 167736 218068
rect 167788 218056 167794 218068
rect 168282 218056 168288 218068
rect 167788 218028 168288 218056
rect 167788 218016 167794 218028
rect 168282 218016 168288 218028
rect 168340 218016 168346 218068
rect 173526 218016 173532 218068
rect 173584 218056 173590 218068
rect 174170 218056 174176 218068
rect 173584 218028 174176 218056
rect 173584 218016 173590 218028
rect 174170 218016 174176 218028
rect 174228 218016 174234 218068
rect 174354 218016 174360 218068
rect 174412 218056 174418 218068
rect 175182 218056 175188 218068
rect 174412 218028 175188 218056
rect 174412 218016 174418 218028
rect 175182 218016 175188 218028
rect 175240 218016 175246 218068
rect 175384 218056 175412 218164
rect 176010 218152 176016 218204
rect 176068 218192 176074 218204
rect 176470 218192 176476 218204
rect 176068 218164 176476 218192
rect 176068 218152 176074 218164
rect 176470 218152 176476 218164
rect 176528 218152 176534 218204
rect 180150 218152 180156 218204
rect 180208 218192 180214 218204
rect 219406 218192 219434 218300
rect 224218 218288 224224 218300
rect 224276 218288 224282 218340
rect 228174 218288 228180 218340
rect 228232 218328 228238 218340
rect 229186 218328 229192 218340
rect 228232 218300 229192 218328
rect 228232 218288 228238 218300
rect 229186 218288 229192 218300
rect 229244 218288 229250 218340
rect 365622 218288 365628 218340
rect 365680 218328 365686 218340
rect 373258 218328 373264 218340
rect 365680 218300 373264 218328
rect 365680 218288 365686 218300
rect 373258 218288 373264 218300
rect 373316 218288 373322 218340
rect 426802 218288 426808 218340
rect 426860 218328 426866 218340
rect 429378 218328 429384 218340
rect 426860 218300 429384 218328
rect 426860 218288 426866 218300
rect 429378 218288 429384 218300
rect 429436 218288 429442 218340
rect 435910 218288 435916 218340
rect 435968 218328 435974 218340
rect 436278 218328 436284 218340
rect 435968 218300 436284 218328
rect 435968 218288 435974 218300
rect 436278 218288 436284 218300
rect 436336 218288 436342 218340
rect 479518 218288 479524 218340
rect 479576 218328 479582 218340
rect 480346 218328 480352 218340
rect 479576 218300 480352 218328
rect 479576 218288 479582 218300
rect 480346 218288 480352 218300
rect 480404 218288 480410 218340
rect 533338 218328 533344 218340
rect 532160 218300 533344 218328
rect 180208 218164 219434 218192
rect 180208 218152 180214 218164
rect 224034 218152 224040 218204
rect 224092 218192 224098 218204
rect 224678 218192 224684 218204
rect 224092 218164 224684 218192
rect 224092 218152 224098 218164
rect 224678 218152 224684 218164
rect 224736 218152 224742 218204
rect 224862 218152 224868 218204
rect 224920 218192 224926 218204
rect 225506 218192 225512 218204
rect 224920 218164 225512 218192
rect 224920 218152 224926 218164
rect 225506 218152 225512 218164
rect 225564 218152 225570 218204
rect 225690 218152 225696 218204
rect 225748 218192 225754 218204
rect 226150 218192 226156 218204
rect 225748 218164 226156 218192
rect 225748 218152 225754 218164
rect 226150 218152 226156 218164
rect 226208 218152 226214 218204
rect 229830 218152 229836 218204
rect 229888 218192 229894 218204
rect 231118 218192 231124 218204
rect 229888 218164 231124 218192
rect 229888 218152 229894 218164
rect 231118 218152 231124 218164
rect 231176 218152 231182 218204
rect 232314 218152 232320 218204
rect 232372 218192 232378 218204
rect 233142 218192 233148 218204
rect 232372 218164 233148 218192
rect 232372 218152 232378 218164
rect 233142 218152 233148 218164
rect 233200 218152 233206 218204
rect 233970 218152 233976 218204
rect 234028 218192 234034 218204
rect 234522 218192 234528 218204
rect 234028 218164 234528 218192
rect 234028 218152 234034 218164
rect 234522 218152 234528 218164
rect 234580 218152 234586 218204
rect 236454 218152 236460 218204
rect 236512 218192 236518 218204
rect 237006 218192 237012 218204
rect 236512 218164 237012 218192
rect 236512 218152 236518 218164
rect 237006 218152 237012 218164
rect 237064 218152 237070 218204
rect 249058 218192 249064 218204
rect 238726 218164 249064 218192
rect 176286 218056 176292 218068
rect 175384 218028 176292 218056
rect 176286 218016 176292 218028
rect 176344 218016 176350 218068
rect 176562 218016 176568 218068
rect 176620 218056 176626 218068
rect 177850 218056 177856 218068
rect 176620 218028 177856 218056
rect 176620 218016 176626 218028
rect 177850 218016 177856 218028
rect 177908 218016 177914 218068
rect 180794 218016 180800 218068
rect 180852 218056 180858 218068
rect 182082 218056 182088 218068
rect 180852 218028 182088 218056
rect 180852 218016 180858 218028
rect 182082 218016 182088 218028
rect 182140 218016 182146 218068
rect 194870 218016 194876 218068
rect 194928 218056 194934 218068
rect 195882 218056 195888 218068
rect 194928 218028 195888 218056
rect 194928 218016 194934 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 198918 218016 198924 218068
rect 198976 218056 198982 218068
rect 200022 218056 200028 218068
rect 198976 218028 200028 218056
rect 198976 218016 198982 218028
rect 200022 218016 200028 218028
rect 200080 218016 200086 218068
rect 200850 218016 200856 218068
rect 200908 218056 200914 218068
rect 201402 218056 201408 218068
rect 200908 218028 201408 218056
rect 200908 218016 200914 218028
rect 201402 218016 201408 218028
rect 201460 218016 201466 218068
rect 203334 218016 203340 218068
rect 203392 218056 203398 218068
rect 203886 218056 203892 218068
rect 203392 218028 203892 218056
rect 203392 218016 203398 218028
rect 203886 218016 203892 218028
rect 203944 218016 203950 218068
rect 204990 218016 204996 218068
rect 205048 218056 205054 218068
rect 206002 218056 206008 218068
rect 205048 218028 206008 218056
rect 205048 218016 205054 218028
rect 206002 218016 206008 218028
rect 206060 218016 206066 218068
rect 209130 218016 209136 218068
rect 209188 218056 209194 218068
rect 209682 218056 209688 218068
rect 209188 218028 209688 218056
rect 209188 218016 209194 218028
rect 209682 218016 209688 218028
rect 209740 218016 209746 218068
rect 215754 218016 215760 218068
rect 215812 218056 215818 218068
rect 216490 218056 216496 218068
rect 215812 218028 216496 218056
rect 215812 218016 215818 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 216674 218016 216680 218068
rect 216732 218056 216738 218068
rect 238726 218056 238754 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 249518 218152 249524 218204
rect 249576 218192 249582 218204
rect 251818 218192 251824 218204
rect 249576 218164 251824 218192
rect 249576 218152 249582 218164
rect 251818 218152 251824 218164
rect 251876 218152 251882 218204
rect 302694 218152 302700 218204
rect 302752 218192 302758 218204
rect 304718 218192 304724 218204
rect 302752 218164 304724 218192
rect 302752 218152 302758 218164
rect 304718 218152 304724 218164
rect 304776 218152 304782 218204
rect 310974 218152 310980 218204
rect 311032 218192 311038 218204
rect 315298 218192 315304 218204
rect 311032 218164 315304 218192
rect 311032 218152 311038 218164
rect 315298 218152 315304 218164
rect 315356 218152 315362 218204
rect 348878 218152 348884 218204
rect 348936 218192 348942 218204
rect 351178 218192 351184 218204
rect 348936 218164 351184 218192
rect 348936 218152 348942 218164
rect 351178 218152 351184 218164
rect 351236 218152 351242 218204
rect 364794 218152 364800 218204
rect 364852 218192 364858 218204
rect 367738 218192 367744 218204
rect 364852 218164 367744 218192
rect 364852 218152 364858 218164
rect 367738 218152 367744 218164
rect 367796 218152 367802 218204
rect 368934 218152 368940 218204
rect 368992 218192 368998 218204
rect 369762 218192 369768 218204
rect 368992 218164 369768 218192
rect 368992 218152 368998 218164
rect 369762 218152 369768 218164
rect 369820 218152 369826 218204
rect 377214 218152 377220 218204
rect 377272 218192 377278 218204
rect 382826 218192 382832 218204
rect 377272 218164 382832 218192
rect 377272 218152 377278 218164
rect 382826 218152 382832 218164
rect 382884 218152 382890 218204
rect 394418 218152 394424 218204
rect 394476 218192 394482 218204
rect 402238 218192 402244 218204
rect 394476 218164 402244 218192
rect 394476 218152 394482 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 422754 218152 422760 218204
rect 422812 218192 422818 218204
rect 425422 218192 425428 218204
rect 422812 218164 425428 218192
rect 422812 218152 422818 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 426066 218152 426072 218204
rect 426124 218192 426130 218204
rect 427906 218192 427912 218204
rect 426124 218164 427912 218192
rect 426124 218152 426130 218164
rect 427906 218152 427912 218164
rect 427964 218152 427970 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 455046 218152 455052 218204
rect 455104 218192 455110 218204
rect 460198 218192 460204 218204
rect 455104 218164 460204 218192
rect 455104 218152 455110 218164
rect 460198 218152 460204 218164
rect 460256 218152 460262 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 465994 218192 466000 218204
rect 462004 218164 466000 218192
rect 462004 218152 462010 218164
rect 465994 218152 466000 218164
rect 466052 218152 466058 218204
rect 509878 218152 509884 218204
rect 509936 218192 509942 218204
rect 510522 218192 510528 218204
rect 509936 218164 510528 218192
rect 509936 218152 509942 218164
rect 510522 218152 510528 218164
rect 510580 218192 510586 218204
rect 532160 218192 532188 218300
rect 533338 218288 533344 218300
rect 533396 218288 533402 218340
rect 533540 218328 533568 218436
rect 534046 218436 546316 218464
rect 534046 218328 534074 218436
rect 546310 218424 546316 218436
rect 546368 218424 546374 218476
rect 546586 218424 546592 218476
rect 546644 218464 546650 218476
rect 563192 218464 563198 218476
rect 546644 218436 563198 218464
rect 546644 218424 546650 218436
rect 563192 218424 563198 218436
rect 563250 218424 563256 218476
rect 572088 218464 572116 218572
rect 572530 218560 572536 218612
rect 572588 218600 572594 218612
rect 584398 218600 584404 218612
rect 572588 218572 584404 218600
rect 572588 218560 572594 218572
rect 584398 218560 584404 218572
rect 584456 218560 584462 218612
rect 573082 218464 573088 218476
rect 572088 218436 573088 218464
rect 573082 218424 573088 218436
rect 573140 218424 573146 218476
rect 574646 218424 574652 218476
rect 574704 218464 574710 218476
rect 575658 218464 575664 218476
rect 574704 218436 575664 218464
rect 574704 218424 574710 218436
rect 575658 218424 575664 218436
rect 575716 218424 575722 218476
rect 582098 218424 582104 218476
rect 582156 218464 582162 218476
rect 582742 218464 582748 218476
rect 582156 218436 582748 218464
rect 582156 218424 582162 218436
rect 582742 218424 582748 218436
rect 582800 218424 582806 218476
rect 570874 218396 570880 218408
rect 563440 218368 570880 218396
rect 533540 218300 534074 218328
rect 534166 218288 534172 218340
rect 534224 218328 534230 218340
rect 534224 218300 538904 218328
rect 534224 218288 534230 218300
rect 538876 218192 538904 218300
rect 539226 218288 539232 218340
rect 539284 218328 539290 218340
rect 563440 218328 563468 218368
rect 570874 218356 570880 218368
rect 570932 218356 570938 218408
rect 571058 218356 571064 218408
rect 571116 218396 571122 218408
rect 571116 218368 572024 218396
rect 571116 218356 571122 218368
rect 539284 218300 563468 218328
rect 571996 218328 572024 218368
rect 601418 218356 601424 218408
rect 601476 218396 601482 218408
rect 607490 218396 607496 218408
rect 601476 218368 607496 218396
rect 601476 218356 601482 218368
rect 607490 218356 607496 218368
rect 607548 218356 607554 218408
rect 573726 218328 573732 218340
rect 571996 218300 573732 218328
rect 539284 218288 539290 218300
rect 573726 218288 573732 218300
rect 573784 218288 573790 218340
rect 573910 218288 573916 218340
rect 573968 218328 573974 218340
rect 577682 218328 577688 218340
rect 573968 218300 577688 218328
rect 573968 218288 573974 218300
rect 577682 218288 577688 218300
rect 577740 218288 577746 218340
rect 578234 218288 578240 218340
rect 578292 218328 578298 218340
rect 582558 218328 582564 218340
rect 578292 218300 582564 218328
rect 578292 218288 578298 218300
rect 582558 218288 582564 218300
rect 582616 218288 582622 218340
rect 592126 218288 592132 218340
rect 592184 218328 592190 218340
rect 597738 218328 597744 218340
rect 592184 218300 597744 218328
rect 592184 218288 592190 218300
rect 597738 218288 597744 218300
rect 597796 218288 597802 218340
rect 563606 218220 563612 218272
rect 563664 218260 563670 218272
rect 564526 218260 564532 218272
rect 563664 218232 564532 218260
rect 563664 218220 563670 218232
rect 564526 218220 564532 218232
rect 564584 218220 564590 218272
rect 564802 218220 564808 218272
rect 564860 218260 564866 218272
rect 571794 218260 571800 218272
rect 564860 218232 571800 218260
rect 564860 218220 564866 218232
rect 571794 218220 571800 218232
rect 571852 218220 571858 218272
rect 543918 218192 543924 218204
rect 510580 218164 532188 218192
rect 532252 218164 538076 218192
rect 538876 218164 543924 218192
rect 510580 218152 510586 218164
rect 216732 218028 238754 218056
rect 216732 218016 216738 218028
rect 242250 218016 242256 218068
rect 242308 218056 242314 218068
rect 242710 218056 242716 218068
rect 242308 218028 242716 218056
rect 242308 218016 242314 218028
rect 242710 218016 242716 218028
rect 242768 218016 242774 218068
rect 244734 218016 244740 218068
rect 244792 218056 244798 218068
rect 247678 218056 247684 218068
rect 244792 218028 247684 218056
rect 244792 218016 244798 218028
rect 247678 218016 247684 218028
rect 247736 218016 247742 218068
rect 248874 218016 248880 218068
rect 248932 218056 248938 218068
rect 249702 218056 249708 218068
rect 248932 218028 249708 218056
rect 248932 218016 248938 218028
rect 249702 218016 249708 218028
rect 249760 218016 249766 218068
rect 250530 218016 250536 218068
rect 250588 218056 250594 218068
rect 251082 218056 251088 218068
rect 250588 218028 251088 218056
rect 250588 218016 250594 218028
rect 251082 218016 251088 218028
rect 251140 218016 251146 218068
rect 258810 218016 258816 218068
rect 258868 218056 258874 218068
rect 259270 218056 259276 218068
rect 258868 218028 259276 218056
rect 258868 218016 258874 218028
rect 259270 218016 259276 218028
rect 259328 218016 259334 218068
rect 262950 218016 262956 218068
rect 263008 218056 263014 218068
rect 263502 218056 263508 218068
rect 263008 218028 263508 218056
rect 263008 218016 263014 218028
rect 263502 218016 263508 218028
rect 263560 218016 263566 218068
rect 265434 218016 265440 218068
rect 265492 218056 265498 218068
rect 266262 218056 266268 218068
rect 265492 218028 266268 218056
rect 265492 218016 265498 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 267090 218016 267096 218068
rect 267148 218056 267154 218068
rect 267550 218056 267556 218068
rect 267148 218028 267556 218056
rect 267148 218016 267154 218028
rect 267550 218016 267556 218028
rect 267608 218016 267614 218068
rect 269574 218016 269580 218068
rect 269632 218056 269638 218068
rect 273898 218056 273904 218068
rect 269632 218028 273904 218056
rect 269632 218016 269638 218028
rect 273898 218016 273904 218028
rect 273956 218016 273962 218068
rect 277854 218016 277860 218068
rect 277912 218056 277918 218068
rect 278406 218056 278412 218068
rect 277912 218028 278412 218056
rect 277912 218016 277918 218028
rect 278406 218016 278412 218028
rect 278464 218016 278470 218068
rect 281994 218016 282000 218068
rect 282052 218056 282058 218068
rect 282638 218056 282644 218068
rect 282052 218028 282644 218056
rect 282052 218016 282058 218028
rect 282638 218016 282644 218028
rect 282696 218016 282702 218068
rect 283650 218016 283656 218068
rect 283708 218056 283714 218068
rect 284110 218056 284116 218068
rect 283708 218028 284116 218056
rect 283708 218016 283714 218028
rect 284110 218016 284116 218028
rect 284168 218016 284174 218068
rect 287790 218016 287796 218068
rect 287848 218056 287854 218068
rect 288250 218056 288256 218068
rect 287848 218028 288256 218056
rect 287848 218016 287854 218028
rect 288250 218016 288256 218028
rect 288308 218016 288314 218068
rect 298554 218016 298560 218068
rect 298612 218056 298618 218068
rect 299198 218056 299204 218068
rect 298612 218028 299204 218056
rect 298612 218016 298618 218028
rect 299198 218016 299204 218028
rect 299256 218016 299262 218068
rect 299382 218016 299388 218068
rect 299440 218056 299446 218068
rect 300302 218056 300308 218068
rect 299440 218028 300308 218056
rect 299440 218016 299446 218028
rect 300302 218016 300308 218028
rect 300360 218016 300366 218068
rect 304350 218016 304356 218068
rect 304408 218056 304414 218068
rect 305638 218056 305644 218068
rect 304408 218028 305644 218056
rect 304408 218016 304414 218028
rect 305638 218016 305644 218028
rect 305696 218016 305702 218068
rect 306834 218016 306840 218068
rect 306892 218056 306898 218068
rect 307662 218056 307668 218068
rect 306892 218028 307668 218056
rect 306892 218016 306898 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 312630 218016 312636 218068
rect 312688 218056 312694 218068
rect 314562 218056 314568 218068
rect 312688 218028 314568 218056
rect 312688 218016 312694 218028
rect 314562 218016 314568 218028
rect 314620 218016 314626 218068
rect 315114 218016 315120 218068
rect 315172 218056 315178 218068
rect 315850 218056 315856 218068
rect 315172 218028 315856 218056
rect 315172 218016 315178 218028
rect 315850 218016 315856 218028
rect 315908 218016 315914 218068
rect 319254 218016 319260 218068
rect 319312 218056 319318 218068
rect 319990 218056 319996 218068
rect 319312 218028 319996 218056
rect 319312 218016 319318 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 325050 218016 325056 218068
rect 325108 218056 325114 218068
rect 325602 218056 325608 218068
rect 325108 218028 325608 218056
rect 325108 218016 325114 218028
rect 325602 218016 325608 218028
rect 325660 218016 325666 218068
rect 329190 218016 329196 218068
rect 329248 218056 329254 218068
rect 330478 218056 330484 218068
rect 329248 218028 330484 218056
rect 329248 218016 329254 218028
rect 330478 218016 330484 218028
rect 330536 218016 330542 218068
rect 330846 218016 330852 218068
rect 330904 218056 330910 218068
rect 333146 218056 333152 218068
rect 330904 218028 333152 218056
rect 330904 218016 330910 218028
rect 333146 218016 333152 218028
rect 333204 218016 333210 218068
rect 333330 218016 333336 218068
rect 333388 218056 333394 218068
rect 333882 218056 333888 218068
rect 333388 218028 333888 218056
rect 333388 218016 333394 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 335814 218016 335820 218068
rect 335872 218056 335878 218068
rect 336458 218056 336464 218068
rect 335872 218028 336464 218056
rect 335872 218016 335878 218028
rect 336458 218016 336464 218028
rect 336516 218016 336522 218068
rect 339954 218016 339960 218068
rect 340012 218056 340018 218068
rect 340690 218056 340696 218068
rect 340012 218028 340696 218056
rect 340012 218016 340018 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 348234 218016 348240 218068
rect 348292 218056 348298 218068
rect 349062 218056 349068 218068
rect 348292 218028 349068 218056
rect 348292 218016 348298 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 354030 218016 354036 218068
rect 354088 218056 354094 218068
rect 354582 218056 354588 218068
rect 354088 218028 354588 218056
rect 354088 218016 354094 218028
rect 354582 218016 354588 218028
rect 354640 218016 354646 218068
rect 356514 218016 356520 218068
rect 356572 218056 356578 218068
rect 357342 218056 357348 218068
rect 356572 218028 357348 218056
rect 356572 218016 356578 218028
rect 357342 218016 357348 218028
rect 357400 218016 357406 218068
rect 358170 218016 358176 218068
rect 358228 218056 358234 218068
rect 359458 218056 359464 218068
rect 358228 218028 359464 218056
rect 358228 218016 358234 218028
rect 359458 218016 359464 218028
rect 359516 218016 359522 218068
rect 366450 218016 366456 218068
rect 366508 218056 366514 218068
rect 366910 218056 366916 218068
rect 366508 218028 366916 218056
rect 366508 218016 366514 218028
rect 366910 218016 366916 218028
rect 366968 218016 366974 218068
rect 369762 218016 369768 218068
rect 369820 218056 369826 218068
rect 370498 218056 370504 218068
rect 369820 218028 370504 218056
rect 369820 218016 369826 218028
rect 370498 218016 370504 218028
rect 370556 218016 370562 218068
rect 374730 218016 374736 218068
rect 374788 218056 374794 218068
rect 375282 218056 375288 218068
rect 374788 218028 375288 218056
rect 374788 218016 374794 218028
rect 375282 218016 375288 218028
rect 375340 218016 375346 218068
rect 378870 218016 378876 218068
rect 378928 218056 378934 218068
rect 379330 218056 379336 218068
rect 378928 218028 379336 218056
rect 378928 218016 378934 218028
rect 379330 218016 379336 218028
rect 379388 218016 379394 218068
rect 381354 218016 381360 218068
rect 381412 218056 381418 218068
rect 381906 218056 381912 218068
rect 381412 218028 381912 218056
rect 381412 218016 381418 218028
rect 381906 218016 381912 218028
rect 381964 218016 381970 218068
rect 385494 218016 385500 218068
rect 385552 218056 385558 218068
rect 386322 218056 386328 218068
rect 385552 218028 386328 218056
rect 385552 218016 385558 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 387150 218016 387156 218068
rect 387208 218056 387214 218068
rect 388438 218056 388444 218068
rect 387208 218028 388444 218056
rect 387208 218016 387214 218028
rect 388438 218016 388444 218028
rect 388496 218016 388502 218068
rect 389634 218016 389640 218068
rect 389692 218056 389698 218068
rect 390278 218056 390284 218068
rect 389692 218028 390284 218056
rect 389692 218016 389698 218028
rect 390278 218016 390284 218028
rect 390336 218016 390342 218068
rect 393774 218016 393780 218068
rect 393832 218056 393838 218068
rect 394602 218056 394608 218068
rect 393832 218028 394608 218056
rect 393832 218016 393838 218028
rect 394602 218016 394608 218028
rect 394660 218016 394666 218068
rect 395430 218016 395436 218068
rect 395488 218056 395494 218068
rect 395982 218056 395988 218068
rect 395488 218028 395988 218056
rect 395488 218016 395494 218028
rect 395982 218016 395988 218028
rect 396040 218016 396046 218068
rect 399570 218016 399576 218068
rect 399628 218056 399634 218068
rect 400030 218056 400036 218068
rect 399628 218028 400036 218056
rect 399628 218016 399634 218028
rect 400030 218016 400036 218028
rect 400088 218016 400094 218068
rect 403526 218016 403532 218068
rect 403584 218056 403590 218068
rect 404262 218056 404268 218068
rect 403584 218028 404268 218056
rect 403584 218016 403590 218028
rect 404262 218016 404268 218028
rect 404320 218016 404326 218068
rect 410334 218016 410340 218068
rect 410392 218056 410398 218068
rect 410886 218056 410892 218068
rect 410392 218028 410892 218056
rect 410392 218016 410398 218028
rect 410886 218016 410892 218028
rect 410944 218016 410950 218068
rect 416130 218016 416136 218068
rect 416188 218056 416194 218068
rect 416682 218056 416688 218068
rect 416188 218028 416688 218056
rect 416188 218016 416194 218028
rect 416682 218016 416688 218028
rect 416740 218016 416746 218068
rect 418614 218016 418620 218068
rect 418672 218056 418678 218068
rect 419442 218056 419448 218068
rect 418672 218028 419448 218056
rect 418672 218016 418678 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 420270 218016 420276 218068
rect 420328 218056 420334 218068
rect 420822 218056 420828 218068
rect 420328 218028 420828 218056
rect 420328 218016 420334 218028
rect 420822 218016 420828 218028
rect 420880 218016 420886 218068
rect 424410 218016 424416 218068
rect 424468 218056 424474 218068
rect 426986 218056 426992 218068
rect 424468 218028 426992 218056
rect 424468 218016 424474 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427722 218016 427728 218068
rect 427780 218056 427786 218068
rect 428458 218056 428464 218068
rect 427780 218028 428464 218056
rect 427780 218016 427786 218028
rect 428458 218016 428464 218028
rect 428516 218016 428522 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430666 218056 430672 218068
rect 429160 218028 430672 218056
rect 429160 218016 429166 218028
rect 430666 218016 430672 218028
rect 430724 218016 430730 218068
rect 432690 218016 432696 218068
rect 432748 218056 432754 218068
rect 433794 218056 433800 218068
rect 432748 218028 433800 218056
rect 432748 218016 432754 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 436830 218016 436836 218068
rect 436888 218056 436894 218068
rect 437474 218056 437480 218068
rect 436888 218028 437480 218056
rect 436888 218016 436894 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438486 218016 438492 218068
rect 438544 218056 438550 218068
rect 438946 218056 438952 218068
rect 438544 218028 438952 218056
rect 438544 218016 438550 218028
rect 438946 218016 438952 218028
rect 439004 218016 439010 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 462958 218016 462964 218068
rect 463016 218056 463022 218068
rect 464430 218056 464436 218068
rect 463016 218028 464436 218056
rect 463016 218016 463022 218028
rect 464430 218016 464436 218028
rect 464488 218016 464494 218068
rect 467098 218016 467104 218068
rect 467156 218056 467162 218068
rect 467834 218056 467840 218068
rect 467156 218028 467840 218056
rect 467156 218016 467162 218028
rect 467834 218016 467840 218028
rect 467892 218016 467898 218068
rect 471698 218016 471704 218068
rect 471756 218056 471762 218068
rect 472618 218056 472624 218068
rect 471756 218028 472624 218056
rect 471756 218016 471762 218028
rect 472618 218016 472624 218028
rect 472676 218016 472682 218068
rect 482830 218016 482836 218068
rect 482888 218056 482894 218068
rect 485038 218056 485044 218068
rect 482888 218028 485044 218056
rect 482888 218016 482894 218028
rect 485038 218016 485044 218028
rect 485096 218016 485102 218068
rect 491386 218016 491392 218068
rect 491444 218056 491450 218068
rect 492306 218056 492312 218068
rect 491444 218028 492312 218056
rect 491444 218016 491450 218028
rect 492306 218016 492312 218028
rect 492364 218056 492370 218068
rect 505094 218056 505100 218068
rect 492364 218028 505100 218056
rect 492364 218016 492370 218028
rect 505094 218016 505100 218028
rect 505152 218016 505158 218068
rect 525242 218016 525248 218068
rect 525300 218056 525306 218068
rect 532252 218056 532280 218164
rect 525300 218028 532280 218056
rect 525300 218016 525306 218028
rect 533338 218016 533344 218068
rect 533396 218056 533402 218068
rect 537846 218056 537852 218068
rect 533396 218028 537852 218056
rect 533396 218016 533402 218028
rect 537846 218016 537852 218028
rect 537904 218016 537910 218068
rect 538048 218056 538076 218164
rect 543918 218152 543924 218164
rect 543976 218152 543982 218204
rect 575014 218152 575020 218204
rect 575072 218192 575078 218204
rect 616138 218192 616144 218204
rect 575072 218164 616144 218192
rect 575072 218152 575078 218164
rect 616138 218152 616144 218164
rect 616196 218152 616202 218204
rect 544102 218084 544108 218136
rect 544160 218124 544166 218136
rect 554222 218124 554228 218136
rect 544160 218096 554228 218124
rect 544160 218084 544166 218096
rect 554222 218084 554228 218096
rect 554280 218084 554286 218136
rect 572898 218124 572904 218136
rect 555344 218096 572904 218124
rect 543688 218056 543694 218068
rect 538048 218028 543694 218056
rect 543688 218016 543694 218028
rect 543746 218016 543752 218068
rect 167012 217920 167040 218016
rect 543826 217948 543832 218000
rect 543884 217988 543890 218000
rect 555344 217988 555372 218096
rect 572898 218084 572904 218096
rect 572956 218084 572962 218136
rect 573100 218096 574876 218124
rect 543884 217960 555372 217988
rect 543884 217948 543890 217960
rect 555694 217948 555700 218000
rect 555752 217988 555758 218000
rect 563606 217988 563612 218000
rect 555752 217960 563612 217988
rect 555752 217948 555758 217960
rect 563606 217948 563612 217960
rect 563664 217948 563670 218000
rect 563790 217948 563796 218000
rect 563848 217988 563854 218000
rect 573100 217988 573128 218096
rect 563848 217960 573128 217988
rect 563848 217948 563854 217960
rect 573266 217948 573272 218000
rect 573324 217988 573330 218000
rect 574646 217988 574652 218000
rect 573324 217960 574652 217988
rect 573324 217948 573330 217960
rect 574646 217948 574652 217960
rect 574704 217948 574710 218000
rect 574848 217988 574876 218096
rect 676398 218084 676404 218136
rect 676456 218124 676462 218136
rect 677594 218124 677600 218136
rect 676456 218096 677600 218124
rect 676456 218084 676462 218096
rect 677594 218084 677600 218096
rect 677652 218084 677658 218136
rect 577682 218016 577688 218068
rect 577740 218056 577746 218068
rect 629386 218056 629392 218068
rect 577740 218028 629392 218056
rect 577740 218016 577746 218028
rect 629386 218016 629392 218028
rect 629444 218016 629450 218068
rect 577314 217988 577320 218000
rect 574848 217960 577320 217988
rect 577314 217948 577320 217960
rect 577372 217948 577378 218000
rect 165908 217892 167040 217920
rect 447134 217812 447140 217864
rect 447192 217852 447198 217864
rect 447778 217852 447784 217864
rect 447192 217824 447784 217852
rect 447192 217812 447198 217824
rect 447778 217812 447784 217824
rect 447836 217812 447842 217864
rect 448606 217812 448612 217864
rect 448664 217852 448670 217864
rect 449434 217852 449440 217864
rect 448664 217824 449440 217852
rect 448664 217812 448670 217824
rect 449434 217812 449440 217824
rect 449492 217812 449498 217864
rect 498194 217812 498200 217864
rect 498252 217852 498258 217864
rect 499114 217852 499120 217864
rect 498252 217824 499120 217852
rect 498252 217812 498258 217824
rect 499114 217812 499120 217824
rect 499172 217812 499178 217864
rect 543182 217812 543188 217864
rect 543240 217852 543246 217864
rect 543240 217824 548564 217852
rect 543240 217812 543246 217824
rect 508038 217744 508044 217796
rect 508096 217784 508102 217796
rect 509510 217784 509516 217796
rect 508096 217756 509516 217784
rect 508096 217744 508102 217756
rect 509510 217744 509516 217756
rect 509568 217744 509574 217796
rect 523770 217744 523776 217796
rect 523828 217784 523834 217796
rect 529106 217784 529112 217796
rect 523828 217756 529112 217784
rect 523828 217744 523834 217756
rect 529106 217744 529112 217756
rect 529164 217744 529170 217796
rect 544102 217716 544108 217728
rect 535288 217688 544108 217716
rect 509418 217540 509424 217592
rect 509476 217580 509482 217592
rect 519170 217580 519176 217592
rect 509476 217552 519176 217580
rect 509476 217540 509482 217552
rect 519170 217540 519176 217552
rect 519228 217540 519234 217592
rect 528278 217540 528284 217592
rect 528336 217580 528342 217592
rect 528336 217552 528554 217580
rect 528336 217540 528342 217552
rect 528526 217376 528554 217552
rect 528646 217540 528652 217592
rect 528704 217580 528710 217592
rect 534258 217580 534264 217592
rect 528704 217552 534264 217580
rect 528704 217540 528710 217552
rect 534258 217540 534264 217552
rect 534316 217540 534322 217592
rect 535288 217376 535316 217688
rect 544102 217676 544108 217688
rect 544160 217676 544166 217728
rect 548536 217716 548564 217824
rect 548886 217812 548892 217864
rect 548944 217852 548950 217864
rect 601510 217852 601516 217864
rect 548944 217824 601516 217852
rect 548944 217812 548950 217824
rect 601510 217812 601516 217824
rect 601568 217812 601574 217864
rect 601970 217812 601976 217864
rect 602028 217852 602034 217864
rect 609146 217852 609152 217864
rect 602028 217824 609152 217852
rect 602028 217812 602034 217824
rect 609146 217812 609152 217824
rect 609204 217812 609210 217864
rect 676674 217812 676680 217864
rect 676732 217852 676738 217864
rect 677042 217852 677048 217864
rect 676732 217824 677048 217852
rect 676732 217812 676738 217824
rect 677042 217812 677048 217824
rect 677100 217812 677106 217864
rect 592126 217716 592132 217728
rect 548536 217688 592132 217716
rect 592126 217676 592132 217688
rect 592184 217676 592190 217728
rect 592310 217676 592316 217728
rect 592368 217716 592374 217728
rect 594242 217716 594248 217728
rect 592368 217688 594248 217716
rect 592368 217676 592374 217688
rect 594242 217676 594248 217688
rect 594300 217676 594306 217728
rect 594426 217676 594432 217728
rect 594484 217716 594490 217728
rect 601326 217716 601332 217728
rect 594484 217688 601332 217716
rect 594484 217676 594490 217688
rect 601326 217676 601332 217688
rect 601384 217676 601390 217728
rect 601694 217676 601700 217728
rect 601752 217716 601758 217728
rect 605834 217716 605840 217728
rect 601752 217688 605840 217716
rect 601752 217676 601758 217688
rect 605834 217676 605840 217688
rect 605892 217676 605898 217728
rect 606202 217676 606208 217728
rect 606260 217716 606266 217728
rect 615678 217716 615684 217728
rect 606260 217688 615684 217716
rect 606260 217676 606266 217688
rect 615678 217676 615684 217688
rect 615736 217676 615742 217728
rect 543458 217540 543464 217592
rect 543516 217580 543522 217592
rect 543826 217580 543832 217592
rect 543516 217552 543832 217580
rect 543516 217540 543522 217552
rect 543826 217540 543832 217552
rect 543884 217540 543890 217592
rect 545758 217540 545764 217592
rect 545816 217580 545822 217592
rect 563790 217580 563796 217592
rect 545816 217552 563796 217580
rect 545816 217540 545822 217552
rect 563790 217540 563796 217552
rect 563848 217540 563854 217592
rect 564526 217540 564532 217592
rect 564584 217580 564590 217592
rect 572254 217580 572260 217592
rect 564584 217552 572260 217580
rect 564584 217540 564590 217552
rect 572254 217540 572260 217552
rect 572312 217540 572318 217592
rect 572806 217540 572812 217592
rect 572864 217580 572870 217592
rect 575382 217580 575388 217592
rect 572864 217552 575388 217580
rect 572864 217540 572870 217552
rect 575382 217540 575388 217552
rect 575440 217540 575446 217592
rect 575658 217540 575664 217592
rect 575716 217580 575722 217592
rect 601648 217580 601654 217592
rect 575716 217552 601654 217580
rect 575716 217540 575722 217552
rect 601648 217540 601654 217552
rect 601706 217540 601712 217592
rect 601786 217540 601792 217592
rect 601844 217580 601850 217592
rect 607306 217580 607312 217592
rect 601844 217552 607312 217580
rect 601844 217540 601850 217552
rect 607306 217540 607312 217552
rect 607364 217540 607370 217592
rect 538490 217404 538496 217456
rect 538548 217444 538554 217456
rect 594426 217444 594432 217456
rect 538548 217416 594432 217444
rect 538548 217404 538554 217416
rect 594426 217404 594432 217416
rect 594484 217404 594490 217456
rect 594610 217404 594616 217456
rect 594668 217444 594674 217456
rect 603994 217444 604000 217456
rect 594668 217416 604000 217444
rect 594668 217404 594674 217416
rect 603994 217404 604000 217416
rect 604052 217404 604058 217456
rect 605650 217404 605656 217456
rect 605708 217444 605714 217456
rect 627914 217444 627920 217456
rect 605708 217416 627920 217444
rect 605708 217404 605714 217416
rect 627914 217404 627920 217416
rect 627972 217404 627978 217456
rect 528526 217348 535316 217376
rect 601510 217308 601516 217320
rect 543706 217280 601516 217308
rect 146708 217200 146714 217252
rect 146766 217240 146772 217252
rect 152458 217240 152464 217252
rect 146766 217212 152464 217240
rect 146766 217200 146772 217212
rect 152458 217200 152464 217212
rect 152516 217200 152522 217252
rect 525932 217200 525938 217252
rect 525990 217240 525996 217252
rect 526530 217240 526536 217252
rect 525990 217212 526536 217240
rect 525990 217200 525996 217212
rect 526530 217200 526536 217212
rect 526588 217240 526594 217252
rect 526588 217212 533384 217240
rect 526588 217200 526594 217212
rect 519078 217064 519084 217116
rect 519136 217104 519142 217116
rect 528462 217104 528468 217116
rect 519136 217076 528468 217104
rect 519136 217064 519142 217076
rect 528462 217064 528468 217076
rect 528520 217064 528526 217116
rect 533356 216968 533384 217212
rect 536006 217200 536012 217252
rect 536064 217240 536070 217252
rect 543706 217240 543734 217280
rect 601510 217268 601516 217280
rect 601568 217268 601574 217320
rect 601694 217308 601700 217320
rect 601666 217268 601700 217308
rect 601752 217268 601758 217320
rect 536064 217212 543734 217240
rect 536064 217200 536070 217212
rect 594610 217172 594616 217184
rect 582346 217144 594616 217172
rect 533706 217064 533712 217116
rect 533764 217104 533770 217116
rect 582346 217104 582374 217144
rect 594610 217132 594616 217144
rect 594668 217132 594674 217184
rect 594794 217132 594800 217184
rect 594852 217172 594858 217184
rect 594852 217144 595392 217172
rect 594852 217132 594858 217144
rect 533764 217076 582374 217104
rect 533764 217064 533770 217076
rect 592126 216996 592132 217048
rect 592184 217036 592190 217048
rect 595162 217036 595168 217048
rect 592184 217008 595168 217036
rect 592184 216996 592190 217008
rect 595162 216996 595168 217008
rect 595220 216996 595226 217048
rect 572990 216968 572996 216980
rect 533356 216940 572996 216968
rect 572990 216928 572996 216940
rect 573048 216928 573054 216980
rect 575566 216968 575572 216980
rect 573284 216940 575572 216968
rect 528554 216792 528560 216844
rect 528612 216832 528618 216844
rect 573284 216832 573312 216940
rect 575566 216928 575572 216940
rect 575624 216928 575630 216980
rect 577314 216928 577320 216980
rect 577372 216968 577378 216980
rect 591942 216968 591948 216980
rect 577372 216940 591948 216968
rect 577372 216928 577378 216940
rect 591942 216928 591948 216940
rect 592000 216928 592006 216980
rect 595364 216968 595392 217144
rect 596634 217064 596640 217116
rect 596692 217104 596698 217116
rect 601666 217104 601694 217268
rect 601970 217200 601976 217252
rect 602028 217240 602034 217252
rect 606202 217240 606208 217252
rect 602028 217212 606208 217240
rect 602028 217200 602034 217212
rect 606202 217200 606208 217212
rect 606260 217200 606266 217252
rect 596692 217076 601694 217104
rect 596692 217064 596698 217076
rect 601786 217064 601792 217116
rect 601844 217104 601850 217116
rect 603074 217104 603080 217116
rect 601844 217076 603080 217104
rect 601844 217064 601850 217076
rect 603074 217064 603080 217076
rect 603132 217064 603138 217116
rect 603258 217064 603264 217116
rect 603316 217104 603322 217116
rect 610618 217104 610624 217116
rect 603316 217076 610624 217104
rect 603316 217064 603322 217076
rect 610618 217064 610624 217076
rect 610676 217064 610682 217116
rect 601142 216968 601148 216980
rect 595364 216940 601148 216968
rect 601142 216928 601148 216940
rect 601200 216928 601206 216980
rect 601510 216928 601516 216980
rect 601568 216968 601574 216980
rect 625246 216968 625252 216980
rect 601568 216940 625252 216968
rect 601568 216928 601574 216940
rect 625246 216928 625252 216940
rect 625304 216928 625310 216980
rect 528612 216804 573312 216832
rect 528612 216792 528618 216804
rect 573450 216792 573456 216844
rect 573508 216832 573514 216844
rect 596634 216832 596640 216844
rect 573508 216804 596640 216832
rect 573508 216792 573514 216804
rect 596634 216792 596640 216804
rect 596692 216792 596698 216844
rect 614482 216832 614488 216844
rect 597572 216804 614488 216832
rect 521286 216656 521292 216708
rect 521344 216696 521350 216708
rect 575014 216696 575020 216708
rect 521344 216668 575020 216696
rect 521344 216656 521350 216668
rect 575014 216656 575020 216668
rect 575072 216656 575078 216708
rect 584398 216656 584404 216708
rect 584456 216696 584462 216708
rect 597572 216696 597600 216804
rect 614482 216792 614488 216804
rect 614540 216792 614546 216844
rect 584456 216668 597600 216696
rect 584456 216656 584462 216668
rect 597738 216656 597744 216708
rect 597796 216696 597802 216708
rect 601648 216696 601654 216708
rect 597796 216668 601654 216696
rect 597796 216656 597802 216668
rect 601648 216656 601654 216668
rect 601706 216656 601712 216708
rect 601786 216656 601792 216708
rect 601844 216696 601850 216708
rect 605098 216696 605104 216708
rect 601844 216668 605104 216696
rect 601844 216656 601850 216668
rect 605098 216656 605104 216668
rect 605156 216656 605162 216708
rect 605834 216656 605840 216708
rect 605892 216696 605898 216708
rect 606754 216696 606760 216708
rect 605892 216668 606760 216696
rect 605892 216656 605898 216668
rect 606754 216656 606760 216668
rect 606812 216656 606818 216708
rect 607490 216656 607496 216708
rect 607548 216696 607554 216708
rect 614114 216696 614120 216708
rect 607548 216668 614120 216696
rect 607548 216656 607554 216668
rect 614114 216656 614120 216668
rect 614172 216656 614178 216708
rect 534074 216520 534080 216572
rect 534132 216560 534138 216572
rect 543642 216560 543648 216572
rect 534132 216532 543648 216560
rect 534132 216520 534138 216532
rect 543642 216520 543648 216532
rect 543700 216520 543706 216572
rect 547782 216520 547788 216572
rect 547840 216560 547846 216572
rect 554590 216560 554596 216572
rect 547840 216532 554596 216560
rect 547840 216520 547846 216532
rect 554590 216520 554596 216532
rect 554648 216520 554654 216572
rect 555050 216520 555056 216572
rect 555108 216560 555114 216572
rect 562686 216560 562692 216572
rect 555108 216532 562692 216560
rect 555108 216520 555114 216532
rect 562686 216520 562692 216532
rect 562744 216520 562750 216572
rect 563330 216520 563336 216572
rect 563388 216560 563394 216572
rect 563388 216532 582374 216560
rect 563388 216520 563394 216532
rect 582346 216492 582374 216532
rect 623314 216492 623320 216504
rect 582346 216464 623320 216492
rect 623314 216452 623320 216464
rect 623372 216452 623378 216504
rect 557074 216384 557080 216436
rect 557132 216424 557138 216436
rect 558546 216424 558552 216436
rect 557132 216396 558552 216424
rect 557132 216384 557138 216396
rect 558546 216384 558552 216396
rect 558604 216384 558610 216436
rect 562502 216384 562508 216436
rect 562560 216424 562566 216436
rect 571058 216424 571064 216436
rect 562560 216396 571064 216424
rect 562560 216384 562566 216396
rect 571058 216384 571064 216396
rect 571116 216384 571122 216436
rect 571242 216384 571248 216436
rect 571300 216424 571306 216436
rect 571300 216396 574048 216424
rect 571300 216384 571306 216396
rect 574020 215948 574048 216396
rect 574646 216316 574652 216368
rect 574704 216356 574710 216368
rect 621106 216356 621112 216368
rect 574704 216328 621112 216356
rect 574704 216316 574710 216328
rect 621106 216316 621112 216328
rect 621164 216316 621170 216368
rect 582558 216180 582564 216232
rect 582616 216220 582622 216232
rect 597554 216220 597560 216232
rect 582616 216192 597560 216220
rect 582616 216180 582622 216192
rect 597554 216180 597560 216192
rect 597612 216180 597618 216232
rect 619634 216084 619640 216096
rect 579586 216056 619640 216084
rect 574646 215948 574652 215960
rect 574020 215920 574652 215948
rect 574646 215908 574652 215920
rect 574704 215908 574710 215960
rect 574094 215772 574100 215824
rect 574152 215812 574158 215824
rect 579586 215812 579614 216056
rect 619634 216044 619640 216056
rect 619692 216044 619698 216096
rect 623038 215908 623044 215960
rect 623096 215948 623102 215960
rect 633802 215948 633808 215960
rect 623096 215920 633808 215948
rect 623096 215908 623102 215920
rect 633802 215908 633808 215920
rect 633860 215908 633866 215960
rect 574152 215784 579614 215812
rect 574152 215772 574158 215784
rect 590102 215568 590108 215620
rect 590160 215608 590166 215620
rect 595714 215608 595720 215620
rect 590160 215580 595720 215608
rect 590160 215568 590166 215580
rect 595714 215568 595720 215580
rect 595772 215568 595778 215620
rect 575382 215432 575388 215484
rect 575440 215472 575446 215484
rect 575440 215444 579614 215472
rect 575440 215432 575446 215444
rect 575198 215296 575204 215348
rect 575256 215336 575262 215348
rect 576394 215336 576400 215348
rect 575256 215308 576400 215336
rect 575256 215296 575262 215308
rect 576394 215296 576400 215308
rect 576452 215296 576458 215348
rect 579586 215268 579614 215444
rect 612274 215268 612280 215280
rect 579586 215240 612280 215268
rect 612274 215228 612280 215240
rect 612332 215228 612338 215280
rect 574278 215092 574284 215144
rect 574336 215132 574342 215144
rect 620002 215132 620008 215144
rect 574336 215104 620008 215132
rect 574336 215092 574342 215104
rect 620002 215092 620008 215104
rect 620060 215092 620066 215144
rect 676214 215092 676220 215144
rect 676272 215132 676278 215144
rect 677226 215132 677232 215144
rect 676272 215104 677232 215132
rect 676272 215092 676278 215104
rect 677226 215092 677232 215104
rect 677284 215092 677290 215144
rect 574830 214956 574836 215008
rect 574888 214996 574894 215008
rect 622394 214996 622400 215008
rect 574888 214968 622400 214996
rect 574888 214956 574894 214968
rect 622394 214956 622400 214968
rect 622452 214956 622458 215008
rect 663518 214888 663524 214940
rect 663576 214928 663582 214940
rect 664438 214928 664444 214940
rect 663576 214900 664444 214928
rect 663576 214888 663582 214900
rect 664438 214888 664444 214900
rect 664496 214888 664502 214940
rect 576026 214820 576032 214872
rect 576084 214860 576090 214872
rect 626074 214860 626080 214872
rect 576084 214832 626080 214860
rect 576084 214820 576090 214832
rect 626074 214820 626080 214832
rect 626132 214820 626138 214872
rect 574462 214684 574468 214736
rect 574520 214724 574526 214736
rect 616690 214724 616696 214736
rect 574520 214696 616696 214724
rect 574520 214684 574526 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 616874 214684 616880 214736
rect 616932 214724 616938 214736
rect 617794 214724 617800 214736
rect 616932 214696 617800 214724
rect 616932 214684 616938 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 658734 214684 658740 214736
rect 658792 214724 658798 214736
rect 661678 214724 661684 214736
rect 658792 214696 661684 214724
rect 658792 214684 658798 214696
rect 661678 214684 661684 214696
rect 661736 214684 661742 214736
rect 574646 214548 574652 214600
rect 574704 214588 574710 214600
rect 628282 214588 628288 214600
rect 574704 214560 628288 214588
rect 574704 214548 574710 214560
rect 628282 214548 628288 214560
rect 628340 214548 628346 214600
rect 631410 214548 631416 214600
rect 631468 214588 631474 214600
rect 632698 214588 632704 214600
rect 631468 214560 632704 214588
rect 631468 214548 631474 214560
rect 632698 214548 632704 214560
rect 632756 214548 632762 214600
rect 656802 214548 656808 214600
rect 656860 214588 656866 214600
rect 658918 214588 658924 214600
rect 656860 214560 658924 214588
rect 656860 214548 656866 214560
rect 658918 214548 658924 214560
rect 658976 214548 658982 214600
rect 662046 214548 662052 214600
rect 662104 214588 662110 214600
rect 663242 214588 663248 214600
rect 662104 214560 663248 214588
rect 662104 214548 662110 214560
rect 663242 214548 663248 214560
rect 663300 214548 663306 214600
rect 608778 214412 608784 214464
rect 608836 214452 608842 214464
rect 609514 214452 609520 214464
rect 608836 214424 609520 214452
rect 608836 214412 608842 214424
rect 609514 214412 609520 214424
rect 609572 214412 609578 214464
rect 611446 214412 611452 214464
rect 611504 214452 611510 214464
rect 611814 214452 611820 214464
rect 611504 214424 611820 214452
rect 611504 214412 611510 214424
rect 611814 214412 611820 214424
rect 611872 214412 611878 214464
rect 616690 214412 616696 214464
rect 616748 214452 616754 214464
rect 624418 214452 624424 214464
rect 616748 214424 624424 214452
rect 616748 214412 616754 214424
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 627730 214140 627736 214192
rect 627788 214180 627794 214192
rect 631042 214180 631048 214192
rect 627788 214152 631048 214180
rect 627788 214140 627794 214152
rect 631042 214140 631048 214152
rect 631100 214140 631106 214192
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 40678 213976 40684 213988
rect 35860 213948 40684 213976
rect 35860 213936 35866 213948
rect 40678 213936 40684 213948
rect 40736 213936 40742 213988
rect 612734 213868 612740 213920
rect 612792 213908 612798 213920
rect 615034 213908 615040 213920
rect 612792 213880 615040 213908
rect 612792 213868 612798 213880
rect 615034 213868 615040 213880
rect 615092 213868 615098 213920
rect 637574 213868 637580 213920
rect 637632 213908 637638 213920
rect 638218 213908 638224 213920
rect 637632 213880 638224 213908
rect 637632 213868 637638 213880
rect 638218 213868 638224 213880
rect 638276 213868 638282 213920
rect 639966 213868 639972 213920
rect 640024 213908 640030 213920
rect 643186 213908 643192 213920
rect 640024 213880 643192 213908
rect 640024 213868 640030 213880
rect 643186 213868 643192 213880
rect 643244 213868 643250 213920
rect 654870 213868 654876 213920
rect 654928 213908 654934 213920
rect 655422 213908 655428 213920
rect 654928 213880 655428 213908
rect 654928 213868 654934 213880
rect 655422 213868 655428 213880
rect 655480 213868 655486 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 576394 213732 576400 213784
rect 576452 213772 576458 213784
rect 598474 213772 598480 213784
rect 576452 213744 598480 213772
rect 576452 213732 576458 213744
rect 598474 213732 598480 213744
rect 598532 213732 598538 213784
rect 638034 213732 638040 213784
rect 638092 213772 638098 213784
rect 640426 213772 640432 213784
rect 638092 213744 640432 213772
rect 638092 213732 638098 213744
rect 640426 213732 640432 213744
rect 640484 213732 640490 213784
rect 644934 213732 644940 213784
rect 644992 213772 644998 213784
rect 646866 213772 646872 213784
rect 644992 213744 646872 213772
rect 644992 213732 644998 213744
rect 646866 213732 646872 213744
rect 646924 213732 646930 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 662966 213772 662972 213784
rect 661000 213744 662972 213772
rect 661000 213732 661006 213744
rect 662966 213732 662972 213744
rect 663024 213732 663030 213784
rect 575014 213596 575020 213648
rect 575072 213636 575078 213648
rect 601234 213636 601240 213648
rect 575072 213608 601240 213636
rect 575072 213596 575078 213608
rect 601234 213596 601240 213608
rect 601292 213596 601298 213648
rect 641622 213596 641628 213648
rect 641680 213636 641686 213648
rect 650638 213636 650644 213648
rect 641680 213608 650644 213636
rect 641680 213596 641686 213608
rect 650638 213596 650644 213608
rect 650696 213596 650702 213648
rect 652018 213596 652024 213648
rect 652076 213636 652082 213648
rect 657998 213636 658004 213648
rect 652076 213608 658004 213636
rect 652076 213596 652082 213608
rect 657998 213596 658004 213608
rect 658056 213596 658062 213648
rect 659562 213596 659568 213648
rect 659620 213636 659626 213648
rect 664898 213636 664904 213648
rect 659620 213608 664904 213636
rect 659620 213596 659626 213608
rect 664898 213596 664904 213608
rect 664956 213596 664962 213648
rect 603074 213528 603080 213580
rect 603132 213568 603138 213580
rect 604546 213568 604552 213580
rect 603132 213540 604552 213568
rect 603132 213528 603138 213540
rect 604546 213528 604552 213540
rect 604604 213528 604610 213580
rect 574094 213460 574100 213512
rect 574152 213500 574158 213512
rect 601786 213500 601792 213512
rect 574152 213472 601792 213500
rect 574152 213460 574158 213472
rect 601786 213460 601792 213472
rect 601844 213460 601850 213512
rect 642174 213460 642180 213512
rect 642232 213500 642238 213512
rect 659378 213500 659384 213512
rect 642232 213472 659384 213500
rect 642232 213460 642238 213472
rect 659378 213460 659384 213472
rect 659436 213460 659442 213512
rect 574094 213324 574100 213376
rect 574152 213364 574158 213376
rect 602338 213364 602344 213376
rect 574152 213336 602344 213364
rect 574152 213324 574158 213336
rect 602338 213324 602344 213336
rect 602396 213324 602402 213376
rect 602522 213324 602528 213376
rect 602580 213364 602586 213376
rect 622762 213364 622768 213376
rect 602580 213336 622768 213364
rect 602580 213324 602586 213336
rect 622762 213324 622768 213336
rect 622820 213324 622826 213376
rect 635550 213324 635556 213376
rect 635608 213364 635614 213376
rect 651834 213364 651840 213376
rect 635608 213336 651840 213364
rect 635608 213324 635614 213336
rect 651834 213324 651840 213336
rect 651892 213324 651898 213376
rect 652846 213324 652852 213376
rect 652904 213364 652910 213376
rect 660206 213364 660212 213376
rect 652904 213336 660212 213364
rect 652904 213324 652910 213336
rect 660206 213324 660212 213336
rect 660264 213324 660270 213376
rect 575566 213188 575572 213240
rect 575624 213228 575630 213240
rect 603074 213228 603080 213240
rect 575624 213200 603080 213228
rect 575624 213188 575630 213200
rect 603074 213188 603080 213200
rect 603132 213188 603138 213240
rect 623958 213188 623964 213240
rect 624016 213228 624022 213240
rect 629938 213228 629944 213240
rect 624016 213200 629944 213228
rect 624016 213188 624022 213200
rect 629938 213188 629944 213200
rect 629996 213188 630002 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 665266 213228 665272 213240
rect 643888 213200 665272 213228
rect 643888 213188 643894 213200
rect 665266 213188 665272 213200
rect 665324 213188 665330 213240
rect 676214 213188 676220 213240
rect 676272 213228 676278 213240
rect 676858 213228 676864 213240
rect 676272 213200 676864 213228
rect 676272 213188 676278 213200
rect 676858 213188 676864 213200
rect 676916 213188 676922 213240
rect 650454 212984 650460 213036
rect 650512 213024 650518 213036
rect 651282 213024 651288 213036
rect 650512 212996 651288 213024
rect 650512 212984 650518 212996
rect 651282 212984 651288 212996
rect 651340 212984 651346 213036
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 632882 212848 632888 212900
rect 632940 212888 632946 212900
rect 634354 212888 634360 212900
rect 632940 212860 634360 212888
rect 632940 212848 632946 212860
rect 634354 212848 634360 212860
rect 634412 212848 634418 212900
rect 636654 212780 636660 212832
rect 636712 212820 636718 212832
rect 639598 212820 639604 212832
rect 636712 212792 639604 212820
rect 636712 212780 636718 212792
rect 639598 212780 639604 212792
rect 639656 212780 639662 212832
rect 578510 211624 578516 211676
rect 578568 211664 578574 211676
rect 580442 211664 580448 211676
rect 578568 211636 580448 211664
rect 578568 211624 578574 211636
rect 580442 211624 580448 211636
rect 580500 211624 580506 211676
rect 612918 211624 612924 211676
rect 612976 211664 612982 211676
rect 613378 211664 613384 211676
rect 612976 211636 613384 211664
rect 612976 211624 612982 211636
rect 613378 211624 613384 211636
rect 613436 211624 613442 211676
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 41690 211188 41696 211200
rect 35860 211160 41696 211188
rect 35860 211148 35866 211160
rect 41690 211148 41696 211160
rect 41748 211148 41754 211200
rect 599210 210060 599216 210112
rect 599268 210100 599274 210112
rect 599578 210100 599584 210112
rect 599268 210072 599584 210100
rect 599268 210060 599274 210072
rect 599578 210060 599584 210072
rect 599636 210060 599642 210112
rect 579246 209788 579252 209840
rect 579304 209828 579310 209840
rect 581730 209828 581736 209840
rect 579304 209800 581736 209828
rect 579304 209788 579310 209800
rect 581730 209788 581736 209800
rect 581788 209788 581794 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 591298 208632 591304 208684
rect 591356 208672 591362 208684
rect 625126 208672 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 652260 209528 654134 209556
rect 652260 209516 652266 209528
rect 654106 209080 654134 209528
rect 667014 209080 667020 209092
rect 654106 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 591356 208644 625154 208672
rect 591356 208632 591362 208644
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 40034 208400 40040 208412
rect 35860 208372 40040 208400
rect 35860 208360 35866 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 580442 207612 580448 207664
rect 580500 207652 580506 207664
rect 589458 207652 589464 207664
rect 580500 207624 589464 207652
rect 580500 207612 580506 207624
rect 589458 207612 589464 207624
rect 589516 207612 589522 207664
rect 581730 206252 581736 206304
rect 581788 206292 581794 206304
rect 589642 206292 589648 206304
rect 581788 206264 589648 206292
rect 581788 206252 581794 206264
rect 589642 206252 589648 206264
rect 589700 206252 589706 206304
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 45462 196596 45468 196648
rect 45520 196636 45526 196648
rect 48590 196636 48596 196648
rect 45520 196608 48596 196636
rect 45520 196596 45526 196608
rect 48590 196596 48596 196608
rect 48648 196596 48654 196648
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 668118 194148 668124 194200
rect 668176 194188 668182 194200
rect 670786 194188 670792 194200
rect 668176 194160 670792 194188
rect 668176 194148 668182 194160
rect 670786 194148 670792 194160
rect 670844 194148 670850 194200
rect 668026 192516 668032 192568
rect 668084 192556 668090 192568
rect 669038 192556 669044 192568
rect 668084 192528 669044 192556
rect 668084 192516 668090 192528
rect 669038 192516 669044 192528
rect 669096 192516 669102 192568
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 669130 189252 669136 189304
rect 669188 189292 669194 189304
rect 670786 189292 670792 189304
rect 669188 189264 670792 189292
rect 669188 189252 669194 189264
rect 670786 189252 670792 189264
rect 670844 189252 670850 189304
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 668026 184356 668032 184408
rect 668084 184396 668090 184408
rect 669590 184396 669596 184408
rect 668084 184368 669596 184396
rect 668084 184356 668090 184368
rect 669590 184356 669596 184368
rect 669648 184356 669654 184408
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 583202 175244 583208 175296
rect 583260 175284 583266 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 583260 175256 586514 175284
rect 583260 175244 583266 175256
rect 667934 174836 667940 174888
rect 667992 174876 667998 174888
rect 669774 174876 669780 174888
rect 667992 174848 669780 174876
rect 667992 174836 667998 174848
rect 669774 174836 669780 174848
rect 669832 174836 669838 174888
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 581638 171096 581644 171148
rect 581696 171136 581702 171148
rect 589458 171136 589464 171148
rect 581696 171108 589464 171136
rect 581696 171096 581702 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 579522 170960 579528 171012
rect 579580 171000 579586 171012
rect 583202 171000 583208 171012
rect 579580 170972 583208 171000
rect 579580 170960 579586 170972
rect 583202 170960 583208 170972
rect 583260 170960 583266 171012
rect 582374 169736 582380 169788
rect 582432 169776 582438 169788
rect 589458 169776 589464 169788
rect 582432 169748 589464 169776
rect 582432 169736 582438 169748
rect 589458 169736 589464 169748
rect 589516 169736 589522 169788
rect 578326 169668 578332 169720
rect 578384 169708 578390 169720
rect 580902 169708 580908 169720
rect 578384 169680 580908 169708
rect 578384 169668 578390 169680
rect 580902 169668 580908 169680
rect 580960 169668 580966 169720
rect 579614 168376 579620 168428
rect 579672 168416 579678 168428
rect 589458 168416 589464 168428
rect 579672 168388 589464 168416
rect 579672 168376 579678 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578970 167152 578976 167204
rect 579028 167192 579034 167204
rect 581638 167192 581644 167204
rect 579028 167164 581644 167192
rect 579028 167152 579034 167164
rect 581638 167152 581644 167164
rect 581696 167152 581702 167204
rect 581638 167016 581644 167068
rect 581696 167056 581702 167068
rect 589458 167056 589464 167068
rect 581696 167028 589464 167056
rect 581696 167016 581702 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 669130 166064 669136 166116
rect 669188 166104 669194 166116
rect 670142 166104 670148 166116
rect 669188 166076 670148 166104
rect 669188 166064 669194 166076
rect 670142 166064 670148 166076
rect 670200 166064 670206 166116
rect 578878 165520 578884 165572
rect 578936 165560 578942 165572
rect 582374 165560 582380 165572
rect 578936 165532 582380 165560
rect 578936 165520 578942 165532
rect 582374 165520 582380 165532
rect 582432 165520 582438 165572
rect 668026 164772 668032 164824
rect 668084 164812 668090 164824
rect 670326 164812 670332 164824
rect 668084 164784 670332 164812
rect 668084 164772 668090 164784
rect 670326 164772 670332 164784
rect 670384 164772 670390 164824
rect 585962 164228 585968 164280
rect 586020 164268 586026 164280
rect 589458 164268 589464 164280
rect 586020 164240 589464 164268
rect 586020 164228 586026 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 584398 162868 584404 162920
rect 584456 162908 584462 162920
rect 589458 162908 589464 162920
rect 584456 162880 589464 162908
rect 584456 162868 584462 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 675846 162800 675852 162852
rect 675904 162840 675910 162852
rect 678238 162840 678244 162852
rect 675904 162812 678244 162840
rect 675904 162800 675910 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 676030 162596 676036 162648
rect 676088 162636 676094 162648
rect 679618 162636 679624 162648
rect 676088 162608 679624 162636
rect 676088 162596 676094 162608
rect 679618 162596 679624 162608
rect 679676 162596 679682 162648
rect 675846 161712 675852 161764
rect 675904 161752 675910 161764
rect 680998 161752 681004 161764
rect 675904 161724 681004 161752
rect 675904 161712 675910 161724
rect 680998 161712 681004 161724
rect 681056 161712 681062 161764
rect 580442 161440 580448 161492
rect 580500 161480 580506 161492
rect 589458 161480 589464 161492
rect 580500 161452 589464 161480
rect 580500 161440 580506 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 582374 160080 582380 160132
rect 582432 160120 582438 160132
rect 589458 160120 589464 160132
rect 582432 160092 589464 160120
rect 582432 160080 582438 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 579246 160012 579252 160064
rect 579304 160052 579310 160064
rect 581638 160052 581644 160064
rect 579304 160024 581644 160052
rect 579304 160012 579310 160024
rect 581638 160012 581644 160024
rect 581696 160012 581702 160064
rect 581822 158788 581828 158840
rect 581880 158828 581886 158840
rect 589458 158828 589464 158840
rect 581880 158800 589464 158828
rect 581880 158788 581886 158800
rect 589458 158788 589464 158800
rect 589516 158788 589522 158840
rect 579154 158652 579160 158704
rect 579212 158692 579218 158704
rect 585962 158692 585968 158704
rect 579212 158664 585968 158692
rect 579212 158652 579218 158664
rect 585962 158652 585968 158664
rect 586020 158652 586026 158704
rect 585778 157360 585784 157412
rect 585836 157400 585842 157412
rect 589458 157400 589464 157412
rect 585836 157372 589464 157400
rect 585836 157360 585842 157372
rect 589458 157360 589464 157372
rect 589516 157360 589522 157412
rect 579522 155864 579528 155916
rect 579580 155904 579586 155916
rect 584398 155904 584404 155916
rect 579580 155876 584404 155904
rect 579580 155864 579586 155876
rect 584398 155864 584404 155876
rect 584456 155864 584462 155916
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 578234 154504 578240 154556
rect 578292 154544 578298 154556
rect 580442 154544 580448 154556
rect 578292 154516 580448 154544
rect 578292 154504 578298 154516
rect 580442 154504 580448 154516
rect 580500 154504 580506 154556
rect 580258 153212 580264 153264
rect 580316 153252 580322 153264
rect 589458 153252 589464 153264
rect 580316 153224 589464 153252
rect 580316 153212 580322 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 582374 152776 582380 152788
rect 578292 152748 582380 152776
rect 578292 152736 578298 152748
rect 582374 152736 582380 152748
rect 582432 152736 582438 152788
rect 583018 151784 583024 151836
rect 583076 151824 583082 151836
rect 589458 151824 589464 151836
rect 583076 151796 589464 151824
rect 583076 151784 583082 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 581822 150600 581828 150612
rect 578936 150572 581828 150600
rect 578936 150560 578942 150572
rect 581822 150560 581828 150572
rect 581880 150560 581886 150612
rect 581638 150424 581644 150476
rect 581696 150464 581702 150476
rect 589458 150464 589464 150476
rect 581696 150436 589464 150464
rect 581696 150424 581702 150436
rect 589458 150424 589464 150436
rect 589516 150424 589522 150476
rect 668670 150220 668676 150272
rect 668728 150260 668734 150272
rect 670786 150260 670792 150272
rect 668728 150232 670792 150260
rect 668728 150220 668734 150232
rect 670786 150220 670792 150232
rect 670844 150220 670850 150272
rect 579522 147364 579528 147416
rect 579580 147404 579586 147416
rect 585778 147404 585784 147416
rect 579580 147376 585784 147404
rect 579580 147364 579586 147376
rect 585778 147364 585784 147376
rect 585836 147364 585842 147416
rect 587342 146276 587348 146328
rect 587400 146316 587406 146328
rect 589366 146316 589372 146328
rect 587400 146288 589372 146316
rect 587400 146276 587406 146288
rect 589366 146276 589372 146288
rect 589424 146276 589430 146328
rect 578878 145528 578884 145580
rect 578936 145568 578942 145580
rect 589182 145568 589188 145580
rect 578936 145540 589188 145568
rect 578936 145528 578942 145540
rect 589182 145528 589188 145540
rect 589240 145528 589246 145580
rect 585778 144916 585784 144968
rect 585836 144956 585842 144968
rect 589458 144956 589464 144968
rect 585836 144928 589464 144956
rect 585836 144916 585842 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 578510 143284 578516 143336
rect 578568 143324 578574 143336
rect 580258 143324 580264 143336
rect 578568 143296 580264 143324
rect 578568 143284 578574 143296
rect 580258 143284 580264 143296
rect 580316 143284 580322 143336
rect 580442 142128 580448 142180
rect 580500 142168 580506 142180
rect 589458 142168 589464 142180
rect 580500 142140 589464 142168
rect 580500 142128 580506 142140
rect 589458 142128 589464 142140
rect 589516 142128 589522 142180
rect 579522 140564 579528 140616
rect 579580 140604 579586 140616
rect 583018 140604 583024 140616
rect 579580 140576 583024 140604
rect 579580 140564 579586 140576
rect 583018 140564 583024 140576
rect 583076 140564 583082 140616
rect 584398 139408 584404 139460
rect 584456 139448 584462 139460
rect 589458 139448 589464 139460
rect 584456 139420 589464 139448
rect 584456 139408 584462 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578694 139340 578700 139392
rect 578752 139380 578758 139392
rect 581638 139380 581644 139392
rect 578752 139352 581644 139380
rect 578752 139340 578758 139352
rect 581638 139340 581644 139352
rect 581696 139340 581702 139392
rect 581638 136620 581644 136672
rect 581696 136660 581702 136672
rect 589458 136660 589464 136672
rect 581696 136632 589464 136660
rect 581696 136620 581702 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 667934 136416 667940 136468
rect 667992 136456 667998 136468
rect 669958 136456 669964 136468
rect 667992 136428 669964 136456
rect 667992 136416 667998 136428
rect 669958 136416 669964 136428
rect 670016 136416 670022 136468
rect 578326 135872 578332 135924
rect 578384 135912 578390 135924
rect 587342 135912 587348 135924
rect 578384 135884 587348 135912
rect 578384 135872 578390 135884
rect 587342 135872 587348 135884
rect 587400 135872 587406 135924
rect 587158 135260 587164 135312
rect 587216 135300 587222 135312
rect 589274 135300 589280 135312
rect 587216 135272 589280 135300
rect 587216 135260 587222 135272
rect 589274 135260 589280 135272
rect 589332 135260 589338 135312
rect 578234 134240 578240 134292
rect 578292 134280 578298 134292
rect 585778 134280 585784 134292
rect 578292 134252 585784 134280
rect 578292 134240 578298 134252
rect 585778 134240 585784 134252
rect 585836 134240 585842 134292
rect 585962 133900 585968 133952
rect 586020 133940 586026 133952
rect 589458 133940 589464 133952
rect 586020 133912 589464 133940
rect 586020 133900 586026 133912
rect 589458 133900 589464 133912
rect 589516 133900 589522 133952
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 579246 133152 579252 133204
rect 579304 133192 579310 133204
rect 589090 133192 589096 133204
rect 579304 133164 589096 133192
rect 579304 133152 579310 133164
rect 589090 133152 589096 133164
rect 589148 133152 589154 133204
rect 582374 131724 582380 131776
rect 582432 131764 582438 131776
rect 589918 131764 589924 131776
rect 582432 131736 589924 131764
rect 582432 131724 582438 131736
rect 589918 131724 589924 131736
rect 589976 131724 589982 131776
rect 579522 129684 579528 129736
rect 579580 129724 579586 129736
rect 582374 129724 582380 129736
rect 579580 129696 582380 129724
rect 579580 129684 579586 129696
rect 582374 129684 582380 129696
rect 582432 129684 582438 129736
rect 583018 128324 583024 128376
rect 583076 128364 583082 128376
rect 589458 128364 589464 128376
rect 583076 128336 589464 128364
rect 583076 128324 583082 128336
rect 589458 128324 589464 128336
rect 589516 128324 589522 128376
rect 578326 128256 578332 128308
rect 578384 128296 578390 128308
rect 580442 128296 580448 128308
rect 578384 128268 580448 128296
rect 578384 128256 578390 128268
rect 580442 128256 580448 128268
rect 580500 128256 580506 128308
rect 580258 126964 580264 127016
rect 580316 127004 580322 127016
rect 589458 127004 589464 127016
rect 580316 126976 589464 127004
rect 580316 126964 580322 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 585778 124176 585784 124228
rect 585836 124216 585842 124228
rect 589458 124216 589464 124228
rect 585836 124188 589464 124216
rect 585836 124176 585842 124188
rect 589458 124176 589464 124188
rect 589516 124176 589522 124228
rect 579246 124108 579252 124160
rect 579304 124148 579310 124160
rect 584398 124148 584404 124160
rect 579304 124120 584404 124148
rect 579304 124108 579310 124120
rect 584398 124108 584404 124120
rect 584456 124108 584462 124160
rect 579246 122816 579252 122868
rect 579304 122856 579310 122868
rect 589458 122856 589464 122868
rect 579304 122828 589464 122856
rect 579304 122816 579310 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 584398 121456 584404 121508
rect 584456 121496 584462 121508
rect 589458 121496 589464 121508
rect 584456 121468 589464 121496
rect 584456 121456 584462 121468
rect 589458 121456 589464 121468
rect 589516 121456 589522 121508
rect 579062 121116 579068 121168
rect 579120 121156 579126 121168
rect 581638 121156 581644 121168
rect 579120 121128 581644 121156
rect 579120 121116 579126 121128
rect 581638 121116 581644 121128
rect 581696 121116 581702 121168
rect 582006 120708 582012 120760
rect 582064 120748 582070 120760
rect 590102 120748 590108 120760
rect 582064 120720 590108 120748
rect 582064 120708 582070 120720
rect 590102 120708 590108 120720
rect 590160 120708 590166 120760
rect 578510 118600 578516 118652
rect 578568 118640 578574 118652
rect 587158 118640 587164 118652
rect 578568 118612 587164 118640
rect 578568 118600 578574 118612
rect 587158 118600 587164 118612
rect 587216 118600 587222 118652
rect 668026 118328 668032 118380
rect 668084 118368 668090 118380
rect 670142 118368 670148 118380
rect 668084 118340 670148 118368
rect 668084 118328 668090 118340
rect 670142 118328 670148 118340
rect 670200 118328 670206 118380
rect 583202 117308 583208 117360
rect 583260 117348 583266 117360
rect 589458 117348 589464 117360
rect 583260 117320 589464 117348
rect 583260 117308 583266 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 682378 117280 682384 117292
rect 675904 117252 682384 117280
rect 675904 117240 675910 117252
rect 682378 117240 682384 117252
rect 682436 117240 682442 117292
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 585962 116940 585968 116952
rect 579580 116912 585968 116940
rect 579580 116900 579586 116912
rect 585962 116900 585968 116912
rect 586020 116900 586026 116952
rect 587802 115948 587808 116000
rect 587860 115988 587866 116000
rect 589458 115988 589464 116000
rect 587860 115960 589464 115988
rect 587860 115948 587866 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 585134 115336 585140 115388
rect 585192 115376 585198 115388
rect 589918 115376 589924 115388
rect 585192 115348 589924 115376
rect 585192 115336 585198 115348
rect 589918 115336 589924 115348
rect 589976 115336 589982 115388
rect 579062 115200 579068 115252
rect 579120 115240 579126 115252
rect 587802 115240 587808 115252
rect 579120 115212 587808 115240
rect 579120 115200 579126 115212
rect 587802 115200 587808 115212
rect 587860 115200 587866 115252
rect 587158 114520 587164 114572
rect 587216 114560 587222 114572
rect 589826 114560 589832 114572
rect 587216 114532 589832 114560
rect 587216 114520 587222 114532
rect 589826 114520 589832 114532
rect 589884 114520 589890 114572
rect 579522 114384 579528 114436
rect 579580 114424 579586 114436
rect 591298 114424 591304 114436
rect 579580 114396 591304 114424
rect 579580 114384 579586 114396
rect 591298 114384 591304 114396
rect 591356 114384 591362 114436
rect 668118 114112 668124 114164
rect 668176 114152 668182 114164
rect 669958 114152 669964 114164
rect 668176 114124 669964 114152
rect 668176 114112 668182 114124
rect 669958 114112 669964 114124
rect 670016 114112 670022 114164
rect 579522 113092 579528 113144
rect 579580 113132 579586 113144
rect 588538 113132 588544 113144
rect 579580 113104 588544 113132
rect 579580 113092 579586 113104
rect 588538 113092 588544 113104
rect 588596 113092 588602 113144
rect 588538 110440 588544 110492
rect 588596 110480 588602 110492
rect 590562 110480 590568 110492
rect 588596 110452 590568 110480
rect 588596 110440 588602 110452
rect 590562 110440 590568 110452
rect 590620 110440 590626 110492
rect 579430 110236 579436 110288
rect 579488 110276 579494 110288
rect 582006 110276 582012 110288
rect 579488 110248 582012 110276
rect 579488 110236 579494 110248
rect 582006 110236 582012 110248
rect 582064 110236 582070 110288
rect 581822 109692 581828 109744
rect 581880 109732 581886 109744
rect 589366 109732 589372 109744
rect 581880 109704 589372 109732
rect 581880 109692 581886 109704
rect 589366 109692 589372 109704
rect 589424 109692 589430 109744
rect 578326 108332 578332 108384
rect 578384 108372 578390 108384
rect 585134 108372 585140 108384
rect 578384 108344 585140 108372
rect 578384 108332 578390 108344
rect 585134 108332 585140 108344
rect 585192 108332 585198 108384
rect 589458 107692 589464 107704
rect 579632 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 579632 107624 579660 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 579660 107624
rect 578936 107584 578942 107596
rect 580626 107040 580632 107092
rect 580684 107080 580690 107092
rect 590102 107080 590108 107092
rect 580684 107052 590108 107080
rect 580684 107040 580690 107052
rect 590102 107040 590108 107052
rect 590160 107040 590166 107092
rect 578326 106904 578332 106956
rect 578384 106944 578390 106956
rect 580258 106944 580264 106956
rect 578384 106916 580264 106944
rect 578384 106904 578390 106916
rect 580258 106904 580264 106916
rect 580316 106904 580322 106956
rect 580442 106904 580448 106956
rect 580500 106944 580506 106956
rect 589642 106944 589648 106956
rect 580500 106916 589648 106944
rect 580500 106904 580506 106916
rect 589642 106904 589648 106916
rect 589700 106904 589706 106956
rect 667198 106156 667204 106208
rect 667256 106196 667262 106208
rect 670694 106196 670700 106208
rect 667256 106168 670700 106196
rect 667256 106156 667262 106168
rect 670694 106156 670700 106168
rect 670752 106156 670758 106208
rect 581638 104864 581644 104916
rect 581696 104904 581702 104916
rect 589458 104904 589464 104916
rect 581696 104876 589464 104904
rect 581696 104864 581702 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 579522 103300 579528 103352
rect 579580 103340 579586 103352
rect 583018 103340 583024 103352
rect 579580 103312 583024 103340
rect 579580 103300 579586 103312
rect 583018 103300 583024 103312
rect 583076 103300 583082 103352
rect 585962 100716 585968 100768
rect 586020 100756 586026 100768
rect 589458 100756 589464 100768
rect 586020 100728 589464 100756
rect 586020 100716 586026 100728
rect 589458 100716 589464 100728
rect 589516 100716 589522 100768
rect 615218 100104 615224 100156
rect 615276 100144 615282 100156
rect 668026 100144 668032 100156
rect 615276 100116 668032 100144
rect 615276 100104 615282 100116
rect 668026 100104 668032 100116
rect 668084 100104 668090 100156
rect 613378 99968 613384 100020
rect 613436 100008 613442 100020
rect 668486 100008 668492 100020
rect 613436 99980 668492 100008
rect 613436 99968 613442 99980
rect 668486 99968 668492 99980
rect 668544 99968 668550 100020
rect 577498 99288 577504 99340
rect 577556 99328 577562 99340
rect 595254 99328 595260 99340
rect 577556 99300 595260 99328
rect 577556 99288 577562 99300
rect 595254 99288 595260 99300
rect 595312 99288 595318 99340
rect 624602 99288 624608 99340
rect 624660 99328 624666 99340
rect 632974 99328 632980 99340
rect 624660 99300 632980 99328
rect 624660 99288 624666 99300
rect 632974 99288 632980 99300
rect 633032 99288 633038 99340
rect 579522 99152 579528 99204
rect 579580 99192 579586 99204
rect 585778 99192 585784 99204
rect 579580 99164 585784 99192
rect 579580 99152 579586 99164
rect 585778 99152 585784 99164
rect 585836 99152 585842 99204
rect 626810 99152 626816 99204
rect 626868 99192 626874 99204
rect 636378 99192 636384 99204
rect 626868 99164 636384 99192
rect 626868 99152 626874 99164
rect 636378 99152 636384 99164
rect 636436 99152 636442 99204
rect 623682 99016 623688 99068
rect 623740 99056 623746 99068
rect 632146 99056 632152 99068
rect 623740 99028 632152 99056
rect 623740 99016 623746 99028
rect 632146 99016 632152 99028
rect 632204 99016 632210 99068
rect 629754 98880 629760 98932
rect 629812 98920 629818 98932
rect 640978 98920 640984 98932
rect 629812 98892 640984 98920
rect 629812 98880 629818 98892
rect 640978 98880 640984 98892
rect 641036 98880 641042 98932
rect 622302 98744 622308 98796
rect 622360 98784 622366 98796
rect 629478 98784 629484 98796
rect 622360 98756 629484 98784
rect 622360 98744 622366 98756
rect 629478 98744 629484 98756
rect 629536 98744 629542 98796
rect 630490 98744 630496 98796
rect 630548 98784 630554 98796
rect 642174 98784 642180 98796
rect 630548 98756 642180 98784
rect 630548 98744 630554 98756
rect 642174 98744 642180 98756
rect 642232 98744 642238 98796
rect 625062 98608 625068 98660
rect 625120 98648 625126 98660
rect 634446 98648 634452 98660
rect 625120 98620 634452 98648
rect 625120 98608 625126 98620
rect 634446 98608 634452 98620
rect 634504 98608 634510 98660
rect 637850 98608 637856 98660
rect 637908 98648 637914 98660
rect 660390 98648 660396 98660
rect 637908 98620 660396 98648
rect 637908 98608 637914 98620
rect 660390 98608 660396 98620
rect 660448 98608 660454 98660
rect 605466 97928 605472 97980
rect 605524 97968 605530 97980
rect 606478 97968 606484 97980
rect 605524 97940 606484 97968
rect 605524 97928 605530 97940
rect 606478 97928 606484 97940
rect 606536 97928 606542 97980
rect 620186 97928 620192 97980
rect 620244 97968 620250 97980
rect 626258 97968 626264 97980
rect 620244 97940 626264 97968
rect 620244 97928 620250 97940
rect 626258 97928 626264 97940
rect 626316 97928 626322 97980
rect 632698 97928 632704 97980
rect 632756 97968 632762 97980
rect 644014 97968 644020 97980
rect 632756 97940 644020 97968
rect 632756 97928 632762 97940
rect 644014 97928 644020 97940
rect 644072 97928 644078 97980
rect 651098 97928 651104 97980
rect 651156 97968 651162 97980
rect 655054 97968 655060 97980
rect 651156 97940 655060 97968
rect 651156 97928 651162 97940
rect 655054 97928 655060 97940
rect 655112 97928 655118 97980
rect 655422 97928 655428 97980
rect 655480 97968 655486 97980
rect 662506 97968 662512 97980
rect 655480 97940 662512 97968
rect 655480 97928 655486 97940
rect 662506 97928 662512 97940
rect 662564 97928 662570 97980
rect 618714 97792 618720 97844
rect 618772 97832 618778 97844
rect 625430 97832 625436 97844
rect 618772 97804 625436 97832
rect 618772 97792 618778 97804
rect 625430 97792 625436 97804
rect 625488 97792 625494 97844
rect 643738 97792 643744 97844
rect 643796 97832 643802 97844
rect 650638 97832 650644 97844
rect 643796 97804 650644 97832
rect 643796 97792 643802 97804
rect 650638 97792 650644 97804
rect 650696 97792 650702 97844
rect 651834 97792 651840 97844
rect 651892 97832 651898 97844
rect 659562 97832 659568 97844
rect 651892 97804 659568 97832
rect 651892 97792 651898 97804
rect 659562 97792 659568 97804
rect 659620 97792 659626 97844
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665542 97832 665548 97844
rect 659988 97804 665548 97832
rect 659988 97792 659994 97804
rect 665542 97792 665548 97804
rect 665600 97792 665606 97844
rect 621658 97656 621664 97708
rect 621716 97696 621722 97708
rect 628374 97696 628380 97708
rect 621716 97668 628380 97696
rect 621716 97656 621722 97668
rect 628374 97656 628380 97668
rect 628432 97656 628438 97708
rect 633342 97656 633348 97708
rect 633400 97696 633406 97708
rect 643462 97696 643468 97708
rect 633400 97668 643468 97696
rect 633400 97656 633406 97668
rect 643462 97656 643468 97668
rect 643520 97656 643526 97708
rect 659194 97656 659200 97708
rect 659252 97696 659258 97708
rect 663886 97696 663892 97708
rect 659252 97668 663892 97696
rect 659252 97656 659258 97668
rect 663886 97656 663892 97668
rect 663944 97656 663950 97708
rect 615034 97520 615040 97572
rect 615092 97560 615098 97572
rect 616138 97560 616144 97572
rect 615092 97532 616144 97560
rect 615092 97520 615098 97532
rect 616138 97520 616144 97532
rect 616196 97520 616202 97572
rect 623130 97520 623136 97572
rect 623188 97560 623194 97572
rect 630674 97560 630680 97572
rect 623188 97532 630680 97560
rect 623188 97520 623194 97532
rect 630674 97520 630680 97532
rect 630732 97520 630738 97572
rect 631962 97520 631968 97572
rect 632020 97560 632026 97572
rect 644934 97560 644940 97572
rect 632020 97532 644940 97560
rect 632020 97520 632026 97532
rect 644934 97520 644940 97532
rect 644992 97520 644998 97572
rect 647142 97520 647148 97572
rect 647200 97560 647206 97572
rect 657998 97560 658004 97572
rect 647200 97532 658004 97560
rect 647200 97520 647206 97532
rect 657998 97520 658004 97532
rect 658056 97520 658062 97572
rect 658182 97520 658188 97572
rect 658240 97560 658246 97572
rect 663058 97560 663064 97572
rect 658240 97532 663064 97560
rect 658240 97520 658246 97532
rect 663058 97520 663064 97532
rect 663116 97520 663122 97572
rect 579522 97452 579528 97504
rect 579580 97492 579586 97504
rect 584398 97492 584404 97504
rect 579580 97464 584404 97492
rect 579580 97452 579586 97464
rect 584398 97452 584404 97464
rect 584456 97452 584462 97504
rect 627546 97384 627552 97436
rect 627604 97424 627610 97436
rect 637574 97424 637580 97436
rect 627604 97396 637580 97424
rect 627604 97384 627610 97396
rect 637574 97384 637580 97396
rect 637632 97384 637638 97436
rect 639874 97424 639880 97436
rect 639524 97396 639880 97424
rect 577498 97248 577504 97300
rect 577556 97288 577562 97300
rect 600406 97288 600412 97300
rect 577556 97260 600412 97288
rect 577556 97248 577562 97260
rect 600406 97248 600412 97260
rect 600464 97248 600470 97300
rect 612642 97248 612648 97300
rect 612700 97288 612706 97300
rect 620278 97288 620284 97300
rect 612700 97260 620284 97288
rect 612700 97248 612706 97260
rect 620278 97248 620284 97260
rect 620336 97248 620342 97300
rect 629018 97248 629024 97300
rect 629076 97288 629082 97300
rect 639524 97288 639552 97396
rect 639874 97384 639880 97396
rect 639932 97384 639938 97436
rect 644290 97384 644296 97436
rect 644348 97424 644354 97436
rect 658826 97424 658832 97436
rect 644348 97396 658832 97424
rect 644348 97384 644354 97396
rect 658826 97384 658832 97396
rect 658884 97384 658890 97436
rect 644750 97288 644756 97300
rect 629076 97260 639552 97288
rect 639616 97260 644756 97288
rect 629076 97248 629082 97260
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 639616 97152 639644 97260
rect 644750 97248 644756 97260
rect 644808 97248 644814 97300
rect 653950 97248 653956 97300
rect 654008 97288 654014 97300
rect 655238 97288 655244 97300
rect 654008 97260 655244 97288
rect 654008 97248 654014 97260
rect 655238 97248 655244 97260
rect 655296 97248 655302 97300
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 634228 97124 639644 97152
rect 634228 97112 634234 97124
rect 643002 97112 643008 97164
rect 643060 97152 643066 97164
rect 643060 97124 644474 97152
rect 643060 97112 643066 97124
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 643738 97016 643744 97028
rect 634780 96988 643744 97016
rect 634780 96976 634786 96988
rect 643738 96976 643744 96988
rect 643796 96976 643802 97028
rect 598934 96908 598940 96960
rect 598992 96948 598998 96960
rect 599670 96948 599676 96960
rect 598992 96920 599676 96948
rect 598992 96908 598998 96920
rect 599670 96908 599676 96920
rect 599728 96908 599734 96960
rect 612090 96908 612096 96960
rect 612148 96948 612154 96960
rect 612642 96948 612648 96960
rect 612148 96920 612648 96948
rect 612148 96908 612154 96920
rect 612642 96908 612648 96920
rect 612700 96908 612706 96960
rect 617242 96908 617248 96960
rect 617300 96948 617306 96960
rect 618162 96948 618168 96960
rect 617300 96920 618168 96948
rect 617300 96908 617306 96920
rect 618162 96908 618168 96920
rect 618220 96908 618226 96960
rect 626074 96840 626080 96892
rect 626132 96880 626138 96892
rect 635274 96880 635280 96892
rect 626132 96852 635280 96880
rect 626132 96840 626138 96852
rect 635274 96840 635280 96852
rect 635332 96840 635338 96892
rect 606202 96772 606208 96824
rect 606260 96812 606266 96824
rect 611998 96812 612004 96824
rect 606260 96784 612004 96812
rect 606260 96772 606266 96784
rect 611998 96772 612004 96784
rect 612056 96772 612062 96824
rect 615770 96772 615776 96824
rect 615828 96812 615834 96824
rect 618898 96812 618904 96824
rect 615828 96784 618904 96812
rect 615828 96772 615834 96784
rect 618898 96772 618904 96784
rect 618956 96772 618962 96824
rect 644446 96812 644474 97124
rect 650362 97112 650368 97164
rect 650420 97152 650426 97164
rect 658274 97152 658280 97164
rect 650420 97124 658280 97152
rect 650420 97112 650426 97124
rect 658274 97112 658280 97124
rect 658332 97112 658338 97164
rect 645210 97044 645216 97096
rect 645268 97084 645274 97096
rect 649258 97084 649264 97096
rect 645268 97056 649264 97084
rect 645268 97044 645274 97056
rect 649258 97044 649264 97056
rect 649316 97044 649322 97096
rect 657998 96976 658004 97028
rect 658056 97016 658062 97028
rect 661954 97016 661960 97028
rect 658056 96988 661960 97016
rect 658056 96976 658062 96988
rect 661954 96976 661960 96988
rect 662012 96976 662018 97028
rect 646682 96908 646688 96960
rect 646740 96948 646746 96960
rect 647878 96948 647884 96960
rect 646740 96920 647884 96948
rect 646740 96908 646746 96920
rect 647878 96908 647884 96920
rect 647936 96908 647942 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 660114 96812 660120 96824
rect 644446 96784 660120 96812
rect 660114 96772 660120 96784
rect 660172 96772 660178 96824
rect 628190 96704 628196 96756
rect 628248 96744 628254 96756
rect 639046 96744 639052 96756
rect 628248 96716 639052 96744
rect 628248 96704 628254 96716
rect 639046 96704 639052 96716
rect 639104 96704 639110 96756
rect 660666 96704 660672 96756
rect 660724 96744 660730 96756
rect 663242 96744 663248 96756
rect 660724 96716 663248 96744
rect 660724 96704 660730 96716
rect 663242 96704 663248 96716
rect 663300 96704 663306 96756
rect 631226 96568 631232 96620
rect 631284 96608 631290 96620
rect 643186 96608 643192 96620
rect 631284 96580 643192 96608
rect 631284 96568 631290 96580
rect 643186 96568 643192 96580
rect 643244 96568 643250 96620
rect 649626 96568 649632 96620
rect 649684 96608 649690 96620
rect 650822 96608 650828 96620
rect 649684 96580 650828 96608
rect 649684 96568 649690 96580
rect 650822 96568 650828 96580
rect 650880 96568 650886 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 665358 96608 665364 96620
rect 652628 96580 665364 96608
rect 652628 96568 652634 96580
rect 665358 96568 665364 96580
rect 665416 96568 665422 96620
rect 640058 96432 640064 96484
rect 640116 96472 640122 96484
rect 647694 96472 647700 96484
rect 640116 96444 647700 96472
rect 640116 96432 640122 96444
rect 647694 96432 647700 96444
rect 647752 96432 647758 96484
rect 648154 96432 648160 96484
rect 648212 96472 648218 96484
rect 652018 96472 652024 96484
rect 648212 96444 652024 96472
rect 648212 96432 648218 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 653858 96472 653864 96484
rect 652220 96444 653864 96472
rect 610618 96296 610624 96348
rect 610676 96336 610682 96348
rect 623038 96336 623044 96348
rect 610676 96308 623044 96336
rect 610676 96296 610682 96308
rect 623038 96296 623044 96308
rect 623096 96296 623102 96348
rect 639322 96296 639328 96348
rect 639380 96336 639386 96348
rect 652220 96336 652248 96444
rect 653858 96432 653864 96444
rect 653916 96432 653922 96484
rect 639380 96308 652248 96336
rect 639380 96296 639386 96308
rect 653306 96296 653312 96348
rect 653364 96336 653370 96348
rect 664162 96336 664168 96348
rect 653364 96308 664168 96336
rect 653364 96296 653370 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 609146 96160 609152 96212
rect 609204 96200 609210 96212
rect 621658 96200 621664 96212
rect 609204 96172 621664 96200
rect 609204 96160 609210 96172
rect 621658 96160 621664 96172
rect 621716 96160 621722 96212
rect 640794 96160 640800 96212
rect 640852 96200 640858 96212
rect 663702 96200 663708 96212
rect 640852 96172 663708 96200
rect 640852 96160 640858 96172
rect 663702 96160 663708 96172
rect 663760 96160 663766 96212
rect 607674 96024 607680 96076
rect 607732 96064 607738 96076
rect 620738 96064 620744 96076
rect 607732 96036 620744 96064
rect 607732 96024 607738 96036
rect 620738 96024 620744 96036
rect 620796 96024 620802 96076
rect 620922 96024 620928 96076
rect 620980 96064 620986 96076
rect 626442 96064 626448 96076
rect 620980 96036 626448 96064
rect 620980 96024 620986 96036
rect 626442 96024 626448 96036
rect 626500 96024 626506 96076
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 665174 96064 665180 96076
rect 641588 96036 665180 96064
rect 641588 96024 641594 96036
rect 665174 96024 665180 96036
rect 665232 96024 665238 96076
rect 594058 95888 594064 95940
rect 594116 95928 594122 95940
rect 601878 95928 601884 95940
rect 594116 95900 601884 95928
rect 594116 95888 594122 95900
rect 601878 95888 601884 95900
rect 601936 95888 601942 95940
rect 613562 95888 613568 95940
rect 613620 95928 613626 95940
rect 613620 95900 625154 95928
rect 613620 95888 613626 95900
rect 625126 95656 625154 95900
rect 635458 95888 635464 95940
rect 635516 95928 635522 95940
rect 646038 95928 646044 95940
rect 635516 95900 646044 95928
rect 635516 95888 635522 95900
rect 646038 95888 646044 95900
rect 646096 95888 646102 95940
rect 647694 95888 647700 95940
rect 647752 95928 647758 95940
rect 653398 95928 653404 95940
rect 647752 95900 653404 95928
rect 647752 95888 647758 95900
rect 653398 95888 653404 95900
rect 653456 95888 653462 95940
rect 664622 95928 664628 95940
rect 654106 95900 664628 95928
rect 638586 95752 638592 95804
rect 638644 95792 638650 95804
rect 642818 95792 642824 95804
rect 638644 95764 642824 95792
rect 638644 95752 638650 95764
rect 642818 95752 642824 95764
rect 642876 95752 642882 95804
rect 648890 95752 648896 95804
rect 648948 95792 648954 95804
rect 654106 95792 654134 95900
rect 664622 95888 664628 95900
rect 664680 95888 664686 95940
rect 648948 95764 654134 95792
rect 648948 95752 648954 95764
rect 646222 95656 646228 95668
rect 625126 95628 646228 95656
rect 646222 95616 646228 95628
rect 646280 95616 646286 95668
rect 642818 95480 642824 95532
rect 642876 95520 642882 95532
rect 648522 95520 648528 95532
rect 642876 95492 648528 95520
rect 642876 95480 642882 95492
rect 648522 95480 648528 95492
rect 648580 95480 648586 95532
rect 642634 95208 642640 95260
rect 642692 95248 642698 95260
rect 644474 95248 644480 95260
rect 642692 95220 644480 95248
rect 642692 95208 642698 95220
rect 644474 95208 644480 95220
rect 644532 95208 644538 95260
rect 578694 95004 578700 95056
rect 578752 95044 578758 95056
rect 580626 95044 580632 95056
rect 578752 95016 580632 95044
rect 578752 95004 578758 95016
rect 580626 95004 580632 95016
rect 580684 95004 580690 95056
rect 616506 94596 616512 94648
rect 616564 94636 616570 94648
rect 625798 94636 625804 94648
rect 616564 94608 625804 94636
rect 616564 94596 616570 94608
rect 625798 94596 625804 94608
rect 625856 94596 625862 94648
rect 608410 94460 608416 94512
rect 608468 94500 608474 94512
rect 624418 94500 624424 94512
rect 608468 94472 624424 94500
rect 608468 94460 608474 94472
rect 624418 94460 624424 94472
rect 624476 94460 624482 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 644474 93780 644480 93832
rect 644532 93820 644538 93832
rect 654870 93820 654876 93832
rect 644532 93792 654876 93820
rect 644532 93780 644538 93792
rect 654870 93780 654876 93792
rect 654928 93780 654934 93832
rect 579522 93236 579528 93288
rect 579580 93276 579586 93288
rect 583202 93276 583208 93288
rect 579580 93248 583208 93276
rect 579580 93236 579586 93248
rect 583202 93236 583208 93248
rect 583260 93236 583266 93288
rect 580258 93100 580264 93152
rect 580316 93140 580322 93152
rect 590102 93140 590108 93152
rect 580316 93112 590108 93140
rect 580316 93100 580322 93112
rect 590102 93100 590108 93112
rect 590160 93100 590166 93152
rect 664438 92488 664444 92540
rect 664496 92528 664502 92540
rect 668302 92528 668308 92540
rect 664496 92500 668308 92528
rect 664496 92488 664502 92500
rect 668302 92488 668308 92500
rect 668360 92488 668366 92540
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 625430 92460 625436 92472
rect 618036 92432 625436 92460
rect 618036 92420 618042 92432
rect 625430 92420 625436 92432
rect 625488 92420 625494 92472
rect 648522 92420 648528 92472
rect 648580 92460 648586 92472
rect 655422 92460 655428 92472
rect 648580 92432 655428 92460
rect 648580 92420 648586 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 617334 91032 617340 91044
rect 611320 91004 617340 91032
rect 611320 90992 611326 91004
rect 617334 90992 617340 91004
rect 617392 90992 617398 91044
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 620738 89632 620744 89684
rect 620796 89672 620802 89684
rect 626442 89672 626448 89684
rect 620796 89644 626448 89672
rect 620796 89632 620802 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 645762 88748 645768 88800
rect 645820 88788 645826 88800
rect 657446 88788 657452 88800
rect 645820 88760 657452 88788
rect 645820 88748 645826 88760
rect 657446 88748 657452 88760
rect 657504 88748 657510 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 579522 88272 579528 88324
rect 579580 88312 579586 88324
rect 587158 88312 587164 88324
rect 579580 88284 587164 88312
rect 579580 88272 579586 88284
rect 587158 88272 587164 88284
rect 587216 88272 587222 88324
rect 607214 88272 607220 88324
rect 607272 88312 607278 88324
rect 626442 88312 626448 88324
rect 607272 88284 626448 88312
rect 607272 88272 607278 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655054 88272 655060 88324
rect 655112 88312 655118 88324
rect 658458 88312 658464 88324
rect 655112 88284 658464 88312
rect 655112 88272 655118 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 617334 88136 617340 88188
rect 617392 88176 617398 88188
rect 625614 88176 625620 88188
rect 617392 88148 625620 88176
rect 617392 88136 617398 88148
rect 625614 88136 625620 88148
rect 625672 88136 625678 88188
rect 647878 87116 647884 87168
rect 647936 87156 647942 87168
rect 657170 87156 657176 87168
rect 647936 87128 657176 87156
rect 647936 87116 647942 87128
rect 657170 87116 657176 87128
rect 657228 87116 657234 87168
rect 649258 86980 649264 87032
rect 649316 87020 649322 87032
rect 660666 87020 660672 87032
rect 649316 86992 660672 87020
rect 649316 86980 649322 86992
rect 660666 86980 660672 86992
rect 660724 86980 660730 87032
rect 650822 86844 650828 86896
rect 650880 86884 650886 86896
rect 658826 86884 658832 86896
rect 650880 86856 658832 86884
rect 650880 86844 650886 86856
rect 658826 86844 658832 86856
rect 658884 86844 658890 86896
rect 659562 86844 659568 86896
rect 659620 86884 659626 86896
rect 663242 86884 663248 86896
rect 659620 86856 663248 86884
rect 659620 86844 659626 86856
rect 663242 86844 663248 86856
rect 663300 86844 663306 86896
rect 652018 86708 652024 86760
rect 652076 86748 652082 86760
rect 662506 86748 662512 86760
rect 652076 86720 662512 86748
rect 652076 86708 652082 86720
rect 662506 86708 662512 86720
rect 662564 86708 662570 86760
rect 578602 86572 578608 86624
rect 578660 86612 578666 86624
rect 580442 86612 580448 86624
rect 578660 86584 580448 86612
rect 578660 86572 578666 86584
rect 580442 86572 580448 86584
rect 580500 86572 580506 86624
rect 650638 86572 650644 86624
rect 650696 86612 650702 86624
rect 661402 86612 661408 86624
rect 650696 86584 661408 86612
rect 650696 86572 650702 86584
rect 661402 86572 661408 86584
rect 661460 86572 661466 86624
rect 623038 86436 623044 86488
rect 623096 86476 623102 86488
rect 626442 86476 626448 86488
rect 623096 86448 626448 86476
rect 623096 86436 623102 86448
rect 626442 86436 626448 86448
rect 626500 86436 626506 86488
rect 653398 86300 653404 86352
rect 653456 86340 653462 86352
rect 660114 86340 660120 86352
rect 653456 86312 660120 86340
rect 653456 86300 653462 86312
rect 660114 86300 660120 86312
rect 660172 86300 660178 86352
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 579246 84124 579252 84176
rect 579304 84164 579310 84176
rect 581822 84164 581828 84176
rect 579304 84136 581828 84164
rect 579304 84124 579310 84136
rect 581822 84124 581828 84136
rect 581880 84124 581886 84176
rect 621658 84124 621664 84176
rect 621716 84164 621722 84176
rect 625614 84164 625620 84176
rect 621716 84136 625620 84164
rect 621716 84124 621722 84136
rect 625614 84124 625620 84136
rect 625672 84124 625678 84176
rect 579246 82764 579252 82816
rect 579304 82804 579310 82816
rect 588538 82804 588544 82816
rect 579304 82776 588544 82804
rect 579304 82764 579310 82776
rect 588538 82764 588544 82776
rect 588596 82764 588602 82816
rect 628650 80928 628656 80980
rect 628708 80968 628714 80980
rect 642450 80968 642456 80980
rect 628708 80940 642456 80968
rect 628708 80928 628714 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 614022 80792 614028 80844
rect 614080 80832 614086 80844
rect 647326 80832 647332 80844
rect 614080 80804 647332 80832
rect 614080 80792 614086 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 578970 80656 578976 80708
rect 579028 80696 579034 80708
rect 589918 80696 589924 80708
rect 579028 80668 589924 80696
rect 579028 80656 579034 80668
rect 589918 80656 589924 80668
rect 589976 80656 589982 80708
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636102 80696 636108 80708
rect 595496 80668 636108 80696
rect 595496 80656 595502 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 579154 80044 579160 80096
rect 579212 80084 579218 80096
rect 585962 80084 585968 80096
rect 579212 80056 585968 80084
rect 579212 80044 579218 80056
rect 585962 80044 585968 80056
rect 586020 80044 586026 80096
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 638862 79472 638868 79484
rect 629260 79444 638868 79472
rect 629260 79432 629266 79444
rect 638862 79432 638868 79444
rect 638920 79432 638926 79484
rect 616138 79296 616144 79348
rect 616196 79336 616202 79348
rect 648982 79336 648988 79348
rect 616196 79308 648988 79336
rect 616196 79296 616202 79308
rect 648982 79296 648988 79308
rect 649040 79296 649046 79348
rect 638862 78276 638868 78328
rect 638920 78316 638926 78328
rect 645302 78316 645308 78328
rect 638920 78288 645308 78316
rect 638920 78276 638926 78288
rect 645302 78276 645308 78288
rect 645360 78276 645366 78328
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 639046 78112 639052 78124
rect 631100 78084 639052 78112
rect 631100 78072 631106 78084
rect 639046 78072 639052 78084
rect 639104 78072 639110 78124
rect 612642 77936 612648 77988
rect 612700 77976 612706 77988
rect 647510 77976 647516 77988
rect 612700 77948 647516 77976
rect 612700 77936 612706 77948
rect 647510 77936 647516 77948
rect 647568 77936 647574 77988
rect 633894 77432 633900 77444
rect 625126 77404 633900 77432
rect 623038 77256 623044 77308
rect 623096 77296 623102 77308
rect 625126 77296 625154 77404
rect 633894 77392 633900 77404
rect 633952 77392 633958 77444
rect 623096 77268 625154 77296
rect 623096 77256 623102 77268
rect 628374 77256 628380 77308
rect 628432 77296 628438 77308
rect 631502 77296 631508 77308
rect 628432 77268 631508 77296
rect 628432 77256 628438 77268
rect 631502 77256 631508 77268
rect 631560 77256 631566 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 649166 76820 649172 76832
rect 620336 76792 649172 76820
rect 620336 76780 620342 76792
rect 649166 76780 649172 76792
rect 649224 76780 649230 76832
rect 611998 76644 612004 76696
rect 612056 76684 612062 76696
rect 647050 76684 647056 76696
rect 612056 76656 647056 76684
rect 612056 76644 612062 76656
rect 647050 76644 647056 76656
rect 647108 76644 647114 76696
rect 606478 76508 606484 76560
rect 606536 76548 606542 76560
rect 662414 76548 662420 76560
rect 606536 76520 662420 76548
rect 606536 76508 606542 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 578878 75896 578884 75948
rect 578936 75936 578942 75948
rect 631042 75936 631048 75948
rect 578936 75908 631048 75936
rect 578936 75896 578942 75908
rect 631042 75896 631048 75908
rect 631100 75896 631106 75948
rect 578694 75420 578700 75472
rect 578752 75460 578758 75472
rect 581638 75460 581644 75472
rect 578752 75432 581644 75460
rect 578752 75420 578758 75432
rect 581638 75420 581644 75432
rect 581696 75420 581702 75472
rect 618898 75148 618904 75200
rect 618956 75188 618962 75200
rect 646866 75188 646872 75200
rect 618956 75160 646872 75188
rect 618956 75148 618962 75160
rect 646866 75148 646872 75160
rect 646924 75148 646930 75200
rect 588538 74808 588544 74860
rect 588596 74848 588602 74860
rect 628006 74848 628012 74860
rect 588596 74820 628012 74848
rect 588596 74808 588602 74820
rect 628006 74808 628012 74820
rect 628064 74808 628070 74860
rect 578510 73108 578516 73160
rect 578568 73148 578574 73160
rect 580258 73148 580264 73160
rect 578568 73120 580264 73148
rect 578568 73108 578574 73120
rect 580258 73108 580264 73120
rect 580316 73108 580322 73160
rect 579522 67600 579528 67652
rect 579580 67640 579586 67652
rect 624418 67640 624424 67652
rect 579580 67612 624424 67640
rect 579580 67600 579586 67612
rect 624418 67600 624424 67612
rect 624476 67600 624482 67652
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 605834 66280 605840 66292
rect 579580 66252 605840 66280
rect 579580 66240 579586 66252
rect 605834 66240 605840 66252
rect 605892 66240 605898 66292
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 613378 64852 613384 64864
rect 579580 64824 613384 64852
rect 579580 64812 579586 64824
rect 613378 64812 613384 64824
rect 613436 64812 613442 64864
rect 578510 62024 578516 62076
rect 578568 62064 578574 62076
rect 664438 62064 664444 62076
rect 578568 62036 664444 62064
rect 578568 62024 578574 62036
rect 664438 62024 664444 62036
rect 664496 62024 664502 62076
rect 579522 60664 579528 60716
rect 579580 60704 579586 60716
rect 614850 60704 614856 60716
rect 579580 60676 614856 60704
rect 579580 60664 579586 60676
rect 614850 60664 614856 60676
rect 614908 60664 614914 60716
rect 581638 59984 581644 60036
rect 581696 60024 581702 60036
rect 603074 60024 603080 60036
rect 581696 59996 603080 60024
rect 581696 59984 581702 59996
rect 603074 59984 603080 59996
rect 603132 59984 603138 60036
rect 580258 58760 580264 58812
rect 580316 58800 580322 58812
rect 601878 58800 601884 58812
rect 580316 58772 601884 58800
rect 580316 58760 580322 58772
rect 601878 58760 601884 58772
rect 601936 58760 601942 58812
rect 577682 58624 577688 58676
rect 577740 58664 577746 58676
rect 604454 58664 604460 58676
rect 577740 58636 604460 58664
rect 577740 58624 577746 58636
rect 604454 58624 604460 58636
rect 604512 58624 604518 58676
rect 605834 58624 605840 58676
rect 605892 58664 605898 58676
rect 663794 58664 663800 58676
rect 605892 58636 663800 58664
rect 605892 58624 605898 58636
rect 663794 58624 663800 58636
rect 663852 58624 663858 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 666554 57916 666560 57928
rect 579580 57888 666560 57916
rect 579580 57876 579586 57888
rect 666554 57876 666560 57888
rect 666612 57876 666618 57928
rect 575474 57196 575480 57248
rect 575532 57236 575538 57248
rect 600314 57236 600320 57248
rect 575532 57208 600320 57236
rect 575532 57196 575538 57208
rect 600314 57196 600320 57208
rect 600372 57196 600378 57248
rect 579522 56516 579528 56568
rect 579580 56556 579586 56568
rect 588538 56556 588544 56568
rect 579580 56528 588544 56556
rect 579580 56516 579586 56528
rect 588538 56516 588544 56528
rect 588596 56516 588602 56568
rect 574922 56108 574928 56160
rect 574980 56148 574986 56160
rect 597922 56148 597928 56160
rect 574980 56120 597928 56148
rect 574980 56108 574986 56120
rect 597922 56108 597928 56120
rect 597980 56108 597986 56160
rect 574554 55972 574560 56024
rect 574612 56012 574618 56024
rect 598934 56012 598940 56024
rect 574612 55984 598940 56012
rect 574612 55972 574618 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 599118 55876 599124 55888
rect 574796 55848 599124 55876
rect 574796 55836 574802 55848
rect 599118 55836 599124 55848
rect 599176 55836 599182 55888
rect 624418 55836 624424 55888
rect 624476 55876 624482 55888
rect 663978 55876 663984 55888
rect 624476 55848 663984 55876
rect 624476 55836 624482 55848
rect 663978 55836 663984 55848
rect 664036 55836 664042 55888
rect 574002 55564 574008 55616
rect 574060 55604 574066 55616
rect 596450 55604 596456 55616
rect 574060 55576 596456 55604
rect 574060 55564 574066 55576
rect 596450 55564 596456 55576
rect 596508 55564 596514 55616
rect 462378 55372 467144 55400
rect 459480 55168 462314 55196
rect 459480 53644 459508 55168
rect 462286 55128 462314 55168
rect 462378 55128 462406 55372
rect 462286 55100 462406 55128
rect 465000 55236 466500 55264
rect 465000 54448 465028 55236
rect 465552 55100 466132 55128
rect 465552 54856 465580 55100
rect 466104 54924 466132 55100
rect 466472 55060 466500 55236
rect 467116 55196 467144 55372
rect 574738 55196 574744 55208
rect 467116 55168 574744 55196
rect 574738 55156 574744 55168
rect 574796 55156 574802 55208
rect 578878 55060 578884 55072
rect 466472 55032 578884 55060
rect 578878 55020 578884 55032
rect 578936 55020 578942 55072
rect 585778 54924 585784 54936
rect 466104 54896 585784 54924
rect 585778 54884 585784 54896
rect 585836 54884 585842 54936
rect 460400 54420 465028 54448
rect 465276 54828 465580 54856
rect 460400 53644 460428 54420
rect 463160 53808 463694 53836
rect 463160 53644 463188 53808
rect 463666 53644 463694 53808
rect 465276 53768 465304 54828
rect 596174 54788 596180 54800
rect 466012 54760 596180 54788
rect 466012 54720 466040 54760
rect 596174 54748 596180 54760
rect 596232 54748 596238 54800
rect 465460 54692 465764 54720
rect 465460 53836 465488 54692
rect 465736 54652 465764 54692
rect 465920 54692 466040 54720
rect 465920 54652 465948 54692
rect 597554 54652 597560 54664
rect 465736 54624 465948 54652
rect 468864 54624 597560 54652
rect 468864 54516 468892 54624
rect 597554 54612 597560 54624
rect 597612 54612 597618 54664
rect 623038 54516 623044 54528
rect 465184 53740 465304 53768
rect 465368 53808 465488 53836
rect 465552 54488 468892 54516
rect 470566 54488 623044 54516
rect 465184 53644 465212 53740
rect 465368 53644 465396 53808
rect 465552 53644 465580 54488
rect 470566 54380 470594 54488
rect 623038 54476 623044 54488
rect 623096 54476 623102 54528
rect 577498 54380 577504 54392
rect 465736 54352 470594 54380
rect 471992 54352 577504 54380
rect 465736 53644 465764 54352
rect 471992 54312 472020 54352
rect 577498 54340 577504 54352
rect 577556 54340 577562 54392
rect 471900 54284 472020 54312
rect 471900 53644 471928 54284
rect 574554 54244 574560 54256
rect 472268 54216 574560 54244
rect 472268 54176 472296 54216
rect 574554 54204 574560 54216
rect 574612 54204 574618 54256
rect 472176 54148 472296 54176
rect 472176 54108 472204 54148
rect 575474 54108 575480 54120
rect 472084 54080 472204 54108
rect 472636 54080 575480 54108
rect 459462 53592 459468 53644
rect 459520 53592 459526 53644
rect 460382 53592 460388 53644
rect 460440 53592 460446 53644
rect 462268 53592 462274 53644
rect 462326 53632 462332 53644
rect 462958 53632 462964 53644
rect 462326 53604 462964 53632
rect 462326 53592 462332 53604
rect 462958 53592 462964 53604
rect 463016 53592 463022 53644
rect 463142 53592 463148 53644
rect 463200 53592 463206 53644
rect 463648 53592 463654 53644
rect 463706 53592 463712 53644
rect 465166 53592 465172 53644
rect 465224 53592 465230 53644
rect 465350 53592 465356 53644
rect 465408 53592 465414 53644
rect 465534 53592 465540 53644
rect 465592 53592 465598 53644
rect 465718 53592 465724 53644
rect 465776 53592 465782 53644
rect 471882 53592 471888 53644
rect 471940 53592 471946 53644
rect 461302 53456 461308 53508
rect 461360 53496 461366 53508
rect 472084 53496 472112 54080
rect 472636 53904 472664 54080
rect 575474 54068 575480 54080
rect 575532 54068 575538 54120
rect 574922 53972 574928 53984
rect 472268 53876 472664 53904
rect 472820 53944 574928 53972
rect 472268 53644 472296 53876
rect 472820 53768 472848 53944
rect 574922 53932 574928 53944
rect 574980 53932 574986 53984
rect 574002 53836 574008 53848
rect 472452 53740 472848 53768
rect 473326 53808 574008 53836
rect 472452 53644 472480 53740
rect 472250 53592 472256 53644
rect 472308 53592 472314 53644
rect 472434 53592 472440 53644
rect 472492 53592 472498 53644
rect 472618 53592 472624 53644
rect 472676 53632 472682 53644
rect 473326 53632 473354 53808
rect 574002 53796 574008 53808
rect 574060 53796 574066 53848
rect 472676 53604 473354 53632
rect 472676 53592 472682 53604
rect 461360 53468 472112 53496
rect 461360 53456 461366 53468
rect 50522 53320 50528 53372
rect 50580 53360 50586 53372
rect 128998 53360 129004 53372
rect 50580 53332 129004 53360
rect 50580 53320 50586 53332
rect 128998 53320 129004 53332
rect 129056 53320 129062 53372
rect 464522 53320 464528 53372
rect 464580 53360 464586 53372
rect 465534 53360 465540 53372
rect 464580 53332 465540 53360
rect 464580 53320 464586 53332
rect 465534 53320 465540 53332
rect 465592 53320 465598 53372
rect 47762 53184 47768 53236
rect 47820 53224 47826 53236
rect 130378 53224 130384 53236
rect 47820 53196 130384 53224
rect 47820 53184 47826 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 463602 53184 463608 53236
rect 463660 53224 463666 53236
rect 472434 53224 472440 53236
rect 463660 53196 472440 53224
rect 463660 53184 463666 53196
rect 472434 53184 472440 53196
rect 472492 53184 472498 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 130562 53088 130568 53100
rect 46256 53060 130568 53088
rect 46256 53048 46262 53060
rect 130562 53048 130568 53060
rect 130620 53048 130626 53100
rect 464982 53048 464988 53100
rect 465040 53088 465046 53100
rect 465350 53088 465356 53100
rect 465040 53060 465356 53088
rect 465040 53048 465046 53060
rect 465350 53048 465356 53060
rect 465408 53048 465414 53100
rect 463740 52776 463746 52828
rect 463798 52816 463804 52828
rect 472618 52816 472624 52828
rect 463798 52788 472624 52816
rect 463798 52776 463804 52788
rect 472618 52776 472624 52788
rect 472676 52776 472682 52828
rect 145374 52436 145380 52488
rect 145432 52476 145438 52488
rect 306006 52476 306012 52488
rect 145432 52448 306012 52476
rect 145432 52436 145438 52448
rect 306006 52436 306012 52448
rect 306064 52436 306070 52488
rect 50706 51960 50712 52012
rect 50764 52000 50770 52012
rect 130746 52000 130752 52012
rect 50764 51972 130752 52000
rect 50764 51960 50770 51972
rect 130746 51960 130752 51972
rect 130804 51960 130810 52012
rect 48958 51824 48964 51876
rect 49016 51864 49022 51876
rect 129458 51864 129464 51876
rect 49016 51836 129464 51864
rect 49016 51824 49022 51836
rect 129458 51824 129464 51836
rect 129516 51824 129522 51876
rect 49142 51688 49148 51740
rect 49200 51728 49206 51740
rect 126882 51728 126888 51740
rect 49200 51700 126888 51728
rect 49200 51688 49206 51700
rect 126882 51688 126888 51700
rect 126940 51688 126946 51740
rect 126882 50736 126888 50788
rect 126940 50776 126946 50788
rect 129274 50776 129280 50788
rect 126940 50748 129280 50776
rect 126940 50736 126946 50748
rect 129274 50736 129280 50748
rect 129332 50736 129338 50788
rect 50338 50464 50344 50516
rect 50396 50504 50402 50516
rect 128630 50504 128636 50516
rect 50396 50476 128636 50504
rect 50396 50464 50402 50476
rect 128630 50464 128636 50476
rect 128688 50464 128694 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 128998 50368 129004 50380
rect 45520 50340 129004 50368
rect 45520 50328 45526 50340
rect 128998 50328 129004 50340
rect 129056 50328 129062 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 128446 49144 128452 49156
rect 51776 49116 128452 49144
rect 51776 49104 51782 49116
rect 128446 49104 128452 49116
rect 128504 49104 128510 49156
rect 47578 48968 47584 49020
rect 47636 49008 47642 49020
rect 129642 49008 129648 49020
rect 47636 48980 129648 49008
rect 47636 48968 47642 48980
rect 129642 48968 129648 48980
rect 129700 48968 129706 49020
rect 128630 48084 128636 48136
rect 128688 48124 128694 48136
rect 132126 48124 132132 48136
rect 128688 48096 132132 48124
rect 128688 48084 128694 48096
rect 132126 48084 132132 48096
rect 132184 48084 132190 48136
rect 129182 47676 129188 47728
rect 129240 47716 129246 47728
rect 131850 47716 131856 47728
rect 129240 47688 131856 47716
rect 129240 47676 129246 47688
rect 131850 47676 131856 47688
rect 131908 47676 131914 47728
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 130856 45064 131146 45076
rect 129608 45048 131146 45064
rect 129608 45036 130884 45048
rect 129608 45024 129614 45036
rect 131316 44964 131376 44992
rect 129734 44888 129740 44940
rect 129792 44928 129798 44940
rect 131316 44928 131344 44964
rect 129792 44900 131344 44928
rect 129792 44888 129798 44900
rect 131592 44792 131620 44894
rect 131546 44764 131620 44792
rect 131730 44796 131790 44824
rect 131546 44740 131574 44764
rect 131500 44724 131574 44740
rect 131408 44712 131574 44724
rect 131408 44696 131528 44712
rect 128446 44616 128452 44668
rect 128504 44656 128510 44668
rect 131408 44656 131436 44696
rect 128504 44628 131436 44656
rect 128504 44616 128510 44628
rect 129366 44480 129372 44532
rect 129424 44520 129430 44532
rect 131730 44520 131758 44796
rect 131960 44724 131988 44726
rect 131868 44696 131988 44724
rect 131868 44600 131896 44696
rect 131850 44548 131856 44600
rect 131908 44548 131914 44600
rect 132236 44520 132264 44642
rect 129424 44492 131758 44520
rect 132144 44500 132264 44520
rect 129424 44480 129430 44492
rect 132126 44448 132132 44500
rect 132184 44492 132264 44500
rect 132184 44448 132190 44492
rect 132420 44464 132448 44558
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 130746 44276 130752 44328
rect 130804 44316 130810 44328
rect 132604 44316 132632 44474
rect 130804 44288 132632 44316
rect 130804 44276 130810 44288
rect 128998 44140 129004 44192
rect 129056 44180 129062 44192
rect 132218 44180 132224 44192
rect 129056 44152 132224 44180
rect 129056 44140 129062 44152
rect 132218 44140 132224 44152
rect 132276 44140 132282 44192
rect 132788 44180 132816 44362
rect 132420 44152 132816 44180
rect 130562 44004 130568 44056
rect 130620 44044 130626 44056
rect 132420 44044 132448 44152
rect 130620 44016 132448 44044
rect 130620 44004 130626 44016
rect 130378 43868 130384 43920
rect 130436 43908 130442 43920
rect 132972 43908 133000 44250
rect 130436 43880 133000 43908
rect 130436 43868 130442 43880
rect 43438 42780 43444 42832
rect 43496 42820 43502 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43496 42792 133184 42820
rect 43496 42780 43502 42792
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 307352 42724 369256 42752
rect 307352 42712 307358 42724
rect 369228 42616 369256 42724
rect 369394 42712 369400 42764
rect 369452 42752 369458 42764
rect 431218 42752 431224 42764
rect 369452 42724 431224 42752
rect 369452 42712 369458 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 464338 42752 464344 42764
rect 456116 42724 464344 42752
rect 456116 42712 456122 42724
rect 464338 42712 464344 42724
rect 464396 42712 464402 42764
rect 427078 42616 427084 42628
rect 369228 42588 427084 42616
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 455874 42576 455880 42628
rect 455932 42616 455938 42628
rect 463970 42616 463976 42628
rect 455932 42588 463976 42616
rect 455932 42576 455938 42588
rect 463970 42576 463976 42588
rect 464028 42576 464034 42628
rect 361758 42440 361764 42492
rect 361816 42480 361822 42492
rect 369394 42480 369400 42492
rect 361816 42452 369400 42480
rect 361816 42440 361822 42452
rect 369394 42440 369400 42452
rect 369452 42440 369458 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 308950 42173 308956 42225
rect 309008 42173 309014 42225
rect 427078 42032 427084 42084
rect 427136 42072 427142 42084
rect 427136 42044 427814 42072
rect 427136 42032 427142 42044
rect 427786 41936 427814 42044
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 455874 41936 455880 41948
rect 427786 41908 455880 41936
rect 455874 41896 455880 41908
rect 455932 41896 455938 41948
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 510344 1007156 510396 1007208
rect 518164 1007156 518216 1007208
rect 431684 1007088 431736 1007140
rect 434628 1007088 434680 1007140
rect 505008 1007020 505060 1007072
rect 515588 1007020 515640 1007072
rect 428004 1006952 428056 1007004
rect 359740 1006884 359792 1006936
rect 374644 1006884 374696 1006936
rect 428372 1006816 428424 1006868
rect 436744 1006816 436796 1006868
rect 145564 1006748 145616 1006800
rect 151728 1006748 151780 1006800
rect 359372 1006748 359424 1006800
rect 369124 1006748 369176 1006800
rect 429200 1006680 429252 1006732
rect 552296 1006952 552348 1007004
rect 568028 1006952 568080 1007004
rect 505376 1006884 505428 1006936
rect 510344 1006884 510396 1006936
rect 510528 1006816 510580 1006868
rect 520924 1006816 520976 1006868
rect 557172 1006748 557224 1006800
rect 565268 1006748 565320 1006800
rect 145748 1006612 145800 1006664
rect 360568 1006612 360620 1006664
rect 371884 1006612 371936 1006664
rect 152096 1006544 152148 1006596
rect 157432 1006544 157484 1006596
rect 166264 1006544 166316 1006596
rect 451832 1006680 451884 1006732
rect 505376 1006612 505428 1006664
rect 514208 1006612 514260 1006664
rect 553124 1006612 553176 1006664
rect 562508 1006612 562560 1006664
rect 469864 1006544 469916 1006596
rect 144184 1006476 144236 1006528
rect 151268 1006476 151320 1006528
rect 551100 1006476 551152 1006528
rect 556620 1006476 556672 1006528
rect 556804 1006476 556856 1006528
rect 564440 1006476 564492 1006528
rect 94688 1006408 94740 1006460
rect 101128 1006408 101180 1006460
rect 158628 1006408 158680 1006460
rect 173164 1006408 173216 1006460
rect 249248 1006408 249300 1006460
rect 255320 1006408 255372 1006460
rect 361396 1006408 361448 1006460
rect 376760 1006408 376812 1006460
rect 422668 1006408 422720 1006460
rect 148508 1006340 148560 1006392
rect 96068 1006272 96120 1006324
rect 101956 1006272 102008 1006324
rect 108488 1006272 108540 1006324
rect 126244 1006272 126296 1006324
rect 144368 1006204 144420 1006256
rect 150900 1006204 150952 1006256
rect 93308 1006136 93360 1006188
rect 99472 1006136 99524 1006188
rect 102968 1006136 103020 1006188
rect 104808 1006136 104860 1006188
rect 106832 1006136 106884 1006188
rect 113824 1006136 113876 1006188
rect 153936 1006272 153988 1006324
rect 158260 1006272 158312 1006324
rect 159456 1006272 159508 1006324
rect 177304 1006272 177356 1006324
rect 249064 1006272 249116 1006324
rect 254124 1006272 254176 1006324
rect 301504 1006272 301556 1006324
rect 306932 1006272 306984 1006324
rect 314660 1006272 314712 1006324
rect 319444 1006272 319496 1006324
rect 354864 1006272 354916 1006324
rect 153752 1006136 153804 1006188
rect 160284 1006136 160336 1006188
rect 164884 1006136 164936 1006188
rect 166264 1006136 166316 1006188
rect 175924 1006136 175976 1006188
rect 210424 1006136 210476 1006188
rect 228364 1006136 228416 1006188
rect 262680 1006136 262732 1006188
rect 279424 1006136 279476 1006188
rect 298744 1006136 298796 1006188
rect 304908 1006136 304960 1006188
rect 355692 1006136 355744 1006188
rect 363604 1006136 363656 1006188
rect 365076 1006136 365128 1006188
rect 367744 1006136 367796 1006188
rect 369124 1006272 369176 1006324
rect 380164 1006272 380216 1006324
rect 373264 1006136 373316 1006188
rect 402244 1006136 402296 1006188
rect 431684 1006272 431736 1006324
rect 436744 1006408 436796 1006460
rect 448520 1006408 448572 1006460
rect 513564 1006408 513616 1006460
rect 519544 1006408 519596 1006460
rect 507860 1006340 507912 1006392
rect 510528 1006340 510580 1006392
rect 555424 1006340 555476 1006392
rect 558828 1006340 558880 1006392
rect 456800 1006272 456852 1006324
rect 506204 1006204 506256 1006256
rect 522304 1006272 522356 1006324
rect 553952 1006204 554004 1006256
rect 571984 1006272 572036 1006324
rect 148876 1006068 148928 1006120
rect 150072 1006068 150124 1006120
rect 93124 1006000 93176 1006052
rect 96068 1006000 96120 1006052
rect 96252 1006000 96304 1006052
rect 98276 1006000 98328 1006052
rect 101404 1006000 101456 1006052
rect 103980 1006000 104032 1006052
rect 106004 1006000 106056 1006052
rect 124864 1006000 124916 1006052
rect 158260 1006000 158312 1006052
rect 171784 1006000 171836 1006052
rect 198188 1006000 198240 1006052
rect 201040 1006000 201092 1006052
rect 208400 1006000 208452 1006052
rect 229744 1006000 229796 1006052
rect 251088 1006000 251140 1006052
rect 252468 1006000 252520 1006052
rect 261852 1006000 261904 1006052
rect 280804 1006000 280856 1006052
rect 298928 1006000 298980 1006052
rect 311808 1006000 311860 1006052
rect 314660 1006000 314712 1006052
rect 320824 1006000 320876 1006052
rect 363420 1006000 363472 1006052
rect 382924 1006000 382976 1006052
rect 400864 1006000 400916 1006052
rect 429200 1006136 429252 1006188
rect 434628 1006136 434680 1006188
rect 471428 1006136 471480 1006188
rect 514208 1006136 514260 1006188
rect 522488 1006136 522540 1006188
rect 562508 1006136 562560 1006188
rect 570604 1006136 570656 1006188
rect 425520 1006000 425572 1006052
rect 429200 1006000 429252 1006052
rect 430028 1006000 430080 1006052
rect 471244 1006000 471296 1006052
rect 496728 1006000 496780 1006052
rect 498844 1006000 498896 1006052
rect 500500 1006000 500552 1006052
rect 513564 1006000 513616 1006052
rect 554320 1006000 554372 1006052
rect 574744 1006000 574796 1006052
rect 509056 1005864 509108 1005916
rect 514024 1005864 514076 1005916
rect 564440 1005864 564492 1005916
rect 567844 1005864 567896 1005916
rect 427544 1005660 427596 1005712
rect 440884 1005660 440936 1005712
rect 428372 1005524 428424 1005576
rect 446404 1005524 446456 1005576
rect 360568 1005388 360620 1005440
rect 378784 1005388 378836 1005440
rect 423496 1005388 423548 1005440
rect 464344 1005388 464396 1005440
rect 555976 1005388 556028 1005440
rect 573364 1005388 573416 1005440
rect 102784 1005252 102836 1005304
rect 108856 1005252 108908 1005304
rect 204904 1005252 204956 1005304
rect 212080 1005252 212132 1005304
rect 357716 1005252 357768 1005304
rect 375380 1005252 375432 1005304
rect 424324 1005252 424376 1005304
rect 465724 1005252 465776 1005304
rect 498844 1005252 498896 1005304
rect 516784 1005252 516836 1005304
rect 149704 1005048 149756 1005100
rect 152924 1005048 152976 1005100
rect 354588 1005048 354640 1005100
rect 356520 1005048 356572 1005100
rect 365076 1005048 365128 1005100
rect 370504 1005048 370556 1005100
rect 551468 1005048 551520 1005100
rect 569224 1005048 569276 1005100
rect 151084 1004912 151136 1004964
rect 153752 1004912 153804 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 263048 1004912 263100 1004964
rect 268384 1004912 268436 1004964
rect 353208 1004912 353260 1004964
rect 355692 1004912 355744 1004964
rect 361396 1004912 361448 1004964
rect 364984 1004912 365036 1004964
rect 422024 1004912 422076 1004964
rect 423496 1004912 423548 1004964
rect 149888 1004776 149940 1004828
rect 152924 1004776 152976 1004828
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 211252 1004776 211304 1004828
rect 215944 1004776 215996 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 362592 1004776 362644 1004828
rect 365168 1004776 365220 1004828
rect 420828 1004776 420880 1004828
rect 422668 1004776 422720 1004828
rect 430856 1004776 430908 1004828
rect 433984 1004912 434036 1004964
rect 498108 1004912 498160 1004964
rect 499672 1004912 499724 1004964
rect 508228 1004912 508280 1004964
rect 511264 1004912 511316 1004964
rect 560852 1004912 560904 1004964
rect 566464 1004912 566516 1004964
rect 432052 1004776 432104 1004828
rect 436744 1004776 436796 1004828
rect 499304 1004776 499356 1004828
rect 501328 1004776 501380 1004828
rect 507032 1004776 507084 1004828
rect 509884 1004776 509936 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 151268 1004640 151320 1004692
rect 154120 1004640 154172 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 430028 1004640 430080 1004692
rect 431960 1004640 432012 1004692
rect 432880 1004640 432932 1004692
rect 438124 1004640 438176 1004692
rect 503352 1004640 503404 1004692
rect 507308 1004640 507360 1004692
rect 508228 1004640 508280 1004692
rect 510620 1004640 510672 1004692
rect 557632 1004640 557684 1004692
rect 559472 1004640 559524 1004692
rect 560852 1004640 560904 1004692
rect 565084 1004640 565136 1004692
rect 422208 1004572 422260 1004624
rect 424324 1004572 424376 1004624
rect 499488 1004572 499540 1004624
rect 500500 1004572 500552 1004624
rect 510068 1004504 510120 1004556
rect 515404 1004504 515456 1004556
rect 425520 1004164 425572 1004216
rect 449164 1004164 449216 1004216
rect 451832 1004164 451884 1004216
rect 467564 1004164 467616 1004216
rect 425152 1004028 425204 1004080
rect 454868 1004028 454920 1004080
rect 456800 1004028 456852 1004080
rect 422208 1003892 422260 1003944
rect 458824 1003892 458876 1003944
rect 502524 1004028 502576 1004080
rect 514668 1004028 514720 1004080
rect 461584 1003892 461636 1003944
rect 499488 1003892 499540 1003944
rect 518348 1003892 518400 1003944
rect 422024 1003484 422076 1003536
rect 423772 1003484 423824 1003536
rect 448520 1003280 448572 1003332
rect 451648 1003280 451700 1003332
rect 97448 1002736 97500 1002788
rect 102324 1002736 102376 1002788
rect 94504 1002600 94556 1002652
rect 100300 1002600 100352 1002652
rect 253480 1002600 253532 1002652
rect 256148 1002600 256200 1002652
rect 100024 1002464 100076 1002516
rect 103152 1002464 103204 1002516
rect 252008 1002464 252060 1002516
rect 255320 1002464 255372 1002516
rect 261024 1002464 261076 1002516
rect 264244 1002464 264296 1002516
rect 558000 1002464 558052 1002516
rect 560944 1002464 560996 1002516
rect 555148 1002396 555200 1002448
rect 557540 1002396 557592 1002448
rect 97264 1002328 97316 1002380
rect 100300 1002328 100352 1002380
rect 107660 1002328 107712 1002380
rect 109500 1002328 109552 1002380
rect 253020 1002328 253072 1002380
rect 256148 1002328 256200 1002380
rect 558828 1002328 558880 1002380
rect 562508 1002328 562560 1002380
rect 98644 1002192 98696 1002244
rect 101956 1002192 102008 1002244
rect 105636 1002192 105688 1002244
rect 107844 1002192 107896 1002244
rect 108028 1002192 108080 1002244
rect 110420 1002192 110472 1002244
rect 155776 1002192 155828 1002244
rect 158720 1002192 158772 1002244
rect 203524 1002192 203576 1002244
rect 206376 1002192 206428 1002244
rect 206744 1002192 206796 1002244
rect 208400 1002192 208452 1002244
rect 210884 1002192 210936 1002244
rect 213184 1002192 213236 1002244
rect 251824 1002192 251876 1002244
rect 254492 1002192 254544 1002244
rect 358544 1002192 358596 1002244
rect 360844 1002192 360896 1002244
rect 423588 1002192 423640 1002244
rect 426348 1002192 426400 1002244
rect 501696 1002192 501748 1002244
rect 504364 1002192 504416 1002244
rect 551928 1002192 551980 1002244
rect 554320 1002192 554372 1002244
rect 558000 1002192 558052 1002244
rect 560300 1002192 560352 1002244
rect 560484 1002192 560536 1002244
rect 563060 1002192 563112 1002244
rect 96068 1002056 96120 1002108
rect 99104 1002056 99156 1002108
rect 100208 1002056 100260 1002108
rect 103152 1002056 103204 1002108
rect 103980 1002056 104032 1002108
rect 106464 1002056 106516 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111800 1002056 111852 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 152464 1002056 152516 1002108
rect 154580 1002056 154632 1002108
rect 205088 1002056 205140 1002108
rect 207204 1002056 207256 1002108
rect 212540 1002056 212592 1002108
rect 214564 1002056 214616 1002108
rect 263508 1002056 263560 1002108
rect 265624 1002056 265676 1002108
rect 300308 1002056 300360 1002108
rect 305276 1002056 305328 1002108
rect 310152 1002056 310204 1002108
rect 311900 1002056 311952 1002108
rect 355784 1002056 355836 1002108
rect 356520 1002056 356572 1002108
rect 504548 1002056 504600 1002108
rect 507124 1002056 507176 1002108
rect 559656 1002056 559708 1002108
rect 561496 1002056 561548 1002108
rect 561680 1002056 561732 1002108
rect 563704 1002056 563756 1002108
rect 95884 1001920 95936 1001972
rect 98276 1001920 98328 1001972
rect 98828 1001920 98880 1001972
rect 101128 1001920 101180 1001972
rect 106004 1001920 106056 1001972
rect 107752 1001920 107804 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 155776 1001920 155828 1001972
rect 157340 1001920 157392 1001972
rect 157800 1001920 157852 1001972
rect 160100 1001920 160152 1001972
rect 202972 1001920 203024 1001972
rect 205548 1001920 205600 1001972
rect 210884 1001920 210936 1001972
rect 212540 1001920 212592 1001972
rect 261024 1001920 261076 1001972
rect 263600 1001920 263652 1001972
rect 263876 1001920 263928 1001972
rect 267004 1001920 267056 1001972
rect 310980 1001920 311032 1001972
rect 313280 1001920 313332 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 360200 1001920 360252 1001972
rect 362224 1001920 362276 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 425704 1001920 425756 1001972
rect 427176 1001920 427228 1001972
rect 433340 1001920 433392 1001972
rect 435364 1001920 435416 1001972
rect 500868 1001920 500920 1001972
rect 501696 1001920 501748 1001972
rect 501880 1001920 501932 1001972
rect 503352 1001920 503404 1001972
rect 504180 1001920 504232 1001972
rect 505744 1001920 505796 1001972
rect 510344 1001920 510396 1001972
rect 512644 1001920 512696 1001972
rect 560024 1001920 560076 1001972
rect 562324 1001920 562376 1001972
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 423772 1001172 423824 1001224
rect 456800 1001172 456852 1001224
rect 498108 1001172 498160 1001224
rect 520372 1001172 520424 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 423588 1000900 423640 1000952
rect 429384 1000900 429436 1000952
rect 298100 1000492 298152 1000544
rect 308956 1000492 309008 1000544
rect 375380 1000492 375432 1000544
rect 383292 1000492 383344 1000544
rect 92756 999744 92808 999796
rect 102968 999744 103020 999796
rect 360844 999744 360896 999796
rect 369860 999744 369912 999796
rect 373264 999064 373316 999116
rect 374644 999064 374696 999116
rect 565268 999064 565320 999116
rect 568212 999064 568264 999116
rect 196624 998996 196676 999048
rect 204352 998996 204404 999048
rect 467564 998860 467616 998912
rect 472624 998860 472676 998912
rect 200764 998724 200816 998776
rect 203892 998724 203944 998776
rect 378784 998724 378836 998776
rect 383568 998724 383620 998776
rect 426532 998656 426584 998708
rect 466460 998656 466512 998708
rect 515588 998656 515640 998708
rect 523868 998656 523920 998708
rect 197820 998588 197872 998640
rect 202696 998588 202748 998640
rect 376760 998588 376812 998640
rect 383476 998588 383528 998640
rect 247224 998520 247276 998572
rect 256976 998520 257028 998572
rect 429384 998520 429436 998572
rect 472440 998520 472492 998572
rect 514668 998520 514720 998572
rect 524052 998520 524104 998572
rect 553124 998520 553176 998572
rect 565820 998520 565872 998572
rect 200948 998452 201000 998504
rect 203892 998452 203944 998504
rect 304264 998452 304316 998504
rect 307300 998452 307352 998504
rect 92388 998384 92440 998436
rect 100208 998384 100260 998436
rect 247408 998384 247460 998436
rect 259000 998384 259052 998436
rect 351828 998384 351880 998436
rect 382280 998384 382332 998436
rect 429200 998384 429252 998436
rect 472256 998384 472308 998436
rect 499304 998384 499356 998436
rect 517520 998384 517572 998436
rect 552296 998384 552348 998436
rect 572720 998384 572772 998436
rect 200212 998316 200264 998368
rect 202972 998316 203024 998368
rect 303068 998316 303120 998368
rect 306104 998316 306156 998368
rect 247040 998248 247092 998300
rect 253664 998248 253716 998300
rect 304448 998180 304500 998232
rect 306932 998180 306984 998232
rect 568028 998180 568080 998232
rect 572904 998180 572956 998232
rect 198004 998112 198056 998164
rect 201868 998112 201920 998164
rect 202144 998112 202196 998164
rect 205548 998112 205600 998164
rect 246764 998112 246816 998164
rect 251088 998112 251140 998164
rect 258172 998112 258224 998164
rect 259460 998112 259512 998164
rect 92572 998044 92624 998096
rect 96252 998044 96304 998096
rect 260196 998044 260248 998096
rect 262864 998044 262916 998096
rect 305644 998044 305696 998096
rect 307760 998044 307812 998096
rect 308404 998044 308456 998096
rect 310612 998044 310664 998096
rect 199384 997976 199436 998028
rect 202696 997976 202748 998028
rect 250444 997976 250496 998028
rect 253296 997976 253348 998028
rect 254584 997976 254636 998028
rect 256516 997976 256568 998028
rect 259828 997908 259880 997960
rect 262220 997908 262272 997960
rect 307208 997908 307260 997960
rect 308956 997908 309008 997960
rect 591304 997908 591356 997960
rect 625804 997908 625856 997960
rect 198372 997840 198424 997892
rect 200672 997840 200724 997892
rect 247684 997840 247736 997892
rect 252468 997840 252520 997892
rect 256332 997840 256384 997892
rect 257344 997840 257396 997892
rect 202328 997772 202380 997824
rect 204720 997772 204772 997824
rect 260196 997772 260248 997824
rect 260932 997772 260984 997824
rect 302884 997772 302936 997824
rect 306104 997772 306156 997824
rect 307024 997772 307076 997824
rect 308128 997772 308180 997824
rect 549168 997772 549220 997824
rect 551468 997772 551520 997824
rect 590844 997772 590896 997824
rect 625620 997772 625672 997824
rect 93492 997704 93544 997756
rect 106464 997704 106516 997756
rect 113824 997704 113876 997756
rect 117136 997704 117188 997756
rect 143724 997704 143776 997756
rect 160100 997704 160152 997756
rect 246580 997704 246632 997756
rect 256332 997704 256384 997756
rect 359464 997704 359516 997756
rect 372344 997704 372396 997756
rect 425704 997704 425756 997756
rect 439688 997704 439740 997756
rect 507308 997704 507360 997756
rect 516876 997704 516928 997756
rect 195244 997636 195296 997688
rect 198372 997636 198424 997688
rect 540888 997636 540940 997688
rect 555424 997636 555476 997688
rect 573364 997636 573416 997688
rect 623688 997636 623740 997688
rect 109500 997568 109552 997620
rect 116216 997568 116268 997620
rect 144184 997500 144236 997552
rect 153936 997568 153988 997620
rect 369860 997568 369912 997620
rect 372528 997568 372580 997620
rect 433984 997568 434036 997620
rect 439872 997568 439924 997620
rect 509884 997568 509936 997620
rect 517060 997568 517112 997620
rect 551928 997500 551980 997552
rect 591304 997500 591356 997552
rect 502340 997432 502392 997484
rect 516692 997432 516744 997484
rect 571984 997364 572036 997416
rect 590568 997364 590620 997416
rect 488908 997296 488960 997348
rect 510620 997296 510672 997348
rect 565820 997296 565872 997348
rect 570236 997296 570288 997348
rect 200212 997228 200264 997280
rect 205088 997228 205140 997280
rect 574744 997228 574796 997280
rect 590844 997228 590896 997280
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 557540 997160 557592 997212
rect 570788 997160 570840 997212
rect 399944 997092 399996 997144
rect 431960 997092 432012 997144
rect 144552 997024 144604 997076
rect 158720 997024 158772 997076
rect 320824 997024 320876 997076
rect 332600 997024 332652 997076
rect 505744 997024 505796 997076
rect 517704 997024 517756 997076
rect 549168 997024 549220 997076
rect 617156 997024 617208 997076
rect 365168 996956 365220 997008
rect 372712 996956 372764 997008
rect 572720 996888 572772 996940
rect 590384 996888 590436 996940
rect 558184 996752 558236 996804
rect 590568 996684 590620 996736
rect 143724 996480 143776 996532
rect 151268 996480 151320 996532
rect 92940 996344 92992 996396
rect 121736 996344 121788 996396
rect 144184 996344 144236 996396
rect 149888 996344 149940 996396
rect 549444 996344 549496 996396
rect 550640 996344 550692 996396
rect 253204 996208 253256 996260
rect 263600 996208 263652 996260
rect 368940 996208 368992 996260
rect 377588 996208 377640 996260
rect 171784 996072 171836 996124
rect 211160 996072 211212 996124
rect 211804 996072 211856 996124
rect 260932 996072 260984 996124
rect 279424 996072 279476 996124
rect 316040 996072 316092 996124
rect 354588 996072 354640 996124
rect 366364 996072 366416 996124
rect 144368 995936 144420 995988
rect 168748 995936 168800 995988
rect 171508 995936 171560 995988
rect 177304 995936 177356 995988
rect 212540 995936 212592 995988
rect 229744 995936 229796 995988
rect 136456 995800 136508 995852
rect 168564 995800 168616 995852
rect 171232 995800 171284 995852
rect 213184 995800 213236 995852
rect 255412 995800 255464 995852
rect 264244 995936 264296 995988
rect 298928 995936 298980 995988
rect 382740 995936 382792 995988
rect 402244 996072 402296 996124
rect 511264 996072 511316 996124
rect 563060 996072 563112 996124
rect 522304 995868 522356 995920
rect 560300 995936 560352 995988
rect 570604 995936 570656 995988
rect 262220 995800 262272 995852
rect 262864 995800 262916 995852
rect 313280 995800 313332 995852
rect 355784 995800 355836 995852
rect 368940 995800 368992 995852
rect 369308 995800 369360 995852
rect 383108 995800 383160 995852
rect 506204 995800 506256 995852
rect 509056 995800 509108 995852
rect 540244 995800 540296 995852
rect 561680 995800 561732 995852
rect 562140 995800 562192 995852
rect 625620 995800 625672 995852
rect 642088 995868 642140 995920
rect 92204 995528 92256 995580
rect 92756 995528 92808 995580
rect 170680 995528 170732 995580
rect 194968 995528 195020 995580
rect 201684 995528 201736 995580
rect 255412 995528 255464 995580
rect 261852 995528 261904 995580
rect 299572 995528 299624 995580
rect 301688 995528 301740 995580
rect 364984 995528 365036 995580
rect 369308 995528 369360 995580
rect 377588 995528 377640 995580
rect 246212 995460 246264 995512
rect 247224 995460 247276 995512
rect 300124 995392 300176 995444
rect 304080 995392 304132 995444
rect 380164 995528 380216 995580
rect 383292 995528 383344 995580
rect 383476 995528 383528 995580
rect 385592 995528 385644 995580
rect 472624 995528 472676 995580
rect 473360 995528 473412 995580
rect 524052 995528 524104 995580
rect 525340 995528 525392 995580
rect 554688 995528 554740 995580
rect 562140 995528 562192 995580
rect 623688 995528 623740 995580
rect 626540 995528 626592 995580
rect 388812 995392 388864 995444
rect 389824 995392 389876 995444
rect 171692 995277 171744 995329
rect 180708 995324 180760 995376
rect 182640 995324 182692 995376
rect 185124 995324 185176 995376
rect 186780 995324 186832 995376
rect 193128 995324 193180 995376
rect 198188 995324 198240 995376
rect 228364 995324 228416 995376
rect 253204 995324 253256 995376
rect 296168 995324 296220 995376
rect 298284 995324 298336 995376
rect 415400 995392 415452 995444
rect 398932 995324 398984 995376
rect 374644 995256 374696 995308
rect 171508 995165 171560 995217
rect 178868 995188 178920 995240
rect 180340 995188 180392 995240
rect 180478 995188 180530 995240
rect 202144 995188 202196 995240
rect 235586 995188 235638 995240
rect 253020 995188 253072 995240
rect 397644 995256 397696 995308
rect 416136 995235 416188 995287
rect 362224 995120 362276 995172
rect 387524 995120 387576 995172
rect 532148 995120 532200 995172
rect 540244 995120 540296 995172
rect 171232 995053 171284 995105
rect 180156 995052 180208 995104
rect 206284 995052 206336 995104
rect 235264 995052 235316 995104
rect 253480 995052 253532 995104
rect 282828 995052 282880 995104
rect 311900 995052 311952 995104
rect 451648 995052 451700 995104
rect 485964 995052 486016 995104
rect 507124 995052 507176 995104
rect 528192 995052 528244 995104
rect 556620 995052 556672 995104
rect 639512 995052 639564 995104
rect 357440 994984 357492 995036
rect 395160 994984 395212 995036
rect 180708 994916 180760 994968
rect 208400 994916 208452 994968
rect 232872 994916 232924 994968
rect 256056 994916 256108 994968
rect 283472 994916 283524 994968
rect 307024 994916 307076 994968
rect 474556 994916 474608 994968
rect 482928 994916 482980 994968
rect 486608 994916 486660 994968
rect 489920 994916 489972 994968
rect 519820 994916 519872 994968
rect 530216 994916 530268 994968
rect 534356 994916 534408 994968
rect 538128 994916 538180 994968
rect 570788 994916 570840 994968
rect 640708 994916 640760 994968
rect 78312 994780 78364 994832
rect 104164 994780 104216 994832
rect 132132 994780 132184 994832
rect 142988 994780 143040 994832
rect 143172 994780 143224 994832
rect 155960 994780 156012 994832
rect 171048 994829 171100 994881
rect 171232 994829 171284 994881
rect 371884 994848 371936 994900
rect 397000 994848 397052 994900
rect 286508 994780 286560 994832
rect 305644 994780 305696 994832
rect 458824 994780 458876 994832
rect 482284 994780 482336 994832
rect 501880 994780 501932 994832
rect 539232 994780 539284 994832
rect 567844 994780 567896 994832
rect 639052 994780 639104 994832
rect 168564 994712 168616 994764
rect 250444 994712 250496 994764
rect 363604 994712 363656 994764
rect 393964 994712 394016 994764
rect 81348 994644 81400 994696
rect 98644 994644 98696 994696
rect 129740 994644 129792 994696
rect 134892 994644 134944 994696
rect 77668 994508 77720 994560
rect 97448 994508 97500 994560
rect 128452 994508 128504 994560
rect 157340 994644 157392 994696
rect 284116 994644 284168 994696
rect 308404 994644 308456 994696
rect 419448 994644 419500 994696
rect 660580 994983 660632 995035
rect 168748 994576 168800 994628
rect 243084 994576 243136 994628
rect 244188 994576 244240 994628
rect 246764 994576 246816 994628
rect 356060 994576 356112 994628
rect 393320 994576 393372 994628
rect 660764 994576 660816 994628
rect 80704 994372 80756 994424
rect 93124 994372 93176 994424
rect 131580 994372 131632 994424
rect 154580 994508 154632 994560
rect 420828 994508 420880 994560
rect 590568 994508 590620 994560
rect 625620 994508 625672 994560
rect 633992 994508 634044 994560
rect 660948 994508 661000 994560
rect 168932 994440 168984 994492
rect 298744 994440 298796 994492
rect 383292 994440 383344 994492
rect 389824 994440 389876 994492
rect 129096 994236 129148 994288
rect 142804 994372 142856 994424
rect 142988 994372 143040 994424
rect 148508 994372 148560 994424
rect 461584 994372 461636 994424
rect 186780 994304 186832 994356
rect 194968 994304 195020 994356
rect 232228 994304 232280 994356
rect 254584 994304 254636 994356
rect 382740 994304 382792 994356
rect 392676 994304 392728 994356
rect 134892 994100 134944 994152
rect 143172 994236 143224 994288
rect 186504 994236 186556 994288
rect 295340 994236 295392 994288
rect 381176 994236 381228 994288
rect 396356 994236 396408 994288
rect 446128 994236 446180 994288
rect 456800 994236 456852 994288
rect 474556 994236 474608 994288
rect 475384 994372 475436 994424
rect 487804 994372 487856 994424
rect 496728 994372 496780 994424
rect 519820 994372 519872 994424
rect 523684 994372 523736 994424
rect 538312 994372 538364 994424
rect 489920 994236 489972 994288
rect 500868 994236 500920 994288
rect 144920 994100 144972 994152
rect 169392 994032 169444 994084
rect 300124 994100 300176 994152
rect 466460 994100 466512 994152
rect 475384 994100 475436 994152
rect 518348 994100 518400 994152
rect 523684 994100 523736 994152
rect 530216 994236 530268 994288
rect 537668 994236 537720 994288
rect 550640 994236 550692 994288
rect 572720 994236 572772 994288
rect 535552 994100 535604 994152
rect 574100 994032 574152 994084
rect 142804 993964 142856 994016
rect 151084 993964 151136 994016
rect 180340 993964 180392 994016
rect 196624 993964 196676 994016
rect 243912 993964 243964 994016
rect 247408 993964 247460 994016
rect 569224 993896 569276 993948
rect 243084 993828 243136 993880
rect 247684 993828 247736 993880
rect 171232 993760 171284 993812
rect 195244 993760 195296 993812
rect 520372 993760 520424 993812
rect 660948 993760 661000 993812
rect 171048 993624 171100 993676
rect 198004 993624 198056 993676
rect 517244 993624 517296 993676
rect 660764 993624 660816 993676
rect 164884 993420 164936 993472
rect 169760 993420 169812 993472
rect 214564 993420 214616 993472
rect 219440 993420 219492 993472
rect 50344 993148 50396 993200
rect 107752 993148 107804 993200
rect 44824 993012 44876 993064
rect 109040 993012 109092 993064
rect 138020 993012 138072 993064
rect 163136 993012 163188 993064
rect 318064 993012 318116 993064
rect 349160 993012 349212 993064
rect 562508 993012 562560 993064
rect 660304 993012 660356 993064
rect 54484 992876 54536 992928
rect 148324 992876 148376 992928
rect 319444 992876 319496 992928
rect 364984 992876 365036 992928
rect 367744 992876 367796 992928
rect 429936 992876 429988 992928
rect 435364 992876 435416 992928
rect 478972 992876 479024 992928
rect 560944 992876 560996 992928
rect 668584 992876 668636 992928
rect 638868 992264 638920 992316
rect 640800 992264 640852 992316
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 51724 991584 51776 991636
rect 110420 991584 110472 991636
rect 55864 991448 55916 991500
rect 146944 991448 146996 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 369124 991448 369176 991500
rect 414112 991448 414164 991500
rect 512644 991448 512696 991500
rect 543832 991448 543884 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 53288 990224 53340 990276
rect 95884 990224 95936 990276
rect 48964 990088 49016 990140
rect 108120 990088 108172 990140
rect 562324 990088 562376 990140
rect 669964 990088 670016 990140
rect 572720 989476 572772 989528
rect 576308 989476 576360 989528
rect 89628 987368 89680 987420
rect 111800 987368 111852 987420
rect 563704 987368 563756 987420
rect 608784 987368 608836 987420
rect 203156 986620 203208 986672
rect 204904 986620 204956 986672
rect 438124 986076 438176 986128
rect 462780 986076 462832 986128
rect 515404 986076 515456 986128
rect 527640 986076 527692 986128
rect 566464 986076 566516 986128
rect 592500 986076 592552 986128
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 370504 985940 370556 985992
rect 397828 985940 397880 985992
rect 436744 985940 436796 985992
rect 495164 985940 495216 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 672724 975672 672776 975724
rect 46204 961868 46256 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952348 36596 952400
rect 41696 952348 41748 952400
rect 33784 951464 33836 951516
rect 41512 951464 41564 951516
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 663064 948064 663116 948116
rect 45560 945956 45612 946008
rect 62120 945956 62172 946008
rect 28724 945276 28776 945328
rect 31760 945276 31812 945328
rect 35808 942556 35860 942608
rect 41604 942556 41656 942608
rect 35808 941196 35860 941248
rect 41420 941196 41472 941248
rect 35808 939768 35860 939820
rect 41604 939768 41656 939820
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 663064 921816 663116 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 665824 909440 665876 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 671344 895636 671396 895688
rect 44088 892712 44140 892764
rect 42938 892270 42990 892322
rect 43076 892202 43128 892254
rect 44088 891896 44140 891948
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 652392 855584 652444 855636
rect 664444 855584 664496 855636
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 651840 841780 651892 841832
rect 669964 841780 670016 841832
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 35808 817028 35860 817080
rect 41696 817028 41748 817080
rect 35808 815600 35860 815652
rect 41420 815600 41472 815652
rect 651472 815600 651524 815652
rect 661684 815600 661736 815652
rect 35808 814240 35860 814292
rect 41604 814240 41656 814292
rect 41328 811452 41380 811504
rect 41696 811452 41748 811504
rect 40592 808528 40644 808580
rect 41604 808528 41656 808580
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 35164 802408 35216 802460
rect 41696 802408 41748 802460
rect 35900 802272 35952 802324
rect 41696 802272 41748 802324
rect 53104 793568 53156 793620
rect 62120 793568 62172 793620
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 652392 775548 652444 775600
rect 668400 775548 668452 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35532 768952 35584 769004
rect 40040 768952 40092 769004
rect 35348 768816 35400 768868
rect 41696 768816 41748 768868
rect 35808 768680 35860 768732
rect 41328 768680 41380 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35532 767320 35584 767372
rect 37924 767320 37976 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 37096 763240 37148 763292
rect 39304 763240 39356 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 672172 761880 672224 761932
rect 672724 761880 672776 761932
rect 31024 759636 31076 759688
rect 39120 759636 39172 759688
rect 37924 759024 37976 759076
rect 41512 759024 41564 759076
rect 35164 758276 35216 758328
rect 41696 758276 41748 758328
rect 676036 757120 676088 757172
rect 676588 757120 676640 757172
rect 675852 754264 675904 754316
rect 683120 754264 683172 754316
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 35808 730056 35860 730108
rect 41696 730056 41748 730108
rect 673368 728560 673420 728612
rect 670700 728424 670752 728476
rect 673368 728288 673420 728340
rect 673368 728084 673420 728136
rect 41328 725908 41380 725960
rect 41696 725908 41748 725960
rect 41328 724480 41380 724532
rect 41696 724480 41748 724532
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 33784 715776 33836 715828
rect 41696 715776 41748 715828
rect 33048 715640 33100 715692
rect 41144 715640 41196 715692
rect 31668 715504 31720 715556
rect 41696 715504 41748 715556
rect 36544 714824 36596 714876
rect 41696 714824 41748 714876
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 651472 709316 651524 709368
rect 664444 709316 664496 709368
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 651472 696940 651524 696992
rect 661868 696940 661920 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 41328 687216 41380 687268
rect 41696 687216 41748 687268
rect 41328 683136 41380 683188
rect 41696 683136 41748 683188
rect 651656 683136 651708 683188
rect 669964 683136 670016 683188
rect 41328 681844 41380 681896
rect 41696 681844 41748 681896
rect 40040 677968 40092 678020
rect 41696 677968 41748 678020
rect 51724 674840 51776 674892
rect 62120 674840 62172 674892
rect 35164 672732 35216 672784
rect 40132 672732 40184 672784
rect 36728 672052 36780 672104
rect 41512 672052 41564 672104
rect 39948 671712 40000 671764
rect 41696 671712 41748 671764
rect 651472 669332 651524 669384
rect 661684 669332 661736 669384
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651472 656888 651524 656940
rect 663064 656888 663116 656940
rect 46204 647844 46256 647896
rect 62120 647844 62172 647896
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639072 35860 639124
rect 40040 639072 40092 639124
rect 35624 638936 35676 638988
rect 41512 638936 41564 638988
rect 35808 637576 35860 637628
rect 40040 637576 40092 637628
rect 35808 636216 35860 636268
rect 41696 636216 41748 636268
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 40040 635876 40092 635928
rect 41696 635876 41748 635928
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651472 629280 651524 629332
rect 667204 629280 667256 629332
rect 675852 626560 675904 626612
rect 676496 626560 676548 626612
rect 673368 623976 673420 624028
rect 673368 623840 673420 623892
rect 50344 623772 50396 623824
rect 62120 623772 62172 623824
rect 672632 620984 672684 621036
rect 673000 620984 673052 621036
rect 672264 618332 672316 618384
rect 672908 618332 672960 618384
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 43812 612892 43864 612944
rect 43720 612688 43772 612740
rect 43996 612552 44048 612604
rect 43582 612280 43634 612332
rect 43720 612280 43772 612332
rect 46020 611872 46072 611924
rect 47952 611668 48004 611720
rect 46940 611464 46992 611516
rect 44155 611260 44207 611312
rect 44379 611056 44431 611108
rect 44272 610920 44324 610972
rect 44502 610716 44554 610768
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 664628 603100 664680 603152
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 41236 594668 41288 594720
rect 41512 594668 41564 594720
rect 676036 591336 676088 591388
rect 682384 591336 682436 591388
rect 652392 590656 652444 590708
rect 658924 590656 658976 590708
rect 40500 589636 40552 589688
rect 41696 589636 41748 589688
rect 33784 585760 33836 585812
rect 39672 585760 39724 585812
rect 37924 585284 37976 585336
rect 41420 585284 41472 585336
rect 36544 585148 36596 585200
rect 40224 585148 40276 585200
rect 51724 583720 51776 583772
rect 62120 583720 62172 583772
rect 651472 576852 651524 576904
rect 666008 576852 666060 576904
rect 651656 563048 651708 563100
rect 659108 563048 659160 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 35808 557540 35860 557592
rect 41512 557540 41564 557592
rect 35808 554752 35860 554804
rect 41696 554752 41748 554804
rect 35808 553528 35860 553580
rect 41420 553528 41472 553580
rect 35624 553392 35676 553444
rect 41696 553392 41748 553444
rect 41236 550740 41288 550792
rect 41696 550740 41748 550792
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 41236 549244 41288 549296
rect 41696 549312 41748 549364
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 675944 547612 675996 547664
rect 678244 547612 678296 547664
rect 31760 547408 31812 547460
rect 37188 547408 37240 547460
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 33784 542988 33836 543040
rect 41512 542988 41564 543040
rect 37188 542308 37240 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669964 536800 670016 536852
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 672724 532108 672776 532160
rect 674012 532108 674064 532160
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 676036 518780 676088 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 675852 503616 675904 503668
rect 681004 503616 681056 503668
rect 675852 499536 675904 499588
rect 679624 499536 679676 499588
rect 652576 494708 652628 494760
rect 665824 494708 665876 494760
rect 675852 492668 675904 492720
rect 683120 492668 683172 492720
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 651472 484440 651524 484492
rect 670148 484372 670200 484424
rect 675852 480360 675904 480412
rect 683120 480360 683172 480412
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 675852 476076 675904 476128
rect 680360 476076 680412 476128
rect 651472 470568 651524 470620
rect 663064 470568 663116 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 676128 457444 676180 457496
rect 676312 457444 676364 457496
rect 676864 457444 676916 457496
rect 676128 457172 676180 457224
rect 652392 456764 652444 456816
rect 667204 456764 667256 456816
rect 673184 456764 673236 456816
rect 675852 456084 675904 456136
rect 677140 456084 677192 456136
rect 673828 456016 673880 456068
rect 673736 455812 673788 455864
rect 673460 455540 673512 455592
rect 673506 455336 673558 455388
rect 672080 455200 672132 455252
rect 673388 455132 673440 455184
rect 673164 454928 673216 454980
rect 673046 454792 673098 454844
rect 672816 454384 672868 454436
rect 672954 454180 673006 454232
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672264 453908 672316 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 671344 430584 671396 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 41328 423784 41380 423836
rect 41696 423784 41748 423836
rect 40960 423172 41012 423224
rect 41604 423172 41656 423224
rect 651840 416780 651892 416832
rect 661684 416780 661736 416832
rect 49148 415420 49200 415472
rect 62120 415420 62172 415472
rect 36544 415352 36596 415404
rect 41696 415352 41748 415404
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 41144 387064 41196 387116
rect 41696 387064 41748 387116
rect 41328 382372 41380 382424
rect 41696 382372 41748 382424
rect 41144 382236 41196 382288
rect 41696 382236 41748 382288
rect 35808 379516 35860 379568
rect 41696 379516 41748 379568
rect 35808 375980 35860 376032
rect 39488 375980 39540 376032
rect 51724 375368 51776 375420
rect 62120 375368 62172 375420
rect 28908 371832 28960 371884
rect 41696 371832 41748 371884
rect 651656 364352 651708 364404
rect 663248 364352 663300 364404
rect 46388 362924 46440 362976
rect 62120 362924 62172 362976
rect 45008 355784 45060 355836
rect 45652 355784 45704 355836
rect 44640 355648 44692 355700
rect 44575 354832 44627 354884
rect 44575 354628 44627 354680
rect 44799 354424 44851 354476
rect 44686 354288 44738 354340
rect 45652 354016 45704 354068
rect 45928 353744 45980 353796
rect 45560 353200 45612 353252
rect 651472 350548 651524 350600
rect 667388 350548 667440 350600
rect 28908 345040 28960 345092
rect 38292 345040 38344 345092
rect 35808 339464 35860 339516
rect 37924 339464 37976 339516
rect 651472 338104 651524 338156
rect 666376 338104 666428 338156
rect 50344 336744 50396 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 666652 324300 666704 324352
rect 53104 310496 53156 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667204 310496 667256 310548
rect 676036 304852 676088 304904
rect 676312 304852 676364 304904
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675852 298052 675904 298104
rect 678980 298052 679032 298104
rect 676036 297032 676088 297084
rect 681004 297032 681056 297084
rect 41328 285064 41380 285116
rect 41696 285064 41748 285116
rect 32404 284928 32456 284980
rect 41696 284928 41748 284980
rect 651472 284316 651524 284368
rect 667572 284316 667624 284368
rect 88340 275952 88392 276004
rect 143356 275952 143408 276004
rect 156880 275952 156932 276004
rect 193864 275952 193916 276004
rect 201776 275952 201828 276004
rect 222108 275952 222160 276004
rect 389180 275952 389232 276004
rect 393320 275952 393372 276004
rect 413100 275952 413152 276004
rect 434720 275952 434772 276004
rect 437480 275952 437532 276004
rect 450084 275952 450136 276004
rect 456800 275952 456852 276004
rect 460664 275952 460716 276004
rect 460848 275952 460900 276004
rect 502064 275952 502116 276004
rect 510252 275952 510304 276004
rect 597836 275952 597888 276004
rect 95424 275816 95476 275868
rect 104808 275816 104860 275868
rect 113180 275816 113232 275868
rect 169944 275816 169996 275868
rect 181720 275816 181772 275868
rect 218888 275816 218940 275868
rect 396356 275816 396408 275868
rect 412272 275816 412324 275868
rect 416412 275816 416464 275868
rect 463056 275816 463108 275868
rect 471152 275816 471204 275868
rect 493784 275816 493836 275868
rect 493968 275816 494020 275868
rect 497372 275816 497424 275868
rect 498200 275816 498252 275868
rect 81256 275680 81308 275732
rect 88984 275680 89036 275732
rect 103704 275680 103756 275732
rect 160100 275680 160152 275732
rect 178132 275680 178184 275732
rect 216864 275680 216916 275732
rect 370504 275680 370556 275732
rect 388628 275680 388680 275732
rect 410064 275680 410116 275732
rect 428832 275680 428884 275732
rect 433156 275680 433208 275732
rect 487896 275680 487948 275732
rect 488080 275680 488132 275732
rect 498752 275680 498804 275732
rect 504180 275816 504232 275868
rect 509148 275816 509200 275868
rect 512184 275816 512236 275868
rect 519820 275816 519872 275868
rect 505652 275680 505704 275732
rect 507124 275680 507176 275732
rect 512736 275680 512788 275732
rect 512920 275680 512972 275732
rect 516232 275680 516284 275732
rect 516784 275680 516836 275732
rect 604920 275816 604972 275868
rect 520188 275680 520240 275732
rect 525524 275680 525576 275732
rect 525892 275680 525944 275732
rect 527272 275680 527324 275732
rect 527732 275680 527784 275732
rect 612004 275680 612056 275732
rect 76472 275544 76524 275596
rect 86868 275544 86920 275596
rect 96620 275544 96672 275596
rect 156604 275544 156656 275596
rect 163964 275544 164016 275596
rect 202144 275544 202196 275596
rect 221924 275544 221976 275596
rect 233884 275544 233936 275596
rect 236092 275544 236144 275596
rect 255504 275544 255556 275596
rect 350724 275544 350776 275596
rect 361396 275544 361448 275596
rect 361580 275544 361632 275596
rect 385040 275544 385092 275596
rect 388076 275544 388128 275596
rect 418160 275544 418212 275596
rect 418344 275544 418396 275596
rect 435916 275544 435968 275596
rect 439504 275544 439556 275596
rect 494980 275544 495032 275596
rect 496820 275544 496872 275596
rect 538220 275544 538272 275596
rect 85948 275408 86000 275460
rect 146760 275408 146812 275460
rect 160468 275408 160520 275460
rect 167736 275408 167788 275460
rect 171048 275408 171100 275460
rect 210424 275408 210476 275460
rect 218336 275408 218388 275460
rect 237380 275408 237432 275460
rect 260932 275408 260984 275460
rect 273536 275408 273588 275460
rect 284576 275408 284628 275460
rect 290096 275408 290148 275460
rect 341524 275408 341576 275460
rect 354312 275408 354364 275460
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 142712 275272 142764 275324
rect 183468 275272 183520 275324
rect 186412 275272 186464 275324
rect 187792 275272 187844 275324
rect 188804 275272 188856 275324
rect 222844 275272 222896 275324
rect 225420 275272 225472 275324
rect 245108 275272 245160 275324
rect 250260 275272 250312 275324
rect 266636 275272 266688 275324
rect 273904 275272 273956 275324
rect 282920 275272 282972 275324
rect 334348 275272 334400 275324
rect 338948 275272 339000 275324
rect 290464 275204 290516 275256
rect 294328 275204 294380 275256
rect 74080 275136 74132 275188
rect 77208 275136 77260 275188
rect 110788 275136 110840 275188
rect 162124 275136 162176 275188
rect 338948 275136 339000 275188
rect 353116 275272 353168 275324
rect 353944 275272 353996 275324
rect 360200 275408 360252 275460
rect 363052 275408 363104 275460
rect 367284 275408 367336 275460
rect 369124 275408 369176 275460
rect 377956 275408 378008 275460
rect 382280 275408 382332 275460
rect 414572 275408 414624 275460
rect 415308 275408 415360 275460
rect 425244 275408 425296 275460
rect 429200 275408 429252 275460
rect 446496 275408 446548 275460
rect 449900 275408 449952 275460
rect 504180 275408 504232 275460
rect 504364 275408 504416 275460
rect 356336 275272 356388 275324
rect 368480 275272 368532 275324
rect 375104 275272 375156 275324
rect 403992 275272 404044 275324
rect 411260 275272 411312 275324
rect 455972 275272 456024 275324
rect 456156 275272 456208 275324
rect 512920 275272 512972 275324
rect 517520 275408 517572 275460
rect 521016 275408 521068 275460
rect 521200 275408 521252 275460
rect 523408 275408 523460 275460
rect 530124 275408 530176 275460
rect 531320 275408 531372 275460
rect 537576 275408 537628 275460
rect 543004 275544 543056 275596
rect 545120 275544 545172 275596
rect 552664 275544 552716 275596
rect 552848 275544 552900 275596
rect 525524 275272 525576 275324
rect 527088 275272 527140 275324
rect 527272 275272 527324 275324
rect 532792 275272 532844 275324
rect 532976 275272 533028 275324
rect 535276 275272 535328 275324
rect 535460 275272 535512 275324
rect 537944 275272 537996 275324
rect 577228 275408 577280 275460
rect 599124 275408 599176 275460
rect 611360 275408 611412 275460
rect 616788 275408 616840 275460
rect 538864 275272 538916 275324
rect 590752 275272 590804 275324
rect 626172 275408 626224 275460
rect 626448 275408 626500 275460
rect 641628 275408 641680 275460
rect 400588 275136 400640 275188
rect 415768 275136 415820 275188
rect 427820 275136 427872 275188
rect 443000 275136 443052 275188
rect 445944 275136 445996 275188
rect 471336 275136 471388 275188
rect 484584 275136 484636 275188
rect 488080 275136 488132 275188
rect 492496 275136 492548 275188
rect 504364 275136 504416 275188
rect 505192 275136 505244 275188
rect 506848 275136 506900 275188
rect 508044 275136 508096 275188
rect 577044 275136 577096 275188
rect 577228 275136 577280 275188
rect 599124 275136 599176 275188
rect 633348 275136 633400 275188
rect 224224 275068 224276 275120
rect 226156 275068 226208 275120
rect 135628 275000 135680 275052
rect 182088 275000 182140 275052
rect 443368 275000 443420 275052
rect 453580 275000 453632 275052
rect 462964 275000 463016 275052
rect 467840 275000 467892 275052
rect 473084 275000 473136 275052
rect 538036 275000 538088 275052
rect 71780 274932 71832 274984
rect 73804 274932 73856 274984
rect 277492 274932 277544 274984
rect 284300 274932 284352 274984
rect 129648 274864 129700 274916
rect 136548 274864 136600 274916
rect 149796 274864 149848 274916
rect 185584 274864 185636 274916
rect 289268 274864 289320 274916
rect 293408 274864 293460 274916
rect 453396 274864 453448 274916
rect 457168 274864 457220 274916
rect 467748 274864 467800 274916
rect 531320 274864 531372 274916
rect 531504 274864 531556 274916
rect 533988 274864 534040 274916
rect 534172 274864 534224 274916
rect 537208 274864 537260 274916
rect 537392 274864 537444 274916
rect 540980 275000 541032 275052
rect 543004 275000 543056 275052
rect 538496 274864 538548 274916
rect 545856 274864 545908 274916
rect 546040 274864 546092 274916
rect 550548 274864 550600 274916
rect 552664 275000 552716 275052
rect 578884 275000 578936 275052
rect 552848 274864 552900 274916
rect 577044 274864 577096 274916
rect 583668 274864 583720 274916
rect 604460 274864 604512 274916
rect 607312 274864 607364 274916
rect 283380 274796 283432 274848
rect 289084 274796 289136 274848
rect 407120 274796 407172 274848
rect 411076 274796 411128 274848
rect 106004 274728 106056 274780
rect 110420 274728 110472 274780
rect 140320 274728 140372 274780
rect 144644 274728 144696 274780
rect 146208 274728 146260 274780
rect 149888 274728 149940 274780
rect 425336 274728 425388 274780
rect 432328 274728 432380 274780
rect 435548 274728 435600 274780
rect 439044 274728 439096 274780
rect 462228 274728 462280 274780
rect 466644 274728 466696 274780
rect 498752 274728 498804 274780
rect 521200 274728 521252 274780
rect 521660 274728 521712 274780
rect 526904 274728 526956 274780
rect 527088 274728 527140 274780
rect 619088 274728 619140 274780
rect 66996 274660 67048 274712
rect 71044 274660 71096 274712
rect 90640 274660 90692 274712
rect 95884 274660 95936 274712
rect 161572 274660 161624 274712
rect 163136 274660 163188 274712
rect 170128 274660 170180 274712
rect 173072 274660 173124 274712
rect 185216 274660 185268 274712
rect 187148 274660 187200 274712
rect 210056 274660 210108 274712
rect 104808 274592 104860 274644
rect 157616 274592 157668 274644
rect 195888 274592 195940 274644
rect 206284 274592 206336 274644
rect 238484 274660 238536 274712
rect 239772 274660 239824 274712
rect 244372 274660 244424 274712
rect 251088 274660 251140 274712
rect 270408 274660 270460 274712
rect 271144 274660 271196 274712
rect 285772 274660 285824 274712
rect 286968 274660 287020 274712
rect 292856 274660 292908 274712
rect 293868 274660 293920 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 298744 274660 298796 274712
rect 300124 274660 300176 274712
rect 321376 274660 321428 274712
rect 328276 274660 328328 274712
rect 331404 274660 331456 274712
rect 335360 274660 335412 274712
rect 360292 274660 360344 274712
rect 363788 274660 363840 274712
rect 367100 274660 367152 274712
rect 369676 274660 369728 274712
rect 386052 274660 386104 274712
rect 389732 274660 389784 274712
rect 404268 274660 404320 274712
rect 407488 274660 407540 274712
rect 409144 274660 409196 274712
rect 409880 274660 409932 274712
rect 488540 274660 488592 274712
rect 492220 274660 492272 274712
rect 494060 274660 494112 274712
rect 498568 274660 498620 274712
rect 619548 274660 619600 274712
rect 623872 274660 623924 274712
rect 410248 274592 410300 274644
rect 437480 274592 437532 274644
rect 440884 274592 440936 274644
rect 486700 274592 486752 274644
rect 498752 274592 498804 274644
rect 571800 274592 571852 274644
rect 121368 274456 121420 274508
rect 176752 274456 176804 274508
rect 182916 274456 182968 274508
rect 199660 274456 199712 274508
rect 237840 274456 237892 274508
rect 362868 274456 362920 274508
rect 386236 274456 386288 274508
rect 395896 274456 395948 274508
rect 413100 274456 413152 274508
rect 427084 274456 427136 274508
rect 477224 274456 477276 274508
rect 101312 274320 101364 274372
rect 160928 274320 160980 274372
rect 187792 274320 187844 274372
rect 220912 274320 220964 274372
rect 237380 274320 237432 274372
rect 243728 274320 243780 274372
rect 384948 274320 385000 274372
rect 419356 274320 419408 274372
rect 424968 274320 425020 274372
rect 474924 274320 474976 274372
rect 476580 274320 476632 274372
rect 491484 274456 491536 274508
rect 492312 274456 492364 274508
rect 496360 274456 496412 274508
rect 496636 274456 496688 274508
rect 577780 274456 577832 274508
rect 585784 274456 585836 274508
rect 477684 274320 477736 274372
rect 528514 274320 528566 274372
rect 528652 274320 528704 274372
rect 538128 274320 538180 274372
rect 538312 274320 538364 274372
rect 586060 274320 586112 274372
rect 601424 274320 601476 274372
rect 82360 274184 82412 274236
rect 145564 274184 145616 274236
rect 160100 274184 160152 274236
rect 164240 274184 164292 274236
rect 176936 274184 176988 274236
rect 214656 274184 214708 274236
rect 220544 274184 220596 274236
rect 240600 274184 240652 274236
rect 342904 274184 342956 274236
rect 347228 274184 347280 274236
rect 366916 274184 366968 274236
rect 389180 274184 389232 274236
rect 390284 274184 390336 274236
rect 426440 274184 426492 274236
rect 438768 274184 438820 274236
rect 496176 274184 496228 274236
rect 496360 274184 496412 274236
rect 498752 274184 498804 274236
rect 501972 274184 502024 274236
rect 84752 274048 84804 274100
rect 148324 274048 148376 274100
rect 158076 274048 158128 274100
rect 200672 274048 200724 274100
rect 206560 274048 206612 274100
rect 235448 274048 235500 274100
rect 239588 274048 239640 274100
rect 258632 274048 258684 274100
rect 346124 274048 346176 274100
rect 362592 274048 362644 274100
rect 377772 274048 377824 274100
rect 408684 274048 408736 274100
rect 413928 274048 413980 274100
rect 456800 274048 456852 274100
rect 459376 274048 459428 274100
rect 523500 274048 523552 274100
rect 523868 274184 523920 274236
rect 602160 274184 602212 274236
rect 602344 274184 602396 274236
rect 608508 274184 608560 274236
rect 528514 274048 528566 274100
rect 528652 274048 528704 274100
rect 619548 274048 619600 274100
rect 77208 273912 77260 273964
rect 143540 273912 143592 273964
rect 145012 273912 145064 273964
rect 192484 273912 192536 273964
rect 193496 273912 193548 273964
rect 226340 273912 226392 273964
rect 234896 273912 234948 273964
rect 255688 273912 255740 273964
rect 256148 273912 256200 273964
rect 270592 273912 270644 273964
rect 271512 273912 271564 273964
rect 280804 273912 280856 273964
rect 331036 273912 331088 273964
rect 342444 273912 342496 273964
rect 360108 273912 360160 273964
rect 383844 273912 383896 273964
rect 385500 273912 385552 273964
rect 395712 273912 395764 273964
rect 405004 273912 405056 273964
rect 444196 273912 444248 273964
rect 451188 273912 451240 273964
rect 513932 273912 513984 273964
rect 514116 273912 514168 273964
rect 523868 273912 523920 273964
rect 524052 273912 524104 273964
rect 613200 273912 613252 273964
rect 123760 273776 123812 273828
rect 177488 273776 177540 273828
rect 406844 273776 406896 273828
rect 410248 273776 410300 273828
rect 428464 273776 428516 273828
rect 458364 273776 458416 273828
rect 465724 273776 465776 273828
rect 482008 273776 482060 273828
rect 491208 273776 491260 273828
rect 570696 273776 570748 273828
rect 280988 273708 281040 273760
rect 287520 273708 287572 273760
rect 134432 273640 134484 273692
rect 185032 273640 185084 273692
rect 457444 273640 457496 273692
rect 484308 273640 484360 273692
rect 487068 273640 487120 273692
rect 563520 273640 563572 273692
rect 570604 273640 570656 273692
rect 587164 273776 587216 273828
rect 613384 273708 613436 273760
rect 615592 273708 615644 273760
rect 144644 273504 144696 273556
rect 187792 273504 187844 273556
rect 475568 273504 475620 273556
rect 477684 273504 477736 273556
rect 482468 273504 482520 273556
rect 558828 273504 558880 273556
rect 481364 273368 481416 273420
rect 556436 273368 556488 273420
rect 347044 273232 347096 273284
rect 349620 273232 349672 273284
rect 350264 273232 350316 273284
rect 356336 273232 356388 273284
rect 114284 273164 114336 273216
rect 169024 273164 169076 273216
rect 104992 273028 105044 273080
rect 163320 273028 163372 273080
rect 167552 273028 167604 273080
rect 184204 273028 184256 273080
rect 187608 273028 187660 273080
rect 211804 273164 211856 273216
rect 419172 273164 419224 273216
rect 462964 273164 463016 273216
rect 473452 273164 473504 273216
rect 496820 273164 496872 273216
rect 500960 273164 501012 273216
rect 581276 273164 581328 273216
rect 211252 273028 211304 273080
rect 220084 273028 220136 273080
rect 397276 273028 397328 273080
rect 418344 273028 418396 273080
rect 426348 273028 426400 273080
rect 478420 273028 478472 273080
rect 485044 273028 485096 273080
rect 492496 273028 492548 273080
rect 493600 273028 493652 273080
rect 574192 273028 574244 273080
rect 580264 273028 580316 273080
rect 640432 273028 640484 273080
rect 78864 272892 78916 272944
rect 138664 272892 138716 272944
rect 141792 272892 141844 272944
rect 189816 272892 189868 272944
rect 191196 272892 191248 272944
rect 224868 272892 224920 272944
rect 288072 272892 288124 272944
rect 290464 272892 290516 272944
rect 373172 272892 373224 272944
rect 382648 272892 382700 272944
rect 391756 272892 391808 272944
rect 410064 272892 410116 272944
rect 412456 272892 412508 272944
rect 453396 272892 453448 272944
rect 458088 272892 458140 272944
rect 521844 272892 521896 272944
rect 94228 272756 94280 272808
rect 156052 272756 156104 272808
rect 180524 272756 180576 272808
rect 217232 272756 217284 272808
rect 228824 272756 228876 272808
rect 249064 272756 249116 272808
rect 352932 272756 352984 272808
rect 372988 272756 373040 272808
rect 380716 272756 380768 272808
rect 396356 272756 396408 272808
rect 403992 272756 404044 272808
rect 429200 272756 429252 272808
rect 434628 272756 434680 272808
rect 488724 272756 488776 272808
rect 496268 272756 496320 272808
rect 528514 272892 528566 272944
rect 528652 272892 528704 272944
rect 611360 272892 611412 272944
rect 87144 272620 87196 272672
rect 152004 272620 152056 272672
rect 168656 272620 168708 272672
rect 208492 272620 208544 272672
rect 217416 272620 217468 272672
rect 242164 272620 242216 272672
rect 242348 272620 242400 272672
rect 259552 272620 259604 272672
rect 333612 272620 333664 272672
rect 344836 272620 344888 272672
rect 368388 272620 368440 272672
rect 393780 272620 393832 272672
rect 393964 272620 394016 272672
rect 406292 272620 406344 272672
rect 408408 272620 408460 272672
rect 452476 272620 452528 272672
rect 453856 272620 453908 272672
rect 516416 272620 516468 272672
rect 516600 272620 516652 272672
rect 606116 272756 606168 272808
rect 524328 272620 524380 272672
rect 527916 272620 527968 272672
rect 528376 272620 528428 272672
rect 614396 272620 614448 272672
rect 77668 272484 77720 272536
rect 145104 272484 145156 272536
rect 152188 272484 152240 272536
rect 197544 272484 197596 272536
rect 199476 272484 199528 272536
rect 230572 272484 230624 272536
rect 231400 272484 231452 272536
rect 252744 272484 252796 272536
rect 252928 272484 252980 272536
rect 267832 272484 267884 272536
rect 268016 272484 268068 272536
rect 278780 272484 278832 272536
rect 279792 272484 279844 272536
rect 287152 272484 287204 272536
rect 322572 272484 322624 272536
rect 330668 272484 330720 272536
rect 338028 272484 338080 272536
rect 351920 272484 351972 272536
rect 358636 272484 358688 272536
rect 380348 272484 380400 272536
rect 382924 272484 382976 272536
rect 413376 272484 413428 272536
rect 415124 272484 415176 272536
rect 461860 272484 461912 272536
rect 463516 272484 463568 272536
rect 528560 272484 528612 272536
rect 529020 272484 529072 272536
rect 538128 272484 538180 272536
rect 538312 272484 538364 272536
rect 632152 272484 632204 272536
rect 127348 272348 127400 272400
rect 179880 272348 179932 272400
rect 451740 272348 451792 272400
rect 139124 272212 139176 272264
rect 141608 272212 141660 272264
rect 143908 272212 143960 272264
rect 190736 272212 190788 272264
rect 447600 272212 447652 272264
rect 470048 272212 470100 272264
rect 471428 272348 471480 272400
rect 485044 272348 485096 272400
rect 488356 272348 488408 272400
rect 567108 272348 567160 272400
rect 578884 272348 578936 272400
rect 594340 272348 594392 272400
rect 153292 272076 153344 272128
rect 171784 272076 171836 272128
rect 463148 272076 463200 272128
rect 471428 272076 471480 272128
rect 487988 272212 488040 272264
rect 565912 272212 565964 272264
rect 480812 272076 480864 272128
rect 483756 272076 483808 272128
rect 560024 272076 560076 272128
rect 470048 271940 470100 271992
rect 473728 271940 473780 271992
rect 478696 271940 478748 271992
rect 552480 271940 552532 271992
rect 552664 271940 552716 271992
rect 580080 271940 580132 271992
rect 110420 271804 110472 271856
rect 164976 271804 165028 271856
rect 175832 271804 175884 271856
rect 207664 271804 207716 271856
rect 214840 271804 214892 271856
rect 221464 271804 221516 271856
rect 222108 271804 222160 271856
rect 232136 271804 232188 271856
rect 381360 271804 381412 271856
rect 399208 271804 399260 271856
rect 411904 271804 411956 271856
rect 438216 271804 438268 271856
rect 443644 271804 443696 271856
rect 500500 271804 500552 271856
rect 500684 271804 500736 271856
rect 508044 271804 508096 271856
rect 508964 271804 509016 271856
rect 596640 271804 596692 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 93032 271668 93084 271720
rect 120724 271668 120776 271720
rect 120908 271668 120960 271720
rect 175280 271668 175332 271720
rect 192300 271668 192352 271720
rect 225512 271668 225564 271720
rect 372528 271668 372580 271720
rect 400404 271668 400456 271720
rect 401324 271668 401376 271720
rect 427820 271668 427872 271720
rect 453304 271668 453356 271720
rect 511540 271668 511592 271720
rect 511908 271668 511960 271720
rect 600228 271668 600280 271720
rect 111984 271532 112036 271584
rect 168380 271532 168432 271584
rect 173440 271532 173492 271584
rect 212632 271532 212684 271584
rect 226156 271532 226208 271584
rect 247224 271532 247276 271584
rect 259736 271532 259788 271584
rect 268384 271532 268436 271584
rect 362224 271532 362276 271584
rect 381176 271532 381228 271584
rect 394332 271532 394384 271584
rect 425336 271532 425388 271584
rect 89720 271396 89772 271448
rect 152648 271396 152700 271448
rect 165160 271396 165212 271448
rect 205732 271396 205784 271448
rect 223580 271396 223632 271448
rect 247408 271396 247460 271448
rect 247868 271396 247920 271448
rect 264336 271396 264388 271448
rect 275100 271396 275152 271448
rect 283472 271396 283524 271448
rect 340604 271396 340656 271448
rect 355140 271396 355192 271448
rect 355324 271396 355376 271448
rect 374368 271396 374420 271448
rect 379428 271396 379480 271448
rect 407120 271396 407172 271448
rect 409788 271396 409840 271448
rect 443368 271532 443420 271584
rect 445668 271532 445720 271584
rect 504548 271532 504600 271584
rect 504732 271532 504784 271584
rect 589372 271532 589424 271584
rect 591304 271532 591356 271584
rect 603724 271532 603776 271584
rect 607864 271532 607916 271584
rect 643928 271532 643980 271584
rect 435364 271396 435416 271448
rect 454500 271396 454552 271448
rect 454684 271396 454736 271448
rect 515128 271396 515180 271448
rect 517336 271396 517388 271448
rect 604460 271396 604512 271448
rect 68192 271260 68244 271312
rect 138480 271260 138532 271312
rect 150992 271260 151044 271312
rect 195980 271260 196032 271312
rect 215944 271260 215996 271312
rect 242072 271260 242124 271312
rect 243176 271260 243228 271312
rect 261024 271260 261076 271312
rect 266820 271260 266872 271312
rect 276664 271260 276716 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 325516 271260 325568 271312
rect 334164 271260 334216 271312
rect 334808 271260 334860 271312
rect 341340 271260 341392 271312
rect 344652 271260 344704 271312
rect 350724 271260 350776 271312
rect 351828 271260 351880 271312
rect 372068 271260 372120 271312
rect 387708 271260 387760 271312
rect 421656 271260 421708 271312
rect 422116 271260 422168 271312
rect 445944 271260 445996 271312
rect 461584 271260 461636 271312
rect 514300 271260 514352 271312
rect 514484 271260 514536 271312
rect 72976 271124 73028 271176
rect 142160 271124 142212 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 208860 271124 208912 271176
rect 237472 271124 237524 271176
rect 240784 271124 240836 271176
rect 259828 271124 259880 271176
rect 262128 271124 262180 271176
rect 274640 271124 274692 271176
rect 276296 271124 276348 271176
rect 284484 271124 284536 271176
rect 328092 271124 328144 271176
rect 337752 271124 337804 271176
rect 342168 271124 342220 271176
rect 356152 271124 356204 271176
rect 364156 271124 364208 271176
rect 386052 271124 386104 271176
rect 431684 271124 431736 271176
rect 484032 271124 484084 271176
rect 484216 271124 484268 271176
rect 519728 271124 519780 271176
rect 519912 271124 519964 271176
rect 523500 271124 523552 271176
rect 523868 271260 523920 271312
rect 610808 271260 610860 271312
rect 621664 271260 621716 271312
rect 636844 271260 636896 271312
rect 538036 271124 538088 271176
rect 538174 271124 538226 271176
rect 625068 271124 625120 271176
rect 356520 271056 356572 271108
rect 359004 271056 359056 271108
rect 128544 270988 128596 271040
rect 181352 270988 181404 271040
rect 190000 270988 190052 271040
rect 216128 270988 216180 271040
rect 389088 270988 389140 271040
rect 415308 270988 415360 271040
rect 439964 270988 440016 271040
rect 493784 270988 493836 271040
rect 499948 270988 500000 271040
rect 500684 270988 500736 271040
rect 507676 270988 507728 271040
rect 593144 270988 593196 271040
rect 130844 270852 130896 270904
rect 182456 270852 182508 270904
rect 200488 270852 200540 270904
rect 224224 270852 224276 270904
rect 416596 270852 416648 270904
rect 463976 270852 464028 270904
rect 464344 270852 464396 270904
rect 519636 270852 519688 270904
rect 520188 270852 520240 270904
rect 523868 270852 523920 270904
rect 526812 270852 526864 270904
rect 621480 270852 621532 270904
rect 137928 270716 137980 270768
rect 187884 270716 187936 270768
rect 418068 270716 418120 270768
rect 462228 270716 462280 270768
rect 464804 270716 464856 270768
rect 484216 270716 484268 270768
rect 484400 270716 484452 270768
rect 485504 270716 485556 270768
rect 489368 270716 489420 270768
rect 551744 270716 551796 270768
rect 116676 270580 116728 270632
rect 151084 270580 151136 270632
rect 237196 270580 237248 270632
rect 115848 270444 115900 270496
rect 171232 270444 171284 270496
rect 172428 270444 172480 270496
rect 209504 270444 209556 270496
rect 233148 270444 233200 270496
rect 237288 270444 237340 270496
rect 400128 270580 400180 270632
rect 435548 270580 435600 270632
rect 437388 270580 437440 270632
rect 471152 270580 471204 270632
rect 474740 270580 474792 270632
rect 538036 270580 538088 270632
rect 538174 270580 538226 270632
rect 591304 270716 591356 270768
rect 110236 270308 110288 270360
rect 167920 270308 167972 270360
rect 173072 270308 173124 270360
rect 210148 270308 210200 270360
rect 213828 270308 213880 270360
rect 240508 270308 240560 270360
rect 249616 270444 249668 270496
rect 253664 270444 253716 270496
rect 291660 270444 291712 270496
rect 295524 270444 295576 270496
rect 297916 270444 297968 270496
rect 299572 270444 299624 270496
rect 299940 270444 299992 270496
rect 300860 270444 300912 270496
rect 359924 270444 359976 270496
rect 376760 270444 376812 270496
rect 377588 270444 377640 270496
rect 391940 270444 391992 270496
rect 396264 270444 396316 270496
rect 423680 270444 423732 270496
rect 429568 270444 429620 270496
rect 480168 270444 480220 270496
rect 480352 270444 480404 270496
rect 485044 270444 485096 270496
rect 486700 270444 486752 270496
rect 494704 270444 494756 270496
rect 494888 270444 494940 270496
rect 560852 270444 560904 270496
rect 252008 270308 252060 270360
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 166908 270172 166960 270224
rect 207388 270172 207440 270224
rect 212448 270172 212500 270224
rect 239956 270172 240008 270224
rect 251088 270172 251140 270224
rect 262312 270308 262364 270360
rect 348424 270308 348476 270360
rect 363052 270308 363104 270360
rect 369400 270308 369452 270360
rect 396080 270308 396132 270360
rect 402060 270308 402112 270360
rect 430580 270308 430632 270360
rect 446956 270308 447008 270360
rect 504916 270308 504968 270360
rect 505054 270308 505106 270360
rect 543188 270308 543240 270360
rect 543372 270308 543424 270360
rect 627920 270308 627972 270360
rect 316960 270240 317012 270292
rect 321560 270240 321612 270292
rect 339316 270240 339368 270292
rect 341524 270240 341576 270292
rect 253848 270172 253900 270224
rect 265072 270172 265124 270224
rect 356704 270172 356756 270224
rect 378140 270172 378192 270224
rect 381544 270172 381596 270224
rect 382280 270172 382332 270224
rect 385684 270172 385736 270224
rect 419540 270172 419592 270224
rect 428280 270172 428332 270224
rect 459560 270172 459612 270224
rect 461860 270172 461912 270224
rect 529204 270172 529256 270224
rect 529664 270172 529716 270224
rect 530768 270172 530820 270224
rect 530952 270172 531004 270224
rect 536104 270172 536156 270224
rect 536288 270172 536340 270224
rect 538036 270172 538088 270224
rect 538174 270172 538226 270224
rect 626632 270172 626684 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 146760 270036 146812 270088
rect 151360 270036 151412 270088
rect 75828 269900 75880 269952
rect 142620 269900 142672 269952
rect 143356 269900 143408 269952
rect 153844 270036 153896 270088
rect 159916 270036 159968 270088
rect 202696 270036 202748 270088
rect 205548 270036 205600 270088
rect 234988 270036 235040 270088
rect 239772 270036 239824 270088
rect 250904 270036 250956 270088
rect 266268 270036 266320 270088
rect 277216 270036 277268 270088
rect 326896 270036 326948 270088
rect 335544 270036 335596 270088
rect 336832 270036 336884 270088
rect 350540 270036 350592 270088
rect 354220 270036 354272 270088
rect 375380 270036 375432 270088
rect 376576 270036 376628 270088
rect 154488 269900 154540 269952
rect 198188 269900 198240 269952
rect 198648 269900 198700 269952
rect 230020 269900 230072 269952
rect 230388 269900 230440 269952
rect 252376 269900 252428 269952
rect 258448 269900 258500 269952
rect 272248 269900 272300 269952
rect 273076 269900 273128 269952
rect 282184 269900 282236 269952
rect 286784 269900 286836 269952
rect 292120 269900 292172 269952
rect 323584 269900 323636 269952
rect 331220 269900 331272 269952
rect 333888 269900 333940 269952
rect 345112 269900 345164 269952
rect 347596 269900 347648 269952
rect 365720 269900 365772 269952
rect 372344 269900 372396 269952
rect 401876 269900 401928 269952
rect 403072 270036 403124 270088
rect 444380 270036 444432 270088
rect 447784 270036 447836 270088
rect 449900 270036 449952 270088
rect 457720 270036 457772 270088
rect 482284 270036 482336 270088
rect 482652 270036 482704 270088
rect 538680 270036 538732 270088
rect 404268 269900 404320 269952
rect 417148 269900 417200 269952
rect 465080 269900 465132 269952
rect 466000 269900 466052 269952
rect 531320 269900 531372 269952
rect 531688 269900 531740 269952
rect 537852 269900 537904 269952
rect 538036 269900 538088 269952
rect 633624 270036 633676 270088
rect 543188 269900 543240 269952
rect 548708 269900 548760 269952
rect 548892 269900 548944 269952
rect 641904 269900 641956 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 139952 269764 140004 269816
rect 181168 269764 181220 269816
rect 182088 269764 182140 269816
rect 186964 269764 187016 269816
rect 187332 269764 187384 269816
rect 191932 269764 191984 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 84108 269628 84160 269680
rect 119804 269628 119856 269680
rect 119068 269492 119120 269544
rect 173716 269628 173768 269680
rect 184756 269628 184808 269680
rect 213828 269628 213880 269680
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 251456 269764 251508 269816
rect 267280 269764 267332 269816
rect 269212 269764 269264 269816
rect 279700 269764 279752 269816
rect 314476 269764 314528 269816
rect 318800 269764 318852 269816
rect 321928 269764 321980 269816
rect 328460 269764 328512 269816
rect 329380 269764 329432 269816
rect 339500 269764 339552 269816
rect 341800 269764 341852 269816
rect 357440 269764 357492 269816
rect 364984 269764 365036 269816
rect 390560 269764 390612 269816
rect 392308 269764 392360 269816
rect 429384 269764 429436 269816
rect 434444 269764 434496 269816
rect 469220 269764 469272 269816
rect 470968 269764 471020 269816
rect 250904 269628 250956 269680
rect 258172 269628 258224 269680
rect 351644 269628 351696 269680
rect 364340 269628 364392 269680
rect 384028 269628 384080 269680
rect 388076 269628 388128 269680
rect 394700 269628 394752 269680
rect 416780 269628 416832 269680
rect 424600 269628 424652 269680
rect 475384 269628 475436 269680
rect 476028 269764 476080 269816
rect 482652 269764 482704 269816
rect 541440 269764 541492 269816
rect 543004 269764 543056 269816
rect 644480 269764 644532 269816
rect 485044 269628 485096 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 187332 269492 187384 269544
rect 208308 269492 208360 269544
rect 230756 269492 230808 269544
rect 390468 269492 390520 269544
rect 118608 269356 118660 269408
rect 166908 269356 166960 269408
rect 335636 269356 335688 269408
rect 343824 269356 343876 269408
rect 401600 269492 401652 269544
rect 426624 269492 426676 269544
rect 427360 269492 427412 269544
rect 475752 269492 475804 269544
rect 402428 269356 402480 269408
rect 419632 269356 419684 269408
rect 468300 269356 468352 269408
rect 469220 269356 469272 269408
rect 489874 269492 489926 269544
rect 490012 269492 490064 269544
rect 494520 269492 494572 269544
rect 494704 269492 494756 269544
rect 504916 269492 504968 269544
rect 505054 269492 505106 269544
rect 545856 269492 545908 269544
rect 546500 269492 546552 269544
rect 548708 269628 548760 269680
rect 564440 269628 564492 269680
rect 553400 269492 553452 269544
rect 558920 269492 558972 269544
rect 572720 269492 572772 269544
rect 136824 269220 136876 269272
rect 182180 269220 182232 269272
rect 264888 269220 264940 269272
rect 269120 269220 269172 269272
rect 295340 269220 295392 269272
rect 297916 269220 297968 269272
rect 420920 269220 420972 269272
rect 448520 269220 448572 269272
rect 450728 269220 450780 269272
rect 471980 269220 472032 269272
rect 474280 269220 474332 269272
rect 479064 269356 479116 269408
rect 479248 269356 479300 269408
rect 480168 269356 480220 269408
rect 480352 269356 480404 269408
rect 476764 269220 476816 269272
rect 538220 269220 538272 269272
rect 538588 269356 538640 269408
rect 543372 269356 543424 269408
rect 543556 269356 543608 269408
rect 545304 269356 545356 269408
rect 541624 269220 541676 269272
rect 545488 269220 545540 269272
rect 541440 269152 541492 269204
rect 545856 269356 545908 269408
rect 548892 269356 548944 269408
rect 549260 269356 549312 269408
rect 568580 269356 568632 269408
rect 557540 269220 557592 269272
rect 282736 269084 282788 269136
rect 288808 269084 288860 269136
rect 294052 269084 294104 269136
rect 297088 269084 297140 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 502616 269084 502668 269136
rect 505008 269084 505060 269136
rect 108948 269016 109000 269068
rect 166264 269016 166316 269068
rect 185584 269016 185636 269068
rect 196900 269016 196952 269068
rect 86868 268880 86920 268932
rect 144736 268880 144788 268932
rect 179328 268880 179380 268932
rect 215944 268880 215996 268932
rect 382372 268880 382424 268932
rect 400588 268880 400640 268932
rect 102508 268744 102560 268796
rect 162952 268744 163004 268796
rect 163136 268744 163188 268796
rect 203524 268744 203576 268796
rect 203984 268744 204036 268796
rect 227720 268744 227772 268796
rect 227904 268744 227956 268796
rect 250720 268744 250772 268796
rect 387340 268744 387392 268796
rect 422300 269016 422352 269068
rect 443920 269016 443972 269068
rect 502340 269016 502392 269068
rect 506112 269016 506164 269068
rect 591028 269016 591080 269068
rect 418988 268880 419040 268932
rect 440240 268880 440292 268932
rect 441160 268880 441212 268932
rect 499580 268880 499632 268932
rect 503260 268880 503312 268932
rect 587900 268880 587952 268932
rect 422300 268744 422352 268796
rect 436100 268744 436152 268796
rect 446128 268744 446180 268796
rect 505192 268744 505244 268796
rect 508228 268744 508280 268796
rect 514024 268744 514076 268796
rect 99288 268608 99340 268660
rect 160468 268608 160520 268660
rect 162768 268608 162820 268660
rect 205180 268608 205232 268660
rect 219532 268608 219584 268660
rect 244924 268608 244976 268660
rect 363052 268608 363104 268660
rect 386420 268608 386472 268660
rect 397644 268608 397696 268660
rect 433340 268608 433392 268660
rect 448612 268608 448664 268660
rect 509332 268608 509384 268660
rect 510712 268608 510764 268660
rect 598848 268744 598900 268796
rect 514944 268608 514996 268660
rect 517520 268608 517572 268660
rect 518440 268608 518492 268660
rect 608692 268608 608744 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 155868 268472 155920 268524
rect 200212 268472 200264 268524
rect 202972 268472 203024 268524
rect 233332 268472 233384 268524
rect 245568 268472 245620 268524
rect 263140 268472 263192 268524
rect 263508 268472 263560 268524
rect 275560 268472 275612 268524
rect 328552 268472 328604 268524
rect 334348 268472 334400 268524
rect 345940 268472 345992 268524
rect 360292 268472 360344 268524
rect 360752 268472 360804 268524
rect 369860 268472 369912 268524
rect 370320 268472 370372 268524
rect 397460 268472 397512 268524
rect 400588 268472 400640 268524
rect 441620 268472 441672 268524
rect 456064 268472 456116 268524
rect 66260 268336 66312 268388
rect 137284 268336 137336 268388
rect 147588 268336 147640 268388
rect 193588 268336 193640 268388
rect 197268 268336 197320 268388
rect 229192 268336 229244 268388
rect 233700 268336 233752 268388
rect 254860 268336 254912 268388
rect 255228 268336 255280 268388
rect 269764 268336 269816 268388
rect 335176 268336 335228 268388
rect 347780 268336 347832 268388
rect 350080 268336 350132 268388
rect 367100 268336 367152 268388
rect 374920 268336 374972 268388
rect 404452 268336 404504 268388
rect 407212 268336 407264 268388
rect 451464 268336 451516 268388
rect 466828 268336 466880 268388
rect 512368 268336 512420 268388
rect 512736 268472 512788 268524
rect 523684 268472 523736 268524
rect 525340 268472 525392 268524
rect 527180 268472 527232 268524
rect 527364 268472 527416 268524
rect 513840 268336 513892 268388
rect 514024 268336 514076 268388
rect 528928 268472 528980 268524
rect 619732 268472 619784 268524
rect 122748 268200 122800 268252
rect 176200 268200 176252 268252
rect 326068 268200 326120 268252
rect 331404 268200 331456 268252
rect 420460 268200 420512 268252
rect 469404 268200 469456 268252
rect 470140 268200 470192 268252
rect 523500 268200 523552 268252
rect 523684 268200 523736 268252
rect 528514 268200 528566 268252
rect 543694 268336 543746 268388
rect 543832 268336 543884 268388
rect 548432 268200 548484 268252
rect 548800 268336 548852 268388
rect 594800 268336 594852 268388
rect 638960 268200 639012 268252
rect 133788 268064 133840 268116
rect 183652 268064 183704 268116
rect 436192 268064 436244 268116
rect 488540 268064 488592 268116
rect 125508 267928 125560 267980
rect 147588 267928 147640 267980
rect 442816 267928 442868 267980
rect 460848 267928 460900 267980
rect 431960 267792 432012 267844
rect 447140 267792 447192 267844
rect 489184 267792 489236 267844
rect 88984 267656 89036 267708
rect 144552 267656 144604 267708
rect 144920 267656 144972 267708
rect 150532 267656 150584 267708
rect 171784 267656 171836 267708
rect 199384 267656 199436 267708
rect 207664 267656 207716 267708
rect 213460 267656 213512 267708
rect 216128 267656 216180 267708
rect 223396 267656 223448 267708
rect 370780 267656 370832 267708
rect 381360 267656 381412 267708
rect 393136 267656 393188 267708
rect 402060 267656 402112 267708
rect 405556 267656 405608 267708
rect 420920 267656 420972 267708
rect 440332 267656 440384 267708
rect 494060 267860 494112 267912
rect 500776 268064 500828 268116
rect 583852 268064 583904 268116
rect 496452 267928 496504 267980
rect 498200 267928 498252 267980
rect 499120 267928 499172 267980
rect 582380 267928 582432 267980
rect 567660 267792 567712 267844
rect 493324 267656 493376 267708
rect 495624 267656 495676 267708
rect 495808 267656 495860 267708
rect 496636 267656 496688 267708
rect 497464 267656 497516 267708
rect 543694 267656 543746 267708
rect 543832 267656 543884 267708
rect 571984 267656 572036 267708
rect 581276 267656 581328 267708
rect 585784 267656 585836 267708
rect 95884 267520 95936 267572
rect 154672 267520 154724 267572
rect 162124 267520 162176 267572
rect 169576 267520 169628 267572
rect 187148 267520 187200 267572
rect 221740 267520 221792 267572
rect 365812 267520 365864 267572
rect 377588 267520 377640 267572
rect 383200 267520 383252 267572
rect 394700 267520 394752 267572
rect 399760 267520 399812 267572
rect 418988 267520 419040 267572
rect 430396 267520 430448 267572
rect 457444 267520 457496 267572
rect 459192 267520 459244 267572
rect 464344 267520 464396 267572
rect 465172 267520 465224 267572
rect 531504 267520 531556 267572
rect 531872 267520 531924 267572
rect 538174 267520 538226 267572
rect 538312 267520 538364 267572
rect 621664 267520 621716 267572
rect 107568 267384 107620 267436
rect 167092 267384 167144 267436
rect 167736 267384 167788 267436
rect 204352 267384 204404 267436
rect 211804 267384 211856 267436
rect 222568 267384 222620 267436
rect 224224 267384 224276 267436
rect 231676 267384 231728 267436
rect 233884 267384 233936 267436
rect 246580 267384 246632 267436
rect 313648 267384 313700 267436
rect 317788 267384 317840 267436
rect 334348 267384 334400 267436
rect 342904 267384 342956 267436
rect 350908 267384 350960 267436
rect 360752 267384 360804 267436
rect 363328 267384 363380 267436
rect 370504 267384 370556 267436
rect 373264 267384 373316 267436
rect 390468 267384 390520 267436
rect 390652 267384 390704 267436
rect 401600 267384 401652 267436
rect 409604 267384 409656 267436
rect 435364 267384 435416 267436
rect 445944 267384 445996 267436
rect 450728 267384 450780 267436
rect 450912 267384 450964 267436
rect 496452 267384 496504 267436
rect 496820 267384 496872 267436
rect 507860 267384 507912 267436
rect 508044 267384 508096 267436
rect 570604 267384 570656 267436
rect 571984 267384 572036 267436
rect 602344 267384 602396 267436
rect 100668 267248 100720 267300
rect 162124 267248 162176 267300
rect 166908 267248 166960 267300
rect 174544 267248 174596 267300
rect 175096 267248 175148 267300
rect 214288 267248 214340 267300
rect 220084 267248 220136 267300
rect 239128 267248 239180 267300
rect 253664 267248 253716 267300
rect 265624 267248 265676 267300
rect 312820 267248 312872 267300
rect 316040 267248 316092 267300
rect 343456 267248 343508 267300
rect 353944 267248 353996 267300
rect 368204 267248 368256 267300
rect 385500 267248 385552 267300
rect 397092 267248 397144 267300
rect 422300 267248 422352 267300
rect 427912 267248 427964 267300
rect 73804 267112 73856 267164
rect 141424 267112 141476 267164
rect 144552 267112 144604 267164
rect 147404 267112 147456 267164
rect 147588 267112 147640 267164
rect 149060 267112 149112 267164
rect 149888 267112 149940 267164
rect 194416 267112 194468 267164
rect 199660 267112 199712 267164
rect 218428 267112 218480 267164
rect 221464 267112 221516 267164
rect 241612 267112 241664 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 336004 267112 336056 267164
rect 347044 267112 347096 267164
rect 355876 267112 355928 267164
rect 369124 267112 369176 267164
rect 375748 267112 375800 267164
rect 393964 267112 394016 267164
rect 404728 267112 404780 267164
rect 431960 267112 432012 267164
rect 432328 267112 432380 267164
rect 440884 267112 440936 267164
rect 71044 266976 71096 267028
rect 138112 266976 138164 267028
rect 141608 266976 141660 267028
rect 184020 266976 184072 267028
rect 184204 266976 184256 267028
rect 132408 266840 132460 266892
rect 184480 266840 184532 266892
rect 193864 266976 193916 267028
rect 201868 266976 201920 267028
rect 227720 266976 227772 267028
rect 234160 266976 234212 267028
rect 237288 266976 237340 267028
rect 254032 266976 254084 267028
rect 271420 266976 271472 267028
rect 276664 266976 276716 267028
rect 278044 266976 278096 267028
rect 286968 266976 287020 267028
rect 291292 266976 291344 267028
rect 324412 266976 324464 267028
rect 332508 266976 332560 267028
rect 353392 266976 353444 267028
rect 355324 266976 355376 267028
rect 378232 266976 378284 267028
rect 409144 266976 409196 267028
rect 421288 266976 421340 267028
rect 422116 266976 422168 267028
rect 422300 266976 422352 267028
rect 445944 266976 445996 267028
rect 449440 267248 449492 267300
rect 453304 267248 453356 267300
rect 455236 267248 455288 267300
rect 511724 267248 511776 267300
rect 519176 267248 519228 267300
rect 528514 267248 528566 267300
rect 528652 267248 528704 267300
rect 613384 267248 613436 267300
rect 450268 267112 450320 267164
rect 507124 267112 507176 267164
rect 507400 267112 507452 267164
rect 512368 267044 512420 267096
rect 514668 267044 514720 267096
rect 514852 267044 514904 267096
rect 516324 267044 516376 267096
rect 516508 267044 516560 267096
rect 517336 267044 517388 267096
rect 517520 267044 517572 267096
rect 518716 267044 518768 267096
rect 451740 266976 451792 267028
rect 454408 266976 454460 267028
rect 459560 266976 459612 267028
rect 460204 266976 460256 267028
rect 487252 266976 487304 267028
rect 487436 266976 487488 267028
rect 209320 266840 209372 266892
rect 209504 266840 209556 266892
rect 210976 266840 211028 266892
rect 257988 266840 258040 266892
rect 271144 266840 271196 266892
rect 280528 266840 280580 266892
rect 316132 266840 316184 266892
rect 320180 266840 320232 266892
rect 331864 266840 331916 266892
rect 335636 266840 335688 266892
rect 342628 266840 342680 266892
rect 356520 266840 356572 266892
rect 359188 266840 359240 266892
rect 373080 266840 373132 266892
rect 388168 266840 388220 266892
rect 396264 266840 396316 266892
rect 402244 266840 402296 266892
rect 405004 266840 405056 266892
rect 412180 266840 412232 266892
rect 428464 266840 428516 266892
rect 435364 266840 435416 266892
rect 439688 266840 439740 266892
rect 441804 266840 441856 266892
rect 447600 266840 447652 266892
rect 452752 266840 452804 266892
rect 455880 266840 455932 266892
rect 461032 266840 461084 266892
rect 470140 266840 470192 266892
rect 471796 266840 471848 266892
rect 475568 266840 475620 266892
rect 477592 266840 477644 266892
rect 489368 266840 489420 266892
rect 492496 266976 492548 267028
rect 500224 266976 500276 267028
rect 502432 266976 502484 267028
rect 504916 266976 504968 267028
rect 495440 266840 495492 266892
rect 495624 266840 495676 266892
rect 509240 266976 509292 267028
rect 506572 266840 506624 266892
rect 507676 266840 507728 266892
rect 507860 266840 507912 266892
rect 518716 266908 518768 266960
rect 518992 267112 519044 267164
rect 581276 267112 581328 267164
rect 581644 267112 581696 267164
rect 622400 267112 622452 267164
rect 518992 266976 519044 267028
rect 520188 266976 520240 267028
rect 523132 266976 523184 267028
rect 524328 266976 524380 267028
rect 524788 266976 524840 267028
rect 525524 266976 525576 267028
rect 527272 266976 527324 267028
rect 528468 266976 528520 267028
rect 528744 266976 528796 267028
rect 540428 266976 540480 267028
rect 540888 266976 540940 267028
rect 629300 266976 629352 267028
rect 120724 266704 120776 266756
rect 156420 266704 156472 266756
rect 156604 266704 156656 266756
rect 159640 266704 159692 266756
rect 169024 266704 169076 266756
rect 172060 266704 172112 266756
rect 184020 266704 184072 266756
rect 189448 266704 189500 266756
rect 206284 266704 206336 266756
rect 228364 266704 228416 266756
rect 240692 266704 240744 266756
rect 245752 266704 245804 266756
rect 249064 266704 249116 266756
rect 251548 266704 251600 266756
rect 265072 266704 265124 266756
rect 268936 266704 268988 266756
rect 320272 266704 320324 266756
rect 327080 266704 327132 266756
rect 355048 266704 355100 266756
rect 359924 266704 359976 266756
rect 398104 266704 398156 266756
rect 411904 266704 411956 266756
rect 413008 266704 413060 266756
rect 428280 266704 428332 266756
rect 428740 266704 428792 266756
rect 465724 266704 465776 266756
rect 138664 266568 138716 266620
rect 119804 266432 119856 266484
rect 144920 266432 144972 266484
rect 149060 266568 149112 266620
rect 179512 266568 179564 266620
rect 213828 266568 213880 266620
rect 220084 266568 220136 266620
rect 245108 266568 245160 266620
rect 249064 266568 249116 266620
rect 358360 266568 358412 266620
rect 362224 266568 362276 266620
rect 422944 266568 422996 266620
rect 441804 266568 441856 266620
rect 441988 266568 442040 266620
rect 443644 266568 443696 266620
rect 444472 266568 444524 266620
rect 445668 266568 445720 266620
rect 445852 266568 445904 266620
rect 450912 266568 450964 266620
rect 451924 266568 451976 266620
rect 454684 266568 454736 266620
rect 456892 266568 456944 266620
rect 458088 266568 458140 266620
rect 458548 266568 458600 266620
rect 459376 266568 459428 266620
rect 459560 266568 459612 266620
rect 461584 266568 461636 266620
rect 145564 266500 145616 266552
rect 148876 266500 148928 266552
rect 269120 266500 269172 266552
rect 276388 266500 276440 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 330208 266500 330260 266552
rect 334808 266500 334860 266552
rect 346768 266500 346820 266552
rect 351644 266500 351696 266552
rect 380532 266500 380584 266552
rect 382924 266500 382976 266552
rect 394792 266500 394844 266552
rect 397644 266500 397696 266552
rect 151084 266432 151136 266484
rect 172888 266432 172940 266484
rect 361672 266432 361724 266484
rect 362776 266432 362828 266484
rect 439688 266432 439740 266484
rect 476580 266704 476632 266756
rect 481732 266704 481784 266756
rect 484860 266704 484912 266756
rect 485044 266704 485096 266756
rect 496820 266704 496872 266756
rect 497004 266704 497056 266756
rect 549260 266704 549312 266756
rect 572168 266840 572220 266892
rect 581644 266840 581696 266892
rect 470140 266568 470192 266620
rect 528744 266568 528796 266620
rect 528928 266568 528980 266620
rect 529848 266568 529900 266620
rect 532240 266568 532292 266620
rect 540244 266568 540296 266620
rect 540428 266568 540480 266620
rect 578884 266704 578936 266756
rect 572168 266568 572220 266620
rect 469312 266432 469364 266484
rect 474740 266432 474792 266484
rect 475936 266432 475988 266484
rect 485044 266432 485096 266484
rect 487252 266432 487304 266484
rect 493324 266432 493376 266484
rect 500224 266432 500276 266484
rect 558920 266432 558972 266484
rect 147220 266364 147272 266416
rect 148324 266364 148376 266416
rect 149704 266364 149756 266416
rect 182180 266364 182232 266416
rect 186136 266364 186188 266416
rect 202144 266364 202196 266416
rect 206836 266364 206888 266416
rect 210424 266364 210476 266416
rect 211804 266364 211856 266416
rect 222844 266364 222896 266416
rect 224224 266364 224276 266416
rect 230756 266364 230808 266416
rect 236644 266364 236696 266416
rect 242256 266364 242308 266416
rect 243268 266364 243320 266416
rect 252008 266364 252060 266416
rect 257344 266364 257396 266416
rect 268384 266364 268436 266416
rect 273076 266364 273128 266416
rect 278596 266364 278648 266416
rect 286324 266364 286376 266416
rect 290464 266364 290516 266416
rect 292948 266364 293000 266416
rect 293868 266364 293920 266416
rect 296260 266364 296312 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 312360 266364 312412 266416
rect 314660 266364 314712 266416
rect 317788 266364 317840 266416
rect 323124 266364 323176 266416
rect 332692 266364 332744 266416
rect 333612 266364 333664 266416
rect 340972 266364 341024 266416
rect 342168 266364 342220 266416
rect 345112 266364 345164 266416
rect 346124 266364 346176 266416
rect 349252 266364 349304 266416
rect 350264 266364 350316 266416
rect 357532 266364 357584 266416
rect 358636 266364 358688 266416
rect 367468 266364 367520 266416
rect 368388 266364 368440 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375104 266364 375156 266416
rect 379888 266364 379940 266416
rect 380716 266364 380768 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412456 266364 412508 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 423772 266364 423824 266416
rect 424968 266364 425020 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 433708 266364 433760 266416
rect 434628 266364 434680 266416
rect 437848 266364 437900 266416
rect 439504 266364 439556 266416
rect 485872 266364 485924 266416
rect 487068 266364 487120 266416
rect 490288 266296 490340 266348
rect 497004 266364 497056 266416
rect 495440 266228 495492 266280
rect 502616 266296 502668 266348
rect 498568 266160 498620 266212
rect 500960 266160 501012 266212
rect 475108 266024 475160 266076
rect 547880 266024 547932 266076
rect 485044 265888 485096 265940
rect 561680 265888 561732 265940
rect 494980 265752 495032 265804
rect 575848 265752 575900 265804
rect 187700 265616 187752 265668
rect 188252 265616 188304 265668
rect 247224 265616 247276 265668
rect 247868 265616 247920 265668
rect 255504 265616 255556 265668
rect 256148 265616 256200 265668
rect 259552 265616 259604 265668
rect 260380 265616 260432 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 480076 265616 480128 265668
rect 554780 265616 554832 265668
rect 558184 265616 558236 265668
rect 647240 265616 647292 265668
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 565084 259428 565136 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 560944 256708 560996 256760
rect 553492 255552 553544 255604
rect 555424 255552 555476 255604
rect 39028 252968 39080 253020
rect 41512 252968 41564 253020
rect 35808 252832 35860 252884
rect 40684 252832 40736 252884
rect 35624 252696 35676 252748
rect 39028 252696 39080 252748
rect 35440 252560 35492 252612
rect 554412 252560 554464 252612
rect 563704 252560 563756 252612
rect 41696 252492 41748 252544
rect 676036 252356 676088 252408
rect 678428 252356 678480 252408
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 35808 251200 35860 251252
rect 36544 251200 36596 251252
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 553860 246304 553912 246356
rect 632704 246304 632756 246356
rect 554412 245624 554464 245676
rect 598204 245624 598256 245676
rect 554504 244264 554556 244316
rect 623044 244264 623096 244316
rect 36544 242836 36596 242888
rect 41696 242836 41748 242888
rect 587164 242156 587216 242208
rect 648620 242156 648672 242208
rect 553952 241476 554004 241528
rect 631324 241476 631376 241528
rect 553860 240116 553912 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 587164 238688 587216 238740
rect 671896 237804 671948 237856
rect 672264 237600 672316 237652
rect 668768 237192 668820 237244
rect 673092 237464 673144 237516
rect 671528 236988 671580 237040
rect 673304 237056 673356 237108
rect 672908 236852 672960 236904
rect 673276 236852 673328 236904
rect 673528 236648 673580 236700
rect 673460 236512 673512 236564
rect 672540 236172 672592 236224
rect 673752 236240 673804 236292
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 671712 236036 671764 236088
rect 673736 235900 673788 235952
rect 672908 235696 672960 235748
rect 669780 235492 669832 235544
rect 668124 235288 668176 235340
rect 598204 235220 598256 235272
rect 633624 235220 633676 235272
rect 674312 234948 674364 235000
rect 672816 234812 672868 234864
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 671344 234540 671396 234592
rect 668400 234404 668452 234456
rect 671896 234404 671948 234456
rect 675852 234540 675904 234592
rect 678244 234540 678296 234592
rect 674748 234472 674800 234524
rect 674886 234268 674938 234320
rect 667940 234064 667992 234116
rect 670792 233860 670844 233912
rect 675236 233860 675288 233912
rect 675852 233792 675904 233844
rect 677784 233792 677836 233844
rect 675852 233520 675904 233572
rect 683488 233520 683540 233572
rect 670608 233452 670660 233504
rect 669596 233316 669648 233368
rect 671344 233316 671396 233368
rect 676036 233248 676088 233300
rect 678428 233248 678480 233300
rect 671344 233180 671396 233232
rect 673092 233180 673144 233232
rect 671160 233044 671212 233096
rect 674840 233044 674892 233096
rect 652024 232500 652076 232552
rect 675484 232500 675536 232552
rect 662328 232364 662380 232416
rect 675852 232364 675904 232416
rect 679256 232364 679308 232416
rect 672264 232296 672316 232348
rect 665088 232160 665140 232212
rect 672264 231956 672316 232008
rect 675180 231752 675232 231804
rect 668216 231548 668268 231600
rect 669412 231548 669464 231600
rect 675070 231548 675122 231600
rect 673460 231480 673512 231532
rect 674748 231480 674800 231532
rect 674956 231276 675008 231328
rect 674840 231208 674892 231260
rect 675852 231208 675904 231260
rect 677600 231208 677652 231260
rect 674732 230936 674784 230988
rect 673276 230800 673328 230852
rect 144644 230528 144696 230580
rect 150532 230528 150584 230580
rect 152188 230528 152240 230580
rect 158260 230664 158312 230716
rect 668952 230664 669004 230716
rect 673460 230664 673512 230716
rect 90364 230392 90416 230444
rect 166080 230528 166132 230580
rect 168196 230528 168248 230580
rect 439320 230528 439372 230580
rect 161112 230392 161164 230444
rect 161296 230392 161348 230444
rect 215208 230392 215260 230444
rect 223396 230392 223448 230444
rect 271880 230392 271932 230444
rect 274180 230392 274232 230444
rect 307944 230392 307996 230444
rect 312544 230392 312596 230444
rect 315672 230392 315724 230444
rect 377404 230392 377456 230444
rect 378784 230392 378836 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443552 230392 443604 230444
rect 468300 230392 468352 230444
rect 469036 230392 469088 230444
rect 526904 230392 526956 230444
rect 537484 230392 537536 230444
rect 674396 230596 674448 230648
rect 674518 230528 674570 230580
rect 404268 230324 404320 230376
rect 412272 230324 412324 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444840 230324 444892 230376
rect 446404 230324 446456 230376
rect 449164 230324 449216 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 476672 230324 476724 230376
rect 479708 230324 479760 230376
rect 480536 230324 480588 230376
rect 481548 230324 481600 230376
rect 483112 230324 483164 230376
rect 484308 230324 484360 230376
rect 490196 230324 490248 230376
rect 491208 230324 491260 230376
rect 492772 230324 492824 230376
rect 493784 230324 493836 230376
rect 494704 230324 494756 230376
rect 496360 230324 496412 230376
rect 499856 230324 499908 230376
rect 501328 230324 501380 230376
rect 505008 230324 505060 230376
rect 505744 230324 505796 230376
rect 516600 230324 516652 230376
rect 517428 230324 517480 230376
rect 520464 230324 520516 230376
rect 521568 230324 521620 230376
rect 669044 230324 669096 230376
rect 673644 230324 673696 230376
rect 118424 230256 118476 230308
rect 189448 230256 189500 230308
rect 190920 230256 190972 230308
rect 111064 230120 111116 230172
rect 184296 230120 184348 230172
rect 88248 229984 88300 230036
rect 166264 229984 166316 230036
rect 166632 229984 166684 230036
rect 181720 229984 181772 230036
rect 184204 229984 184256 230036
rect 191288 230120 191340 230172
rect 196992 230256 197044 230308
rect 202328 230120 202380 230172
rect 205364 230256 205416 230308
rect 256424 230256 256476 230308
rect 261392 230256 261444 230308
rect 297640 230256 297692 230308
rect 302884 230256 302936 230308
rect 305368 230256 305420 230308
rect 307852 230256 307904 230308
rect 323400 230256 323452 230308
rect 497924 230256 497976 230308
rect 408868 230188 408920 230240
rect 410984 230188 411036 230240
rect 447048 230188 447100 230240
rect 449900 230188 449952 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 454132 230188 454184 230240
rect 455236 230188 455288 230240
rect 470876 230188 470928 230240
rect 471888 230188 471940 230240
rect 475384 230188 475436 230240
rect 479064 230188 479116 230240
rect 532700 230256 532752 230308
rect 547144 230256 547196 230308
rect 504364 230188 504416 230240
rect 511448 230188 511500 230240
rect 516784 230188 516836 230240
rect 521108 230188 521160 230240
rect 530308 230188 530360 230240
rect 674396 230392 674448 230444
rect 251272 230120 251324 230172
rect 276848 230120 276900 230172
rect 313096 230120 313148 230172
rect 315304 230120 315356 230172
rect 340144 230120 340196 230172
rect 488264 230120 488316 230172
rect 533528 230120 533580 230172
rect 543924 230120 543976 230172
rect 555424 230120 555476 230172
rect 571340 230120 571392 230172
rect 345664 230052 345716 230104
rect 353024 230052 353076 230104
rect 444472 230052 444524 230104
rect 447600 230052 447652 230104
rect 499580 230052 499632 230104
rect 673598 230052 673650 230104
rect 190276 229984 190328 230036
rect 246120 229984 246172 230036
rect 251732 229984 251784 230036
rect 292488 229984 292540 230036
rect 296996 229984 297048 230036
rect 302516 229984 302568 230036
rect 305644 229984 305696 230036
rect 334992 229984 335044 230036
rect 380440 229984 380492 230036
rect 389088 229984 389140 230036
rect 410892 229984 410944 230036
rect 417424 229984 417476 230036
rect 467012 229984 467064 230036
rect 474004 229984 474056 230036
rect 484768 229984 484820 230036
rect 74448 229848 74500 229900
rect 155960 229848 156012 229900
rect 156604 229848 156656 229900
rect 176568 229848 176620 229900
rect 177580 229848 177632 229900
rect 67548 229712 67600 229764
rect 144644 229712 144696 229764
rect 144828 229712 144880 229764
rect 140044 229576 140096 229628
rect 146944 229576 146996 229628
rect 148784 229712 148836 229764
rect 151912 229712 151964 229764
rect 152372 229712 152424 229764
rect 190920 229712 190972 229764
rect 191288 229848 191340 229900
rect 240968 229848 241020 229900
rect 245660 229848 245712 229900
rect 287336 229848 287388 229900
rect 300124 229848 300176 229900
rect 329840 229848 329892 229900
rect 334256 229848 334308 229900
rect 345296 229848 345348 229900
rect 352564 229848 352616 229900
rect 358176 229848 358228 229900
rect 364156 229848 364208 229900
rect 381360 229848 381412 229900
rect 384304 229848 384356 229900
rect 394240 229848 394292 229900
rect 469588 229848 469640 229900
rect 476856 229848 476908 229900
rect 481824 229848 481876 229900
rect 489920 229848 489972 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 235816 229712 235868 229764
rect 236920 229712 236972 229764
rect 282184 229712 282236 229764
rect 285312 229712 285364 229764
rect 318248 229712 318300 229764
rect 324044 229712 324096 229764
rect 350448 229712 350500 229764
rect 210056 229576 210108 229628
rect 210240 229576 210292 229628
rect 261576 229576 261628 229628
rect 350540 229576 350592 229628
rect 371056 229712 371108 229764
rect 370964 229576 371016 229628
rect 386512 229712 386564 229764
rect 386972 229712 387024 229764
rect 396816 229712 396868 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 412456 229712 412508 229764
rect 419356 229712 419408 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 468852 229712 468904 229764
rect 475384 229712 475436 229764
rect 479248 229712 479300 229764
rect 487160 229712 487212 229764
rect 477960 229576 478012 229628
rect 478512 229576 478564 229628
rect 490840 229984 490892 230036
rect 493968 229984 494020 230036
rect 505928 229984 505980 230036
rect 515772 229984 515824 230036
rect 517244 229984 517296 230036
rect 522304 229984 522356 230036
rect 523040 229984 523092 230036
rect 534816 229984 534868 230036
rect 538496 229984 538548 230036
rect 559564 229984 559616 230036
rect 673736 229916 673788 229968
rect 495992 229848 496044 229900
rect 510620 229848 510672 229900
rect 513380 229848 513432 229900
rect 525064 229848 525116 229900
rect 528836 229848 528888 229900
rect 533528 229848 533580 229900
rect 534632 229848 534684 229900
rect 555240 229848 555292 229900
rect 675852 229848 675904 229900
rect 677232 229848 677284 229900
rect 494336 229712 494388 229764
rect 509884 229712 509936 229764
rect 525248 229712 525300 229764
rect 528928 229712 528980 229764
rect 536564 229712 536616 229764
rect 562324 229712 562376 229764
rect 669412 229712 669464 229764
rect 670516 229712 670568 229764
rect 497464 229576 497516 229628
rect 503720 229576 503772 229628
rect 508504 229576 508556 229628
rect 515312 229576 515364 229628
rect 526076 229576 526128 229628
rect 530768 229576 530820 229628
rect 540244 229576 540296 229628
rect 666836 229576 666888 229628
rect 131120 229440 131172 229492
rect 197176 229440 197228 229492
rect 203892 229440 203944 229492
rect 205364 229440 205416 229492
rect 231124 229440 231176 229492
rect 277032 229440 277084 229492
rect 509516 229440 509568 229492
rect 518164 229440 518216 229492
rect 519176 229440 519228 229492
rect 527824 229440 527876 229492
rect 673414 229440 673466 229492
rect 436100 229372 436152 229424
rect 436744 229372 436796 229424
rect 448980 229372 449032 229424
rect 451372 229372 451424 229424
rect 122932 229304 122984 229356
rect 179144 229304 179196 229356
rect 182088 229304 182140 229356
rect 230664 229304 230716 229356
rect 453488 229304 453540 229356
rect 455788 229304 455840 229356
rect 358084 229236 358136 229288
rect 360752 229236 360804 229288
rect 360936 229236 360988 229288
rect 363328 229236 363380 229288
rect 419448 229236 419500 229288
rect 424508 229236 424560 229288
rect 450268 229236 450320 229288
rect 451832 229236 451884 229288
rect 479892 229236 479944 229288
rect 482284 229236 482336 229288
rect 501788 229236 501840 229288
rect 507124 229236 507176 229288
rect 673736 229236 673788 229288
rect 92480 229168 92532 229220
rect 146300 229168 146352 229220
rect 146944 229168 146996 229220
rect 153384 229168 153436 229220
rect 153844 229168 153896 229220
rect 163688 229168 163740 229220
rect 163872 229168 163924 229220
rect 166632 229168 166684 229220
rect 167644 229168 167696 229220
rect 220360 229168 220412 229220
rect 476028 229168 476080 229220
rect 478696 229168 478748 229220
rect 378968 229100 379020 229152
rect 383936 229100 383988 229152
rect 102048 229032 102100 229084
rect 175280 229032 175332 229084
rect 175648 229032 175700 229084
rect 97908 228896 97960 228948
rect 82084 228624 82136 228676
rect 108120 228760 108172 228812
rect 108488 228896 108540 228948
rect 170956 228896 171008 228948
rect 173900 228896 173952 228948
rect 174084 228896 174136 228948
rect 171600 228760 171652 228812
rect 181260 228760 181312 228812
rect 96528 228624 96580 228676
rect 172060 228624 172112 228676
rect 172244 228624 172296 228676
rect 179788 228624 179840 228676
rect 181720 229032 181772 229084
rect 190552 229032 190604 229084
rect 191380 229032 191432 229084
rect 194600 229032 194652 229084
rect 195704 229032 195756 229084
rect 250628 229032 250680 229084
rect 259276 229032 259328 229084
rect 298284 229032 298336 229084
rect 413744 229032 413796 229084
rect 420000 229100 420052 229152
rect 420184 229100 420236 229152
rect 421932 229100 421984 229152
rect 424324 229100 424376 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 519820 229032 519872 229084
rect 543188 229032 543240 229084
rect 673388 229032 673440 229084
rect 675852 229032 675904 229084
rect 676220 229032 676272 229084
rect 181904 228896 181956 228948
rect 190920 228760 190972 228812
rect 192208 228896 192260 228948
rect 241612 228896 241664 228948
rect 251088 228896 251140 228948
rect 291200 228896 291252 228948
rect 319812 228896 319864 228948
rect 345940 228896 345992 228948
rect 349988 228896 350040 228948
rect 369124 228896 369176 228948
rect 517888 228896 517940 228948
rect 540060 228896 540112 228948
rect 212632 228760 212684 228812
rect 219164 228760 219216 228812
rect 224040 228760 224092 228812
rect 231308 228760 231360 228812
rect 246212 228760 246264 228812
rect 253848 228760 253900 228812
rect 255044 228760 255096 228812
rect 295708 228760 295760 228812
rect 318064 228760 318116 228812
rect 344652 228760 344704 228812
rect 346124 228760 346176 228812
rect 366180 228760 366232 228812
rect 373816 228760 373868 228812
rect 387248 228760 387300 228812
rect 401324 228760 401376 228812
rect 408408 228760 408460 228812
rect 487160 228760 487212 228812
rect 489920 228760 489972 228812
rect 493968 228760 494020 228812
rect 505928 228760 505980 228812
rect 507124 228760 507176 228812
rect 519728 228760 519780 228812
rect 526260 228760 526312 228812
rect 551192 228760 551244 228812
rect 673506 228692 673558 228744
rect 62764 228488 62816 228540
rect 140780 228488 140832 228540
rect 140964 228488 141016 228540
rect 156420 228488 156472 228540
rect 65984 228352 66036 228404
rect 150164 228352 150216 228404
rect 150348 228352 150400 228404
rect 204720 228488 204772 228540
rect 204904 228488 204956 228540
rect 156972 228352 157024 228404
rect 157432 228352 157484 228404
rect 157800 228352 157852 228404
rect 212172 228352 212224 228404
rect 212632 228488 212684 228540
rect 237196 228624 237248 228676
rect 239404 228624 239456 228676
rect 284116 228624 284168 228676
rect 292396 228624 292448 228676
rect 326620 228624 326672 228676
rect 333244 228624 333296 228676
rect 355600 228624 355652 228676
rect 222752 228352 222804 228404
rect 224040 228352 224092 228404
rect 267372 228488 267424 228540
rect 267556 228488 267608 228540
rect 307300 228488 307352 228540
rect 307668 228488 307720 228540
rect 335636 228488 335688 228540
rect 336648 228488 336700 228540
rect 358820 228488 358872 228540
rect 225696 228352 225748 228404
rect 273812 228352 273864 228404
rect 283932 228352 283984 228404
rect 320180 228352 320232 228404
rect 326804 228352 326856 228404
rect 351092 228352 351144 228404
rect 355324 228352 355376 228404
rect 369768 228624 369820 228676
rect 376484 228624 376536 228676
rect 389732 228624 389784 228676
rect 390284 228624 390336 228676
rect 400036 228624 400088 228676
rect 411076 228624 411128 228676
rect 416136 228624 416188 228676
rect 479708 228624 479760 228676
rect 487436 228624 487488 228676
rect 495348 228624 495400 228676
rect 511448 228624 511500 228676
rect 528192 228624 528244 228676
rect 553676 228624 553728 228676
rect 672724 228556 672776 228608
rect 672908 228556 672960 228608
rect 366916 228488 366968 228540
rect 382004 228488 382056 228540
rect 362868 228352 362920 228404
rect 379428 228352 379480 228404
rect 381912 228352 381964 228404
rect 392860 228488 392912 228540
rect 393044 228488 393096 228540
rect 391848 228352 391900 228404
rect 400036 228488 400088 228540
rect 407764 228488 407816 228540
rect 482468 228488 482520 228540
rect 494704 228488 494756 228540
rect 502432 228488 502484 228540
rect 520924 228488 520976 228540
rect 531412 228488 531464 228540
rect 558184 228488 558236 228540
rect 673388 228488 673440 228540
rect 672264 228420 672316 228472
rect 108120 228216 108172 228268
rect 140964 228216 141016 228268
rect 141148 228216 141200 228268
rect 190920 228216 190972 228268
rect 106188 228080 106240 228132
rect 108488 228080 108540 228132
rect 113088 228080 113140 228132
rect 181076 228080 181128 228132
rect 181260 228080 181312 228132
rect 204904 228216 204956 228268
rect 122748 227944 122800 227996
rect 181720 227944 181772 227996
rect 181904 227944 181956 227996
rect 184940 227944 184992 227996
rect 190920 227944 190972 227996
rect 201040 228080 201092 228132
rect 201408 228080 201460 228132
rect 252560 228216 252612 228268
rect 277124 228216 277176 228268
rect 311808 228216 311860 228268
rect 402612 228352 402664 228404
rect 409604 228352 409656 228404
rect 415492 228352 415544 228404
rect 486976 228352 487028 228404
rect 501696 228352 501748 228404
rect 506296 228352 506348 228404
rect 526536 228352 526588 228404
rect 537852 228352 537904 228404
rect 566188 228352 566240 228404
rect 403900 228216 403952 228268
rect 478696 228216 478748 228268
rect 487068 228216 487120 228268
rect 512092 228216 512144 228268
rect 533528 228216 533580 228268
rect 671344 228216 671396 228268
rect 205456 228080 205508 228132
rect 257068 228080 257120 228132
rect 288072 228080 288124 228132
rect 321468 228080 321520 228132
rect 671896 228012 671948 228064
rect 198004 227944 198056 227996
rect 204536 227944 204588 227996
rect 212172 227944 212224 227996
rect 218428 227944 218480 227996
rect 222752 227944 222804 227996
rect 226156 227944 226208 227996
rect 133788 227808 133840 227860
rect 200396 227808 200448 227860
rect 204720 227808 204772 227860
rect 210700 227808 210752 227860
rect 226156 227808 226208 227860
rect 272524 227944 272576 227996
rect 369124 227876 369176 227928
rect 375564 227876 375616 227928
rect 407764 227876 407816 227928
rect 411628 227876 411680 227928
rect 471520 227876 471572 227928
rect 479248 227876 479300 227928
rect 242532 227740 242584 227792
rect 245660 227740 245712 227792
rect 255964 227740 256016 227792
rect 259000 227740 259052 227792
rect 366272 227740 366324 227792
rect 372988 227740 373040 227792
rect 393964 227740 394016 227792
rect 395528 227740 395580 227792
rect 396724 227740 396776 227792
rect 397460 227740 397512 227792
rect 402244 227740 402296 227792
rect 403256 227740 403308 227792
rect 404084 227740 404136 227792
rect 408868 227740 408920 227792
rect 409144 227740 409196 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416596 227740 416648 227792
rect 420644 227740 420696 227792
rect 475016 227740 475068 227792
rect 482836 227740 482888 227792
rect 510620 227740 510672 227792
rect 513012 227740 513064 227792
rect 663708 227740 663760 227792
rect 665272 227740 665324 227792
rect 672954 227740 673006 227792
rect 109868 227672 109920 227724
rect 182364 227672 182416 227724
rect 184572 227672 184624 227724
rect 187516 227672 187568 227724
rect 191748 227672 191800 227724
rect 270316 227672 270368 227724
rect 306656 227672 306708 227724
rect 321376 227672 321428 227724
rect 346584 227672 346636 227724
rect 528928 227672 528980 227724
rect 549904 227672 549956 227724
rect 248052 227604 248104 227656
rect 670516 227604 670568 227656
rect 100668 227536 100720 227588
rect 174636 227536 174688 227588
rect 179328 227536 179380 227588
rect 236460 227536 236512 227588
rect 252284 227536 252336 227588
rect 293132 227536 293184 227588
rect 299204 227536 299256 227588
rect 328552 227536 328604 227588
rect 359464 227536 359516 227588
rect 374920 227536 374972 227588
rect 465908 227536 465960 227588
rect 469864 227536 469916 227588
rect 518532 227536 518584 227588
rect 541624 227536 541676 227588
rect 560944 227536 560996 227588
rect 567660 227536 567712 227588
rect 89628 227400 89680 227452
rect 159640 227400 159692 227452
rect 160008 227400 160060 227452
rect 166908 227400 166960 227452
rect 86684 227264 86736 227316
rect 164332 227264 164384 227316
rect 165344 227264 165396 227316
rect 175004 227400 175056 227452
rect 231952 227400 232004 227452
rect 248144 227400 248196 227452
rect 291844 227400 291896 227452
rect 293684 227400 293736 227452
rect 325332 227400 325384 227452
rect 340604 227400 340656 227452
rect 361396 227400 361448 227452
rect 227444 227264 227496 227316
rect 75828 227128 75880 227180
rect 151728 227128 151780 227180
rect 152280 227128 152332 227180
rect 156512 227128 156564 227180
rect 57704 226992 57756 227044
rect 135260 226992 135312 227044
rect 135444 226992 135496 227044
rect 168840 227128 168892 227180
rect 169484 227128 169536 227180
rect 228732 227128 228784 227180
rect 156972 226992 157024 227044
rect 213276 226992 213328 227044
rect 226984 226992 227036 227044
rect 233240 227264 233292 227316
rect 234528 227264 234580 227316
rect 278320 227264 278372 227316
rect 280804 227264 280856 227316
rect 312084 227264 312136 227316
rect 326344 227264 326396 227316
rect 352380 227264 352432 227316
rect 361304 227264 361356 227316
rect 377220 227400 377272 227452
rect 362224 227264 362276 227316
rect 372344 227264 372396 227316
rect 373264 227264 373316 227316
rect 383292 227400 383344 227452
rect 515956 227400 516008 227452
rect 538496 227400 538548 227452
rect 672264 227332 672316 227384
rect 382832 227264 382884 227316
rect 391664 227264 391716 227316
rect 395988 227264 396040 227316
rect 406476 227264 406528 227316
rect 485044 227264 485096 227316
rect 498844 227264 498896 227316
rect 501328 227264 501380 227316
rect 517796 227264 517848 227316
rect 521752 227264 521804 227316
rect 545764 227264 545816 227316
rect 672724 227332 672776 227384
rect 235724 227128 235776 227180
rect 280252 227128 280304 227180
rect 296168 227128 296220 227180
rect 329196 227128 329248 227180
rect 329748 227128 329800 227180
rect 353668 227128 353720 227180
rect 354588 227128 354640 227180
rect 373632 227128 373684 227180
rect 382096 227128 382148 227180
rect 396172 227128 396224 227180
rect 498568 227128 498620 227180
rect 516048 227128 516100 227180
rect 533988 227128 534040 227180
rect 561496 227128 561548 227180
rect 229054 226992 229106 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 106924 226856 106976 226908
rect 125784 226856 125836 226908
rect 121368 226720 121420 226772
rect 190460 226856 190512 226908
rect 200028 226856 200080 226908
rect 252008 226856 252060 226908
rect 272524 226856 272576 226908
rect 284760 226856 284812 226908
rect 308588 226856 308640 226908
rect 336280 226992 336332 227044
rect 336464 226992 336516 227044
rect 360108 226992 360160 227044
rect 369768 226992 369820 227044
rect 385868 226992 385920 227044
rect 386328 226992 386380 227044
rect 398748 226992 398800 227044
rect 472164 226992 472216 227044
rect 480812 226992 480864 227044
rect 481180 226992 481232 227044
rect 493968 226992 494020 227044
rect 497280 226992 497332 227044
rect 513840 226992 513892 227044
rect 514024 226992 514076 227044
rect 536104 226992 536156 227044
rect 537208 226992 537260 227044
rect 565360 226992 565412 227044
rect 670516 226992 670568 227044
rect 355508 226856 355560 226908
rect 362224 226856 362276 226908
rect 398748 226856 398800 226908
rect 408684 226856 408736 226908
rect 671896 226788 671948 226840
rect 119804 226584 119856 226636
rect 190092 226720 190144 226772
rect 195888 226720 195940 226772
rect 199292 226720 199344 226772
rect 212356 226720 212408 226772
rect 262220 226720 262272 226772
rect 125784 226448 125836 226500
rect 135444 226584 135496 226636
rect 135628 226584 135680 226636
rect 129648 226448 129700 226500
rect 137192 226448 137244 226500
rect 137560 226584 137612 226636
rect 197360 226584 197412 226636
rect 222016 226584 222068 226636
rect 269948 226584 270000 226636
rect 142114 226448 142166 226500
rect 142252 226448 142304 226500
rect 205180 226448 205232 226500
rect 213184 226448 213236 226500
rect 217784 226448 217836 226500
rect 221832 226448 221884 226500
rect 229008 226448 229060 226500
rect 232504 226448 232556 226500
rect 266728 226448 266780 226500
rect 291844 226380 291896 226432
rect 295064 226380 295116 226432
rect 672156 226448 672208 226500
rect 83464 226244 83516 226296
rect 154212 226244 154264 226296
rect 69664 226108 69716 226160
rect 143540 226108 143592 226160
rect 146944 226108 146996 226160
rect 166954 226312 167006 226364
rect 221004 226312 221056 226364
rect 490104 226312 490156 226364
rect 494888 226312 494940 226364
rect 671896 226312 671948 226364
rect 161940 226244 161992 226296
rect 162308 226244 162360 226296
rect 166816 226244 166868 226296
rect 222476 226244 222528 226296
rect 225512 226244 225564 226296
rect 228916 226244 228968 226296
rect 275100 226244 275152 226296
rect 278412 226244 278464 226296
rect 315028 226244 315080 226296
rect 317328 226244 317380 226296
rect 334256 226244 334308 226296
rect 672034 226244 672086 226296
rect 154764 226108 154816 226160
rect 157432 226108 157484 226160
rect 157616 226108 157668 226160
rect 215852 226108 215904 226160
rect 216496 226108 216548 226160
rect 264796 226108 264848 226160
rect 266268 226108 266320 226160
rect 303436 226108 303488 226160
rect 325608 226108 325660 226160
rect 349160 226108 349212 226160
rect 514668 226108 514720 226160
rect 535460 226108 535512 226160
rect 667848 226040 667900 226092
rect 93768 225972 93820 226024
rect 161572 225972 161624 226024
rect 161940 225972 161992 226024
rect 171048 225972 171100 226024
rect 171232 225972 171284 226024
rect 186412 225972 186464 226024
rect 186596 225972 186648 226024
rect 224224 225972 224276 226024
rect 94964 225836 95016 225888
rect 166816 225836 166868 225888
rect 166954 225836 167006 225888
rect 64788 225700 64840 225752
rect 92480 225700 92532 225752
rect 108304 225700 108356 225752
rect 171048 225700 171100 225752
rect 171232 225700 171284 225752
rect 175924 225700 175976 225752
rect 176292 225836 176344 225888
rect 176614 225836 176666 225888
rect 176752 225836 176804 225888
rect 181076 225836 181128 225888
rect 181628 225836 181680 225888
rect 183284 225836 183336 225888
rect 186136 225836 186188 225888
rect 186274 225836 186326 225888
rect 233884 225972 233936 226024
rect 243544 225972 243596 226024
rect 248696 225972 248748 226024
rect 267556 225972 267608 226024
rect 304080 225972 304132 226024
rect 313096 225972 313148 226024
rect 340788 225972 340840 226024
rect 181444 225700 181496 225752
rect 184572 225700 184624 225752
rect 187056 225700 187108 225752
rect 239036 225836 239088 225888
rect 249708 225836 249760 225888
rect 290556 225836 290608 225888
rect 295248 225836 295300 225888
rect 325976 225836 326028 225888
rect 340144 225836 340196 225888
rect 347872 225972 347924 226024
rect 349068 225972 349120 226024
rect 367192 225972 367244 226024
rect 501144 225972 501196 226024
rect 347044 225836 347096 225888
rect 365904 225836 365956 225888
rect 367744 225836 367796 225888
rect 379612 225836 379664 225888
rect 488908 225836 488960 225888
rect 502984 225836 503036 225888
rect 458640 225768 458692 225820
rect 462596 225768 462648 225820
rect 61384 225564 61436 225616
rect 136824 225564 136876 225616
rect 137008 225564 137060 225616
rect 146944 225564 146996 225616
rect 147404 225564 147456 225616
rect 204076 225564 204128 225616
rect 204904 225564 204956 225616
rect 222476 225564 222528 225616
rect 224224 225564 224276 225616
rect 242900 225700 242952 225752
rect 257804 225700 257856 225752
rect 299572 225700 299624 225752
rect 304908 225700 304960 225752
rect 333704 225700 333756 225752
rect 335084 225700 335136 225752
rect 356888 225700 356940 225752
rect 379336 225700 379388 225752
rect 393596 225700 393648 225752
rect 394608 225700 394660 225752
rect 404544 225700 404596 225752
rect 487620 225700 487672 225752
rect 501512 225700 501564 225752
rect 524328 225972 524380 226024
rect 547880 225972 547932 226024
rect 508872 225836 508924 225888
rect 528928 225836 528980 225888
rect 530124 225836 530176 225888
rect 556160 225836 556212 225888
rect 519360 225700 519412 225752
rect 527548 225700 527600 225752
rect 553308 225700 553360 225752
rect 556804 225700 556856 225752
rect 570696 225700 570748 225752
rect 671820 225700 671872 225752
rect 671344 225632 671396 225684
rect 234344 225564 234396 225616
rect 281540 225564 281592 225616
rect 285496 225564 285548 225616
rect 318892 225564 318944 225616
rect 322664 225564 322716 225616
rect 349804 225564 349856 225616
rect 351184 225564 351236 225616
rect 370412 225564 370464 225616
rect 372344 225564 372396 225616
rect 388076 225564 388128 225616
rect 388444 225564 388496 225616
rect 399392 225564 399444 225616
rect 467656 225564 467708 225616
rect 476672 225564 476724 225616
rect 477316 225564 477368 225616
rect 488540 225564 488592 225616
rect 494152 225564 494204 225616
rect 509700 225564 509752 225616
rect 510160 225564 510212 225616
rect 530584 225564 530636 225616
rect 535920 225564 535972 225616
rect 564716 225564 564768 225616
rect 103244 225428 103296 225480
rect 108304 225428 108356 225480
rect 105728 225292 105780 225344
rect 127440 225428 127492 225480
rect 117228 225292 117280 225344
rect 181444 225428 181496 225480
rect 181628 225428 181680 225480
rect 185584 225428 185636 225480
rect 187700 225428 187752 225480
rect 190552 225428 190604 225480
rect 190736 225428 190788 225480
rect 242256 225428 242308 225480
rect 667020 225428 667072 225480
rect 127440 225156 127492 225208
rect 137008 225292 137060 225344
rect 128084 225156 128136 225208
rect 142114 225292 142166 225344
rect 142252 225292 142304 225344
rect 202972 225292 203024 225344
rect 204076 225292 204128 225344
rect 207756 225292 207808 225344
rect 208124 225292 208176 225344
rect 260932 225292 260984 225344
rect 463148 225224 463200 225276
rect 467104 225224 467156 225276
rect 670516 225224 670568 225276
rect 126888 225020 126940 225072
rect 187700 225156 187752 225208
rect 188068 225156 188120 225208
rect 195888 225156 195940 225208
rect 199384 225156 199436 225208
rect 204904 225156 204956 225208
rect 205088 225156 205140 225208
rect 254492 225156 254544 225208
rect 137468 225020 137520 225072
rect 141516 225020 141568 225072
rect 141884 225020 141936 225072
rect 116860 224884 116912 224936
rect 122932 224884 122984 224936
rect 126520 224884 126572 224936
rect 142068 224884 142120 224936
rect 142436 225020 142488 225072
rect 162308 225020 162360 225072
rect 162768 225020 162820 225072
rect 166540 225020 166592 225072
rect 166724 225020 166776 225072
rect 169024 225020 169076 225072
rect 169208 225020 169260 225072
rect 170864 225020 170916 225072
rect 171048 225020 171100 225072
rect 223580 225020 223632 225072
rect 224684 225020 224736 225072
rect 270592 225020 270644 225072
rect 671252 225020 671304 225072
rect 275652 224952 275704 225004
rect 276848 224952 276900 225004
rect 282828 224952 282880 225004
rect 285312 224952 285364 225004
rect 209412 224884 209464 224936
rect 209688 224884 209740 224936
rect 259644 224884 259696 224936
rect 264244 224884 264296 224936
rect 269304 224884 269356 224936
rect 288256 224884 288308 224936
rect 322388 224884 322440 224936
rect 407028 224884 407080 224936
rect 414848 224884 414900 224936
rect 426440 224884 426492 224936
rect 426992 224884 427044 224936
rect 118608 224748 118660 224800
rect 181260 224748 181312 224800
rect 115664 224612 115716 224664
rect 187056 224748 187108 224800
rect 187516 224748 187568 224800
rect 190736 224748 190788 224800
rect 194324 224748 194376 224800
rect 247408 224748 247460 224800
rect 282644 224748 282696 224800
rect 316316 224748 316368 224800
rect 515772 224748 515824 224800
rect 525248 224748 525300 224800
rect 526076 224748 526128 224800
rect 537116 224748 537168 224800
rect 460572 224680 460624 224732
rect 462964 224680 463016 224732
rect 671252 224680 671304 224732
rect 181812 224612 181864 224664
rect 191380 224612 191432 224664
rect 192484 224612 192536 224664
rect 194508 224612 194560 224664
rect 195704 224612 195756 224664
rect 248880 224612 248932 224664
rect 249064 224612 249116 224664
rect 263876 224612 263928 224664
rect 271328 224612 271380 224664
rect 309876 224612 309928 224664
rect 315856 224612 315908 224664
rect 341432 224612 341484 224664
rect 344928 224612 344980 224664
rect 364616 224612 364668 224664
rect 486608 224612 486660 224664
rect 500408 224612 500460 224664
rect 508228 224612 508280 224664
rect 528008 224612 528060 224664
rect 670516 224612 670568 224664
rect 60648 224476 60700 224528
rect 103612 224476 103664 224528
rect 108948 224476 109000 224528
rect 183652 224476 183704 224528
rect 184020 224476 184072 224528
rect 233700 224476 233752 224528
rect 233884 224476 233936 224528
rect 246764 224476 246816 224528
rect 247684 224476 247736 224528
rect 289268 224476 289320 224528
rect 319996 224476 320048 224528
rect 347228 224476 347280 224528
rect 491484 224476 491536 224528
rect 506480 224476 506532 224528
rect 510804 224476 510856 224528
rect 531780 224476 531832 224528
rect 532056 224476 532108 224528
rect 558920 224476 558972 224528
rect 670608 224408 670660 224460
rect 82544 224340 82596 224392
rect 126520 224340 126572 224392
rect 126704 224340 126756 224392
rect 131120 224340 131172 224392
rect 131304 224340 131356 224392
rect 193956 224340 194008 224392
rect 194140 224340 194192 224392
rect 204904 224340 204956 224392
rect 205088 224340 205140 224392
rect 255780 224340 255832 224392
rect 262128 224340 262180 224392
rect 300860 224340 300912 224392
rect 303436 224340 303488 224392
rect 333060 224340 333112 224392
rect 333888 224340 333940 224392
rect 356244 224340 356296 224392
rect 357348 224340 357400 224392
rect 374276 224340 374328 224392
rect 375288 224340 375340 224392
rect 387800 224340 387852 224392
rect 456156 224340 456208 224392
rect 459652 224340 459704 224392
rect 479064 224340 479116 224392
rect 485780 224340 485832 224392
rect 499212 224340 499264 224392
rect 516416 224340 516468 224392
rect 525616 224340 525668 224392
rect 550640 224340 550692 224392
rect 59268 224204 59320 224256
rect 141608 224204 141660 224256
rect 142068 224204 142120 224256
rect 157294 224204 157346 224256
rect 157432 224204 157484 224256
rect 170956 224204 171008 224256
rect 171094 224204 171146 224256
rect 186872 224204 186924 224256
rect 187056 224204 187108 224256
rect 188804 224204 188856 224256
rect 188988 224204 189040 224256
rect 243820 224204 243872 224256
rect 246948 224204 247000 224256
rect 288624 224204 288676 224256
rect 289544 224204 289596 224256
rect 307852 224204 307904 224256
rect 308956 224204 309008 224256
rect 339500 224204 339552 224256
rect 341892 224204 341944 224256
rect 364800 224204 364852 224256
rect 364984 224204 365036 224256
rect 378140 224204 378192 224256
rect 388904 224204 388956 224256
rect 400956 224204 401008 224256
rect 416412 224204 416464 224256
rect 422208 224204 422260 224256
rect 451372 224204 451424 224256
rect 452016 224204 452068 224256
rect 462412 224204 462464 224256
rect 469680 224204 469732 224256
rect 470232 224204 470284 224256
rect 479524 224204 479576 224256
rect 483756 224204 483808 224256
rect 497280 224204 497332 224256
rect 513196 224204 513248 224256
rect 534448 224204 534500 224256
rect 535276 224204 535328 224256
rect 563980 224204 564032 224256
rect 423588 224136 423640 224188
rect 424324 224136 424376 224188
rect 667020 224136 667072 224188
rect 104808 224068 104860 224120
rect 116860 224068 116912 224120
rect 117044 224068 117096 224120
rect 118424 224068 118476 224120
rect 122288 224068 122340 224120
rect 131304 224068 131356 224120
rect 131488 224068 131540 224120
rect 192484 224068 192536 224120
rect 192668 224068 192720 224120
rect 194140 224068 194192 224120
rect 194508 224068 194560 224120
rect 196532 224068 196584 224120
rect 201224 224068 201276 224120
rect 204720 224068 204772 224120
rect 204904 224068 204956 224120
rect 233884 224068 233936 224120
rect 76472 223932 76524 223984
rect 141424 223932 141476 223984
rect 141608 223932 141660 223984
rect 145196 223932 145248 223984
rect 145380 223932 145432 223984
rect 147220 223932 147272 223984
rect 147680 223932 147732 223984
rect 154580 223932 154632 223984
rect 156880 223932 156932 223984
rect 217048 223932 217100 223984
rect 217232 223932 217284 223984
rect 228088 223932 228140 223984
rect 231584 223932 231636 223984
rect 278964 224068 279016 224120
rect 286968 224068 287020 224120
rect 319536 224068 319588 224120
rect 238668 223932 238720 223984
rect 282460 223932 282512 223984
rect 125140 223796 125192 223848
rect 131488 223796 131540 223848
rect 134984 223796 135036 223848
rect 204260 223796 204312 223848
rect 205272 223796 205324 223848
rect 212816 223796 212868 223848
rect 215944 223796 215996 223848
rect 222936 223796 222988 223848
rect 233700 223796 233752 223848
rect 239680 223796 239732 223848
rect 242716 223796 242768 223848
rect 285036 223796 285088 223848
rect 132224 223660 132276 223712
rect 201684 223660 201736 223712
rect 88064 223524 88116 223576
rect 164976 223524 165028 223576
rect 166264 223524 166316 223576
rect 168104 223524 168156 223576
rect 168288 223524 168340 223576
rect 226800 223524 226852 223576
rect 268844 223524 268896 223576
rect 297824 223524 297876 223576
rect 300124 223524 300176 223576
rect 563704 223592 563756 223644
rect 571248 223592 571300 223644
rect 306012 223524 306064 223576
rect 329012 223524 329064 223576
rect 342720 223524 342772 223576
rect 457996 223524 458048 223576
rect 460204 223524 460256 223576
rect 473452 223524 473504 223576
rect 475752 223524 475804 223576
rect 499580 223524 499632 223576
rect 503168 223524 503220 223576
rect 81348 223388 81400 223440
rect 157248 223388 157300 223440
rect 157432 223388 157484 223440
rect 159824 223388 159876 223440
rect 161112 223388 161164 223440
rect 162308 223388 162360 223440
rect 164148 223388 164200 223440
rect 224040 223388 224092 223440
rect 260564 223388 260616 223440
rect 298928 223388 298980 223440
rect 301964 223388 302016 223440
rect 331128 223388 331180 223440
rect 516784 223388 516836 223440
rect 532148 223388 532200 223440
rect 543924 223388 543976 223440
rect 554872 223388 554924 223440
rect 96712 223252 96764 223304
rect 117964 223252 118016 223304
rect 118148 223252 118200 223304
rect 166264 223252 166316 223304
rect 168104 223252 168156 223304
rect 185768 223252 185820 223304
rect 186044 223252 186096 223304
rect 192208 223252 192260 223304
rect 192484 223252 192536 223304
rect 196072 223252 196124 223304
rect 204076 223252 204128 223304
rect 254860 223252 254912 223304
rect 264704 223252 264756 223304
rect 304724 223252 304776 223304
rect 306104 223252 306156 223304
rect 336924 223252 336976 223304
rect 343364 223252 343416 223304
rect 363972 223252 364024 223304
rect 506940 223252 506992 223304
rect 526352 223252 526404 223304
rect 530308 223252 530360 223304
rect 544936 223252 544988 223304
rect 78404 223116 78456 223168
rect 152280 223116 152332 223168
rect 152464 223116 152516 223168
rect 166264 223116 166316 223168
rect 166448 223116 166500 223168
rect 222292 223116 222344 223168
rect 224224 223116 224276 223168
rect 238392 223116 238444 223168
rect 245568 223116 245620 223168
rect 287612 223116 287664 223168
rect 291108 223116 291160 223168
rect 323676 223116 323728 223168
rect 330484 223116 330536 223168
rect 354956 223116 355008 223168
rect 357164 223116 357216 223168
rect 376208 223116 376260 223168
rect 522672 223116 522724 223168
rect 546776 223116 546828 223168
rect 92388 222980 92440 223032
rect 96712 222980 96764 223032
rect 98644 222980 98696 223032
rect 166080 222980 166132 223032
rect 166816 222980 166868 223032
rect 181628 222980 181680 223032
rect 181812 222980 181864 223032
rect 234804 222980 234856 223032
rect 235264 222980 235316 223032
rect 243268 222980 243320 223032
rect 250904 222980 250956 223032
rect 294420 222980 294472 223032
rect 300308 222980 300360 223032
rect 331312 222980 331364 223032
rect 337936 222980 337988 223032
rect 359188 222980 359240 223032
rect 370504 222980 370556 223032
rect 384580 222980 384632 223032
rect 387708 222980 387760 223032
rect 398104 222980 398156 223032
rect 478328 222980 478380 223032
rect 485044 222980 485096 223032
rect 485596 222980 485648 223032
rect 498200 222980 498252 223032
rect 503352 222980 503404 223032
rect 521936 222980 521988 223032
rect 523684 222980 523736 223032
rect 548156 222980 548208 223032
rect 570328 222980 570380 223032
rect 575388 222980 575440 223032
rect 56508 222844 56560 222896
rect 137100 222844 137152 222896
rect 137284 222844 137336 222896
rect 152464 222844 152516 222896
rect 154488 222844 154540 222896
rect 212172 222844 212224 222896
rect 85488 222708 85540 222760
rect 162124 222708 162176 222760
rect 162308 222708 162360 222760
rect 168104 222708 168156 222760
rect 166816 222640 166868 222692
rect 89168 222572 89220 222624
rect 98644 222572 98696 222624
rect 99104 222572 99156 222624
rect 166080 222572 166132 222624
rect 167000 222572 167052 222624
rect 174820 222572 174872 222624
rect 175004 222572 175056 222624
rect 181260 222572 181312 222624
rect 181628 222708 181680 222760
rect 196072 222708 196124 222760
rect 203708 222708 203760 222760
rect 221648 222844 221700 222896
rect 233148 222844 233200 222896
rect 277676 222844 277728 222896
rect 284116 222844 284168 222896
rect 316684 222844 316736 222896
rect 316868 222844 316920 222896
rect 343180 222844 343232 222896
rect 347504 222844 347556 222896
rect 368480 222844 368532 222896
rect 375104 222844 375156 222896
rect 391020 222844 391072 222896
rect 397184 222844 397236 222896
rect 407212 222844 407264 222896
rect 408408 222844 408460 222896
rect 416780 222844 416832 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 466736 222844 466788 222896
rect 467472 222844 467524 222896
rect 473452 222844 473504 222896
rect 474740 222844 474792 222896
rect 484860 222844 484912 222896
rect 489552 222844 489604 222896
rect 503996 222844 504048 222896
rect 504640 222844 504692 222896
rect 523776 222844 523828 222896
rect 533712 222844 533764 222896
rect 560668 222844 560720 222896
rect 562968 222844 563020 222896
rect 571432 222844 571484 222896
rect 571892 222844 571944 222896
rect 192024 222572 192076 222624
rect 213828 222708 213880 222760
rect 262864 222708 262916 222760
rect 263508 222708 263560 222760
rect 296996 222708 297048 222760
rect 563980 222640 564032 222692
rect 574652 222640 574704 222692
rect 205088 222572 205140 222624
rect 208768 222572 208820 222624
rect 209504 222572 209556 222624
rect 210240 222572 210292 222624
rect 210884 222572 210936 222624
rect 260288 222572 260340 222624
rect 117964 222436 118016 222488
rect 137284 222436 137336 222488
rect 137468 222436 137520 222488
rect 151360 222436 151412 222488
rect 152280 222436 152332 222488
rect 157064 222436 157116 222488
rect 157248 222436 157300 222488
rect 219716 222436 219768 222488
rect 220084 222436 220136 222488
rect 268660 222436 268712 222488
rect 555240 222368 555292 222420
rect 562140 222368 562192 222420
rect 572260 222504 572312 222556
rect 565084 222368 565136 222420
rect 568672 222368 568724 222420
rect 570144 222368 570196 222420
rect 574468 222368 574520 222420
rect 112904 222300 112956 222352
rect 118148 222300 118200 222352
rect 133604 222300 133656 222352
rect 136916 222300 136968 222352
rect 137100 222300 137152 222352
rect 142620 222300 142672 222352
rect 145012 222300 145064 222352
rect 143448 222232 143500 222284
rect 144828 222232 144880 222284
rect 203708 222300 203760 222352
rect 207480 222300 207532 222352
rect 212172 222300 212224 222352
rect 216220 222300 216272 222352
rect 220728 222300 220780 222352
rect 268016 222300 268068 222352
rect 203524 222232 203576 222284
rect 171140 222164 171192 222216
rect 482836 222164 482888 222216
rect 593972 222232 594024 222284
rect 596640 222232 596692 222284
rect 95700 221960 95752 222012
rect 117964 222096 118016 222148
rect 118148 222096 118200 222148
rect 171324 222096 171376 222148
rect 177396 222096 177448 222148
rect 177580 222096 177632 222148
rect 179972 222096 180024 222148
rect 180156 222096 180208 222148
rect 104624 221960 104676 222012
rect 171048 221960 171100 222012
rect 71688 221824 71740 221876
rect 142804 221824 142856 221876
rect 143172 221824 143224 221876
rect 172980 221960 173032 222012
rect 176292 221960 176344 222012
rect 181444 221960 181496 222012
rect 181812 222096 181864 222148
rect 240140 222096 240192 222148
rect 256332 222096 256384 222148
rect 261208 222096 261260 222148
rect 261392 222096 261444 222148
rect 301688 222096 301740 222148
rect 331680 222096 331732 222148
rect 353944 222096 353996 222148
rect 462136 222096 462188 222148
rect 468484 222096 468536 222148
rect 471888 222096 471940 222148
rect 477592 222096 477644 222148
rect 547144 222096 547196 222148
rect 558000 222096 558052 222148
rect 558184 222096 558236 222148
rect 562876 222096 562928 222148
rect 237380 221960 237432 222012
rect 243912 221960 243964 222012
rect 285680 221960 285732 222012
rect 310152 221960 310204 222012
rect 338120 221960 338172 222012
rect 517612 221960 517664 222012
rect 518532 221960 518584 222012
rect 562692 221960 562744 222012
rect 424968 221892 425020 221944
rect 429200 221892 429252 221944
rect 564900 222096 564952 222148
rect 565360 222096 565412 222148
rect 596824 222096 596876 222148
rect 600412 222096 600464 222148
rect 563520 221960 563572 222012
rect 591948 221960 592000 222012
rect 592132 221960 592184 222012
rect 599124 221960 599176 222012
rect 599308 221960 599360 222012
rect 600596 221960 600648 222012
rect 171416 221824 171468 221876
rect 229652 221824 229704 221876
rect 237288 221824 237340 221876
rect 280436 221824 280488 221876
rect 285680 221824 285732 221876
rect 286324 221824 286376 221876
rect 304724 221824 304776 221876
rect 334072 221824 334124 221876
rect 505744 221824 505796 221876
rect 523960 221824 524012 221876
rect 529848 221824 529900 221876
rect 555700 221824 555752 221876
rect 559564 221824 559616 221876
rect 563336 221824 563388 221876
rect 609980 221824 610032 221876
rect 68376 221688 68428 221740
rect 147496 221688 147548 221740
rect 61752 221552 61804 221604
rect 137284 221552 137336 221604
rect 137468 221552 137520 221604
rect 64604 221416 64656 221468
rect 138572 221416 138624 221468
rect 138756 221416 138808 221468
rect 142436 221416 142488 221468
rect 142804 221552 142856 221604
rect 147312 221552 147364 221604
rect 161756 221688 161808 221740
rect 224408 221688 224460 221740
rect 230388 221688 230440 221740
rect 275192 221688 275244 221740
rect 275376 221688 275428 221740
rect 310888 221688 310940 221740
rect 311532 221688 311584 221740
rect 338396 221688 338448 221740
rect 143172 221416 143224 221468
rect 145380 221416 145432 221468
rect 204904 221552 204956 221604
rect 205088 221552 205140 221604
rect 148784 221416 148836 221468
rect 211988 221416 212040 221468
rect 214932 221552 214984 221604
rect 265716 221552 265768 221604
rect 267740 221552 267792 221604
rect 273996 221552 274048 221604
rect 278228 221552 278280 221604
rect 313280 221552 313332 221604
rect 314568 221552 314620 221604
rect 341616 221688 341668 221740
rect 359832 221688 359884 221740
rect 376852 221688 376904 221740
rect 496176 221688 496228 221740
rect 513564 221688 513616 221740
rect 527824 221688 527876 221740
rect 542452 221688 542504 221740
rect 553216 221688 553268 221740
rect 608968 221688 609020 221740
rect 341616 221552 341668 221604
rect 361580 221552 361632 221604
rect 378048 221552 378100 221604
rect 390008 221552 390060 221604
rect 456708 221552 456760 221604
rect 461768 221552 461820 221604
rect 484308 221552 484360 221604
rect 495808 221552 495860 221604
rect 500040 221552 500092 221604
rect 517612 221552 517664 221604
rect 518164 221552 518216 221604
rect 530032 221552 530084 221604
rect 534816 221552 534868 221604
rect 547420 221552 547472 221604
rect 552664 221552 552716 221604
rect 553676 221552 553728 221604
rect 553860 221552 553912 221604
rect 557080 221552 557132 221604
rect 558000 221552 558052 221604
rect 559840 221552 559892 221604
rect 563152 221552 563204 221604
rect 563704 221552 563756 221604
rect 608784 221552 608836 221604
rect 232136 221416 232188 221468
rect 241244 221416 241296 221468
rect 285680 221416 285732 221468
rect 286048 221416 286100 221468
rect 289912 221416 289964 221468
rect 290280 221416 290332 221468
rect 321744 221416 321796 221468
rect 339132 221416 339184 221468
rect 362040 221416 362092 221468
rect 362316 221416 362368 221468
rect 380256 221416 380308 221468
rect 391296 221416 391348 221468
rect 400404 221416 400456 221468
rect 405372 221416 405424 221468
rect 414204 221416 414256 221468
rect 452568 221416 452620 221468
rect 456708 221416 456760 221468
rect 484032 221416 484084 221468
rect 538680 221416 538732 221468
rect 540060 221416 540112 221468
rect 540888 221416 540940 221468
rect 606024 221416 606076 221468
rect 114468 221280 114520 221332
rect 178316 221280 178368 221332
rect 178500 221280 178552 221332
rect 180156 221280 180208 221332
rect 181444 221280 181496 221332
rect 195244 221280 195296 221332
rect 195428 221280 195480 221332
rect 245108 221280 245160 221332
rect 273720 221280 273772 221332
rect 309232 221280 309284 221332
rect 525064 221280 525116 221332
rect 535092 221280 535144 221332
rect 543556 221280 543608 221332
rect 547880 221212 547932 221264
rect 549076 221212 549128 221264
rect 550640 221212 550692 221264
rect 607772 221212 607824 221264
rect 117964 221144 118016 221196
rect 137100 221144 137152 221196
rect 137284 221144 137336 221196
rect 144000 221144 144052 221196
rect 144184 221144 144236 221196
rect 203248 221144 203300 221196
rect 108120 221008 108172 221060
rect 118148 221008 118200 221060
rect 128820 221008 128872 221060
rect 195060 221008 195112 221060
rect 195244 221008 195296 221060
rect 205088 221144 205140 221196
rect 206008 221144 206060 221196
rect 258080 221144 258132 221196
rect 530584 221076 530636 221128
rect 603448 221076 603500 221128
rect 204904 221008 204956 221060
rect 211620 221008 211672 221060
rect 211988 221008 212040 221060
rect 214288 221008 214340 221060
rect 227352 221008 227404 221060
rect 272708 221008 272760 221060
rect 415124 221008 415176 221060
rect 420184 221008 420236 221060
rect 516048 220940 516100 220992
rect 596640 220940 596692 220992
rect 107936 220872 107988 220924
rect 97724 220736 97776 220788
rect 118056 220872 118108 220924
rect 187884 220872 187936 220924
rect 188436 220872 188488 220924
rect 195428 220872 195480 220924
rect 137284 220736 137336 220788
rect 137468 220736 137520 220788
rect 194876 220736 194928 220788
rect 195060 220736 195112 220788
rect 198924 220872 198976 220924
rect 203248 220872 203300 220924
rect 206468 220872 206520 220924
rect 596824 220872 596876 220924
rect 611636 220872 611688 220924
rect 420644 220804 420696 220856
rect 423772 220804 423824 220856
rect 466092 220804 466144 220856
rect 471704 220804 471756 220856
rect 513564 220804 513616 220856
rect 592132 220804 592184 220856
rect 196072 220736 196124 220788
rect 197820 220736 197872 220788
rect 198372 220736 198424 220788
rect 252744 220736 252796 220788
rect 257160 220736 257212 220788
rect 295892 220736 295944 220788
rect 306380 220736 306432 220788
rect 320364 220736 320416 220788
rect 328828 220736 328880 220788
rect 331956 220736 332008 220788
rect 414480 220736 414532 220788
rect 418252 220736 418304 220788
rect 455236 220736 455288 220788
rect 458548 220736 458600 220788
rect 474004 220736 474056 220788
rect 475108 220736 475160 220788
rect 475384 220736 475436 220788
rect 476120 220736 476172 220788
rect 476856 220736 476908 220788
rect 478420 220736 478472 220788
rect 592316 220736 592368 220788
rect 601516 220736 601568 220788
rect 601700 220736 601752 220788
rect 617524 220736 617576 220788
rect 91560 220600 91612 220652
rect 107936 220600 107988 220652
rect 465724 220668 465776 220720
rect 469312 220668 469364 220720
rect 172704 220600 172756 220652
rect 177488 220600 177540 220652
rect 182640 220600 182692 220652
rect 183468 220600 183520 220652
rect 184204 220600 184256 220652
rect 184388 220600 184440 220652
rect 234068 220600 234120 220652
rect 253848 220600 253900 220652
rect 293408 220600 293460 220652
rect 296996 220600 297048 220652
rect 310704 220600 310756 220652
rect 311716 220600 311768 220652
rect 327264 220600 327316 220652
rect 508504 220600 508556 220652
rect 522672 220600 522724 220652
rect 522856 220600 522908 220652
rect 532884 220600 532936 220652
rect 533344 220600 533396 220652
rect 618812 220600 618864 220652
rect 83280 220464 83332 220516
rect 76656 220328 76708 220380
rect 150624 220328 150676 220380
rect 152648 220464 152700 220516
rect 167184 220464 167236 220516
rect 171048 220464 171100 220516
rect 229284 220464 229336 220516
rect 240600 220464 240652 220516
rect 283012 220464 283064 220516
rect 296628 220464 296680 220516
rect 327448 220464 327500 220516
rect 328184 220464 328236 220516
rect 351368 220464 351420 220516
rect 371148 220464 371200 220516
rect 385224 220464 385276 220516
rect 432236 220464 432288 220516
rect 434812 220464 434864 220516
rect 496360 220464 496412 220516
rect 157616 220328 157668 220380
rect 157800 220328 157852 220380
rect 218612 220328 218664 220380
rect 229192 220328 229244 220380
rect 276112 220328 276164 220380
rect 281172 220328 281224 220380
rect 317512 220328 317564 220380
rect 323400 220328 323452 220380
rect 348148 220328 348200 220380
rect 353208 220328 353260 220380
rect 371424 220328 371476 220380
rect 473268 220328 473320 220380
rect 481732 220328 481784 220380
rect 482284 220328 482336 220380
rect 491392 220328 491444 220380
rect 492588 220328 492640 220380
rect 507400 220328 507452 220380
rect 66720 220192 66772 220244
rect 147220 220192 147272 220244
rect 203248 220192 203300 220244
rect 63408 220056 63460 220108
rect 141056 220056 141108 220108
rect 141240 220056 141292 220108
rect 147634 220056 147686 220108
rect 211344 220192 211396 220244
rect 211620 220192 211672 220244
rect 263048 220192 263100 220244
rect 263324 220192 263376 220244
rect 301044 220192 301096 220244
rect 318432 220192 318484 220244
rect 343732 220192 343784 220244
rect 345848 220192 345900 220244
rect 367376 220192 367428 220244
rect 368112 220192 368164 220244
rect 382464 220192 382516 220244
rect 383016 220192 383068 220244
rect 394792 220192 394844 220244
rect 397920 220192 397972 220244
rect 405832 220192 405884 220244
rect 459468 220192 459520 220244
rect 465172 220192 465224 220244
rect 469036 220192 469088 220244
rect 474280 220192 474332 220244
rect 478604 220192 478656 220244
rect 489184 220192 489236 220244
rect 491208 220192 491260 220244
rect 515220 220464 515272 220516
rect 601332 220464 601384 220516
rect 601976 220464 602028 220516
rect 613292 220464 613344 220516
rect 507768 220328 507820 220380
rect 527272 220328 527324 220380
rect 530032 220328 530084 220380
rect 532700 220328 532752 220380
rect 532884 220328 532936 220380
rect 534034 220328 534086 220380
rect 534172 220328 534224 220380
rect 620468 220328 620520 220380
rect 111432 219920 111484 219972
rect 177488 219920 177540 219972
rect 177672 219920 177724 219972
rect 184388 219920 184440 219972
rect 190920 219920 190972 219972
rect 244464 220056 244516 220108
rect 254676 220056 254728 220108
rect 296812 220056 296864 220108
rect 300124 220056 300176 220108
rect 330024 220056 330076 220108
rect 332508 220056 332560 220108
rect 357532 220056 357584 220108
rect 360660 220056 360712 220108
rect 377404 220056 377456 220108
rect 390468 220056 390520 220108
rect 401692 220056 401744 220108
rect 421932 220056 421984 220108
rect 426808 220056 426860 220108
rect 481548 220056 481600 220108
rect 492772 220056 492824 220108
rect 510988 220192 511040 220244
rect 582748 220192 582800 220244
rect 582932 220192 582984 220244
rect 591672 220192 591724 220244
rect 592500 220192 592552 220244
rect 601516 220192 601568 220244
rect 601700 220192 601752 220244
rect 612924 220192 612976 220244
rect 505192 220056 505244 220108
rect 521568 220056 521620 220108
rect 543372 220056 543424 220108
rect 548340 220056 548392 220108
rect 572628 220056 572680 220108
rect 627092 220056 627144 220108
rect 647332 220056 647384 220108
rect 652760 220056 652812 220108
rect 124680 219784 124732 219836
rect 193496 219784 193548 219836
rect 197268 219784 197320 219836
rect 249892 219920 249944 219972
rect 280068 219920 280120 219972
rect 313924 219920 313976 219972
rect 493784 219920 493836 219972
rect 508228 219920 508280 219972
rect 522672 219920 522724 219972
rect 533344 219920 533396 219972
rect 534080 219920 534132 219972
rect 537300 219920 537352 219972
rect 537484 219852 537536 219904
rect 548524 219988 548576 220040
rect 553860 219988 553912 220040
rect 554044 219988 554096 220040
rect 562876 219988 562928 220040
rect 563244 219988 563296 220040
rect 572076 219988 572128 220040
rect 592040 219920 592092 219972
rect 543740 219852 543792 219904
rect 572628 219852 572680 219904
rect 572812 219852 572864 219904
rect 582196 219852 582248 219904
rect 582380 219852 582432 219904
rect 591856 219852 591908 219904
rect 621572 219852 621624 219904
rect 207480 219784 207532 219836
rect 257344 219784 257396 219836
rect 293868 219784 293920 219836
rect 299940 219784 299992 219836
rect 504364 219784 504416 219836
rect 515220 219784 515272 219836
rect 517428 219716 517480 219768
rect 539048 219716 539100 219768
rect 540244 219716 540296 219768
rect 548524 219716 548576 219768
rect 549904 219716 549956 219768
rect 553216 219716 553268 219768
rect 553354 219716 553406 219768
rect 570512 219716 570564 219768
rect 574836 219716 574888 219768
rect 623780 219716 623832 219768
rect 137284 219648 137336 219700
rect 152648 219648 152700 219700
rect 153108 219648 153160 219700
rect 214104 219648 214156 219700
rect 217416 219648 217468 219700
rect 265164 219648 265216 219700
rect 273076 219580 273128 219632
rect 279240 219580 279292 219632
rect 464988 219580 465040 219632
rect 471980 219580 472032 219632
rect 497280 219580 497332 219632
rect 562876 219580 562928 219632
rect 563060 219580 563112 219632
rect 625436 219580 625488 219632
rect 131028 219512 131080 219564
rect 137468 219512 137520 219564
rect 137928 219512 137980 219564
rect 203064 219512 203116 219564
rect 203248 219512 203300 219564
rect 205824 219512 205876 219564
rect 406200 219512 406252 219564
rect 412732 219512 412784 219564
rect 80796 219376 80848 219428
rect 90364 219376 90416 219428
rect 90732 219376 90784 219428
rect 106924 219376 106976 219428
rect 117872 219376 117924 219428
rect 123484 219376 123536 219428
rect 132776 219376 132828 219428
rect 140044 219376 140096 219428
rect 142804 219376 142856 219428
rect 198004 219376 198056 219428
rect 199844 219376 199896 219428
rect 204720 219376 204772 219428
rect 213000 219376 213052 219428
rect 217232 219376 217284 219428
rect 217968 219376 218020 219428
rect 220084 219376 220136 219428
rect 224040 219376 224092 219428
rect 232504 219376 232556 219428
rect 232964 219376 233016 219428
rect 93216 219240 93268 219292
rect 93768 219240 93820 219292
rect 108304 219240 108356 219292
rect 149980 219240 150032 219292
rect 150164 219240 150216 219292
rect 161296 219240 161348 219292
rect 85304 219104 85356 219156
rect 117872 219104 117924 219156
rect 123852 219104 123904 219156
rect 127072 219104 127124 219156
rect 130476 219104 130528 219156
rect 169024 219240 169076 219292
rect 169208 219240 169260 219292
rect 162308 219104 162360 219156
rect 180984 219104 181036 219156
rect 182640 219240 182692 219292
rect 183284 219240 183336 219292
rect 183652 219240 183704 219292
rect 226984 219240 227036 219292
rect 238116 219240 238168 219292
rect 239404 219240 239456 219292
rect 246396 219376 246448 219428
rect 286048 219376 286100 219428
rect 291660 219376 291712 219428
rect 324688 219376 324740 219428
rect 273076 219240 273128 219292
rect 325424 219240 325476 219292
rect 326344 219240 326396 219292
rect 327540 219240 327592 219292
rect 345572 219376 345624 219428
rect 352380 219376 352432 219428
rect 344100 219240 344152 219292
rect 347044 219240 347096 219292
rect 199384 219104 199436 219156
rect 204720 219104 204772 219156
rect 246212 219104 246264 219156
rect 262680 219104 262732 219156
rect 291844 219104 291896 219156
rect 70860 218968 70912 219020
rect 132776 218968 132828 219020
rect 132960 218968 133012 219020
rect 133788 218968 133840 219020
rect 137100 218968 137152 219020
rect 142804 218968 142856 219020
rect 143172 218968 143224 219020
rect 62580 218832 62632 218884
rect 76472 218832 76524 218884
rect 83924 218832 83976 218884
rect 60096 218696 60148 218748
rect 69664 218696 69716 218748
rect 77208 218696 77260 218748
rect 143632 218832 143684 218884
rect 146208 218832 146260 218884
rect 152464 218968 152516 219020
rect 204904 218968 204956 219020
rect 206652 218968 206704 219020
rect 255964 218968 256016 219020
rect 259092 218968 259144 219020
rect 293868 218968 293920 219020
rect 294420 218968 294472 219020
rect 311716 219104 311768 219156
rect 315672 219104 315724 219156
rect 318064 219104 318116 219156
rect 320916 219104 320968 219156
rect 340144 219104 340196 219156
rect 354404 219104 354456 219156
rect 355508 219104 355560 219156
rect 417792 219376 417844 219428
rect 421012 219444 421064 219496
rect 428280 219376 428332 219428
rect 432052 219512 432104 219564
rect 430212 219376 430264 219428
rect 432696 219376 432748 219428
rect 435088 219376 435140 219428
rect 437020 219444 437072 219496
rect 493968 219444 494020 219496
rect 613108 219444 613160 219496
rect 613292 219444 613344 219496
rect 628104 219444 628156 219496
rect 535460 219308 535512 219360
rect 536380 219308 536432 219360
rect 537300 219308 537352 219360
rect 539692 219308 539744 219360
rect 543372 219308 543424 219360
rect 544292 219308 544344 219360
rect 358728 219240 358780 219292
rect 364984 219240 365036 219292
rect 383568 219240 383620 219292
rect 387064 219240 387116 219292
rect 475752 219240 475804 219292
rect 482560 219240 482612 219292
rect 546316 219240 546368 219292
rect 553492 219240 553544 219292
rect 513012 219172 513064 219224
rect 519176 219172 519228 219224
rect 562508 219308 562560 219360
rect 562876 219308 562928 219360
rect 563244 219308 563296 219360
rect 563428 219308 563480 219360
rect 573180 219308 573232 219360
rect 573456 219308 573508 219360
rect 574836 219308 574888 219360
rect 582196 219308 582248 219360
rect 582380 219308 582432 219360
rect 591856 219308 591908 219360
rect 592316 219308 592368 219360
rect 366272 219104 366324 219156
rect 373080 219104 373132 219156
rect 373816 219104 373868 219156
rect 407580 219104 407632 219156
rect 411904 219104 411956 219156
rect 419264 219104 419316 219156
rect 422668 219104 422720 219156
rect 507216 219104 507268 219156
rect 509516 219104 509568 219156
rect 537116 219104 537168 219156
rect 539232 219104 539284 219156
rect 543740 219104 543792 219156
rect 553952 219172 554004 219224
rect 563612 219172 563664 219224
rect 570144 219172 570196 219224
rect 572352 219172 572404 219224
rect 582932 219172 582984 219224
rect 591672 219172 591724 219224
rect 592500 219172 592552 219224
rect 601516 219172 601568 219224
rect 601700 219172 601752 219224
rect 571432 219104 571484 219156
rect 300768 218968 300820 219020
rect 328828 218968 328880 219020
rect 333704 218968 333756 219020
rect 352564 218968 352616 219020
rect 355692 218968 355744 219020
rect 369124 218968 369176 219020
rect 373724 218968 373776 219020
rect 380164 218968 380216 219020
rect 384672 218968 384724 219020
rect 393964 218968 394016 219020
rect 402060 218968 402112 219020
rect 407764 218968 407816 219020
rect 460204 218968 460256 219020
rect 461124 218968 461176 219020
rect 532148 218968 532200 219020
rect 532608 218968 532660 219020
rect 538864 218968 538916 219020
rect 542452 218968 542504 219020
rect 546592 218968 546644 219020
rect 546960 218968 547012 219020
rect 552848 218968 552900 219020
rect 553492 218968 553544 219020
rect 509516 218900 509568 218952
rect 518716 218900 518768 218952
rect 162308 218832 162360 218884
rect 162492 218832 162544 218884
rect 215944 218832 215996 218884
rect 216312 218832 216364 218884
rect 224040 218832 224092 218884
rect 225972 218832 226024 218884
rect 93768 218560 93820 218612
rect 140228 218560 140280 218612
rect 140412 218560 140464 218612
rect 142620 218560 142672 218612
rect 149336 218696 149388 218748
rect 149520 218696 149572 218748
rect 150348 218696 150400 218748
rect 148508 218560 148560 218612
rect 149980 218560 150032 218612
rect 156328 218696 156380 218748
rect 156972 218696 157024 218748
rect 161940 218696 161992 218748
rect 151176 218560 151228 218612
rect 153108 218560 153160 218612
rect 153660 218560 153712 218612
rect 213184 218696 213236 218748
rect 219900 218696 219952 218748
rect 264244 218696 264296 218748
rect 162308 218560 162360 218612
rect 163964 218560 164016 218612
rect 165620 218560 165672 218612
rect 166816 218560 166868 218612
rect 167000 218560 167052 218612
rect 169208 218560 169260 218612
rect 170220 218560 170272 218612
rect 180800 218560 180852 218612
rect 180984 218560 181036 218612
rect 192484 218560 192536 218612
rect 193128 218560 193180 218612
rect 243544 218560 243596 218612
rect 253020 218560 253072 218612
rect 262680 218560 262732 218612
rect 274548 218832 274600 218884
rect 280804 218832 280856 218884
rect 280988 218832 281040 218884
rect 312544 218832 312596 218884
rect 314292 218832 314344 218884
rect 329012 218832 329064 218884
rect 337476 218832 337528 218884
rect 358084 218832 358136 218884
rect 366732 218832 366784 218884
rect 378692 218832 378744 218884
rect 386144 218832 386196 218884
rect 396724 218832 396776 218884
rect 402704 218832 402756 218884
rect 409144 218832 409196 218884
rect 411996 218832 412048 218884
rect 412456 218832 412508 218884
rect 485044 218832 485096 218884
rect 490656 218832 490708 218884
rect 266084 218696 266136 218748
rect 302884 218696 302936 218748
rect 307484 218696 307536 218748
rect 337108 218696 337160 218748
rect 340512 218696 340564 218748
rect 360844 218696 360896 218748
rect 379152 218696 379204 218748
rect 392124 218696 392176 218748
rect 395804 218696 395856 218748
rect 404544 218696 404596 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 509240 218628 509292 218680
rect 518854 218628 518906 218680
rect 527272 218628 527324 218680
rect 531964 218900 532016 218952
rect 537852 218832 537904 218884
rect 543924 218832 543976 218884
rect 544108 218832 544160 218884
rect 553768 218832 553820 218884
rect 554228 218968 554280 219020
rect 562876 218832 562928 218884
rect 528652 218764 528704 218816
rect 534264 218764 534316 218816
rect 572352 219036 572404 219088
rect 572996 219036 573048 219088
rect 571800 218900 571852 218952
rect 572536 218900 572588 218952
rect 573180 218900 573232 218952
rect 575020 218900 575072 218952
rect 605656 218832 605708 218884
rect 267740 218560 267792 218612
rect 272892 218560 272944 218612
rect 296996 218560 297048 218612
rect 351552 218560 351604 218612
rect 355324 218560 355376 218612
rect 546960 218696 547012 218748
rect 547144 218696 547196 218748
rect 552664 218696 552716 218748
rect 553262 218696 553314 218748
rect 570328 218696 570380 218748
rect 575388 218696 575440 218748
rect 597468 218696 597520 218748
rect 469864 218492 469916 218544
rect 470968 218492 471020 218544
rect 518716 218492 518768 218544
rect 538864 218560 538916 218612
rect 100484 218424 100536 218476
rect 108304 218424 108356 218476
rect 126336 218424 126388 218476
rect 126888 218424 126940 218476
rect 127072 218424 127124 218476
rect 174176 218424 174228 218476
rect 174360 218424 174412 218476
rect 183652 218424 183704 218476
rect 186780 218424 186832 218476
rect 235264 218424 235316 218476
rect 239772 218424 239824 218476
rect 272524 218424 272576 218476
rect 279516 218424 279568 218476
rect 280988 218424 281040 218476
rect 286140 218424 286192 218476
rect 306380 218424 306432 218476
rect 380532 218424 380584 218476
rect 384304 218424 384356 218476
rect 531964 218424 532016 218476
rect 450544 218356 450596 218408
rect 453580 218356 453632 218408
rect 519084 218356 519136 218408
rect 528560 218356 528612 218408
rect 75644 218288 75696 218340
rect 83464 218288 83516 218340
rect 107292 218288 107344 218340
rect 157984 218288 158036 218340
rect 56324 218152 56376 218204
rect 62764 218152 62816 218204
rect 79784 218152 79836 218204
rect 82084 218152 82136 218204
rect 113916 218152 113968 218204
rect 161572 218288 161624 218340
rect 161940 218288 161992 218340
rect 165160 218288 165212 218340
rect 213000 218288 213052 218340
rect 213276 218288 213328 218340
rect 216680 218288 216732 218340
rect 159824 218152 159876 218204
rect 162492 218152 162544 218204
rect 163596 218152 163648 218204
rect 55956 218016 56008 218068
rect 56508 218016 56560 218068
rect 58440 218016 58492 218068
rect 61384 218016 61436 218068
rect 64236 218016 64288 218068
rect 64788 218016 64840 218068
rect 72516 218016 72568 218068
rect 73068 218016 73120 218068
rect 75000 218016 75052 218068
rect 75828 218016 75880 218068
rect 79140 218016 79192 218068
rect 79968 218016 80020 218068
rect 84936 218016 84988 218068
rect 85488 218016 85540 218068
rect 87420 218016 87472 218068
rect 88248 218016 88300 218068
rect 97356 218016 97408 218068
rect 97908 218016 97960 218068
rect 99840 218016 99892 218068
rect 100668 218016 100720 218068
rect 101496 218016 101548 218068
rect 102048 218016 102100 218068
rect 103980 218016 104032 218068
rect 104808 218016 104860 218068
rect 110328 218016 110380 218068
rect 111064 218016 111116 218068
rect 112260 218016 112312 218068
rect 112904 218016 112956 218068
rect 116400 218016 116452 218068
rect 117228 218016 117280 218068
rect 120540 218016 120592 218068
rect 159456 218016 159508 218068
rect 160008 218016 160060 218068
rect 165620 218016 165672 218068
rect 166816 218152 166868 218204
rect 168104 218152 168156 218204
rect 170864 218152 170916 218204
rect 171876 218152 171928 218204
rect 166080 218084 166132 218136
rect 166540 218084 166592 218136
rect 167000 218016 167052 218068
rect 167736 218016 167788 218068
rect 168288 218016 168340 218068
rect 173532 218016 173584 218068
rect 174176 218016 174228 218068
rect 174360 218016 174412 218068
rect 175188 218016 175240 218068
rect 176016 218152 176068 218204
rect 176476 218152 176528 218204
rect 180156 218152 180208 218204
rect 224224 218288 224276 218340
rect 228180 218288 228232 218340
rect 229192 218288 229244 218340
rect 365628 218288 365680 218340
rect 373264 218288 373316 218340
rect 426808 218288 426860 218340
rect 429384 218288 429436 218340
rect 435916 218288 435968 218340
rect 436284 218288 436336 218340
rect 479524 218288 479576 218340
rect 480352 218288 480404 218340
rect 224040 218152 224092 218204
rect 224684 218152 224736 218204
rect 224868 218152 224920 218204
rect 225512 218152 225564 218204
rect 225696 218152 225748 218204
rect 226156 218152 226208 218204
rect 229836 218152 229888 218204
rect 231124 218152 231176 218204
rect 232320 218152 232372 218204
rect 233148 218152 233200 218204
rect 233976 218152 234028 218204
rect 234528 218152 234580 218204
rect 236460 218152 236512 218204
rect 237012 218152 237064 218204
rect 176292 218016 176344 218068
rect 176568 218016 176620 218068
rect 177856 218016 177908 218068
rect 180800 218016 180852 218068
rect 182088 218016 182140 218068
rect 194876 218016 194928 218068
rect 195888 218016 195940 218068
rect 198924 218016 198976 218068
rect 200028 218016 200080 218068
rect 200856 218016 200908 218068
rect 201408 218016 201460 218068
rect 203340 218016 203392 218068
rect 203892 218016 203944 218068
rect 204996 218016 205048 218068
rect 206008 218016 206060 218068
rect 209136 218016 209188 218068
rect 209688 218016 209740 218068
rect 215760 218016 215812 218068
rect 216496 218016 216548 218068
rect 216680 218016 216732 218068
rect 249064 218152 249116 218204
rect 249524 218152 249576 218204
rect 251824 218152 251876 218204
rect 302700 218152 302752 218204
rect 304724 218152 304776 218204
rect 310980 218152 311032 218204
rect 315304 218152 315356 218204
rect 348884 218152 348936 218204
rect 351184 218152 351236 218204
rect 364800 218152 364852 218204
rect 367744 218152 367796 218204
rect 368940 218152 368992 218204
rect 369768 218152 369820 218204
rect 377220 218152 377272 218204
rect 382832 218152 382884 218204
rect 394424 218152 394476 218204
rect 402244 218152 402296 218204
rect 422760 218152 422812 218204
rect 425428 218152 425480 218204
rect 426072 218152 426124 218204
rect 427912 218152 427964 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 455052 218152 455104 218204
rect 460204 218152 460256 218204
rect 461952 218152 462004 218204
rect 466000 218152 466052 218204
rect 509884 218152 509936 218204
rect 510528 218152 510580 218204
rect 533344 218288 533396 218340
rect 546316 218424 546368 218476
rect 546592 218424 546644 218476
rect 563198 218424 563250 218476
rect 572536 218560 572588 218612
rect 584404 218560 584456 218612
rect 573088 218424 573140 218476
rect 574652 218424 574704 218476
rect 575664 218424 575716 218476
rect 582104 218424 582156 218476
rect 582748 218424 582800 218476
rect 534172 218288 534224 218340
rect 539232 218288 539284 218340
rect 570880 218356 570932 218408
rect 571064 218356 571116 218408
rect 601424 218356 601476 218408
rect 607496 218356 607548 218408
rect 573732 218288 573784 218340
rect 573916 218288 573968 218340
rect 577688 218288 577740 218340
rect 578240 218288 578292 218340
rect 582564 218288 582616 218340
rect 592132 218288 592184 218340
rect 597744 218288 597796 218340
rect 563612 218220 563664 218272
rect 564532 218220 564584 218272
rect 564808 218220 564860 218272
rect 571800 218220 571852 218272
rect 242256 218016 242308 218068
rect 242716 218016 242768 218068
rect 244740 218016 244792 218068
rect 247684 218016 247736 218068
rect 248880 218016 248932 218068
rect 249708 218016 249760 218068
rect 250536 218016 250588 218068
rect 251088 218016 251140 218068
rect 258816 218016 258868 218068
rect 259276 218016 259328 218068
rect 262956 218016 263008 218068
rect 263508 218016 263560 218068
rect 265440 218016 265492 218068
rect 266268 218016 266320 218068
rect 267096 218016 267148 218068
rect 267556 218016 267608 218068
rect 269580 218016 269632 218068
rect 273904 218016 273956 218068
rect 277860 218016 277912 218068
rect 278412 218016 278464 218068
rect 282000 218016 282052 218068
rect 282644 218016 282696 218068
rect 283656 218016 283708 218068
rect 284116 218016 284168 218068
rect 287796 218016 287848 218068
rect 288256 218016 288308 218068
rect 298560 218016 298612 218068
rect 299204 218016 299256 218068
rect 299388 218016 299440 218068
rect 300308 218016 300360 218068
rect 304356 218016 304408 218068
rect 305644 218016 305696 218068
rect 306840 218016 306892 218068
rect 307668 218016 307720 218068
rect 312636 218016 312688 218068
rect 314568 218016 314620 218068
rect 315120 218016 315172 218068
rect 315856 218016 315908 218068
rect 319260 218016 319312 218068
rect 319996 218016 320048 218068
rect 325056 218016 325108 218068
rect 325608 218016 325660 218068
rect 329196 218016 329248 218068
rect 330484 218016 330536 218068
rect 330852 218016 330904 218068
rect 333152 218016 333204 218068
rect 333336 218016 333388 218068
rect 333888 218016 333940 218068
rect 335820 218016 335872 218068
rect 336464 218016 336516 218068
rect 339960 218016 340012 218068
rect 340696 218016 340748 218068
rect 348240 218016 348292 218068
rect 349068 218016 349120 218068
rect 354036 218016 354088 218068
rect 354588 218016 354640 218068
rect 356520 218016 356572 218068
rect 357348 218016 357400 218068
rect 358176 218016 358228 218068
rect 359464 218016 359516 218068
rect 366456 218016 366508 218068
rect 366916 218016 366968 218068
rect 369768 218016 369820 218068
rect 370504 218016 370556 218068
rect 374736 218016 374788 218068
rect 375288 218016 375340 218068
rect 378876 218016 378928 218068
rect 379336 218016 379388 218068
rect 381360 218016 381412 218068
rect 381912 218016 381964 218068
rect 385500 218016 385552 218068
rect 386328 218016 386380 218068
rect 387156 218016 387208 218068
rect 388444 218016 388496 218068
rect 389640 218016 389692 218068
rect 390284 218016 390336 218068
rect 393780 218016 393832 218068
rect 394608 218016 394660 218068
rect 395436 218016 395488 218068
rect 395988 218016 396040 218068
rect 399576 218016 399628 218068
rect 400036 218016 400088 218068
rect 403532 218016 403584 218068
rect 404268 218016 404320 218068
rect 410340 218016 410392 218068
rect 410892 218016 410944 218068
rect 416136 218016 416188 218068
rect 416688 218016 416740 218068
rect 418620 218016 418672 218068
rect 419448 218016 419500 218068
rect 420276 218016 420328 218068
rect 420828 218016 420880 218068
rect 424416 218016 424468 218068
rect 426992 218016 427044 218068
rect 427728 218016 427780 218068
rect 428464 218016 428516 218068
rect 429108 218016 429160 218068
rect 430672 218016 430724 218068
rect 432696 218016 432748 218068
rect 433800 218016 433852 218068
rect 436836 218016 436888 218068
rect 437480 218016 437532 218068
rect 438492 218016 438544 218068
rect 438952 218016 439004 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 462964 218016 463016 218068
rect 464436 218016 464488 218068
rect 467104 218016 467156 218068
rect 467840 218016 467892 218068
rect 471704 218016 471756 218068
rect 472624 218016 472676 218068
rect 482836 218016 482888 218068
rect 485044 218016 485096 218068
rect 491392 218016 491444 218068
rect 492312 218016 492364 218068
rect 505100 218016 505152 218068
rect 525248 218016 525300 218068
rect 533344 218016 533396 218068
rect 537852 218016 537904 218068
rect 543924 218152 543976 218204
rect 575020 218152 575072 218204
rect 616144 218152 616196 218204
rect 544108 218084 544160 218136
rect 554228 218084 554280 218136
rect 543694 218016 543746 218068
rect 543832 217948 543884 218000
rect 572904 218084 572956 218136
rect 555700 217948 555752 218000
rect 563612 217948 563664 218000
rect 563796 217948 563848 218000
rect 573272 217948 573324 218000
rect 574652 217948 574704 218000
rect 676404 218084 676456 218136
rect 677600 218084 677652 218136
rect 577688 218016 577740 218068
rect 629392 218016 629444 218068
rect 577320 217948 577372 218000
rect 447140 217812 447192 217864
rect 447784 217812 447836 217864
rect 448612 217812 448664 217864
rect 449440 217812 449492 217864
rect 498200 217812 498252 217864
rect 499120 217812 499172 217864
rect 543188 217812 543240 217864
rect 508044 217744 508096 217796
rect 509516 217744 509568 217796
rect 523776 217744 523828 217796
rect 529112 217744 529164 217796
rect 509424 217540 509476 217592
rect 519176 217540 519228 217592
rect 528284 217540 528336 217592
rect 528652 217540 528704 217592
rect 534264 217540 534316 217592
rect 544108 217676 544160 217728
rect 548892 217812 548944 217864
rect 601516 217812 601568 217864
rect 601976 217812 602028 217864
rect 609152 217812 609204 217864
rect 676680 217812 676732 217864
rect 677048 217812 677100 217864
rect 592132 217676 592184 217728
rect 592316 217676 592368 217728
rect 594248 217676 594300 217728
rect 594432 217676 594484 217728
rect 601332 217676 601384 217728
rect 601700 217676 601752 217728
rect 605840 217676 605892 217728
rect 606208 217676 606260 217728
rect 615684 217676 615736 217728
rect 543464 217540 543516 217592
rect 543832 217540 543884 217592
rect 545764 217540 545816 217592
rect 563796 217540 563848 217592
rect 564532 217540 564584 217592
rect 572260 217540 572312 217592
rect 572812 217540 572864 217592
rect 575388 217540 575440 217592
rect 575664 217540 575716 217592
rect 601654 217540 601706 217592
rect 601792 217540 601844 217592
rect 607312 217540 607364 217592
rect 538496 217404 538548 217456
rect 594432 217404 594484 217456
rect 594616 217404 594668 217456
rect 604000 217404 604052 217456
rect 605656 217404 605708 217456
rect 627920 217404 627972 217456
rect 146714 217200 146766 217252
rect 152464 217200 152516 217252
rect 525938 217200 525990 217252
rect 526536 217200 526588 217252
rect 519084 217064 519136 217116
rect 528468 217064 528520 217116
rect 536012 217200 536064 217252
rect 601516 217268 601568 217320
rect 601700 217268 601752 217320
rect 533712 217064 533764 217116
rect 594616 217132 594668 217184
rect 594800 217132 594852 217184
rect 592132 216996 592184 217048
rect 595168 216996 595220 217048
rect 572996 216928 573048 216980
rect 528560 216792 528612 216844
rect 575572 216928 575624 216980
rect 577320 216928 577372 216980
rect 591948 216928 592000 216980
rect 596640 217064 596692 217116
rect 601976 217200 602028 217252
rect 606208 217200 606260 217252
rect 601792 217064 601844 217116
rect 603080 217064 603132 217116
rect 603264 217064 603316 217116
rect 610624 217064 610676 217116
rect 601148 216928 601200 216980
rect 601516 216928 601568 216980
rect 625252 216928 625304 216980
rect 573456 216792 573508 216844
rect 596640 216792 596692 216844
rect 521292 216656 521344 216708
rect 575020 216656 575072 216708
rect 584404 216656 584456 216708
rect 614488 216792 614540 216844
rect 597744 216656 597796 216708
rect 601654 216656 601706 216708
rect 601792 216656 601844 216708
rect 605104 216656 605156 216708
rect 605840 216656 605892 216708
rect 606760 216656 606812 216708
rect 607496 216656 607548 216708
rect 614120 216656 614172 216708
rect 534080 216520 534132 216572
rect 543648 216520 543700 216572
rect 547788 216520 547840 216572
rect 554596 216520 554648 216572
rect 555056 216520 555108 216572
rect 562692 216520 562744 216572
rect 563336 216520 563388 216572
rect 623320 216452 623372 216504
rect 557080 216384 557132 216436
rect 558552 216384 558604 216436
rect 562508 216384 562560 216436
rect 571064 216384 571116 216436
rect 571248 216384 571300 216436
rect 574652 216316 574704 216368
rect 621112 216316 621164 216368
rect 582564 216180 582616 216232
rect 597560 216180 597612 216232
rect 574652 215908 574704 215960
rect 574100 215772 574152 215824
rect 619640 216044 619692 216096
rect 623044 215908 623096 215960
rect 633808 215908 633860 215960
rect 590108 215568 590160 215620
rect 595720 215568 595772 215620
rect 575388 215432 575440 215484
rect 575204 215296 575256 215348
rect 576400 215296 576452 215348
rect 612280 215228 612332 215280
rect 574284 215092 574336 215144
rect 620008 215092 620060 215144
rect 676220 215092 676272 215144
rect 677232 215092 677284 215144
rect 574836 214956 574888 215008
rect 622400 214956 622452 215008
rect 663524 214888 663576 214940
rect 664444 214888 664496 214940
rect 576032 214820 576084 214872
rect 626080 214820 626132 214872
rect 574468 214684 574520 214736
rect 616696 214684 616748 214736
rect 616880 214684 616932 214736
rect 617800 214684 617852 214736
rect 658740 214684 658792 214736
rect 661684 214684 661736 214736
rect 574652 214548 574704 214600
rect 628288 214548 628340 214600
rect 631416 214548 631468 214600
rect 632704 214548 632756 214600
rect 656808 214548 656860 214600
rect 658924 214548 658976 214600
rect 662052 214548 662104 214600
rect 663248 214548 663300 214600
rect 608784 214412 608836 214464
rect 609520 214412 609572 214464
rect 611452 214412 611504 214464
rect 611820 214412 611872 214464
rect 616696 214412 616748 214464
rect 624424 214412 624476 214464
rect 627736 214140 627788 214192
rect 631048 214140 631100 214192
rect 35808 213936 35860 213988
rect 40684 213936 40736 213988
rect 612740 213868 612792 213920
rect 615040 213868 615092 213920
rect 637580 213868 637632 213920
rect 638224 213868 638276 213920
rect 639972 213868 640024 213920
rect 643192 213868 643244 213920
rect 654876 213868 654928 213920
rect 655428 213868 655480 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 576400 213732 576452 213784
rect 598480 213732 598532 213784
rect 638040 213732 638092 213784
rect 640432 213732 640484 213784
rect 644940 213732 644992 213784
rect 646872 213732 646924 213784
rect 660948 213732 661000 213784
rect 662972 213732 663024 213784
rect 575020 213596 575072 213648
rect 601240 213596 601292 213648
rect 641628 213596 641680 213648
rect 650644 213596 650696 213648
rect 652024 213596 652076 213648
rect 658004 213596 658056 213648
rect 659568 213596 659620 213648
rect 664904 213596 664956 213648
rect 603080 213528 603132 213580
rect 604552 213528 604604 213580
rect 574100 213460 574152 213512
rect 601792 213460 601844 213512
rect 642180 213460 642232 213512
rect 659384 213460 659436 213512
rect 574100 213324 574152 213376
rect 602344 213324 602396 213376
rect 602528 213324 602580 213376
rect 622768 213324 622820 213376
rect 635556 213324 635608 213376
rect 651840 213324 651892 213376
rect 652852 213324 652904 213376
rect 660212 213324 660264 213376
rect 575572 213188 575624 213240
rect 603080 213188 603132 213240
rect 623964 213188 624016 213240
rect 629944 213188 629996 213240
rect 643836 213188 643888 213240
rect 665272 213188 665324 213240
rect 676220 213188 676272 213240
rect 676864 213188 676916 213240
rect 650460 212984 650512 213036
rect 651288 212984 651340 213036
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 632888 212848 632940 212900
rect 634360 212848 634412 212900
rect 636660 212780 636712 212832
rect 639604 212780 639656 212832
rect 578516 211624 578568 211676
rect 580448 211624 580500 211676
rect 612924 211624 612976 211676
rect 613384 211624 613436 211676
rect 35808 211148 35860 211200
rect 41696 211148 41748 211200
rect 599216 210060 599268 210112
rect 599584 210060 599636 210112
rect 579252 209788 579304 209840
rect 581736 209788 581788 209840
rect 591304 208632 591356 208684
rect 632152 209516 632204 209568
rect 652208 209516 652260 209568
rect 667020 209040 667072 209092
rect 35808 208360 35860 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 580448 207612 580500 207664
rect 589464 207612 589516 207664
rect 581736 206252 581788 206304
rect 589648 206252 589700 206304
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 45468 196596 45520 196648
rect 48596 196596 48648 196648
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 668124 194148 668176 194200
rect 670792 194148 670844 194200
rect 668032 192516 668084 192568
rect 669044 192516 669096 192568
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 669136 189252 669188 189304
rect 670792 189252 670844 189304
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 668032 184356 668084 184408
rect 669596 184356 669648 184408
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 583208 175244 583260 175296
rect 589464 175312 589516 175364
rect 667940 174836 667992 174888
rect 669780 174836 669832 174888
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 581644 171096 581696 171148
rect 589464 171096 589516 171148
rect 579528 170960 579580 171012
rect 583208 170960 583260 171012
rect 582380 169736 582432 169788
rect 589464 169736 589516 169788
rect 578332 169668 578384 169720
rect 580908 169668 580960 169720
rect 579620 168376 579672 168428
rect 589464 168376 589516 168428
rect 578976 167152 579028 167204
rect 581644 167152 581696 167204
rect 581644 167016 581696 167068
rect 589464 167016 589516 167068
rect 669136 166064 669188 166116
rect 670148 166064 670200 166116
rect 578884 165520 578936 165572
rect 582380 165520 582432 165572
rect 668032 164772 668084 164824
rect 670332 164772 670384 164824
rect 585968 164228 586020 164280
rect 589464 164228 589516 164280
rect 584404 162868 584456 162920
rect 589464 162868 589516 162920
rect 675852 162800 675904 162852
rect 678244 162800 678296 162852
rect 676036 162596 676088 162648
rect 679624 162596 679676 162648
rect 675852 161712 675904 161764
rect 681004 161712 681056 161764
rect 580448 161440 580500 161492
rect 589464 161440 589516 161492
rect 582380 160080 582432 160132
rect 589464 160080 589516 160132
rect 579252 160012 579304 160064
rect 581644 160012 581696 160064
rect 581828 158788 581880 158840
rect 589464 158788 589516 158840
rect 579160 158652 579212 158704
rect 585968 158652 586020 158704
rect 585784 157360 585836 157412
rect 589464 157360 589516 157412
rect 579528 155864 579580 155916
rect 584404 155864 584456 155916
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 578240 154504 578292 154556
rect 580448 154504 580500 154556
rect 580264 153212 580316 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 582380 152736 582432 152788
rect 583024 151784 583076 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 581828 150560 581880 150612
rect 581644 150424 581696 150476
rect 589464 150424 589516 150476
rect 668676 150220 668728 150272
rect 670792 150220 670844 150272
rect 579528 147364 579580 147416
rect 585784 147364 585836 147416
rect 587348 146276 587400 146328
rect 589372 146276 589424 146328
rect 578884 145528 578936 145580
rect 589188 145528 589240 145580
rect 585784 144916 585836 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 578516 143284 578568 143336
rect 580264 143284 580316 143336
rect 580448 142128 580500 142180
rect 589464 142128 589516 142180
rect 579528 140564 579580 140616
rect 583024 140564 583076 140616
rect 584404 139408 584456 139460
rect 589464 139408 589516 139460
rect 578700 139340 578752 139392
rect 581644 139340 581696 139392
rect 581644 136620 581696 136672
rect 589464 136620 589516 136672
rect 667940 136416 667992 136468
rect 669964 136416 670016 136468
rect 578332 135872 578384 135924
rect 587348 135872 587400 135924
rect 587164 135260 587216 135312
rect 589280 135260 589332 135312
rect 578240 134240 578292 134292
rect 585784 134240 585836 134292
rect 585968 133900 586020 133952
rect 589464 133900 589516 133952
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 579252 133152 579304 133204
rect 589096 133152 589148 133204
rect 582380 131724 582432 131776
rect 589924 131724 589976 131776
rect 579528 129684 579580 129736
rect 582380 129684 582432 129736
rect 583024 128324 583076 128376
rect 589464 128324 589516 128376
rect 578332 128256 578384 128308
rect 580448 128256 580500 128308
rect 580264 126964 580316 127016
rect 589464 126964 589516 127016
rect 585784 124176 585836 124228
rect 589464 124176 589516 124228
rect 579252 124108 579304 124160
rect 584404 124108 584456 124160
rect 579252 122816 579304 122868
rect 589464 122816 589516 122868
rect 584404 121456 584456 121508
rect 589464 121456 589516 121508
rect 579068 121116 579120 121168
rect 581644 121116 581696 121168
rect 582012 120708 582064 120760
rect 590108 120708 590160 120760
rect 578516 118600 578568 118652
rect 587164 118600 587216 118652
rect 668032 118328 668084 118380
rect 670148 118328 670200 118380
rect 583208 117308 583260 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 682384 117240 682436 117292
rect 579528 116900 579580 116952
rect 585968 116900 586020 116952
rect 587808 115948 587860 116000
rect 589464 115948 589516 116000
rect 585140 115336 585192 115388
rect 589924 115336 589976 115388
rect 579068 115200 579120 115252
rect 587808 115200 587860 115252
rect 587164 114520 587216 114572
rect 589832 114520 589884 114572
rect 579528 114384 579580 114436
rect 591304 114384 591356 114436
rect 668124 114112 668176 114164
rect 669964 114112 670016 114164
rect 579528 113092 579580 113144
rect 588544 113092 588596 113144
rect 588544 110440 588596 110492
rect 590568 110440 590620 110492
rect 579436 110236 579488 110288
rect 582012 110236 582064 110288
rect 581828 109692 581880 109744
rect 589372 109692 589424 109744
rect 578332 108332 578384 108384
rect 585140 108332 585192 108384
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 580632 107040 580684 107092
rect 590108 107040 590160 107092
rect 578332 106904 578384 106956
rect 580264 106904 580316 106956
rect 580448 106904 580500 106956
rect 589648 106904 589700 106956
rect 667204 106156 667256 106208
rect 670700 106156 670752 106208
rect 581644 104864 581696 104916
rect 589464 104864 589516 104916
rect 579528 103300 579580 103352
rect 583024 103300 583076 103352
rect 585968 100716 586020 100768
rect 589464 100716 589516 100768
rect 615224 100104 615276 100156
rect 668032 100104 668084 100156
rect 613384 99968 613436 100020
rect 668492 99968 668544 100020
rect 577504 99288 577556 99340
rect 595260 99288 595312 99340
rect 624608 99288 624660 99340
rect 632980 99288 633032 99340
rect 579528 99152 579580 99204
rect 585784 99152 585836 99204
rect 626816 99152 626868 99204
rect 636384 99152 636436 99204
rect 623688 99016 623740 99068
rect 632152 99016 632204 99068
rect 629760 98880 629812 98932
rect 640984 98880 641036 98932
rect 622308 98744 622360 98796
rect 629484 98744 629536 98796
rect 630496 98744 630548 98796
rect 642180 98744 642232 98796
rect 625068 98608 625120 98660
rect 634452 98608 634504 98660
rect 637856 98608 637908 98660
rect 660396 98608 660448 98660
rect 605472 97928 605524 97980
rect 606484 97928 606536 97980
rect 620192 97928 620244 97980
rect 626264 97928 626316 97980
rect 632704 97928 632756 97980
rect 644020 97928 644072 97980
rect 651104 97928 651156 97980
rect 655060 97928 655112 97980
rect 655428 97928 655480 97980
rect 662512 97928 662564 97980
rect 618720 97792 618772 97844
rect 625436 97792 625488 97844
rect 643744 97792 643796 97844
rect 650644 97792 650696 97844
rect 651840 97792 651892 97844
rect 659568 97792 659620 97844
rect 659936 97792 659988 97844
rect 665548 97792 665600 97844
rect 621664 97656 621716 97708
rect 628380 97656 628432 97708
rect 633348 97656 633400 97708
rect 643468 97656 643520 97708
rect 659200 97656 659252 97708
rect 663892 97656 663944 97708
rect 615040 97520 615092 97572
rect 616144 97520 616196 97572
rect 623136 97520 623188 97572
rect 630680 97520 630732 97572
rect 631968 97520 632020 97572
rect 644940 97520 644992 97572
rect 647148 97520 647200 97572
rect 658004 97520 658056 97572
rect 658188 97520 658240 97572
rect 663064 97520 663116 97572
rect 579528 97452 579580 97504
rect 584404 97452 584456 97504
rect 627552 97384 627604 97436
rect 637580 97384 637632 97436
rect 577504 97248 577556 97300
rect 600412 97248 600464 97300
rect 612648 97248 612700 97300
rect 620284 97248 620336 97300
rect 629024 97248 629076 97300
rect 639880 97384 639932 97436
rect 644296 97384 644348 97436
rect 658832 97384 658884 97436
rect 634176 97112 634228 97164
rect 644756 97248 644808 97300
rect 653956 97248 654008 97300
rect 655244 97248 655296 97300
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 643008 97112 643060 97164
rect 634728 96976 634780 97028
rect 643744 96976 643796 97028
rect 598940 96908 598992 96960
rect 599676 96908 599728 96960
rect 612096 96908 612148 96960
rect 612648 96908 612700 96960
rect 617248 96908 617300 96960
rect 618168 96908 618220 96960
rect 626080 96840 626132 96892
rect 635280 96840 635332 96892
rect 606208 96772 606260 96824
rect 612004 96772 612056 96824
rect 615776 96772 615828 96824
rect 618904 96772 618956 96824
rect 650368 97112 650420 97164
rect 658280 97112 658332 97164
rect 645216 97044 645268 97096
rect 649264 97044 649316 97096
rect 658004 96976 658056 97028
rect 661960 96976 662012 97028
rect 646688 96908 646740 96960
rect 647884 96908 647936 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 660120 96772 660172 96824
rect 628196 96704 628248 96756
rect 639052 96704 639104 96756
rect 660672 96704 660724 96756
rect 663248 96704 663300 96756
rect 631232 96568 631284 96620
rect 643192 96568 643244 96620
rect 649632 96568 649684 96620
rect 650828 96568 650880 96620
rect 652576 96568 652628 96620
rect 665364 96568 665416 96620
rect 640064 96432 640116 96484
rect 647700 96432 647752 96484
rect 648160 96432 648212 96484
rect 652024 96432 652076 96484
rect 610624 96296 610676 96348
rect 623044 96296 623096 96348
rect 639328 96296 639380 96348
rect 653864 96432 653916 96484
rect 653312 96296 653364 96348
rect 664168 96296 664220 96348
rect 609152 96160 609204 96212
rect 621664 96160 621716 96212
rect 640800 96160 640852 96212
rect 663708 96160 663760 96212
rect 607680 96024 607732 96076
rect 620744 96024 620796 96076
rect 620928 96024 620980 96076
rect 626448 96024 626500 96076
rect 641536 96024 641588 96076
rect 665180 96024 665232 96076
rect 594064 95888 594116 95940
rect 601884 95888 601936 95940
rect 613568 95888 613620 95940
rect 635464 95888 635516 95940
rect 646044 95888 646096 95940
rect 647700 95888 647752 95940
rect 653404 95888 653456 95940
rect 638592 95752 638644 95804
rect 642824 95752 642876 95804
rect 648896 95752 648948 95804
rect 664628 95888 664680 95940
rect 646228 95616 646280 95668
rect 642824 95480 642876 95532
rect 648528 95480 648580 95532
rect 642640 95208 642692 95260
rect 644480 95208 644532 95260
rect 578700 95004 578752 95056
rect 580632 95004 580684 95056
rect 616512 94596 616564 94648
rect 625804 94596 625856 94648
rect 608416 94460 608468 94512
rect 624424 94460 624476 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 644480 93780 644532 93832
rect 654876 93780 654928 93832
rect 579528 93236 579580 93288
rect 583208 93236 583260 93288
rect 580264 93100 580316 93152
rect 590108 93100 590160 93152
rect 664444 92488 664496 92540
rect 668308 92488 668360 92540
rect 617984 92420 618036 92472
rect 625436 92420 625488 92472
rect 648528 92420 648580 92472
rect 655428 92420 655480 92472
rect 611268 90992 611320 91044
rect 617340 90992 617392 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 620744 89632 620796 89684
rect 626448 89632 626500 89684
rect 645768 88748 645820 88800
rect 657452 88748 657504 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 579528 88272 579580 88324
rect 587164 88272 587216 88324
rect 607220 88272 607272 88324
rect 626448 88272 626500 88324
rect 655060 88272 655112 88324
rect 658464 88272 658516 88324
rect 617340 88136 617392 88188
rect 625620 88136 625672 88188
rect 647884 87116 647936 87168
rect 657176 87116 657228 87168
rect 649264 86980 649316 87032
rect 660672 86980 660724 87032
rect 650828 86844 650880 86896
rect 658832 86844 658884 86896
rect 659568 86844 659620 86896
rect 663248 86844 663300 86896
rect 652024 86708 652076 86760
rect 662512 86708 662564 86760
rect 578608 86572 578660 86624
rect 580448 86572 580500 86624
rect 650644 86572 650696 86624
rect 661408 86572 661460 86624
rect 623044 86436 623096 86488
rect 626448 86436 626500 86488
rect 653404 86300 653456 86352
rect 660120 86300 660172 86352
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 579252 84124 579304 84176
rect 581828 84124 581880 84176
rect 621664 84124 621716 84176
rect 625620 84124 625672 84176
rect 579252 82764 579304 82816
rect 588544 82764 588596 82816
rect 628656 80928 628708 80980
rect 642456 80928 642508 80980
rect 614028 80792 614080 80844
rect 647332 80792 647384 80844
rect 578976 80656 579028 80708
rect 589924 80656 589976 80708
rect 595444 80656 595496 80708
rect 636108 80656 636160 80708
rect 579160 80044 579212 80096
rect 585968 80044 586020 80096
rect 629208 79432 629260 79484
rect 638868 79432 638920 79484
rect 616144 79296 616196 79348
rect 648988 79296 649040 79348
rect 638868 78276 638920 78328
rect 645308 78276 645360 78328
rect 631048 78072 631100 78124
rect 639052 78072 639104 78124
rect 612648 77936 612700 77988
rect 647516 77936 647568 77988
rect 623044 77256 623096 77308
rect 633900 77392 633952 77444
rect 628380 77256 628432 77308
rect 631508 77256 631560 77308
rect 620284 76780 620336 76832
rect 649172 76780 649224 76832
rect 612004 76644 612056 76696
rect 647056 76644 647108 76696
rect 606484 76508 606536 76560
rect 662420 76508 662472 76560
rect 578884 75896 578936 75948
rect 631048 75896 631100 75948
rect 578700 75420 578752 75472
rect 581644 75420 581696 75472
rect 618904 75148 618956 75200
rect 646872 75148 646924 75200
rect 588544 74808 588596 74860
rect 628012 74808 628064 74860
rect 578516 73108 578568 73160
rect 580264 73108 580316 73160
rect 579528 67600 579580 67652
rect 624424 67600 624476 67652
rect 579528 66240 579580 66292
rect 605840 66240 605892 66292
rect 579528 64812 579580 64864
rect 613384 64812 613436 64864
rect 578516 62024 578568 62076
rect 664444 62024 664496 62076
rect 579528 60664 579580 60716
rect 614856 60664 614908 60716
rect 581644 59984 581696 60036
rect 603080 59984 603132 60036
rect 580264 58760 580316 58812
rect 601884 58760 601936 58812
rect 577688 58624 577740 58676
rect 604460 58624 604512 58676
rect 605840 58624 605892 58676
rect 663800 58624 663852 58676
rect 579528 57876 579580 57928
rect 666560 57876 666612 57928
rect 575480 57196 575532 57248
rect 600320 57196 600372 57248
rect 579528 56516 579580 56568
rect 588544 56516 588596 56568
rect 574928 56108 574980 56160
rect 597928 56108 597980 56160
rect 574560 55972 574612 56024
rect 598940 55972 598992 56024
rect 574744 55836 574796 55888
rect 599124 55836 599176 55888
rect 624424 55836 624476 55888
rect 663984 55836 664036 55888
rect 574008 55564 574060 55616
rect 596456 55564 596508 55616
rect 574744 55156 574796 55208
rect 578884 55020 578936 55072
rect 585784 54884 585836 54936
rect 596180 54748 596232 54800
rect 597560 54612 597612 54664
rect 623044 54476 623096 54528
rect 577504 54340 577556 54392
rect 574560 54204 574612 54256
rect 459468 53592 459520 53644
rect 460388 53592 460440 53644
rect 462274 53592 462326 53644
rect 462964 53592 463016 53644
rect 463148 53592 463200 53644
rect 463654 53592 463706 53644
rect 465172 53592 465224 53644
rect 465356 53592 465408 53644
rect 465540 53592 465592 53644
rect 465724 53592 465776 53644
rect 471888 53592 471940 53644
rect 461308 53456 461360 53508
rect 575480 54068 575532 54120
rect 574928 53932 574980 53984
rect 472256 53592 472308 53644
rect 472440 53592 472492 53644
rect 472624 53592 472676 53644
rect 574008 53796 574060 53848
rect 50528 53320 50580 53372
rect 129004 53320 129056 53372
rect 464528 53320 464580 53372
rect 465540 53320 465592 53372
rect 47768 53184 47820 53236
rect 130384 53184 130436 53236
rect 463608 53184 463660 53236
rect 472440 53184 472492 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 46204 53048 46256 53100
rect 130568 53048 130620 53100
rect 464988 53048 465040 53100
rect 465356 53048 465408 53100
rect 463746 52776 463798 52828
rect 472624 52776 472676 52828
rect 145380 52436 145432 52488
rect 306012 52436 306064 52488
rect 50712 51960 50764 52012
rect 130752 51960 130804 52012
rect 48964 51824 49016 51876
rect 129464 51824 129516 51876
rect 49148 51688 49200 51740
rect 126888 51688 126940 51740
rect 126888 50736 126940 50788
rect 129280 50736 129332 50788
rect 50344 50464 50396 50516
rect 128636 50464 128688 50516
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 129004 50328 129056 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 51724 49104 51776 49156
rect 128452 49104 128504 49156
rect 47584 48968 47636 49020
rect 129648 48968 129700 49020
rect 128636 48084 128688 48136
rect 132132 48084 132184 48136
rect 129188 47676 129240 47728
rect 131856 47676 131908 47728
rect 129556 45024 129608 45076
rect 129740 44888 129792 44940
rect 128452 44616 128504 44668
rect 129372 44480 129424 44532
rect 131856 44548 131908 44600
rect 132132 44448 132184 44500
rect 132408 44412 132460 44464
rect 130752 44276 130804 44328
rect 129004 44140 129056 44192
rect 132224 44140 132276 44192
rect 130568 44004 130620 44056
rect 130384 43868 130436 43920
rect 43444 42780 43496 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 307300 42712 307352 42764
rect 369400 42712 369452 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 464344 42712 464396 42764
rect 427084 42576 427136 42628
rect 455880 42576 455932 42628
rect 463976 42576 464028 42628
rect 361764 42440 361816 42492
rect 369400 42440 369452 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 308956 42173 309008 42225
rect 427084 42032 427136 42084
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 455880 41896 455932 41948
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 510344 1007208 510396 1007214
rect 431682 1007176 431738 1007185
rect 510344 1007150 510396 1007156
rect 518164 1007208 518216 1007214
rect 518164 1007150 518216 1007156
rect 431682 1007111 431684 1007120
rect 431736 1007111 431738 1007120
rect 434628 1007140 434680 1007146
rect 431684 1007082 431736 1007088
rect 434628 1007082 434680 1007088
rect 428002 1007040 428058 1007049
rect 428002 1006975 428004 1006984
rect 428056 1006975 428058 1006984
rect 428004 1006946 428056 1006952
rect 359740 1006936 359792 1006942
rect 359738 1006904 359740 1006913
rect 374644 1006936 374696 1006942
rect 359792 1006904 359794 1006913
rect 374644 1006878 374696 1006884
rect 428370 1006904 428426 1006913
rect 359738 1006839 359794 1006848
rect 145564 1006800 145616 1006806
rect 145564 1006742 145616 1006748
rect 151728 1006800 151780 1006806
rect 359372 1006800 359424 1006806
rect 151728 1006742 151780 1006748
rect 359370 1006768 359372 1006777
rect 369124 1006800 369176 1006806
rect 359424 1006768 359426 1006777
rect 144184 1006528 144236 1006534
rect 101126 1006496 101182 1006505
rect 94688 1006460 94740 1006466
rect 144184 1006470 144236 1006476
rect 101126 1006431 101128 1006440
rect 94688 1006402 94740 1006408
rect 101180 1006431 101182 1006440
rect 101128 1006402 101180 1006408
rect 93308 1006188 93360 1006194
rect 93308 1006130 93360 1006136
rect 93124 1006052 93176 1006058
rect 93124 1005994 93176 1006000
rect 92756 999796 92808 999802
rect 92756 999738 92808 999744
rect 92388 998436 92440 998442
rect 92388 998378 92440 998384
rect 80426 995752 80482 995761
rect 80178 995710 80426 995738
rect 85946 995752 86002 995761
rect 85698 995710 85946 995738
rect 80426 995687 80482 995696
rect 86590 995752 86646 995761
rect 86342 995710 86590 995738
rect 85946 995687 86002 995696
rect 87878 995752 87934 995761
rect 87538 995710 87878 995738
rect 86590 995687 86646 995696
rect 92400 995738 92428 998378
rect 92572 998096 92624 998102
rect 92572 998038 92624 998044
rect 87878 995687 87934 995696
rect 92032 995710 92428 995738
rect 88982 995480 89038 995489
rect 77036 995081 77064 995452
rect 77022 995072 77078 995081
rect 77022 995007 77078 995016
rect 77680 994566 77708 995452
rect 78324 994838 78352 995452
rect 78312 994832 78364 994838
rect 78312 994774 78364 994780
rect 77668 994560 77720 994566
rect 77668 994502 77720 994508
rect 80716 994430 80744 995452
rect 81360 994702 81388 995452
rect 82004 994809 82032 995452
rect 81990 994800 82046 994809
rect 81990 994735 82046 994744
rect 81348 994696 81400 994702
rect 81348 994638 81400 994644
rect 80704 994424 80756 994430
rect 80704 994366 80756 994372
rect 84488 994265 84516 995452
rect 85054 995438 85344 995466
rect 88734 995438 88982 995466
rect 85316 994537 85344 995438
rect 90270 995480 90326 995489
rect 89378 995438 89852 995466
rect 90022 995438 90270 995466
rect 88982 995415 89038 995424
rect 89824 995194 89852 995438
rect 91218 995438 91692 995466
rect 90270 995415 90326 995424
rect 91664 995330 91692 995438
rect 92032 995330 92060 995710
rect 92204 995580 92256 995586
rect 92204 995522 92256 995528
rect 91664 995302 92060 995330
rect 92216 995194 92244 995522
rect 92584 995489 92612 998038
rect 92768 995586 92796 999738
rect 92938 996976 92994 996985
rect 92938 996911 92994 996920
rect 92952 996402 92980 996911
rect 92940 996396 92992 996402
rect 92940 996338 92992 996344
rect 92756 995580 92808 995586
rect 92756 995522 92808 995528
rect 92570 995480 92626 995489
rect 92570 995415 92626 995424
rect 89824 995166 92244 995194
rect 85302 994528 85358 994537
rect 85302 994463 85358 994472
rect 93136 994430 93164 1005994
rect 93320 996033 93348 1006130
rect 94504 1002652 94556 1002658
rect 94504 1002594 94556 1002600
rect 93492 997756 93544 997762
rect 93492 997698 93544 997704
rect 93504 997257 93532 997698
rect 93490 997248 93546 997257
rect 93490 997183 93546 997192
rect 94516 996985 94544 1002594
rect 93582 996976 93638 996985
rect 93582 996911 93638 996920
rect 94502 996976 94558 996985
rect 94502 996911 94558 996920
rect 93306 996024 93362 996033
rect 93306 995959 93362 995968
rect 93596 994537 93624 996911
rect 94700 996033 94728 1006402
rect 101954 1006360 102010 1006369
rect 96068 1006324 96120 1006330
rect 101954 1006295 101956 1006304
rect 96068 1006266 96120 1006272
rect 102008 1006295 102010 1006304
rect 108486 1006360 108542 1006369
rect 108486 1006295 108488 1006304
rect 101956 1006266 102008 1006272
rect 108540 1006295 108542 1006304
rect 126244 1006324 126296 1006330
rect 108488 1006266 108540 1006272
rect 126244 1006266 126296 1006272
rect 96080 1006058 96108 1006266
rect 99470 1006224 99526 1006233
rect 104806 1006224 104862 1006233
rect 99470 1006159 99472 1006168
rect 99524 1006159 99526 1006168
rect 102968 1006188 103020 1006194
rect 99472 1006130 99524 1006136
rect 104806 1006159 104808 1006168
rect 102968 1006130 103020 1006136
rect 104860 1006159 104862 1006168
rect 106830 1006224 106886 1006233
rect 106830 1006159 106832 1006168
rect 104808 1006130 104860 1006136
rect 106884 1006159 106886 1006168
rect 113824 1006188 113876 1006194
rect 106832 1006130 106884 1006136
rect 113824 1006130 113876 1006136
rect 98274 1006088 98330 1006097
rect 96068 1006052 96120 1006058
rect 96068 1005994 96120 1006000
rect 96252 1006052 96304 1006058
rect 98274 1006023 98276 1006032
rect 96252 1005994 96304 1006000
rect 98328 1006023 98330 1006032
rect 101404 1006052 101456 1006058
rect 98276 1005994 98328 1006000
rect 101404 1005994 101456 1006000
rect 96068 1002108 96120 1002114
rect 96068 1002050 96120 1002056
rect 95884 1001972 95936 1001978
rect 95884 1001914 95936 1001920
rect 94686 996024 94742 996033
rect 94686 995959 94742 995968
rect 93582 994528 93638 994537
rect 93582 994463 93638 994472
rect 93124 994424 93176 994430
rect 93124 994366 93176 994372
rect 84474 994256 84530 994265
rect 84474 994191 84530 994200
rect 50344 993200 50396 993206
rect 50344 993142 50396 993148
rect 44824 993064 44876 993070
rect 44824 993006 44876 993012
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 969218 42196 969272
rect 42260 969258 42564 969286
rect 42260 969218 42288 969258
rect 42168 969190 42288 969218
rect 42536 968810 42564 969258
rect 42536 968782 42840 968810
rect 42168 967609 42196 968048
rect 42154 967600 42210 967609
rect 42154 967535 42210 967544
rect 42614 967600 42670 967609
rect 42614 967535 42670 967544
rect 41800 967201 41828 967405
rect 41786 967192 41842 967201
rect 41786 967127 41842 967136
rect 42154 967192 42210 967201
rect 42154 967127 42210 967136
rect 42168 966756 42196 967127
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42444 963937 42472 964362
rect 42430 963928 42486 963937
rect 42430 963863 42486 963872
rect 42182 963711 42472 963739
rect 42444 963393 42472 963711
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42430 963112 42486 963121
rect 42182 963070 42430 963098
rect 42430 963047 42486 963056
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 41786 959103 41842 959112
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 41800 957817 41828 958188
rect 41786 957808 41842 957817
rect 41786 957743 41842 957752
rect 42182 956338 42288 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 41800 954689 41828 955060
rect 41786 954680 41842 954689
rect 41786 954615 41842 954624
rect 41786 954408 41842 954417
rect 41786 954343 41842 954352
rect 35162 952912 35218 952921
rect 35162 952847 35218 952856
rect 33784 951516 33836 951522
rect 33784 951458 33836 951464
rect 31758 946656 31814 946665
rect 31758 946591 31814 946600
rect 31772 945334 31800 946591
rect 28724 945328 28776 945334
rect 28724 945270 28776 945276
rect 31760 945328 31812 945334
rect 31760 945270 31812 945276
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28736 942721 28764 945270
rect 28722 942712 28778 942721
rect 28722 942647 28778 942656
rect 33796 938233 33824 951458
rect 33782 938224 33838 938233
rect 33782 938159 33838 938168
rect 35176 937825 35204 952847
rect 41800 952626 41828 954343
rect 41524 952598 41828 952626
rect 37922 952504 37978 952513
rect 37922 952439 37978 952448
rect 36544 952400 36596 952406
rect 36544 952342 36596 952348
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35820 942614 35848 943055
rect 35808 942608 35860 942614
rect 35808 942550 35860 942556
rect 35806 941896 35862 941905
rect 35806 941831 35862 941840
rect 35820 941254 35848 941831
rect 35808 941248 35860 941254
rect 35808 941190 35860 941196
rect 35806 940264 35862 940273
rect 35806 940199 35862 940208
rect 35820 939826 35848 940199
rect 35808 939820 35860 939826
rect 35808 939762 35860 939768
rect 36556 939049 36584 952342
rect 36542 939040 36598 939049
rect 36542 938975 36598 938984
rect 37936 938641 37964 952439
rect 39302 952232 39358 952241
rect 39302 952167 39358 952176
rect 37922 938632 37978 938641
rect 37922 938567 37978 938576
rect 35162 937816 35218 937825
rect 35162 937751 35218 937760
rect 39316 937417 39344 952167
rect 40038 951688 40094 951697
rect 40038 951623 40094 951632
rect 39762 943800 39818 943809
rect 39762 943735 39818 943744
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 39776 935785 39804 943735
rect 39762 935776 39818 935785
rect 39762 935711 39818 935720
rect 40052 934561 40080 951623
rect 41524 951522 41552 952598
rect 42260 952490 42288 956338
rect 41708 952462 42288 952490
rect 41708 952406 41736 952462
rect 41696 952400 41748 952406
rect 41696 952342 41748 952348
rect 41512 951516 41564 951522
rect 41512 951458 41564 951464
rect 42628 949454 42656 967535
rect 42536 949426 42656 949454
rect 41604 942608 41656 942614
rect 41656 942556 41828 942562
rect 41604 942550 41828 942556
rect 41616 942534 41828 942550
rect 41420 941248 41472 941254
rect 41420 941190 41472 941196
rect 40038 934552 40094 934561
rect 40038 934487 40094 934496
rect 41432 911713 41460 941190
rect 41604 939820 41656 939826
rect 41604 939762 41656 939768
rect 41616 911985 41644 939762
rect 41800 935649 41828 942534
rect 42062 940672 42118 940681
rect 42062 940607 42118 940616
rect 42076 939865 42104 940607
rect 42062 939856 42118 939865
rect 42062 939791 42118 939800
rect 42536 939794 42564 949426
rect 42352 939766 42564 939794
rect 41786 935640 41842 935649
rect 41786 935575 41842 935584
rect 42352 932929 42380 939766
rect 42812 937009 42840 968782
rect 43456 967201 43484 975666
rect 43442 967192 43498 967201
rect 43442 967127 43498 967136
rect 43442 964744 43498 964753
rect 43442 964679 43498 964688
rect 43258 963928 43314 963937
rect 43258 963863 43314 963872
rect 43074 963384 43130 963393
rect 43074 963319 43130 963328
rect 42798 937000 42854 937009
rect 42798 936935 42854 936944
rect 43088 934969 43116 963319
rect 43074 934960 43130 934969
rect 43074 934895 43130 934904
rect 43272 933745 43300 963863
rect 43456 935377 43484 964679
rect 44270 963112 44326 963121
rect 44270 963047 44326 963056
rect 43442 935368 43498 935377
rect 43442 935303 43498 935312
rect 44284 934153 44312 963047
rect 44454 958760 44510 958769
rect 44454 958695 44510 958704
rect 44468 936329 44496 958695
rect 44836 941497 44864 993006
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 46204 961920 46256 961926
rect 46204 961862 46256 961868
rect 46216 946665 46244 961862
rect 46202 946656 46258 946665
rect 46202 946591 46258 946600
rect 45560 946008 45612 946014
rect 45560 945950 45612 945956
rect 45572 943537 45600 945950
rect 45558 943528 45614 943537
rect 45558 943463 45614 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44638 941080 44694 941089
rect 44638 941015 44694 941024
rect 44454 936320 44510 936329
rect 44454 936255 44510 936264
rect 44270 934144 44326 934153
rect 44270 934079 44326 934088
rect 43258 933736 43314 933745
rect 43258 933671 43314 933680
rect 43626 933328 43682 933337
rect 43626 933263 43682 933272
rect 42338 932920 42394 932929
rect 42338 932855 42394 932864
rect 41602 911976 41658 911985
rect 41602 911911 41658 911920
rect 41418 911704 41474 911713
rect 41418 911639 41474 911648
rect 42936 892528 42992 892537
rect 42936 892463 42992 892472
rect 42950 892328 42978 892463
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43074 892256 43130 892265
rect 43074 892191 43130 892200
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817086 35848 817255
rect 35808 817080 35860 817086
rect 35808 817022 35860 817028
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 815658 35848 816439
rect 41432 815658 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815810 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815782 41644 815810
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 41420 815652 41472 815658
rect 41420 815594 41472 815600
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814298 35848 814807
rect 41616 814298 41644 815782
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41604 814292 41656 814298
rect 41604 814234 41656 814240
rect 41326 812832 41382 812841
rect 41326 812767 41382 812776
rect 40958 812424 41014 812433
rect 40958 812359 41014 812368
rect 35162 811608 35218 811617
rect 35162 811543 35218 811552
rect 35176 802466 35204 811543
rect 35898 811200 35954 811209
rect 35898 811135 35954 811144
rect 35164 802460 35216 802466
rect 35164 802402 35216 802408
rect 35912 802330 35940 811135
rect 40592 808580 40644 808586
rect 40592 808522 40644 808528
rect 40604 805361 40632 808522
rect 40774 808344 40830 808353
rect 40774 808279 40830 808288
rect 40590 805352 40646 805361
rect 40590 805287 40646 805296
rect 40788 805089 40816 808279
rect 40774 805080 40830 805089
rect 40774 805015 40830 805024
rect 40972 804545 41000 812359
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 41156 804817 41184 811951
rect 41340 811510 41368 812767
rect 41328 811504 41380 811510
rect 41328 811446 41380 811452
rect 41696 811504 41748 811510
rect 41748 811452 42380 811458
rect 41696 811446 42380 811452
rect 41708 811430 42380 811446
rect 41970 809160 42026 809169
rect 41970 809095 42026 809104
rect 41786 808752 41842 808761
rect 41616 808710 41786 808738
rect 41616 808586 41644 808710
rect 41786 808687 41842 808696
rect 41604 808580 41656 808586
rect 41604 808522 41656 808528
rect 41984 805497 42012 809095
rect 42154 806712 42210 806721
rect 42154 806647 42210 806656
rect 41970 805488 42026 805497
rect 41970 805423 42026 805432
rect 41142 804808 41198 804817
rect 41142 804743 41198 804752
rect 40958 804536 41014 804545
rect 40958 804471 41014 804480
rect 41694 802496 41750 802505
rect 41694 802431 41696 802440
rect 41748 802431 41750 802440
rect 41696 802402 41748 802408
rect 35900 802324 35952 802330
rect 35900 802266 35952 802272
rect 41696 802324 41748 802330
rect 41696 802266 41748 802272
rect 41708 802210 41736 802266
rect 41708 802182 41828 802210
rect 41800 800329 41828 802182
rect 41786 800320 41842 800329
rect 42168 800306 42196 806647
rect 42168 800278 42288 800306
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798266 42288 800278
rect 42182 798238 42288 798266
rect 42352 797619 42380 811430
rect 43074 810792 43130 810801
rect 43074 810727 43130 810736
rect 42798 809976 42854 809985
rect 42798 809911 42854 809920
rect 42522 802496 42578 802505
rect 42578 802454 42748 802482
rect 42522 802431 42578 802440
rect 42522 799232 42578 799241
rect 42522 799167 42578 799176
rect 42182 797591 42380 797619
rect 42536 797042 42564 799167
rect 42720 799082 42748 802454
rect 42352 797014 42564 797042
rect 42628 799054 42748 799082
rect 42352 796974 42380 797014
rect 42182 796946 42380 796974
rect 42430 796784 42486 796793
rect 42430 796719 42486 796728
rect 42154 796240 42210 796249
rect 42154 796175 42210 796184
rect 42168 795765 42196 796175
rect 42444 794594 42472 796719
rect 42182 794566 42472 794594
rect 42430 794336 42486 794345
rect 42430 794271 42486 794280
rect 41786 794200 41842 794209
rect 41786 794135 41842 794144
rect 41800 793900 41828 794135
rect 42444 793302 42472 794271
rect 42182 793274 42472 793302
rect 42628 792758 42656 799054
rect 42182 792730 42656 792758
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42812 792282 42840 809911
rect 42168 790622 42288 790650
rect 42628 792254 42840 792282
rect 42168 790228 42196 790622
rect 42628 789834 42656 792254
rect 42890 790800 42946 790809
rect 42890 790735 42946 790744
rect 42904 790650 42932 790735
rect 42260 789806 42656 789834
rect 42720 790622 42932 790650
rect 42260 789630 42288 789806
rect 42182 789602 42288 789630
rect 42720 789018 42748 790622
rect 42168 788990 42288 789018
rect 42168 788936 42196 788990
rect 42260 788950 42288 788990
rect 42536 788990 42748 789018
rect 42536 788950 42564 788990
rect 42260 788922 42564 788950
rect 42522 788760 42578 788769
rect 42522 788695 42578 788704
rect 41786 788624 41842 788633
rect 41786 788559 41842 788568
rect 41800 788392 41828 788559
rect 42536 788474 42564 788695
rect 42706 788624 42762 788633
rect 42706 788559 42762 788568
rect 42536 788446 42656 788474
rect 42430 788352 42486 788361
rect 42430 788287 42486 788296
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42260 786978 42288 788151
rect 42168 786950 42288 786978
rect 42168 786556 42196 786950
rect 42444 785958 42472 788287
rect 42628 788202 42656 788446
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42536 788174 42656 788202
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 788174
rect 42182 785250 42564 785278
rect 42720 779714 42748 788559
rect 43088 788361 43116 810727
rect 43442 809568 43498 809577
rect 43442 809503 43498 809512
rect 43258 807528 43314 807537
rect 43258 807463 43314 807472
rect 43074 788352 43130 788361
rect 43074 788287 43130 788296
rect 41708 779686 42748 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 772886 35848 773463
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768874 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35532 768984
rect 35584 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 40040 769004 40092 769010
rect 35532 768946 35584 768952
rect 35348 768868 35400 768874
rect 35348 768810 35400 768816
rect 35820 768738 35848 768975
rect 40040 768946 40092 768952
rect 35808 768732 35860 768738
rect 35808 768674 35860 768680
rect 31022 768224 31078 768233
rect 31022 768159 31078 768168
rect 31036 759694 31064 768159
rect 35530 767816 35586 767825
rect 35530 767751 35586 767760
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35544 767378 35572 767751
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35532 767372 35584 767378
rect 35532 767314 35584 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 31024 759688 31076 759694
rect 31024 759630 31076 759636
rect 35176 758334 35204 766935
rect 35164 758328 35216 758334
rect 35164 758270 35216 758276
rect 36556 757761 36584 767450
rect 37924 767372 37976 767378
rect 37924 767314 37976 767320
rect 37094 763328 37150 763337
rect 37094 763263 37096 763272
rect 37148 763263 37150 763272
rect 37096 763234 37148 763240
rect 37936 759082 37964 767314
rect 40052 764561 40080 768946
rect 41696 768868 41748 768874
rect 41696 768810 41748 768816
rect 41328 768732 41380 768738
rect 41328 768674 41380 768680
rect 41340 765785 41368 768674
rect 41326 765776 41382 765785
rect 41326 765711 41382 765720
rect 40038 764552 40094 764561
rect 40038 764487 40094 764496
rect 39304 763292 39356 763298
rect 39304 763234 39356 763240
rect 39120 759688 39172 759694
rect 39120 759630 39172 759636
rect 37924 759076 37976 759082
rect 37924 759018 37976 759024
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 39132 757353 39160 759630
rect 39316 758033 39344 763234
rect 41512 759076 41564 759082
rect 41512 759018 41564 759024
rect 39302 758024 39358 758033
rect 39302 757959 39358 757968
rect 41524 757602 41552 759018
rect 41708 758849 41736 768810
rect 42890 766320 42946 766329
rect 42890 766255 42946 766264
rect 42706 765776 42762 765785
rect 42706 765711 42762 765720
rect 41694 758840 41750 758849
rect 41694 758775 41750 758784
rect 42246 758840 42302 758849
rect 42246 758775 42302 758784
rect 41696 758328 41748 758334
rect 41694 758296 41696 758305
rect 41748 758296 41750 758305
rect 41694 758231 41750 758240
rect 42260 758146 42288 758775
rect 42430 758296 42486 758305
rect 42486 758254 42656 758282
rect 42430 758231 42486 758240
rect 42260 758118 42472 758146
rect 42246 758024 42302 758033
rect 42246 757959 42302 757968
rect 41524 757574 41828 757602
rect 39118 757344 39174 757353
rect 39118 757279 39174 757288
rect 41800 757081 41828 757574
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 41878 756664 41934 756673
rect 41878 756599 41934 756608
rect 41892 756226 41920 756599
rect 42168 755018 42196 755072
rect 42260 755018 42288 757959
rect 42168 754990 42288 755018
rect 42444 754882 42472 758118
rect 42260 754854 42472 754882
rect 42260 754406 42288 754854
rect 42430 754488 42486 754497
rect 42430 754423 42486 754432
rect 42182 754378 42288 754406
rect 41970 754080 42026 754089
rect 41970 754015 42026 754024
rect 41984 753780 42012 754015
rect 42246 753944 42302 753953
rect 42246 753879 42302 753888
rect 42260 752570 42288 753879
rect 42182 752542 42288 752570
rect 42246 752176 42302 752185
rect 42246 752111 42302 752120
rect 42062 751768 42118 751777
rect 42062 751703 42118 751712
rect 42076 751369 42104 751703
rect 41786 751088 41842 751097
rect 41786 751023 41842 751032
rect 41800 750720 41828 751023
rect 42168 749986 42196 750108
rect 42260 749986 42288 752111
rect 42168 749958 42288 749986
rect 42168 749550 42380 749578
rect 42168 749529 42196 749550
rect 42352 749543 42380 749550
rect 42444 749543 42472 754423
rect 42352 749515 42472 749543
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 747062 42288 749391
rect 42430 749320 42486 749329
rect 42430 749255 42486 749264
rect 42182 747034 42288 747062
rect 42444 746594 42472 749255
rect 42076 746566 42472 746594
rect 42076 746401 42104 746566
rect 42628 745770 42656 758254
rect 42720 754338 42748 765711
rect 42720 754310 42840 754338
rect 42812 754066 42840 754310
rect 42182 745742 42656 745770
rect 42720 754038 42840 754066
rect 42720 745226 42748 754038
rect 42904 753953 42932 766255
rect 43074 763056 43130 763065
rect 43074 762991 43130 763000
rect 42890 753944 42946 753953
rect 42890 753879 42946 753888
rect 42890 753536 42946 753545
rect 42890 753471 42946 753480
rect 42904 751777 42932 753471
rect 42890 751768 42946 751777
rect 42890 751703 42946 751712
rect 42182 745198 42748 745226
rect 42430 745104 42486 745113
rect 42430 745039 42486 745048
rect 42246 744832 42302 744841
rect 42246 744767 42302 744776
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42260 743050 42288 744767
rect 42168 743022 42288 743050
rect 42168 742696 42196 743022
rect 42444 742098 42472 745039
rect 42706 743064 42762 743073
rect 42706 742999 42762 743008
rect 42182 742070 42472 742098
rect 42720 736934 42748 742999
rect 41708 736906 42748 736934
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35820 730114 35848 730895
rect 41708 730114 41736 736906
rect 35808 730108 35860 730114
rect 35808 730050 35860 730056
rect 41696 730108 41748 730114
rect 41696 730050 41748 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41142 726064 41198 726073
rect 41142 725999 41198 726008
rect 33782 725248 33838 725257
rect 33782 725183 33838 725192
rect 33046 724024 33102 724033
rect 33046 723959 33102 723968
rect 31666 723208 31722 723217
rect 31666 723143 31722 723152
rect 31680 715562 31708 723143
rect 33060 715698 33088 723959
rect 33796 715834 33824 725183
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 33784 715828 33836 715834
rect 33784 715770 33836 715776
rect 33048 715692 33100 715698
rect 33048 715634 33100 715640
rect 31668 715556 31720 715562
rect 31668 715498 31720 715504
rect 36556 714882 36584 724775
rect 40682 724432 40738 724441
rect 40682 724367 40738 724376
rect 36544 714876 36596 714882
rect 36544 714818 36596 714824
rect 40696 714785 40724 724367
rect 41156 721777 41184 725999
rect 41340 725966 41368 726407
rect 41328 725960 41380 725966
rect 41328 725902 41380 725908
rect 41696 725960 41748 725966
rect 41748 725908 41920 725914
rect 41696 725902 41920 725908
rect 41708 725886 41920 725902
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724538 41368 725591
rect 41328 724532 41380 724538
rect 41328 724474 41380 724480
rect 41696 724532 41748 724538
rect 41892 724514 41920 725886
rect 41892 724486 42380 724514
rect 41696 724474 41748 724480
rect 41142 721768 41198 721777
rect 41142 721703 41198 721712
rect 41708 719681 41736 724474
rect 41878 722392 41934 722401
rect 41878 722327 41934 722336
rect 41694 719672 41750 719681
rect 41694 719607 41750 719616
rect 41892 718593 41920 722327
rect 42154 720352 42210 720361
rect 42154 720287 42210 720296
rect 42168 720202 42196 720287
rect 42168 720174 42288 720202
rect 41878 718584 41934 718593
rect 41878 718519 41934 718528
rect 41142 715864 41198 715873
rect 41142 715799 41198 715808
rect 41694 715864 41750 715873
rect 41694 715799 41696 715808
rect 41156 715698 41184 715799
rect 41748 715799 41750 715808
rect 41696 715770 41748 715776
rect 41144 715692 41196 715698
rect 41144 715634 41196 715640
rect 41696 715556 41748 715562
rect 41748 715516 41920 715544
rect 41696 715498 41748 715504
rect 41696 714876 41748 714882
rect 41892 714854 41920 715516
rect 41892 714826 42012 714854
rect 41696 714818 41748 714824
rect 40682 714776 40738 714785
rect 41708 714762 41736 714818
rect 41708 714734 41828 714762
rect 40682 714711 40738 714720
rect 41800 714490 41828 714734
rect 41984 714649 42012 714826
rect 41970 714640 42026 714649
rect 42260 714626 42288 720174
rect 42352 719522 42380 724486
rect 42522 719672 42578 719681
rect 42522 719607 42578 719616
rect 42352 719494 42472 719522
rect 42260 714598 42380 714626
rect 41970 714575 42026 714584
rect 41800 714462 42288 714490
rect 42260 713062 42288 714462
rect 42182 713034 42288 713062
rect 42352 712314 42380 714598
rect 42168 712286 42380 712314
rect 42168 711824 42196 712286
rect 42444 711498 42472 719494
rect 42536 715714 42564 719607
rect 42706 715864 42762 715873
rect 42706 715799 42762 715808
rect 42536 715686 42656 715714
rect 42260 711470 42472 711498
rect 42260 711226 42288 711470
rect 42182 711198 42288 711226
rect 42246 711104 42302 711113
rect 42246 711039 42302 711048
rect 42260 710575 42288 711039
rect 42182 710547 42288 710575
rect 41970 709880 42026 709889
rect 41970 709815 42026 709824
rect 41984 709376 42012 709815
rect 42246 709200 42302 709209
rect 42246 709135 42302 709144
rect 41786 708520 41842 708529
rect 41786 708455 41842 708464
rect 41800 708152 41828 708455
rect 42260 707554 42288 709135
rect 42182 707526 42288 707554
rect 42628 707282 42656 715686
rect 42536 707254 42656 707282
rect 41800 706761 41828 706860
rect 41786 706752 41842 706761
rect 41786 706687 41842 706696
rect 42154 706752 42210 706761
rect 42154 706687 42210 706696
rect 42168 706316 42196 706687
rect 42246 705528 42302 705537
rect 42246 705463 42302 705472
rect 41786 704304 41842 704313
rect 41786 704239 41842 704248
rect 41800 703868 41828 704239
rect 42260 703338 42288 705463
rect 42168 703310 42288 703338
rect 42168 703188 42196 703310
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 42536 702046 42564 707254
rect 42720 706761 42748 715799
rect 42890 715592 42946 715601
rect 42890 715527 42946 715536
rect 42706 706752 42762 706761
rect 42706 706687 42762 706696
rect 42904 705194 42932 715527
rect 42720 705166 42932 705194
rect 42720 703089 42748 705166
rect 42706 703080 42762 703089
rect 42706 703015 42762 703024
rect 42168 701978 42196 702032
rect 42352 702018 42564 702046
rect 42352 701978 42380 702018
rect 42168 701950 42380 701978
rect 42338 701856 42394 701865
rect 42338 701791 42394 701800
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42352 699530 42380 701791
rect 42614 701584 42670 701593
rect 42614 701519 42670 701528
rect 42182 699502 42380 699530
rect 42628 698918 42656 701519
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 41694 697912 41750 697921
rect 41694 697847 41750 697856
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 41326 687712 41382 687721
rect 41326 687647 41382 687656
rect 35622 687304 35678 687313
rect 41340 687274 41368 687647
rect 41708 687274 41736 697847
rect 35622 687239 35678 687248
rect 41328 687268 41380 687274
rect 41328 687210 41380 687216
rect 41696 687268 41748 687274
rect 41696 687210 41748 687216
rect 41326 683224 41382 683233
rect 41326 683159 41328 683168
rect 41380 683159 41382 683168
rect 41696 683188 41748 683194
rect 41328 683130 41380 683136
rect 41696 683130 41748 683136
rect 41326 682408 41382 682417
rect 41326 682343 41382 682352
rect 40038 682000 40094 682009
rect 40038 681935 40094 681944
rect 36726 681592 36782 681601
rect 36726 681527 36782 681536
rect 36542 681184 36598 681193
rect 36542 681119 36598 681128
rect 35162 680776 35218 680785
rect 35162 680711 35218 680720
rect 35176 672790 35204 680711
rect 35164 672784 35216 672790
rect 35164 672726 35216 672732
rect 36556 670993 36584 681119
rect 36740 672110 36768 681527
rect 40052 678026 40080 681935
rect 41340 681902 41368 682343
rect 41708 681986 41736 683130
rect 41708 681958 42012 681986
rect 41328 681896 41380 681902
rect 41696 681896 41748 681902
rect 41328 681838 41380 681844
rect 41694 681864 41696 681873
rect 41748 681864 41750 681873
rect 41694 681799 41750 681808
rect 41984 678974 42012 681958
rect 42614 681864 42670 681873
rect 42614 681799 42670 681808
rect 42628 678974 42656 681799
rect 42798 679960 42854 679969
rect 42798 679895 42854 679904
rect 42812 678974 42840 679895
rect 41984 678946 42380 678974
rect 42628 678946 42748 678974
rect 42812 678946 43024 678974
rect 40040 678020 40092 678026
rect 40040 677962 40092 677968
rect 41696 678020 41748 678026
rect 41696 677962 41748 677968
rect 41708 677385 41736 677962
rect 41694 677376 41750 677385
rect 41694 677311 41750 677320
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 36728 672104 36780 672110
rect 36728 672046 36780 672052
rect 39960 671770 39988 677039
rect 40132 672784 40184 672790
rect 40132 672726 40184 672732
rect 39948 671764 40000 671770
rect 39948 671706 40000 671712
rect 40144 671265 40172 672726
rect 41512 672104 41564 672110
rect 41512 672046 41564 672052
rect 41524 671514 41552 672046
rect 42352 671786 42380 678946
rect 42720 677498 42748 678946
rect 42536 677470 42748 677498
rect 41696 671764 41748 671770
rect 42352 671758 42472 671786
rect 41696 671706 41748 671712
rect 41708 671650 41736 671706
rect 41708 671622 42380 671650
rect 41524 671486 42288 671514
rect 40130 671256 40186 671265
rect 40130 671191 40186 671200
rect 36542 670984 36598 670993
rect 36542 670919 36598 670928
rect 42168 669746 42196 669868
rect 42260 669746 42288 671486
rect 42168 669718 42288 669746
rect 42352 668658 42380 671622
rect 42182 668630 42380 668658
rect 42444 668114 42472 671758
rect 42352 668086 42472 668114
rect 42352 668046 42380 668086
rect 42168 667978 42196 668032
rect 42260 668018 42380 668046
rect 42260 667978 42288 668018
rect 42536 667978 42564 677470
rect 42706 677376 42762 677385
rect 42706 677311 42762 677320
rect 42720 676214 42748 677311
rect 42996 676214 43024 678946
rect 42720 676186 42840 676214
rect 42168 667950 42288 667978
rect 42444 667950 42564 667978
rect 42246 667856 42302 667865
rect 42246 667791 42302 667800
rect 42260 667366 42288 667791
rect 42444 667706 42472 667950
rect 42812 667706 42840 676186
rect 42444 667678 42656 667706
rect 42430 667584 42486 667593
rect 42430 667519 42486 667528
rect 42182 667338 42288 667366
rect 42246 667176 42302 667185
rect 42246 667111 42302 667120
rect 42260 666554 42288 667111
rect 42168 666526 42288 666554
rect 42168 666165 42196 666526
rect 42246 666088 42302 666097
rect 42246 666023 42302 666032
rect 41786 665408 41842 665417
rect 41786 665343 41842 665352
rect 41800 664972 41828 665343
rect 42260 664339 42288 666023
rect 42182 664311 42288 664339
rect 41970 664048 42026 664057
rect 41970 663983 42026 663992
rect 41984 663680 42012 663983
rect 42154 663504 42210 663513
rect 42154 663439 42210 663448
rect 42168 663136 42196 663439
rect 42246 662960 42302 662969
rect 42444 662946 42472 667519
rect 42628 666554 42656 667678
rect 42720 667678 42840 667706
rect 42904 676186 43024 676214
rect 42720 667026 42748 667678
rect 42904 667185 42932 676186
rect 42890 667176 42946 667185
rect 42890 667111 42946 667120
rect 42720 666998 42932 667026
rect 42628 666526 42840 666554
rect 42812 663626 42840 666526
rect 42720 663598 42840 663626
rect 42444 662918 42564 662946
rect 42246 662895 42302 662904
rect 42260 662810 42288 662895
rect 42260 662782 42472 662810
rect 42246 662688 42302 662697
rect 42246 662623 42302 662632
rect 42260 661042 42288 662623
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42444 660022 42472 662782
rect 42182 659994 42472 660022
rect 42536 659371 42564 662918
rect 42182 659343 42564 659371
rect 42720 659002 42748 663598
rect 42904 663513 42932 666998
rect 42890 663504 42946 663513
rect 42890 663439 42946 663448
rect 42536 658974 42748 659002
rect 42168 658838 42288 658866
rect 42168 658784 42196 658838
rect 42260 658798 42288 658838
rect 42536 658798 42564 658974
rect 42260 658770 42564 658798
rect 42614 658608 42670 658617
rect 42614 658543 42670 658552
rect 42430 658336 42486 658345
rect 42430 658271 42486 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42444 656350 42472 658271
rect 42182 656322 42472 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42628 655670 42656 658543
rect 42260 655642 42656 655670
rect 35806 646776 35862 646785
rect 35806 646711 35862 646720
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35820 644745 35848 646711
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35622 639840 35678 639849
rect 35622 639775 35678 639784
rect 35636 638994 35664 639775
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35820 639130 35848 639367
rect 35808 639124 35860 639130
rect 35808 639066 35860 639072
rect 40040 639124 40092 639130
rect 40040 639066 40092 639072
rect 35624 638988 35676 638994
rect 35624 638930 35676 638936
rect 40052 638625 40080 639066
rect 41512 638988 41564 638994
rect 41512 638930 41564 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 40038 638616 40094 638625
rect 40038 638551 40094 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 35820 637634 35848 638551
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 40040 637628 40092 637634
rect 40040 637570 40092 637576
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35820 636274 35848 636511
rect 35808 636268 35860 636274
rect 35808 636210 35860 636216
rect 40052 635934 40080 637570
rect 40040 635928 40092 635934
rect 40040 635870 40092 635876
rect 41524 634814 41552 638930
rect 41786 638208 41842 638217
rect 41786 638143 41842 638152
rect 41800 637605 41828 638143
rect 41786 637596 41842 637605
rect 41786 637531 41842 637540
rect 41696 636268 41748 636274
rect 41696 636210 41748 636216
rect 41708 636018 41736 636210
rect 41708 635990 42656 636018
rect 41696 635928 41748 635934
rect 41748 635876 42564 635882
rect 41696 635870 42564 635876
rect 41708 635854 42564 635870
rect 41524 634786 42472 634814
rect 42246 633856 42302 633865
rect 42246 633791 42302 633800
rect 42260 630674 42288 633791
rect 42260 630646 42380 630674
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625478 42380 630646
rect 42182 625450 42380 625478
rect 42444 625274 42472 634786
rect 42076 625246 42472 625274
rect 42076 624784 42104 625246
rect 42246 625016 42302 625025
rect 42536 625002 42564 635854
rect 42628 634814 42656 635990
rect 42798 635760 42854 635769
rect 42798 635695 42854 635704
rect 42628 634786 42748 634814
rect 42302 624974 42564 625002
rect 42246 624951 42302 624960
rect 42062 624472 42118 624481
rect 42062 624407 42118 624416
rect 42076 624172 42104 624407
rect 42168 623070 42288 623098
rect 42168 622948 42196 623070
rect 42260 622962 42288 623070
rect 42720 622962 42748 634786
rect 42260 622934 42748 622962
rect 41786 622160 41842 622169
rect 41786 622095 41842 622104
rect 41800 621792 41828 622095
rect 42154 621616 42210 621625
rect 42154 621551 42210 621560
rect 42168 621112 42196 621551
rect 42062 620800 42118 620809
rect 42062 620735 42118 620744
rect 42076 620500 42104 620735
rect 41970 620256 42026 620265
rect 41970 620191 42026 620200
rect 41984 619956 42012 620191
rect 42812 619698 42840 635695
rect 42260 619670 42840 619698
rect 42260 617454 42288 619670
rect 42430 619304 42486 619313
rect 42430 619239 42486 619248
rect 42182 617426 42288 617454
rect 42444 616842 42472 619239
rect 42614 619032 42670 619041
rect 42614 618967 42670 618976
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42628 616162 42656 618967
rect 42182 616134 42656 616162
rect 42246 616040 42302 616049
rect 42246 615975 42302 615984
rect 41786 615768 41842 615777
rect 41786 615703 41842 615712
rect 41800 615604 41828 615703
rect 42260 613782 42288 615975
rect 42890 615632 42946 615641
rect 42890 615567 42946 615576
rect 42904 615494 42932 615567
rect 42182 613754 42288 613782
rect 42628 615466 42932 615494
rect 42628 613170 42656 615466
rect 42536 613142 42656 613170
rect 42536 613135 42564 613142
rect 42182 613107 42564 613135
rect 41786 612776 41842 612785
rect 41786 612711 41842 612720
rect 41800 612476 41828 612711
rect 43088 612377 43116 762991
rect 43272 630674 43300 807463
rect 43456 796249 43484 809503
rect 43442 796240 43498 796249
rect 43442 796175 43498 796184
rect 43442 633448 43498 633457
rect 43442 633383 43498 633392
rect 43272 630646 43392 630674
rect 43364 612898 43392 630646
rect 43456 615494 43484 633383
rect 43456 615466 43576 615494
rect 43364 612870 43484 612898
rect 43074 612368 43130 612377
rect 43456 612354 43484 612870
rect 43548 612490 43576 615466
rect 43640 612762 43668 933263
rect 43810 932104 43866 932113
rect 43810 932039 43866 932048
rect 43824 612950 43852 932039
rect 44086 892800 44142 892809
rect 44086 892735 44088 892744
rect 44140 892735 44142 892744
rect 44088 892706 44140 892712
rect 44086 891984 44142 891993
rect 44086 891919 44088 891928
rect 44140 891919 44142 891928
rect 44088 891890 44140 891896
rect 44454 816096 44510 816105
rect 44454 816031 44510 816040
rect 44270 810384 44326 810393
rect 44270 810319 44326 810328
rect 43994 806304 44050 806313
rect 43994 806239 44050 806248
rect 43812 612944 43864 612950
rect 43812 612886 43864 612892
rect 43640 612746 43760 612762
rect 43640 612740 43772 612746
rect 43640 612734 43720 612740
rect 43720 612682 43772 612688
rect 44008 612610 44036 806239
rect 44284 790809 44312 810319
rect 44270 790800 44326 790809
rect 44270 790735 44326 790744
rect 44468 773265 44496 816031
rect 44652 815697 44680 941015
rect 47596 891993 47624 991714
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 48976 940137 49004 990082
rect 48962 940128 49018 940137
rect 48962 940063 49018 940072
rect 50356 939865 50384 993142
rect 54484 992928 54536 992934
rect 54484 992870 54536 992876
rect 51724 991636 51776 991642
rect 51724 991578 51776 991584
rect 51736 942313 51764 991578
rect 53288 990276 53340 990282
rect 53288 990218 53340 990224
rect 51722 942304 51778 942313
rect 51722 942239 51778 942248
rect 50342 939856 50398 939865
rect 50342 939791 50398 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44638 815688 44694 815697
rect 44638 815623 44694 815632
rect 45006 815280 45062 815289
rect 45006 815215 45062 815224
rect 44638 814464 44694 814473
rect 44638 814399 44694 814408
rect 44454 773256 44510 773265
rect 44454 773191 44510 773200
rect 44454 772848 44510 772857
rect 44454 772783 44510 772792
rect 44270 772032 44326 772041
rect 44270 771967 44326 771976
rect 44284 729337 44312 771967
rect 44468 730153 44496 772783
rect 44652 771633 44680 814399
rect 44822 813648 44878 813657
rect 44822 813583 44878 813592
rect 44638 771624 44694 771633
rect 44638 771559 44694 771568
rect 44836 771474 44864 813583
rect 45020 772449 45048 815215
rect 45190 807936 45246 807945
rect 45190 807871 45246 807880
rect 45204 796793 45232 807871
rect 45190 796784 45246 796793
rect 45190 796719 45246 796728
rect 45006 772440 45062 772449
rect 45006 772375 45062 772384
rect 44652 771446 44864 771474
rect 44652 770817 44680 771446
rect 44822 771216 44878 771225
rect 44822 771151 44878 771160
rect 44638 770808 44694 770817
rect 44638 770743 44694 770752
rect 44638 770400 44694 770409
rect 44638 770335 44694 770344
rect 44454 730144 44510 730153
rect 44454 730079 44510 730088
rect 44270 729328 44326 729337
rect 44270 729263 44326 729272
rect 44454 728920 44510 728929
rect 44454 728855 44510 728864
rect 44270 728104 44326 728113
rect 44270 728039 44326 728048
rect 44284 685273 44312 728039
rect 44468 686089 44496 728855
rect 44652 727705 44680 770335
rect 44836 728521 44864 771151
rect 45098 766728 45154 766737
rect 45098 766663 45154 766672
rect 45112 749329 45140 766663
rect 45282 764824 45338 764833
rect 45282 764759 45338 764768
rect 45296 753545 45324 764759
rect 46018 764280 46074 764289
rect 46018 764215 46074 764224
rect 45282 753536 45338 753545
rect 45282 753471 45338 753480
rect 45098 749320 45154 749329
rect 45098 749255 45154 749264
rect 45006 729736 45062 729745
rect 45006 729671 45062 729680
rect 44822 728512 44878 728521
rect 44822 728447 44878 728456
rect 44638 727696 44694 727705
rect 44638 727631 44694 727640
rect 44638 727424 44694 727433
rect 44638 727359 44694 727368
rect 44454 686080 44510 686089
rect 44454 686015 44510 686024
rect 44270 685264 44326 685273
rect 44270 685199 44326 685208
rect 44362 684856 44418 684865
rect 44362 684791 44418 684800
rect 44178 679552 44234 679561
rect 44178 679487 44234 679496
rect 44192 666641 44220 679487
rect 44178 666632 44234 666641
rect 44178 666567 44234 666576
rect 44376 642297 44404 684791
rect 44652 684457 44680 727359
rect 44822 722800 44878 722809
rect 44822 722735 44878 722744
rect 44836 709481 44864 722735
rect 44822 709472 44878 709481
rect 44822 709407 44878 709416
rect 45020 686905 45048 729671
rect 45190 723616 45246 723625
rect 45190 723551 45246 723560
rect 45204 705537 45232 723551
rect 45190 705528 45246 705537
rect 45190 705463 45246 705472
rect 45006 686896 45062 686905
rect 45006 686831 45062 686840
rect 44822 686488 44878 686497
rect 44822 686423 44878 686432
rect 44638 684448 44694 684457
rect 44638 684383 44694 684392
rect 44546 680368 44602 680377
rect 44546 680303 44602 680312
rect 44560 662969 44588 680303
rect 44546 662960 44602 662969
rect 44546 662895 44602 662904
rect 44836 643657 44864 686423
rect 45006 685672 45062 685681
rect 45006 685607 45062 685616
rect 44822 643648 44878 643657
rect 44822 643583 44878 643592
rect 44638 643376 44694 643385
rect 44638 643311 44694 643320
rect 44362 642288 44418 642297
rect 44362 642223 44418 642232
rect 44178 635352 44234 635361
rect 44178 635287 44234 635296
rect 44192 620809 44220 635287
rect 44362 634536 44418 634545
rect 44362 634471 44418 634480
rect 44178 620800 44234 620809
rect 44178 620735 44234 620744
rect 44376 615494 44404 634471
rect 44376 615466 44588 615494
rect 44178 614136 44234 614145
rect 44178 614071 44234 614080
rect 43996 612604 44048 612610
rect 43996 612546 44048 612552
rect 43548 612462 43944 612490
rect 43718 612368 43774 612377
rect 43456 612338 43622 612354
rect 43456 612332 43634 612338
rect 43456 612326 43582 612332
rect 43074 612303 43130 612312
rect 43718 612303 43720 612312
rect 43582 612274 43634 612280
rect 43772 612303 43774 612312
rect 43720 612274 43772 612280
rect 43916 611130 43944 612462
rect 44192 611674 44220 614071
rect 44167 611646 44220 611674
rect 44167 611318 44195 611646
rect 44155 611312 44207 611318
rect 44155 611254 44207 611260
rect 43916 611114 44419 611130
rect 43916 611108 44431 611114
rect 43916 611102 44379 611108
rect 44379 611050 44431 611056
rect 44270 611008 44326 611017
rect 44560 610994 44588 615466
rect 44270 610943 44272 610952
rect 44324 610943 44326 610952
rect 44514 610966 44588 610994
rect 44272 610914 44324 610920
rect 44514 610774 44542 610966
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 44652 600545 44680 643311
rect 45020 643113 45048 685607
rect 45374 684040 45430 684049
rect 45374 683975 45430 683984
rect 45006 643104 45062 643113
rect 45006 643039 45062 643048
rect 44822 642560 44878 642569
rect 44822 642495 44878 642504
rect 44638 600536 44694 600545
rect 44638 600471 44694 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 42430 596864 42486 596873
rect 42430 596799 42486 596808
rect 41234 596048 41290 596057
rect 41234 595983 41290 595992
rect 33782 595640 33838 595649
rect 33782 595575 33838 595584
rect 32402 594824 32458 594833
rect 32402 594759 32458 594768
rect 32416 585721 32444 594759
rect 33796 585818 33824 595575
rect 36542 595232 36598 595241
rect 36542 595167 36598 595176
rect 33784 585812 33836 585818
rect 33784 585754 33836 585760
rect 32402 585712 32458 585721
rect 32402 585647 32458 585656
rect 36556 585206 36584 595167
rect 41248 594726 41276 595983
rect 41236 594720 41288 594726
rect 41236 594662 41288 594668
rect 41512 594720 41564 594726
rect 41512 594662 41564 594668
rect 37922 594416 37978 594425
rect 37922 594351 37978 594360
rect 37936 585342 37964 594351
rect 40682 593600 40738 593609
rect 40682 593535 40738 593544
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 585993 39988 590679
rect 40500 589688 40552 589694
rect 40498 589656 40500 589665
rect 40552 589656 40554 589665
rect 40498 589591 40554 589600
rect 39946 585984 40002 585993
rect 39946 585919 40002 585928
rect 39672 585812 39724 585818
rect 39672 585754 39724 585760
rect 37924 585336 37976 585342
rect 39684 585313 39712 585754
rect 37924 585278 37976 585284
rect 39670 585304 39726 585313
rect 39670 585239 39726 585248
rect 36544 585200 36596 585206
rect 36544 585142 36596 585148
rect 40224 585200 40276 585206
rect 40224 585142 40276 585148
rect 40236 585041 40264 585142
rect 40222 585032 40278 585041
rect 40222 584967 40278 584976
rect 40696 584633 40724 593535
rect 41524 585993 41552 594662
rect 42062 593192 42118 593201
rect 42062 593127 42118 593136
rect 41878 592784 41934 592793
rect 41878 592719 41934 592728
rect 41892 589778 41920 592719
rect 41708 589750 41920 589778
rect 41708 589694 41736 589750
rect 41696 589688 41748 589694
rect 41696 589630 41748 589636
rect 42076 589393 42104 593127
rect 42062 589384 42118 589393
rect 42062 589319 42118 589328
rect 41510 585984 41566 585993
rect 41510 585919 41566 585928
rect 41420 585336 41472 585342
rect 41420 585278 41472 585284
rect 41432 584633 41460 585278
rect 42246 585032 42302 585041
rect 42246 584967 42302 584976
rect 40682 584624 40738 584633
rect 40682 584559 40738 584568
rect 41418 584624 41474 584633
rect 41418 584559 41474 584568
rect 42260 583454 42288 584967
rect 42182 583426 42288 583454
rect 41786 582584 41842 582593
rect 41786 582519 41842 582528
rect 41800 582249 41828 582519
rect 42444 581890 42472 596799
rect 42798 594008 42854 594017
rect 42798 593943 42854 593952
rect 42812 587894 42840 593943
rect 42812 587866 42932 587894
rect 42706 585984 42762 585993
rect 42706 585919 42762 585928
rect 42352 581862 42472 581890
rect 42352 581618 42380 581862
rect 42182 581590 42380 581618
rect 42246 581496 42302 581505
rect 42246 581431 42302 581440
rect 42260 580975 42288 581431
rect 42182 580947 42288 580975
rect 42430 580680 42486 580689
rect 42430 580615 42486 580624
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42062 580136 42118 580145
rect 42118 580094 42288 580122
rect 42062 580071 42118 580080
rect 42062 578912 42118 578921
rect 42062 578847 42118 578856
rect 42076 578544 42104 578847
rect 42260 578377 42288 580094
rect 42444 578558 42472 580615
rect 42444 578530 42564 578558
rect 42246 578368 42302 578377
rect 42246 578303 42302 578312
rect 42536 578218 42564 578530
rect 42720 578234 42748 585919
rect 42168 578190 42564 578218
rect 42628 578206 42748 578234
rect 42168 577932 42196 578190
rect 42246 577824 42302 577833
rect 42246 577759 42302 577768
rect 42260 577295 42288 577759
rect 42628 577402 42656 578206
rect 42182 577267 42288 577295
rect 42352 577374 42656 577402
rect 42352 576994 42380 577374
rect 42352 576966 42472 576994
rect 42246 576872 42302 576881
rect 42246 576807 42302 576816
rect 41984 576609 42012 576708
rect 41970 576600 42026 576609
rect 41970 576535 42026 576544
rect 42260 574274 42288 576807
rect 42182 574246 42288 574274
rect 42154 574152 42210 574161
rect 42154 574087 42210 574096
rect 42168 573580 42196 574087
rect 42444 573730 42472 576966
rect 42904 574161 42932 587866
rect 42996 579614 43024 596935
rect 44454 591968 44510 591977
rect 44454 591903 44510 591912
rect 43442 590336 43498 590345
rect 43442 590271 43498 590280
rect 42996 579586 43208 579614
rect 42890 574152 42946 574161
rect 42890 574087 42946 574096
rect 42352 573702 42472 573730
rect 41970 573200 42026 573209
rect 41970 573135 42026 573144
rect 41984 572968 42012 573135
rect 42352 572438 42380 573702
rect 42168 572370 42196 572424
rect 42260 572410 42380 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42430 571704 42486 571713
rect 42430 571639 42486 571648
rect 42246 571432 42302 571441
rect 42246 571367 42302 571376
rect 42062 571024 42118 571033
rect 42062 570959 42118 570968
rect 42076 570588 42104 570959
rect 42260 569922 42288 571367
rect 42182 569894 42288 569922
rect 42444 569310 42472 571639
rect 43180 569954 43208 579586
rect 42168 569242 42196 569296
rect 42260 569282 42472 569310
rect 42996 569926 43208 569954
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42246 569120 42302 569129
rect 42246 569055 42302 569064
rect 42260 563054 42288 569055
rect 41524 563026 42288 563054
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 41524 557598 41552 563026
rect 42062 558512 42118 558521
rect 42062 558447 42118 558456
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 41512 557592 41564 557598
rect 42076 557569 42104 558447
rect 41512 557534 41564 557540
rect 42062 557560 42118 557569
rect 42996 557534 43024 569926
rect 42062 557495 42118 557504
rect 42812 557506 43024 557534
rect 35806 554840 35862 554849
rect 42812 554826 42840 557506
rect 41708 554810 42840 554826
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 41696 554804 42840 554810
rect 35808 554746 35860 554752
rect 41748 554798 42840 554804
rect 41696 554746 41748 554752
rect 35622 554024 35678 554033
rect 35622 553959 35678 553968
rect 35636 553450 35664 553959
rect 35806 553616 35862 553625
rect 35806 553551 35808 553560
rect 35860 553551 35862 553560
rect 41420 553580 41472 553586
rect 35808 553522 35860 553528
rect 41420 553522 41472 553528
rect 35624 553444 35676 553450
rect 35624 553386 35676 553392
rect 41432 553394 41460 553522
rect 41696 553444 41748 553450
rect 41432 553366 41552 553394
rect 41748 553392 41828 553394
rect 41696 553386 41828 553392
rect 41708 553366 41828 553386
rect 40866 553208 40922 553217
rect 40866 553143 40922 553152
rect 33782 551984 33838 551993
rect 33782 551919 33838 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 33796 543046 33824 551919
rect 40880 549794 40908 553143
rect 41234 551168 41290 551177
rect 41234 551103 41290 551112
rect 41248 550798 41276 551103
rect 41236 550792 41288 550798
rect 41236 550734 41288 550740
rect 40880 549766 41092 549794
rect 37188 547460 37240 547466
rect 37188 547402 37240 547408
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 37200 542366 37228 547402
rect 41064 546802 41092 549766
rect 41234 549536 41290 549545
rect 41234 549471 41290 549480
rect 41248 549302 41276 549471
rect 41236 549296 41288 549302
rect 41236 549238 41288 549244
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41064 546774 41368 546802
rect 41340 546417 41368 546774
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 41524 543734 41552 553366
rect 41800 553217 41828 553366
rect 41786 553208 41842 553217
rect 41786 553143 41842 553152
rect 43166 552392 43222 552401
rect 43166 552327 43222 552336
rect 41696 550792 41748 550798
rect 41748 550752 42840 550780
rect 41696 550734 41748 550740
rect 42062 550352 42118 550361
rect 42062 550287 42118 550296
rect 41878 549944 41934 549953
rect 41878 549879 41934 549888
rect 41694 549400 41750 549409
rect 41694 549335 41696 549344
rect 41748 549335 41750 549344
rect 41696 549306 41748 549312
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 41892 545465 41920 549879
rect 42076 545737 42104 550287
rect 42062 545728 42118 545737
rect 42062 545663 42118 545672
rect 41878 545456 41934 545465
rect 41878 545391 41934 545400
rect 41524 543706 42472 543734
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 37188 542360 37240 542366
rect 37188 542302 37240 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538778 42472 543706
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42076 538750 42472 538778
rect 42076 538424 42104 538750
rect 42246 538248 42302 538257
rect 42246 538183 42302 538192
rect 42062 537976 42118 537985
rect 42062 537911 42118 537920
rect 42076 537744 42104 537911
rect 42168 536466 42196 536588
rect 42260 536466 42288 538183
rect 42628 537985 42656 540223
rect 42614 537976 42670 537985
rect 42614 537911 42670 537920
rect 42168 536438 42288 536466
rect 42168 535265 42196 535364
rect 42154 535256 42210 535265
rect 42154 535191 42210 535200
rect 41786 534984 41842 534993
rect 41786 534919 41842 534928
rect 41800 534752 41828 534919
rect 42154 534440 42210 534449
rect 42154 534375 42210 534384
rect 42168 534072 42196 534375
rect 42154 533896 42210 533905
rect 42154 533831 42210 533840
rect 42168 533528 42196 533831
rect 42246 533216 42302 533225
rect 42246 533151 42302 533160
rect 42260 531162 42288 533151
rect 42812 532930 42840 550752
rect 42982 549400 43038 549409
rect 42982 549335 43038 549344
rect 42996 533225 43024 549335
rect 43180 533905 43208 552327
rect 43166 533896 43222 533905
rect 43166 533831 43222 533840
rect 42982 533216 43038 533225
rect 42982 533151 43038 533160
rect 42720 532902 42840 532930
rect 42522 532808 42578 532817
rect 42522 532743 42578 532752
rect 42168 531134 42288 531162
rect 42168 531045 42196 531134
rect 42536 530890 42564 532743
rect 42352 530862 42564 530890
rect 42352 530754 42380 530862
rect 42260 530726 42380 530754
rect 42260 530414 42288 530726
rect 42522 530632 42578 530641
rect 42182 530386 42288 530414
rect 42352 530590 42522 530618
rect 42154 530088 42210 530097
rect 42154 530023 42210 530032
rect 42168 529757 42196 530023
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42352 527626 42380 530590
rect 42522 530567 42578 530576
rect 42720 530097 42748 532902
rect 42706 530088 42762 530097
rect 42706 530023 42762 530032
rect 42614 529680 42670 529689
rect 42614 529615 42670 529624
rect 42168 527598 42380 527626
rect 42168 527340 42196 527598
rect 42628 526742 42656 529615
rect 42890 529136 42946 529145
rect 42182 526714 42656 526742
rect 42720 529094 42890 529122
rect 42720 526091 42748 529094
rect 42890 529071 42946 529080
rect 42182 526063 42748 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 40958 426048 41014 426057
rect 40958 425983 41014 425992
rect 40774 425640 40830 425649
rect 40774 425575 40830 425584
rect 36542 424416 36598 424425
rect 36542 424351 36598 424360
rect 36556 415410 36584 424351
rect 40498 421968 40554 421977
rect 40498 421903 40554 421912
rect 40512 418713 40540 421903
rect 40788 418849 40816 425575
rect 40972 423230 41000 425983
rect 41326 424008 41382 424017
rect 41326 423943 41382 423952
rect 41340 423842 41368 423943
rect 41328 423836 41380 423842
rect 41328 423778 41380 423784
rect 41696 423836 41748 423842
rect 41748 423796 42840 423824
rect 41696 423778 41748 423784
rect 40960 423224 41012 423230
rect 40960 423166 41012 423172
rect 41604 423224 41656 423230
rect 41656 423172 42012 423178
rect 41604 423166 42012 423172
rect 41616 423150 42012 423166
rect 41786 423056 41842 423065
rect 41786 422991 41842 423000
rect 41800 422249 41828 422991
rect 41786 422240 41842 422249
rect 41786 422175 41842 422184
rect 41786 421560 41842 421569
rect 41786 421495 41842 421504
rect 40774 418840 40830 418849
rect 40774 418775 40830 418784
rect 40498 418704 40554 418713
rect 40498 418639 40554 418648
rect 41800 418305 41828 421495
rect 41786 418296 41842 418305
rect 41786 418231 41842 418240
rect 41984 418154 42012 423150
rect 42154 422784 42210 422793
rect 42154 422719 42210 422728
rect 42168 418577 42196 422719
rect 42522 419928 42578 419937
rect 42522 419863 42578 419872
rect 42154 418568 42210 418577
rect 42154 418503 42210 418512
rect 41984 418126 42380 418154
rect 36544 415404 36596 415410
rect 36544 415346 36596 415352
rect 41696 415404 41748 415410
rect 41696 415346 41748 415352
rect 41708 415290 41736 415346
rect 41708 415262 42288 415290
rect 42260 413114 42288 415262
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42352 411074 42380 418126
rect 42536 411913 42564 419863
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42380 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42430 407144 42486 407153
rect 42182 407102 42430 407130
rect 42430 407079 42486 407088
rect 42430 406872 42486 406881
rect 42430 406807 42486 406816
rect 42444 406518 42472 406807
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42182 402138 42472 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42444 400217 42472 402138
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423796
rect 43074 422240 43130 422249
rect 43074 422175 43130 422184
rect 43088 402937 43116 422175
rect 43258 421152 43314 421161
rect 43258 421087 43314 421096
rect 43272 407833 43300 421087
rect 43258 407824 43314 407833
rect 43258 407759 43314 407768
rect 43074 402928 43130 402937
rect 43074 402863 43130 402872
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41340 387654 41552 387682
rect 41142 387152 41198 387161
rect 41142 387087 41144 387096
rect 41196 387087 41198 387096
rect 41144 387058 41196 387064
rect 41340 386753 41368 387654
rect 41524 386753 41552 387654
rect 41708 387122 41920 387138
rect 41696 387116 41920 387122
rect 41748 387110 41920 387116
rect 41696 387058 41748 387064
rect 41892 387025 41920 387110
rect 41878 387016 41934 387025
rect 41878 386951 41934 386960
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 41142 383072 41198 383081
rect 41142 383007 41198 383016
rect 41156 382294 41184 383007
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41696 382424 41748 382430
rect 41748 382384 41920 382412
rect 41696 382366 41748 382372
rect 41144 382288 41196 382294
rect 40038 382256 40094 382265
rect 41696 382288 41748 382294
rect 41144 382230 41196 382236
rect 41694 382256 41696 382265
rect 41748 382256 41750 382265
rect 40038 382191 40094 382200
rect 41694 382191 41750 382200
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 35820 379409 35848 379510
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 40052 376553 40080 382191
rect 40774 381440 40830 381449
rect 40774 381375 40830 381384
rect 40788 378593 40816 381375
rect 41326 381032 41382 381041
rect 41326 380967 41382 380976
rect 40774 378584 40830 378593
rect 40774 378519 40830 378528
rect 41340 377777 41368 380967
rect 41696 379568 41748 379574
rect 41696 379510 41748 379516
rect 41892 379514 41920 382384
rect 42798 382256 42854 382265
rect 42798 382191 42854 382200
rect 41708 379409 41736 379510
rect 41892 379486 42564 379514
rect 41694 379400 41750 379409
rect 41694 379335 41750 379344
rect 41326 377768 41382 377777
rect 41326 377703 41382 377712
rect 42338 377768 42394 377777
rect 42338 377703 42394 377712
rect 42352 376754 42380 377703
rect 42352 376726 42472 376754
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 40038 376544 40094 376553
rect 40038 376479 40094 376488
rect 28906 376136 28962 376145
rect 28906 376071 28962 376080
rect 28920 371890 28948 376071
rect 35820 376038 35848 376479
rect 35808 376032 35860 376038
rect 35808 375974 35860 375980
rect 39488 376032 39540 376038
rect 39488 375974 39540 375980
rect 39500 375737 39528 375974
rect 39486 375728 39542 375737
rect 39486 375663 39542 375672
rect 41694 371920 41750 371929
rect 28908 371884 28960 371890
rect 41694 371855 41696 371864
rect 28908 371826 28960 371832
rect 41748 371855 41750 371864
rect 41696 371826 41748 371832
rect 42444 369458 42472 376726
rect 42182 369430 42472 369458
rect 41786 368656 41842 368665
rect 41786 368591 41842 368600
rect 41800 368249 41828 368591
rect 42536 367622 42564 379486
rect 42182 367594 42564 367622
rect 42430 367024 42486 367033
rect 42182 366968 42430 366975
rect 42182 366959 42486 366968
rect 42182 366947 42472 366959
rect 42430 365800 42486 365809
rect 42182 365758 42430 365786
rect 42430 365735 42486 365744
rect 41800 364313 41828 364548
rect 41786 364304 41842 364313
rect 41786 364239 41842 364248
rect 42182 363922 42472 363950
rect 41786 363624 41842 363633
rect 41786 363559 41842 363568
rect 41800 363256 41828 363559
rect 41786 362944 41842 362953
rect 41786 362879 41842 362888
rect 41800 362712 41828 362879
rect 42444 361593 42472 363922
rect 42430 361584 42486 361593
rect 42430 361519 42486 361528
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 42182 358958 42472 358986
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42444 357377 42472 358958
rect 42430 357368 42486 357377
rect 42430 357303 42486 357312
rect 42812 356674 42840 382191
rect 43456 379514 43484 590271
rect 44468 578921 44496 591903
rect 44454 578912 44510 578921
rect 44454 578847 44510 578856
rect 44652 557297 44680 600063
rect 44836 599729 44864 642495
rect 45388 641481 45416 683975
rect 45650 677920 45706 677929
rect 45650 677855 45706 677864
rect 45374 641472 45430 641481
rect 45374 641407 45430 641416
rect 45190 641200 45246 641209
rect 45190 641135 45246 641144
rect 45006 640928 45062 640937
rect 45006 640863 45062 640872
rect 44822 599720 44878 599729
rect 44822 599655 44878 599664
rect 44822 599312 44878 599321
rect 44822 599247 44878 599256
rect 44638 557288 44694 557297
rect 44638 557223 44694 557232
rect 44836 556481 44864 599247
rect 45020 598097 45048 640863
rect 45204 598913 45232 641135
rect 45664 611017 45692 677855
rect 45834 637800 45890 637809
rect 45834 637735 45890 637744
rect 45848 615641 45876 637735
rect 45834 615632 45890 615641
rect 45834 615567 45890 615576
rect 46032 611930 46060 764215
rect 46216 756401 46244 870810
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 46202 756392 46258 756401
rect 46202 756327 46258 756336
rect 46938 721168 46994 721177
rect 46938 721103 46994 721112
rect 46204 647896 46256 647902
rect 46204 647838 46256 647844
rect 46020 611924 46072 611930
rect 46020 611866 46072 611872
rect 45650 611008 45706 611017
rect 45650 610943 45706 610952
rect 46216 600953 46244 647838
rect 46386 636984 46442 636993
rect 46386 636919 46442 636928
rect 46400 619313 46428 636919
rect 46386 619304 46442 619313
rect 46386 619239 46442 619248
rect 46952 611522 46980 721103
rect 47596 712201 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47858 719944 47914 719953
rect 47858 719879 47914 719888
rect 47582 712192 47638 712201
rect 47582 712127 47638 712136
rect 47674 676696 47730 676705
rect 47674 676631 47730 676640
rect 47688 669314 47716 676631
rect 47688 669286 47808 669314
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47214 638208 47270 638217
rect 47214 638143 47270 638152
rect 47228 619041 47256 638143
rect 47398 636440 47454 636449
rect 47398 636375 47454 636384
rect 47412 621625 47440 636375
rect 47398 621616 47454 621625
rect 47398 621551 47454 621560
rect 47214 619032 47270 619041
rect 47214 618967 47270 618976
rect 46940 611516 46992 611522
rect 46940 611458 46992 611464
rect 46202 600944 46258 600953
rect 46202 600879 46258 600888
rect 45190 598904 45246 598913
rect 45190 598839 45246 598848
rect 45190 598496 45246 598505
rect 45190 598431 45246 598440
rect 45006 598088 45062 598097
rect 45006 598023 45062 598032
rect 45204 582374 45232 598431
rect 47596 582457 47624 662390
rect 47780 614145 47808 669286
rect 47872 634814 47900 719879
rect 48976 669361 49004 767314
rect 50356 730561 50384 805938
rect 53116 799377 53144 923238
rect 53300 892265 53328 990218
rect 54496 892537 54524 992870
rect 55864 991500 55916 991506
rect 55864 991442 55916 991448
rect 55876 892809 55904 991442
rect 95896 990282 95924 1001914
rect 96080 991778 96108 1002050
rect 96264 998102 96292 1005994
rect 97448 1002788 97500 1002794
rect 97448 1002730 97500 1002736
rect 97264 1002380 97316 1002386
rect 97264 1002322 97316 1002328
rect 96252 998096 96304 998102
rect 96252 998038 96304 998044
rect 97276 994809 97304 1002322
rect 97262 994800 97318 994809
rect 97262 994735 97318 994744
rect 97460 994566 97488 1002730
rect 100298 1002688 100354 1002697
rect 100298 1002623 100300 1002632
rect 100352 1002623 100354 1002632
rect 100300 1002594 100352 1002600
rect 100024 1002516 100076 1002522
rect 100024 1002458 100076 1002464
rect 98644 1002244 98696 1002250
rect 98644 1002186 98696 1002192
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 98656 994702 98684 1002186
rect 99102 1002144 99158 1002153
rect 99102 1002079 99104 1002088
rect 99156 1002079 99158 1002088
rect 99104 1002050 99156 1002056
rect 98828 1001972 98880 1001978
rect 98828 1001914 98880 1001920
rect 98840 995761 98868 1001914
rect 98826 995752 98882 995761
rect 98826 995687 98882 995696
rect 98644 994696 98696 994702
rect 98644 994638 98696 994644
rect 97448 994560 97500 994566
rect 100036 994537 100064 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100300 1002322 100352 1002328
rect 100208 1002108 100260 1002114
rect 100208 1002050 100260 1002056
rect 100220 998442 100248 1002050
rect 101126 1002008 101182 1002017
rect 101126 1001943 101128 1001952
rect 101180 1001943 101182 1001952
rect 101128 1001914 101180 1001920
rect 100208 998436 100260 998442
rect 100208 998378 100260 998384
rect 101416 995081 101444 1005994
rect 102784 1005304 102836 1005310
rect 102784 1005246 102836 1005252
rect 102322 1002824 102378 1002833
rect 102322 1002759 102324 1002768
rect 102376 1002759 102378 1002768
rect 102324 1002730 102376 1002736
rect 101954 1002280 102010 1002289
rect 101954 1002215 101956 1002224
rect 102008 1002215 102010 1002224
rect 101956 1002186 102008 1002192
rect 101402 995072 101458 995081
rect 101402 995007 101458 995016
rect 97448 994502 97500 994508
rect 100022 994528 100078 994537
rect 100022 994463 100078 994472
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 990276 95936 990282
rect 95884 990218 95936 990224
rect 89628 987420 89680 987426
rect 89628 987362 89680 987368
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 987362
rect 102796 985998 102824 1005246
rect 102980 999802 103008 1006130
rect 103978 1006088 104034 1006097
rect 103978 1006023 103980 1006032
rect 104032 1006023 104034 1006032
rect 106002 1006088 106058 1006097
rect 106002 1006023 106004 1006032
rect 103980 1005994 104032 1006000
rect 106056 1006023 106058 1006032
rect 106004 1005994 106056 1006000
rect 108856 1005304 108908 1005310
rect 108854 1005272 108856 1005281
rect 108908 1005272 108910 1005281
rect 108854 1005207 108910 1005216
rect 108486 1004728 108542 1004737
rect 106188 1004692 106240 1004698
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 103150 1002552 103206 1002561
rect 103150 1002487 103152 1002496
rect 103204 1002487 103206 1002496
rect 103152 1002458 103204 1002464
rect 105634 1002280 105690 1002289
rect 105634 1002215 105636 1002224
rect 105688 1002215 105690 1002224
rect 105636 1002186 105688 1002192
rect 103150 1002144 103206 1002153
rect 103150 1002079 103152 1002088
rect 103204 1002079 103206 1002088
rect 103978 1002144 104034 1002153
rect 103978 1002079 103980 1002088
rect 103152 1002050 103204 1002056
rect 104032 1002079 104034 1002088
rect 103980 1002050 104032 1002056
rect 104806 1002008 104862 1002017
rect 104176 1001966 104806 1001994
rect 102968 999796 103020 999802
rect 102968 999738 103020 999744
rect 104176 994838 104204 1001966
rect 104806 1001943 104862 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 104164 994832 104216 994838
rect 104164 994774 104216 994780
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1004634
rect 107658 1002416 107714 1002425
rect 107658 1002351 107660 1002360
rect 107712 1002351 107714 1002360
rect 109500 1002380 109552 1002386
rect 107660 1002322 107712 1002328
rect 109500 1002322 109552 1002328
rect 108026 1002280 108082 1002289
rect 107844 1002244 107896 1002250
rect 108026 1002215 108028 1002224
rect 107844 1002186 107896 1002192
rect 108080 1002215 108082 1002224
rect 108028 1002186 108080 1002192
rect 106830 1002144 106886 1002153
rect 106464 1002108 106516 1002114
rect 106830 1002079 106832 1002088
rect 106464 1002050 106516 1002056
rect 106884 1002079 106886 1002088
rect 107856 1002096 107884 1002186
rect 109040 1002108 109092 1002114
rect 107856 1002068 108160 1002096
rect 106832 1002050 106884 1002056
rect 106476 997762 106504 1002050
rect 107752 1001972 107804 1001978
rect 107752 1001914 107804 1001920
rect 106464 997756 106516 997762
rect 106464 997698 106516 997704
rect 107764 993206 107792 1001914
rect 107752 993200 107804 993206
rect 107752 993142 107804 993148
rect 108132 990146 108160 1002068
rect 109040 1002050 109092 1002056
rect 109052 993070 109080 1002050
rect 109512 997626 109540 1002322
rect 110420 1002244 110472 1002250
rect 110420 1002186 110472 1002192
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 997620 109552 997626
rect 109500 997562 109552 997568
rect 109040 993064 109092 993070
rect 109040 993006 109092 993012
rect 110432 991642 110460 1002186
rect 111800 1002108 111852 1002114
rect 111800 1002050 111852 1002056
rect 110420 991636 110472 991642
rect 110420 991578 110472 991584
rect 108120 990140 108172 990146
rect 108120 990082 108172 990088
rect 111812 987426 111840 1002050
rect 113836 997762 113864 1006130
rect 124864 1006052 124916 1006058
rect 124864 1005994 124916 1006000
rect 113824 997756 113876 997762
rect 113824 997698 113876 997704
rect 117136 997756 117188 997762
rect 117136 997698 117188 997704
rect 116216 997620 116268 997626
rect 116216 997562 116268 997568
rect 116228 996985 116256 997562
rect 117148 997257 117176 997698
rect 117134 997248 117190 997257
rect 117134 997183 117190 997192
rect 116214 996976 116270 996985
rect 116214 996911 116270 996920
rect 121736 996396 121788 996402
rect 121736 996338 121788 996344
rect 111800 987420 111852 987426
rect 111800 987362 111852 987368
rect 105846 983606 106228 983634
rect 121748 983634 121776 996338
rect 124876 995081 124904 1005994
rect 126256 996169 126284 1006266
rect 143998 1000648 144054 1000657
rect 143998 1000583 144054 1000592
rect 143724 997756 143776 997762
rect 143724 997698 143776 997704
rect 143736 997257 143764 997698
rect 143722 997248 143778 997257
rect 143722 997183 143778 997192
rect 143724 996532 143776 996538
rect 143724 996474 143776 996480
rect 126242 996160 126298 996169
rect 126242 996095 126298 996104
rect 136468 995858 136496 995860
rect 136456 995852 136508 995858
rect 136456 995794 136508 995800
rect 138018 995752 138074 995761
rect 137770 995710 138018 995738
rect 141790 995752 141846 995761
rect 141450 995710 141790 995738
rect 138018 995687 138074 995696
rect 143736 995738 143764 996474
rect 144012 995761 144040 1000583
rect 144196 997754 144224 1006470
rect 144368 1006256 144420 1006262
rect 144368 1006198 144420 1006204
rect 144380 997754 144408 1006198
rect 144196 997726 144316 997754
rect 144380 997726 144776 997754
rect 144288 997642 144316 997726
rect 144288 997614 144408 997642
rect 144184 997552 144236 997558
rect 144184 997494 144236 997500
rect 144196 996985 144224 997494
rect 144182 996976 144238 996985
rect 144182 996911 144238 996920
rect 144184 996396 144236 996402
rect 144184 996338 144236 996344
rect 141790 995687 141846 995696
rect 143460 995710 143764 995738
rect 143998 995752 144054 995761
rect 137374 995480 137430 995489
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994566 128492 995452
rect 128452 994560 128504 994566
rect 128452 994502 128504 994508
rect 129108 994294 129136 995452
rect 129752 994702 129780 995452
rect 129740 994696 129792 994702
rect 129740 994638 129792 994644
rect 131592 994430 131620 995452
rect 132144 994838 132172 995452
rect 132802 995438 133184 995466
rect 132132 994832 132184 994838
rect 132132 994774 132184 994780
rect 133156 994537 133184 995438
rect 133432 994809 133460 995452
rect 133418 994800 133474 994809
rect 133418 994735 133474 994744
rect 134892 994696 134944 994702
rect 134892 994638 134944 994644
rect 133142 994528 133198 994537
rect 133142 994463 133198 994472
rect 131580 994424 131632 994430
rect 131580 994366 131632 994372
rect 129096 994288 129148 994294
rect 129096 994230 129148 994236
rect 134904 994158 134932 994638
rect 135916 994265 135944 995452
rect 137126 995438 137374 995466
rect 137374 995415 137430 995424
rect 138952 994809 138980 995452
rect 140162 995438 140544 995466
rect 140516 995353 140544 995438
rect 140502 995344 140558 995353
rect 140502 995279 140558 995288
rect 138754 994800 138810 994809
rect 138754 994735 138810 994744
rect 138938 994800 138994 994809
rect 138938 994735 138994 994744
rect 135902 994256 135958 994265
rect 135902 994191 135958 994200
rect 134892 994152 134944 994158
rect 134892 994094 134944 994100
rect 138768 993993 138796 994735
rect 140792 994537 140820 995452
rect 142646 995438 143028 995466
rect 143000 995330 143028 995438
rect 143460 995330 143488 995710
rect 143998 995687 144054 995696
rect 143000 995302 143488 995330
rect 142988 994832 143040 994838
rect 142988 994774 143040 994780
rect 143172 994832 143224 994838
rect 144196 994809 144224 996338
rect 144380 995994 144408 997614
rect 144552 997076 144604 997082
rect 144552 997018 144604 997024
rect 144368 995988 144420 995994
rect 144368 995930 144420 995936
rect 143172 994774 143224 994780
rect 144182 994800 144238 994809
rect 140594 994528 140650 994537
rect 140594 994463 140650 994472
rect 140778 994528 140834 994537
rect 140778 994463 140834 994472
rect 138754 993984 138810 993993
rect 138754 993919 138810 993928
rect 140608 993721 140636 994463
rect 143000 994430 143028 994774
rect 142804 994424 142856 994430
rect 142804 994366 142856 994372
rect 142988 994424 143040 994430
rect 142988 994366 143040 994372
rect 142816 994022 142844 994366
rect 143184 994294 143212 994774
rect 144182 994735 144238 994744
rect 144564 994537 144592 997018
rect 144748 996033 144776 997726
rect 144734 996024 144790 996033
rect 144734 995959 144790 995968
rect 144918 995344 144974 995353
rect 144918 995279 144974 995288
rect 144550 994528 144606 994537
rect 144550 994463 144606 994472
rect 143172 994288 143224 994294
rect 143172 994230 143224 994236
rect 144932 994158 144960 995279
rect 144920 994152 144972 994158
rect 144920 994094 144972 994100
rect 142804 994016 142856 994022
rect 145576 993993 145604 1006742
rect 145748 1006664 145800 1006670
rect 145748 1006606 145800 1006612
rect 145760 996577 145788 1006606
rect 151268 1006528 151320 1006534
rect 151266 1006496 151268 1006505
rect 151740 1006505 151768 1006742
rect 369124 1006742 369176 1006748
rect 359370 1006703 359426 1006712
rect 360568 1006664 360620 1006670
rect 152094 1006632 152150 1006641
rect 152094 1006567 152096 1006576
rect 152148 1006567 152150 1006576
rect 157430 1006632 157486 1006641
rect 360566 1006632 360568 1006641
rect 360620 1006632 360622 1006641
rect 157430 1006567 157432 1006576
rect 152096 1006538 152148 1006544
rect 157484 1006567 157486 1006576
rect 166264 1006596 166316 1006602
rect 157432 1006538 157484 1006544
rect 360566 1006567 360622 1006576
rect 166264 1006538 166316 1006544
rect 151320 1006496 151322 1006505
rect 151266 1006431 151322 1006440
rect 151726 1006496 151782 1006505
rect 151726 1006431 151782 1006440
rect 158626 1006496 158682 1006505
rect 158626 1006431 158628 1006440
rect 158680 1006431 158682 1006440
rect 158628 1006402 158680 1006408
rect 148508 1006392 148560 1006398
rect 148508 1006334 148560 1006340
rect 158258 1006360 158314 1006369
rect 147126 1006088 147182 1006097
rect 147126 1006023 147182 1006032
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145746 996568 145802 996577
rect 145746 996503 145802 996512
rect 142804 993958 142856 993964
rect 145562 993984 145618 993993
rect 145562 993919 145618 993928
rect 140594 993712 140650 993721
rect 140594 993647 140650 993656
rect 138020 993064 138072 993070
rect 138020 993006 138072 993012
rect 138032 983634 138060 993006
rect 146956 991506 146984 1001914
rect 147140 1000657 147168 1006023
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 147126 1000648 147182 1000657
rect 147126 1000583 147182 1000592
rect 148336 992934 148364 1002050
rect 148520 994430 148548 1006334
rect 153936 1006324 153988 1006330
rect 158258 1006295 158260 1006304
rect 153936 1006266 153988 1006272
rect 158312 1006295 158314 1006304
rect 159454 1006360 159510 1006369
rect 159454 1006295 159456 1006304
rect 158260 1006266 158312 1006272
rect 159508 1006295 159510 1006304
rect 159456 1006266 159508 1006272
rect 150900 1006256 150952 1006262
rect 150898 1006224 150900 1006233
rect 150952 1006224 150954 1006233
rect 150898 1006159 150954 1006168
rect 153750 1006224 153806 1006233
rect 153750 1006159 153752 1006168
rect 153804 1006159 153806 1006168
rect 153752 1006130 153804 1006136
rect 148876 1006120 148928 1006126
rect 148874 1006088 148876 1006097
rect 150072 1006120 150124 1006126
rect 148928 1006088 148930 1006097
rect 148874 1006023 148930 1006032
rect 150070 1006088 150072 1006097
rect 150124 1006088 150126 1006097
rect 150070 1006023 150126 1006032
rect 152922 1005136 152978 1005145
rect 149704 1005100 149756 1005106
rect 152922 1005071 152924 1005080
rect 149704 1005042 149756 1005048
rect 152976 1005071 152978 1005080
rect 152924 1005042 152976 1005048
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 148508 994424 148560 994430
rect 148508 994366 148560 994372
rect 149716 993721 149744 1005042
rect 153750 1005000 153806 1005009
rect 151084 1004964 151136 1004970
rect 153750 1004935 153752 1004944
rect 151084 1004906 151136 1004912
rect 153804 1004935 153806 1004944
rect 153752 1004906 153804 1004912
rect 149888 1004828 149940 1004834
rect 149888 1004770 149940 1004776
rect 149900 996402 149928 1004770
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 149888 996396 149940 996402
rect 149888 996338 149940 996344
rect 151096 994022 151124 1004906
rect 152922 1004864 152978 1004873
rect 152922 1004799 152924 1004808
rect 152976 1004799 152978 1004808
rect 152924 1004770 152976 1004776
rect 151268 1004692 151320 1004698
rect 151268 1004634 151320 1004640
rect 151280 996538 151308 1004634
rect 152464 1002108 152516 1002114
rect 152464 1002050 152516 1002056
rect 151268 996532 151320 996538
rect 151268 996474 151320 996480
rect 152476 994265 152504 1002050
rect 153948 997626 153976 1006266
rect 160282 1006224 160338 1006233
rect 166276 1006194 166304 1006538
rect 255318 1006496 255374 1006505
rect 173164 1006460 173216 1006466
rect 173164 1006402 173216 1006408
rect 249248 1006460 249300 1006466
rect 255318 1006431 255320 1006440
rect 249248 1006402 249300 1006408
rect 255372 1006431 255374 1006440
rect 361394 1006496 361450 1006505
rect 361394 1006431 361396 1006440
rect 255320 1006402 255372 1006408
rect 361448 1006431 361450 1006440
rect 361396 1006402 361448 1006408
rect 160282 1006159 160284 1006168
rect 160336 1006159 160338 1006168
rect 164884 1006188 164936 1006194
rect 160284 1006130 160336 1006136
rect 164884 1006130 164936 1006136
rect 166264 1006188 166316 1006194
rect 166264 1006130 166316 1006136
rect 158258 1006088 158314 1006097
rect 158258 1006023 158260 1006032
rect 158312 1006023 158314 1006032
rect 158260 1005994 158312 1006000
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 160704 1004799 160706 1004808
rect 163136 1004828 163188 1004834
rect 160652 1004770 160704 1004776
rect 163136 1004770 163188 1004776
rect 154118 1004728 154174 1004737
rect 154118 1004663 154120 1004672
rect 154172 1004663 154174 1004672
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 154120 1004634 154172 1004640
rect 161164 1004663 161166 1004672
rect 162952 1004692 163004 1004698
rect 161112 1004634 161164 1004640
rect 162952 1004634 163004 1004640
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 158720 1002244 158772 1002250
rect 155776 1002186 155828 1002192
rect 158720 1002186 158772 1002192
rect 154578 1002144 154634 1002153
rect 154578 1002079 154580 1002088
rect 154632 1002079 154634 1002088
rect 154580 1002050 154632 1002056
rect 154946 1002008 155002 1002017
rect 154592 1001966 154946 1001994
rect 153936 997620 153988 997626
rect 153936 997562 153988 997568
rect 154302 995752 154358 995761
rect 154302 995687 154358 995696
rect 154316 995081 154344 995687
rect 154302 995072 154358 995081
rect 154302 995007 154358 995016
rect 154592 994566 154620 1001966
rect 154946 1001943 155002 1001952
rect 155774 1002008 155830 1002017
rect 156602 1002008 156658 1002017
rect 155774 1001943 155776 1001952
rect 155828 1001943 155830 1001952
rect 155972 1001966 156602 1001994
rect 155776 1001914 155828 1001920
rect 155972 994838 156000 1001966
rect 157798 1002008 157854 1002017
rect 156602 1001943 156658 1001952
rect 157340 1001972 157392 1001978
rect 157798 1001943 157800 1001952
rect 157340 1001914 157392 1001920
rect 157852 1001943 157854 1001952
rect 157800 1001914 157852 1001920
rect 155960 994832 156012 994838
rect 155960 994774 156012 994780
rect 157352 994702 157380 1001914
rect 158732 997082 158760 1002186
rect 160100 1001972 160152 1001978
rect 160100 1001914 160152 1001920
rect 160112 997762 160140 1001914
rect 160100 997756 160152 997762
rect 160100 997698 160152 997704
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 158720 997076 158772 997082
rect 158720 997018 158772 997024
rect 157340 994696 157392 994702
rect 157340 994638 157392 994644
rect 154580 994560 154632 994566
rect 154580 994502 154632 994508
rect 152462 994256 152518 994265
rect 152462 994191 152518 994200
rect 151084 994016 151136 994022
rect 151084 993958 151136 993964
rect 149702 993712 149758 993721
rect 149702 993647 149758 993656
rect 148324 992928 148376 992934
rect 148324 992870 148376 992876
rect 146944 991500 146996 991506
rect 146944 991442 146996 991448
rect 160756 985726 160784 997154
rect 163148 993070 163176 1004770
rect 164896 993478 164924 1006130
rect 171784 1006052 171836 1006058
rect 171784 1005994 171836 1006000
rect 171796 996130 171824 1005994
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 168748 995988 168800 995994
rect 168748 995930 168800 995936
rect 171508 995988 171560 995994
rect 171508 995930 171560 995936
rect 168564 995852 168616 995858
rect 168564 995794 168616 995800
rect 168576 994770 168604 995794
rect 168564 994764 168616 994770
rect 168564 994706 168616 994712
rect 168760 994634 168788 995930
rect 171232 995852 171284 995858
rect 171232 995794 171284 995800
rect 170680 995580 170732 995586
rect 170680 995522 170732 995528
rect 168930 995344 168986 995353
rect 168930 995279 168986 995288
rect 168748 994628 168800 994634
rect 168748 994570 168800 994576
rect 168944 994498 168972 995279
rect 170692 995081 170720 995522
rect 171244 995111 171272 995794
rect 171520 995223 171548 995930
rect 171690 995344 171746 995353
rect 171690 995279 171692 995288
rect 171744 995279 171746 995288
rect 171692 995271 171744 995277
rect 171508 995217 171560 995223
rect 171508 995159 171560 995165
rect 171232 995105 171284 995111
rect 169390 995072 169446 995081
rect 169390 995007 169446 995016
rect 170678 995072 170734 995081
rect 173176 995081 173204 1006402
rect 177304 1006324 177356 1006330
rect 177304 1006266 177356 1006272
rect 249064 1006324 249116 1006330
rect 249064 1006266 249116 1006272
rect 175924 1006188 175976 1006194
rect 175924 1006130 175976 1006136
rect 175936 995761 175964 1006130
rect 177316 995994 177344 1006266
rect 210422 1006224 210478 1006233
rect 210422 1006159 210424 1006168
rect 210476 1006159 210478 1006168
rect 228364 1006188 228416 1006194
rect 210424 1006130 210476 1006136
rect 228364 1006130 228416 1006136
rect 201038 1006088 201094 1006097
rect 198188 1006052 198240 1006058
rect 201038 1006023 201040 1006032
rect 198188 1005994 198240 1006000
rect 201092 1006023 201094 1006032
rect 208398 1006088 208454 1006097
rect 208398 1006023 208400 1006032
rect 201040 1005994 201092 1006000
rect 208452 1006023 208454 1006032
rect 208400 1005994 208452 1006000
rect 196624 999048 196676 999054
rect 196624 998990 196676 998996
rect 195058 998336 195114 998345
rect 195058 998271 195114 998280
rect 178866 996432 178922 996441
rect 178866 996367 178922 996376
rect 177304 995988 177356 995994
rect 177304 995930 177356 995936
rect 175922 995752 175978 995761
rect 175922 995687 175978 995696
rect 178880 995246 178908 996367
rect 195072 995761 195100 998271
rect 195244 997688 195296 997694
rect 195244 997630 195296 997636
rect 188066 995752 188122 995761
rect 187864 995710 188066 995738
rect 189446 995752 189502 995761
rect 189152 995710 189446 995738
rect 188066 995687 188122 995696
rect 191746 995752 191802 995761
rect 191544 995710 191746 995738
rect 189446 995687 189502 995696
rect 192482 995752 192538 995761
rect 192188 995710 192482 995738
rect 191746 995687 191802 995696
rect 194322 995752 194378 995761
rect 194028 995710 194322 995738
rect 192482 995687 192538 995696
rect 194322 995687 194378 995696
rect 195058 995752 195114 995761
rect 195058 995687 195114 995696
rect 194968 995580 195020 995586
rect 194968 995522 195020 995528
rect 183834 995480 183890 995489
rect 179860 995438 180196 995466
rect 178868 995240 178920 995246
rect 178868 995182 178920 995188
rect 180168 995110 180196 995438
rect 180490 995246 180518 995452
rect 181148 995438 181484 995466
rect 180708 995376 180760 995382
rect 180708 995318 180760 995324
rect 180340 995240 180392 995246
rect 180340 995182 180392 995188
rect 180478 995240 180530 995246
rect 180478 995182 180530 995188
rect 180156 995104 180208 995110
rect 171232 995047 171284 995053
rect 173162 995072 173218 995081
rect 170678 995007 170734 995016
rect 180156 995046 180208 995052
rect 173162 995007 173218 995016
rect 168932 994492 168984 994498
rect 168932 994434 168984 994440
rect 169404 994090 169432 995007
rect 171048 994881 171100 994887
rect 171048 994823 171100 994829
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 169392 994084 169444 994090
rect 169392 994026 169444 994032
rect 171060 993682 171088 994823
rect 171244 993818 171272 994823
rect 180352 994022 180380 995182
rect 180720 994974 180748 995318
rect 180708 994968 180760 994974
rect 180708 994910 180760 994916
rect 181456 994809 181484 995438
rect 182652 995438 182988 995466
rect 183540 995438 183834 995466
rect 182652 995382 182680 995438
rect 183834 995415 183890 995424
rect 184032 995438 184184 995466
rect 184828 995438 185164 995466
rect 187312 995438 187648 995466
rect 188508 995438 188844 995466
rect 190348 995438 190408 995466
rect 192832 995438 193168 995466
rect 182640 995376 182692 995382
rect 182640 995318 182692 995324
rect 183650 995344 183706 995353
rect 184032 995330 184060 995438
rect 185136 995382 185164 995438
rect 183706 995302 184060 995330
rect 185124 995376 185176 995382
rect 185124 995318 185176 995324
rect 186780 995376 186832 995382
rect 186780 995318 186832 995324
rect 183650 995279 183706 995288
rect 181442 994800 181498 994809
rect 181442 994735 181498 994744
rect 186792 994362 186820 995318
rect 187620 994537 187648 995438
rect 187606 994528 187662 994537
rect 187606 994463 187662 994472
rect 186780 994356 186832 994362
rect 186780 994298 186832 994304
rect 186504 994288 186556 994294
rect 186504 994230 186556 994236
rect 180340 994016 180392 994022
rect 180340 993958 180392 993964
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 171048 993676 171100 993682
rect 171048 993618 171100 993624
rect 164884 993472 164936 993478
rect 164884 993414 164936 993420
rect 169760 993472 169812 993478
rect 169760 993414 169812 993420
rect 163136 993064 163188 993070
rect 163136 993006 163188 993012
rect 169772 992234 169800 993414
rect 169772 992206 170352 992234
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 121748 983606 122130 983634
rect 138032 983606 138322 983634
rect 154500 983620 154528 985662
rect 170324 983634 170352 992206
rect 186516 983634 186544 994230
rect 188816 993993 188844 995438
rect 190380 994265 190408 995438
rect 193140 995382 193168 995438
rect 193128 995376 193180 995382
rect 193128 995318 193180 995324
rect 194980 994362 195008 995522
rect 194968 994356 195020 994362
rect 194968 994298 195020 994304
rect 190366 994256 190422 994265
rect 190366 994191 190422 994200
rect 188802 993984 188858 993993
rect 188802 993919 188858 993928
rect 195256 993818 195284 997630
rect 196636 994022 196664 998990
rect 197820 998640 197872 998646
rect 197820 998582 197872 998588
rect 197832 996985 197860 998582
rect 198004 998164 198056 998170
rect 198004 998106 198056 998112
rect 197818 996976 197874 996985
rect 197818 996911 197874 996920
rect 196624 994016 196676 994022
rect 196624 993958 196676 993964
rect 195244 993812 195296 993818
rect 195244 993754 195296 993760
rect 198016 993682 198044 998106
rect 198200 995382 198228 1005994
rect 204904 1005304 204956 1005310
rect 212080 1005304 212132 1005310
rect 204904 1005246 204956 1005252
rect 212078 1005272 212080 1005281
rect 212132 1005272 212134 1005281
rect 203524 1002244 203576 1002250
rect 203524 1002186 203576 1002192
rect 202972 1001972 203024 1001978
rect 202972 1001914 203024 1001920
rect 200764 998776 200816 998782
rect 200764 998718 200816 998724
rect 200212 998368 200264 998374
rect 200210 998336 200212 998345
rect 200264 998336 200266 998345
rect 200210 998271 200266 998280
rect 200776 998050 200804 998718
rect 202696 998640 202748 998646
rect 202694 998608 202696 998617
rect 202748 998608 202750 998617
rect 202694 998543 202750 998552
rect 200948 998504 201000 998510
rect 200948 998446 201000 998452
rect 199384 998028 199436 998034
rect 200776 998022 200896 998050
rect 199384 997970 199436 997976
rect 198372 997892 198424 997898
rect 198372 997834 198424 997840
rect 198384 997694 198412 997834
rect 198372 997688 198424 997694
rect 198372 997630 198424 997636
rect 199396 996033 199424 997970
rect 200670 997928 200726 997937
rect 200670 997863 200672 997872
rect 200724 997863 200726 997872
rect 200672 997834 200724 997840
rect 200868 997754 200896 998022
rect 200776 997726 200896 997754
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 199382 996024 199438 996033
rect 199382 995959 199438 995968
rect 198188 995376 198240 995382
rect 198188 995318 198240 995324
rect 200776 993993 200804 997726
rect 200960 994265 200988 998446
rect 202984 998374 203012 1001914
rect 202972 998368 203024 998374
rect 202972 998310 203024 998316
rect 201866 998200 201922 998209
rect 201866 998135 201868 998144
rect 201920 998135 201922 998144
rect 202144 998164 202196 998170
rect 201868 998106 201920 998112
rect 202144 998106 202196 998112
rect 201682 995616 201738 995625
rect 201682 995551 201684 995560
rect 201736 995551 201738 995560
rect 201684 995522 201736 995528
rect 202156 995246 202184 998106
rect 202694 998064 202750 998073
rect 202694 997999 202696 998008
rect 202748 997999 202750 998008
rect 202696 997970 202748 997976
rect 202328 997824 202380 997830
rect 202328 997766 202380 997772
rect 202340 995897 202368 997766
rect 202326 995888 202382 995897
rect 202326 995823 202382 995832
rect 202144 995240 202196 995246
rect 202144 995182 202196 995188
rect 203536 994537 203564 1002186
rect 204352 999048 204404 999054
rect 204350 999016 204352 999025
rect 204404 999016 204406 999025
rect 204350 998951 204406 998960
rect 203892 998776 203944 998782
rect 203890 998744 203892 998753
rect 203944 998744 203946 998753
rect 203890 998679 203946 998688
rect 203892 998504 203944 998510
rect 203890 998472 203892 998481
rect 203944 998472 203946 998481
rect 203890 998407 203946 998416
rect 204720 997824 204772 997830
rect 204718 997792 204720 997801
rect 204772 997792 204774 997801
rect 204718 997727 204774 997736
rect 203522 994528 203578 994537
rect 203522 994463 203578 994472
rect 200946 994256 201002 994265
rect 200946 994191 201002 994200
rect 200762 993984 200818 993993
rect 200762 993919 200818 993928
rect 198004 993676 198056 993682
rect 198004 993618 198056 993624
rect 204916 986678 204944 1005246
rect 212078 1005207 212134 1005216
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 211250 1004864 211306 1004873
rect 211250 1004799 211252 1004808
rect 211304 1004799 211306 1004808
rect 211252 1004770 211304 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 211160 1004692 211212 1004698
rect 209228 1004634 209280 1004640
rect 211160 1004634 211212 1004640
rect 206374 1002280 206430 1002289
rect 206374 1002215 206376 1002224
rect 206428 1002215 206430 1002224
rect 206742 1002280 206798 1002289
rect 210882 1002280 210938 1002289
rect 206742 1002215 206744 1002224
rect 206376 1002186 206428 1002192
rect 206796 1002215 206798 1002224
rect 208400 1002244 208452 1002250
rect 206744 1002186 206796 1002192
rect 210882 1002215 210884 1002224
rect 208400 1002186 208452 1002192
rect 210936 1002215 210938 1002224
rect 210884 1002186 210936 1002192
rect 207202 1002144 207258 1002153
rect 205088 1002108 205140 1002114
rect 207202 1002079 207204 1002088
rect 205088 1002050 205140 1002056
rect 207256 1002079 207258 1002088
rect 207204 1002050 207256 1002056
rect 205100 997286 205128 1002050
rect 205546 1002008 205602 1002017
rect 206742 1002008 206798 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 206296 1001966 206742 1001994
rect 205548 1001914 205600 1001920
rect 205546 998200 205602 998209
rect 205546 998135 205548 998144
rect 205600 998135 205602 998144
rect 205548 998106 205600 998112
rect 205088 997280 205140 997286
rect 205088 997222 205140 997228
rect 206296 995110 206324 1001966
rect 207570 1002008 207626 1002017
rect 206742 1001943 206798 1001952
rect 207032 1001966 207570 1001994
rect 206284 995104 206336 995110
rect 206284 995046 206336 995052
rect 207032 994809 207060 1001966
rect 207570 1001943 207626 1001952
rect 208412 994974 208440 1002186
rect 210882 1002008 210938 1002017
rect 210882 1001943 210884 1001952
rect 210936 1001943 210938 1001952
rect 210884 1001914 210936 1001920
rect 211172 996130 211200 1004634
rect 211816 996130 211844 1004906
rect 215944 1004828 215996 1004834
rect 215944 1004770 215996 1004776
rect 213184 1002244 213236 1002250
rect 213184 1002186 213236 1002192
rect 212538 1002144 212594 1002153
rect 212538 1002079 212540 1002088
rect 212592 1002079 212594 1002088
rect 212540 1002050 212592 1002056
rect 212540 1001972 212592 1001978
rect 212540 1001914 212592 1001920
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211804 996124 211856 996130
rect 211804 996066 211856 996072
rect 212552 995994 212580 1001914
rect 212540 995988 212592 995994
rect 212540 995930 212592 995936
rect 213196 995858 213224 1002186
rect 214564 1002108 214616 1002114
rect 214564 1002050 214616 1002056
rect 213184 995852 213236 995858
rect 213184 995794 213236 995800
rect 208400 994968 208452 994974
rect 208400 994910 208452 994916
rect 207018 994800 207074 994809
rect 207018 994735 207074 994744
rect 214576 993478 214604 1002050
rect 214564 993472 214616 993478
rect 214564 993414 214616 993420
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 204904 986672 204956 986678
rect 204904 986614 204956 986620
rect 170324 983606 170798 983634
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1004770
rect 228376 995382 228404 1006130
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 229756 995994 229784 1005994
rect 247224 998572 247276 998578
rect 247224 998514 247276 998520
rect 247040 998300 247092 998306
rect 247040 998242 247092 998248
rect 246764 998164 246816 998170
rect 246764 998106 246816 998112
rect 246580 997756 246632 997762
rect 246580 997698 246632 997704
rect 246592 996441 246620 997698
rect 246578 996432 246634 996441
rect 246578 996367 246634 996376
rect 229744 995988 229796 995994
rect 229744 995930 229796 995936
rect 240874 995752 240930 995761
rect 240580 995710 240874 995738
rect 240874 995687 240930 995696
rect 236550 995616 236606 995625
rect 236256 995574 236550 995602
rect 236550 995551 236606 995560
rect 246212 995512 246264 995518
rect 242070 995480 242126 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 234416 995438 234568 995466
rect 234968 995438 235304 995466
rect 228364 995376 228416 995382
rect 228364 995318 228416 995324
rect 231596 994809 231624 995438
rect 231582 994800 231638 994809
rect 231582 994735 231638 994744
rect 232240 994362 232268 995438
rect 232884 994974 232912 995438
rect 232872 994968 232924 994974
rect 232872 994910 232924 994916
rect 232228 994356 232280 994362
rect 232228 994298 232280 994304
rect 234540 993993 234568 995438
rect 235276 995110 235304 995438
rect 235598 995246 235626 995452
rect 238588 995438 238740 995466
rect 239292 995438 239628 995466
rect 238588 995353 238616 995438
rect 238574 995344 238630 995353
rect 238574 995279 238630 995288
rect 235586 995240 235638 995246
rect 235586 995182 235638 995188
rect 235264 995104 235316 995110
rect 235264 995046 235316 995052
rect 234526 993984 234582 993993
rect 234526 993919 234582 993928
rect 239600 993721 239628 995438
rect 239922 995217 239950 995452
rect 241776 995438 242070 995466
rect 242972 995438 243308 995466
rect 243616 995438 243952 995466
rect 242070 995415 242126 995424
rect 239908 995208 239964 995217
rect 239908 995143 239964 995152
rect 243084 994628 243136 994634
rect 243084 994570 243136 994576
rect 243096 993886 243124 994570
rect 243280 994537 243308 995438
rect 243266 994528 243322 994537
rect 243266 994463 243322 994472
rect 243542 994528 243598 994537
rect 243542 994463 243598 994472
rect 243556 993993 243584 994463
rect 243924 994022 243952 995438
rect 244200 995438 244260 995466
rect 245456 995438 245884 995466
rect 246212 995454 246264 995460
rect 244200 994634 244228 995438
rect 245856 995330 245884 995438
rect 246224 995330 246252 995454
rect 245856 995302 246252 995330
rect 246776 994634 246804 998106
rect 247052 995761 247080 998242
rect 247038 995752 247094 995761
rect 247038 995687 247094 995696
rect 247236 995518 247264 998514
rect 247408 998436 247460 998442
rect 247408 998378 247460 998384
rect 247224 995512 247276 995518
rect 247224 995454 247276 995460
rect 244188 994628 244240 994634
rect 244188 994570 244240 994576
rect 246764 994628 246816 994634
rect 246764 994570 246816 994576
rect 247420 994022 247448 998378
rect 247684 997892 247736 997898
rect 247684 997834 247736 997840
rect 243912 994016 243964 994022
rect 243542 993984 243598 993993
rect 243912 993958 243964 993964
rect 247408 994016 247460 994022
rect 247408 993958 247460 993964
rect 243542 993919 243598 993928
rect 247696 993886 247724 997834
rect 248142 996024 248198 996033
rect 248142 995959 248198 995968
rect 248156 995058 248184 995959
rect 248326 995072 248382 995081
rect 248156 995030 248326 995058
rect 248326 995007 248382 995016
rect 249076 993993 249104 1006266
rect 249260 996033 249288 1006402
rect 254122 1006360 254178 1006369
rect 306930 1006360 306986 1006369
rect 254122 1006295 254124 1006304
rect 254176 1006295 254178 1006304
rect 301504 1006324 301556 1006330
rect 254124 1006266 254176 1006272
rect 306930 1006295 306932 1006304
rect 301504 1006266 301556 1006272
rect 306984 1006295 306986 1006304
rect 314658 1006360 314714 1006369
rect 369136 1006330 369164 1006742
rect 371884 1006664 371936 1006670
rect 371884 1006606 371936 1006612
rect 314658 1006295 314660 1006304
rect 306932 1006266 306984 1006272
rect 314712 1006295 314714 1006304
rect 319444 1006324 319496 1006330
rect 314660 1006266 314712 1006272
rect 319444 1006266 319496 1006272
rect 354864 1006324 354916 1006330
rect 354864 1006266 354916 1006272
rect 369124 1006324 369176 1006330
rect 369124 1006266 369176 1006272
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 262732 1006159 262734 1006168
rect 279424 1006188 279476 1006194
rect 262680 1006130 262732 1006136
rect 279424 1006130 279476 1006136
rect 298744 1006188 298796 1006194
rect 298744 1006130 298796 1006136
rect 252466 1006088 252522 1006097
rect 251088 1006052 251140 1006058
rect 252466 1006023 252468 1006032
rect 251088 1005994 251140 1006000
rect 252520 1006023 252522 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 252468 1005994 252520 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 251100 998170 251128 1005994
rect 263046 1005000 263102 1005009
rect 263046 1004935 263048 1004944
rect 263100 1004935 263102 1004944
rect 268384 1004964 268436 1004970
rect 263048 1004906 263100 1004912
rect 268384 1004906 268436 1004912
rect 256146 1002688 256202 1002697
rect 253480 1002652 253532 1002658
rect 256146 1002623 256148 1002632
rect 253480 1002594 253532 1002600
rect 256200 1002623 256202 1002632
rect 256148 1002594 256200 1002600
rect 252008 1002516 252060 1002522
rect 252008 1002458 252060 1002464
rect 251824 1002244 251876 1002250
rect 251824 1002186 251876 1002192
rect 251088 998164 251140 998170
rect 251088 998106 251140 998112
rect 250444 998028 250496 998034
rect 250444 997970 250496 997976
rect 249246 996024 249302 996033
rect 249246 995959 249302 995968
rect 250456 994770 250484 997970
rect 251836 995081 251864 1002186
rect 252020 995353 252048 1002458
rect 253020 1002380 253072 1002386
rect 253020 1002322 253072 1002328
rect 252466 997928 252522 997937
rect 252466 997863 252468 997872
rect 252520 997863 252522 997872
rect 252468 997834 252520 997840
rect 252006 995344 252062 995353
rect 252006 995279 252062 995288
rect 253032 995246 253060 1002322
rect 253294 998064 253350 998073
rect 253294 997999 253296 998008
rect 253348 997999 253350 998008
rect 253296 997970 253348 997976
rect 253204 996260 253256 996266
rect 253204 996202 253256 996208
rect 253216 995382 253244 996202
rect 253204 995376 253256 995382
rect 253204 995318 253256 995324
rect 253020 995240 253072 995246
rect 253020 995182 253072 995188
rect 253492 995110 253520 1002594
rect 255318 1002552 255374 1002561
rect 255318 1002487 255320 1002496
rect 255372 1002487 255374 1002496
rect 261022 1002552 261078 1002561
rect 261022 1002487 261024 1002496
rect 255320 1002458 255372 1002464
rect 261076 1002487 261078 1002496
rect 264244 1002516 264296 1002522
rect 261024 1002458 261076 1002464
rect 264244 1002458 264296 1002464
rect 256146 1002416 256202 1002425
rect 256146 1002351 256148 1002360
rect 256200 1002351 256202 1002360
rect 256148 1002322 256200 1002328
rect 254490 1002280 254546 1002289
rect 254490 1002215 254492 1002224
rect 254544 1002215 254546 1002224
rect 254492 1002186 254544 1002192
rect 263506 1002144 263562 1002153
rect 263506 1002079 263508 1002088
rect 263560 1002079 263562 1002088
rect 263508 1002050 263560 1002056
rect 261022 1002008 261078 1002017
rect 263874 1002008 263930 1002017
rect 261022 1001943 261024 1001952
rect 261076 1001943 261078 1001952
rect 263600 1001972 263652 1001978
rect 261024 1001914 261076 1001920
rect 263874 1001943 263876 1001952
rect 263600 1001914 263652 1001920
rect 263928 1001943 263930 1001952
rect 263876 1001914 263928 1001920
rect 256974 998608 257030 998617
rect 256974 998543 256976 998552
rect 257028 998543 257030 998552
rect 256976 998514 257028 998520
rect 258998 998472 259054 998481
rect 258998 998407 259000 998416
rect 259052 998407 259054 998416
rect 259000 998378 259052 998384
rect 253662 998336 253718 998345
rect 253662 998271 253664 998280
rect 253716 998271 253718 998280
rect 253664 998242 253716 998248
rect 258170 998200 258226 998209
rect 258170 998135 258172 998144
rect 258224 998135 258226 998144
rect 259460 998164 259512 998170
rect 258172 998106 258224 998112
rect 259460 998106 259512 998112
rect 256514 998064 256570 998073
rect 254584 998028 254636 998034
rect 256514 997999 256516 998008
rect 254584 997970 254636 997976
rect 256568 997999 256570 998008
rect 256516 997970 256568 997976
rect 253480 995104 253532 995110
rect 251822 995072 251878 995081
rect 253480 995046 253532 995052
rect 251822 995007 251878 995016
rect 250444 994764 250496 994770
rect 250444 994706 250496 994712
rect 254596 994362 254624 997970
rect 257342 997928 257398 997937
rect 256332 997892 256384 997898
rect 257342 997863 257344 997872
rect 256332 997834 256384 997840
rect 257396 997863 257398 997872
rect 257344 997834 257396 997840
rect 256344 997762 256372 997834
rect 256332 997756 256384 997762
rect 256332 997698 256384 997704
rect 255412 995852 255464 995858
rect 255412 995794 255464 995800
rect 255424 995586 255452 995794
rect 255778 995616 255834 995625
rect 255412 995580 255464 995586
rect 255778 995551 255834 995560
rect 255412 995522 255464 995528
rect 255792 994809 255820 995551
rect 256054 995344 256110 995353
rect 256054 995279 256110 995288
rect 256068 994974 256096 995279
rect 256056 994968 256108 994974
rect 256056 994910 256108 994916
rect 255778 994800 255834 994809
rect 255778 994735 255834 994744
rect 259472 994537 259500 998106
rect 260196 998096 260248 998102
rect 260194 998064 260196 998073
rect 262864 998096 262916 998102
rect 260248 998064 260250 998073
rect 262864 998038 262916 998044
rect 260194 997999 260250 998008
rect 259828 997960 259880 997966
rect 259826 997928 259828 997937
rect 262220 997960 262272 997966
rect 259880 997928 259882 997937
rect 262220 997902 262272 997908
rect 259826 997863 259882 997872
rect 260196 997824 260248 997830
rect 260194 997792 260196 997801
rect 260932 997824 260984 997830
rect 260248 997792 260250 997801
rect 260932 997766 260984 997772
rect 261850 997792 261906 997801
rect 260194 997727 260250 997736
rect 260944 996130 260972 997766
rect 261850 997727 261906 997736
rect 260932 996124 260984 996130
rect 260932 996066 260984 996072
rect 261864 995586 261892 997727
rect 262232 995858 262260 997902
rect 262876 995858 262904 998038
rect 263612 996266 263640 1001914
rect 263600 996260 263652 996266
rect 263600 996202 263652 996208
rect 264256 995994 264284 1002458
rect 265624 1002108 265676 1002114
rect 265624 1002050 265676 1002056
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 262220 995852 262272 995858
rect 262220 995794 262272 995800
rect 262864 995852 262916 995858
rect 262864 995794 262916 995800
rect 261852 995580 261904 995586
rect 261852 995522 261904 995528
rect 259458 994528 259514 994537
rect 259458 994463 259514 994472
rect 254584 994356 254636 994362
rect 254584 994298 254636 994304
rect 251454 994256 251510 994265
rect 251454 994191 251510 994200
rect 249062 993984 249118 993993
rect 249062 993919 249118 993928
rect 243084 993880 243136 993886
rect 243084 993822 243136 993828
rect 247684 993880 247736 993886
rect 247684 993822 247736 993828
rect 239586 993712 239642 993721
rect 239586 993647 239642 993656
rect 219440 993472 219492 993478
rect 219440 993414 219492 993420
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 993414
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 994191
rect 265636 990894 265664 1002050
rect 267004 1001972 267056 1001978
rect 267004 1001914 267056 1001920
rect 267016 991506 267044 1001914
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1004906
rect 279436 996130 279464 1006130
rect 280804 1006052 280856 1006058
rect 280804 1005994 280856 1006000
rect 279424 996124 279476 996130
rect 279424 996066 279476 996072
rect 280816 995081 280844 1005994
rect 298100 1000544 298152 1000550
rect 298100 1000486 298152 1000492
rect 287978 995752 288034 995761
rect 287822 995710 287978 995738
rect 290554 995752 290610 995761
rect 290306 995710 290554 995738
rect 287978 995687 288034 995696
rect 291106 995752 291162 995761
rect 290858 995710 291106 995738
rect 290554 995687 290610 995696
rect 293590 995752 293646 995761
rect 293342 995710 293590 995738
rect 291106 995687 291162 995696
rect 298112 995738 298140 1000486
rect 298282 997248 298338 997257
rect 298282 997183 298338 997192
rect 293590 995687 293646 995696
rect 297836 995710 298140 995738
rect 282840 995110 282868 995452
rect 282828 995104 282880 995110
rect 280802 995072 280858 995081
rect 282828 995046 282880 995052
rect 280802 995007 280858 995016
rect 283484 994974 283512 995452
rect 283472 994968 283524 994974
rect 283472 994910 283524 994916
rect 284128 994702 284156 995452
rect 285968 994809 285996 995452
rect 286520 994838 286548 995452
rect 286508 994832 286560 994838
rect 285954 994800 286010 994809
rect 286508 994774 286560 994780
rect 285954 994735 286010 994744
rect 284116 994696 284168 994702
rect 284116 994638 284168 994644
rect 287164 994537 287192 995452
rect 291502 995438 291792 995466
rect 291764 995353 291792 995438
rect 291948 995438 292146 995466
rect 294538 995438 295104 995466
rect 295182 995438 295564 995466
rect 295826 995438 296208 995466
rect 297022 995438 297404 995466
rect 291382 995344 291438 995353
rect 291750 995344 291806 995353
rect 291438 995302 291608 995330
rect 291382 995279 291438 995288
rect 291580 995194 291608 995302
rect 291750 995279 291806 995288
rect 291948 995194 291976 995438
rect 291580 995166 291976 995194
rect 295076 995058 295104 995438
rect 295076 995030 295380 995058
rect 287150 994528 287206 994537
rect 287150 994463 287206 994472
rect 295352 994294 295380 995030
rect 295340 994288 295392 994294
rect 295340 994230 295392 994236
rect 295536 993993 295564 995438
rect 296180 995382 296208 995438
rect 296168 995376 296220 995382
rect 296168 995318 296220 995324
rect 297376 995330 297404 995438
rect 297836 995330 297864 995710
rect 298296 995382 298324 997183
rect 297376 995302 297864 995330
rect 298284 995376 298336 995382
rect 298284 995318 298336 995324
rect 298756 994498 298784 1006130
rect 298928 1006052 298980 1006058
rect 298928 1005994 298980 1006000
rect 298940 995994 298968 1005994
rect 300308 1002108 300360 1002114
rect 300308 1002050 300360 1002056
rect 300320 996713 300348 1002050
rect 300306 996704 300362 996713
rect 300306 996639 300362 996648
rect 298928 995988 298980 995994
rect 298928 995930 298980 995936
rect 299570 995752 299626 995761
rect 299570 995687 299626 995696
rect 299584 995586 299612 995687
rect 299572 995580 299624 995586
rect 299572 995522 299624 995528
rect 300124 995444 300176 995450
rect 300124 995386 300176 995392
rect 298744 994492 298796 994498
rect 298744 994434 298796 994440
rect 300136 994158 300164 995386
rect 301516 995353 301544 1006266
rect 304906 1006224 304962 1006233
rect 304906 1006159 304908 1006168
rect 304960 1006159 304962 1006168
rect 304908 1006130 304960 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 304078 1006088 304134 1006097
rect 303306 1006046 304078 1006074
rect 303250 1006023 303306 1006032
rect 304078 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311808 1006032
rect 301700 997257 301728 1006023
rect 311860 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 314658 1006023 314660 1006032
rect 311808 1005994 311860 1006000
rect 314712 1006023 314714 1006032
rect 314660 1005994 314712 1006000
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 305274 1002144 305330 1002153
rect 305274 1002079 305276 1002088
rect 305328 1002079 305330 1002088
rect 310150 1002144 310206 1002153
rect 310150 1002079 310152 1002088
rect 305276 1002050 305328 1002056
rect 310204 1002079 310206 1002088
rect 311900 1002108 311952 1002114
rect 310152 1002050 310204 1002056
rect 311900 1002050 311952 1002056
rect 310978 1002008 311034 1002017
rect 310978 1001943 310980 1001952
rect 311032 1001943 311034 1001952
rect 310980 1001914 311032 1001920
rect 308956 1000544 309008 1000550
rect 308954 1000512 308956 1000521
rect 309008 1000512 309010 1000521
rect 308954 1000447 309010 1000456
rect 304264 998504 304316 998510
rect 307300 998504 307352 998510
rect 304264 998446 304316 998452
rect 307298 998472 307300 998481
rect 307352 998472 307354 998481
rect 303068 998368 303120 998374
rect 303068 998310 303120 998316
rect 302884 997824 302936 997830
rect 302884 997766 302936 997772
rect 301686 997248 301742 997257
rect 301686 997183 301742 997192
rect 302896 995625 302924 997766
rect 303080 996985 303108 998310
rect 303066 996976 303122 996985
rect 303066 996911 303122 996920
rect 304078 996160 304134 996169
rect 304078 996095 304134 996104
rect 302882 995616 302938 995625
rect 301688 995580 301740 995586
rect 302882 995551 302938 995560
rect 301688 995522 301740 995528
rect 301700 995353 301728 995522
rect 304092 995450 304120 996095
rect 304080 995444 304132 995450
rect 304080 995386 304132 995392
rect 301502 995344 301558 995353
rect 301502 995279 301558 995288
rect 301686 995344 301742 995353
rect 301686 995279 301742 995288
rect 304276 994537 304304 998446
rect 307298 998407 307354 998416
rect 306104 998368 306156 998374
rect 306102 998336 306104 998345
rect 306156 998336 306158 998345
rect 306102 998271 306158 998280
rect 304448 998232 304500 998238
rect 306932 998232 306984 998238
rect 304448 998174 304500 998180
rect 306930 998200 306932 998209
rect 306984 998200 306986 998209
rect 304460 995353 304488 998174
rect 306930 998135 306986 998144
rect 305644 998096 305696 998102
rect 307760 998096 307812 998102
rect 305644 998038 305696 998044
rect 307758 998064 307760 998073
rect 308404 998096 308456 998102
rect 307812 998064 307814 998073
rect 304446 995344 304502 995353
rect 304446 995279 304502 995288
rect 305656 994838 305684 998038
rect 310612 998096 310664 998102
rect 308404 998038 308456 998044
rect 310610 998064 310612 998073
rect 310664 998064 310666 998073
rect 307758 997999 307814 998008
rect 307208 997960 307260 997966
rect 307208 997902 307260 997908
rect 306104 997824 306156 997830
rect 306102 997792 306104 997801
rect 307024 997824 307076 997830
rect 306156 997792 306158 997801
rect 307024 997766 307076 997772
rect 306102 997727 306158 997736
rect 307036 994974 307064 997766
rect 307220 995353 307248 997902
rect 308128 997824 308180 997830
rect 308126 997792 308128 997801
rect 308180 997792 308182 997801
rect 308126 997727 308182 997736
rect 307206 995344 307262 995353
rect 307206 995279 307262 995288
rect 307024 994968 307076 994974
rect 307024 994910 307076 994916
rect 305644 994832 305696 994838
rect 305644 994774 305696 994780
rect 308416 994702 308444 998038
rect 310610 997999 310666 998008
rect 308956 997960 309008 997966
rect 308954 997928 308956 997937
rect 309008 997928 309010 997937
rect 308954 997863 309010 997872
rect 309782 997792 309838 997801
rect 309152 997736 309782 997754
rect 310610 997792 310666 997801
rect 309152 997727 309838 997736
rect 310532 997736 310610 997754
rect 310532 997727 310666 997736
rect 309152 997726 309824 997727
rect 310532 997726 310652 997727
rect 309152 994809 309180 997726
rect 309138 994800 309194 994809
rect 309138 994735 309194 994744
rect 308404 994696 308456 994702
rect 308404 994638 308456 994644
rect 304262 994528 304318 994537
rect 304262 994463 304318 994472
rect 300124 994152 300176 994158
rect 300124 994094 300176 994100
rect 310532 993993 310560 997726
rect 311912 995110 311940 1002050
rect 313280 1001972 313332 1001978
rect 313280 1001914 313332 1001920
rect 313292 995858 313320 1001914
rect 316052 996130 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 313280 995852 313332 995858
rect 313280 995794 313332 995800
rect 311900 995104 311952 995110
rect 311900 995046 311952 995052
rect 316406 994256 316462 994265
rect 316406 994191 316462 994200
rect 295522 993984 295578 993993
rect 295522 993919 295578 993928
rect 310518 993984 310574 993993
rect 310518 993919 310574 993928
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994191
rect 318076 993070 318104 1004634
rect 318064 993064 318116 993070
rect 318064 993006 318116 993012
rect 319456 992934 319484 1006266
rect 354876 1006097 354904 1006266
rect 355690 1006224 355746 1006233
rect 365074 1006224 365130 1006233
rect 355690 1006159 355692 1006168
rect 355744 1006159 355746 1006168
rect 363604 1006188 363656 1006194
rect 355692 1006130 355744 1006136
rect 365074 1006159 365076 1006168
rect 363604 1006130 363656 1006136
rect 365128 1006159 365130 1006168
rect 367744 1006188 367796 1006194
rect 365076 1006130 365128 1006136
rect 367744 1006130 367796 1006136
rect 354862 1006088 354918 1006097
rect 320824 1006052 320876 1006058
rect 354862 1006023 354918 1006032
rect 363418 1006088 363474 1006097
rect 363418 1006023 363420 1006032
rect 320824 1005994 320876 1006000
rect 363472 1006023 363474 1006032
rect 363420 1005994 363472 1006000
rect 320836 997082 320864 1005994
rect 360568 1005440 360620 1005446
rect 360566 1005408 360568 1005417
rect 360620 1005408 360622 1005417
rect 360566 1005343 360622 1005352
rect 357716 1005304 357768 1005310
rect 357714 1005272 357716 1005281
rect 357768 1005272 357770 1005281
rect 357714 1005207 357770 1005216
rect 356518 1005136 356574 1005145
rect 354588 1005100 354640 1005106
rect 356518 1005071 356520 1005080
rect 354588 1005042 354640 1005048
rect 356572 1005071 356574 1005080
rect 356520 1005042 356572 1005048
rect 353208 1004964 353260 1004970
rect 353208 1004906 353260 1004912
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998442 351868 1001914
rect 353220 1001230 353248 1004906
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998436 351880 998442
rect 351828 998378 351880 998384
rect 320824 997076 320876 997082
rect 320824 997018 320876 997024
rect 332600 997076 332652 997082
rect 332600 997018 332652 997024
rect 319444 992928 319496 992934
rect 319444 992870 319496 992876
rect 332612 983634 332640 997018
rect 354600 996130 354628 1005042
rect 355690 1005000 355746 1005009
rect 355690 1004935 355692 1004944
rect 355744 1004935 355746 1004944
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 355692 1004906 355744 1004912
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 358542 1002280 358598 1002289
rect 358542 1002215 358544 1002224
rect 358596 1002215 358598 1002224
rect 360844 1002244 360896 1002250
rect 358544 1002186 358596 1002192
rect 360844 1002186 360896 1002192
rect 356518 1002144 356574 1002153
rect 355784 1002108 355836 1002114
rect 356518 1002079 356520 1002088
rect 355784 1002050 355836 1002056
rect 356572 1002079 356574 1002088
rect 356520 1002050 356572 1002056
rect 354588 996124 354640 996130
rect 354588 996066 354640 996072
rect 355796 995858 355824 1002050
rect 356886 1002008 356942 1002017
rect 356072 1001966 356886 1001994
rect 355784 995852 355836 995858
rect 355784 995794 355836 995800
rect 356072 994634 356100 1001966
rect 357714 1002008 357770 1002017
rect 356886 1001943 356942 1001952
rect 357452 1001966 357714 1001994
rect 357452 995042 357480 1001966
rect 357714 1001943 357770 1001952
rect 358542 1002008 358598 1002017
rect 360198 1002008 360254 1002017
rect 358598 1001966 359504 1001994
rect 358542 1001943 358598 1001952
rect 359476 997762 359504 1001966
rect 360198 1001943 360200 1001952
rect 360252 1001943 360254 1001952
rect 360200 1001914 360252 1001920
rect 360856 999802 360884 1002186
rect 362224 1001972 362276 1001978
rect 362224 1001914 362276 1001920
rect 360844 999796 360896 999802
rect 360844 999738 360896 999744
rect 359464 997756 359516 997762
rect 359464 997698 359516 997704
rect 362236 995178 362264 1001914
rect 362224 995172 362276 995178
rect 362224 995114 362276 995120
rect 357440 995036 357492 995042
rect 357440 994978 357492 994984
rect 363616 994770 363644 1006130
rect 365074 1005136 365130 1005145
rect 365074 1005071 365076 1005080
rect 365128 1005071 365130 1005080
rect 365076 1005042 365128 1005048
rect 364984 1004964 365036 1004970
rect 364984 1004906 365036 1004912
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 364996 995586 365024 1004906
rect 365168 1004828 365220 1004834
rect 365168 1004770 365220 1004776
rect 365180 997014 365208 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365168 997008 365220 997014
rect 365168 996950 365220 996956
rect 366376 996130 366404 1004634
rect 366364 996124 366416 996130
rect 366364 996066 366416 996072
rect 364984 995580 365036 995586
rect 364984 995522 365036 995528
rect 363604 994764 363656 994770
rect 363604 994706 363656 994712
rect 356060 994628 356112 994634
rect 356060 994570 356112 994576
rect 349160 993064 349212 993070
rect 349160 993006 349212 993012
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 993006
rect 367756 992934 367784 1006130
rect 370504 1005100 370556 1005106
rect 370504 1005042 370556 1005048
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 368940 996260 368992 996266
rect 368940 996202 368992 996208
rect 368952 995858 368980 996202
rect 368940 995852 368992 995858
rect 368940 995794 368992 995800
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 367744 992928 367796 992934
rect 367744 992870 367796 992876
rect 364996 983634 365024 992870
rect 369136 991506 369164 1001914
rect 369860 999796 369912 999802
rect 369860 999738 369912 999744
rect 369872 997626 369900 999738
rect 369860 997620 369912 997626
rect 369860 997562 369912 997568
rect 369308 995852 369360 995858
rect 369308 995794 369360 995800
rect 369320 995586 369348 995794
rect 369308 995580 369360 995586
rect 369308 995522 369360 995528
rect 369124 991500 369176 991506
rect 369124 991442 369176 991448
rect 370516 985998 370544 1005042
rect 371896 994906 371924 1006606
rect 373264 1006188 373316 1006194
rect 373264 1006130 373316 1006136
rect 373276 999122 373304 1006130
rect 374656 1001894 374684 1006878
rect 428370 1006839 428372 1006848
rect 428424 1006839 428426 1006848
rect 428372 1006810 428424 1006816
rect 429198 1006768 429254 1006777
rect 429198 1006703 429200 1006712
rect 429252 1006703 429254 1006712
rect 429200 1006674 429252 1006680
rect 376760 1006460 376812 1006466
rect 376760 1006402 376812 1006408
rect 422668 1006460 422720 1006466
rect 422668 1006402 422720 1006408
rect 375380 1005304 375432 1005310
rect 375380 1005246 375432 1005252
rect 374656 1001866 374868 1001894
rect 373264 999116 373316 999122
rect 373264 999058 373316 999064
rect 374644 999116 374696 999122
rect 374644 999058 374696 999064
rect 372344 997756 372396 997762
rect 372344 997698 372396 997704
rect 372356 996441 372384 997698
rect 372528 997620 372580 997626
rect 372528 997562 372580 997568
rect 372540 996713 372568 997562
rect 372712 997008 372764 997014
rect 372710 996976 372712 996985
rect 372764 996976 372766 996985
rect 372710 996911 372766 996920
rect 372526 996704 372582 996713
rect 372526 996639 372582 996648
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 374656 995314 374684 999058
rect 374644 995308 374696 995314
rect 374644 995250 374696 995256
rect 371884 994900 371936 994906
rect 371884 994842 371936 994848
rect 374840 994809 374868 1001866
rect 375392 1000550 375420 1005246
rect 375380 1000544 375432 1000550
rect 375380 1000486 375432 1000492
rect 376772 998646 376800 1006402
rect 380164 1006324 380216 1006330
rect 380164 1006266 380216 1006272
rect 378784 1005440 378836 1005446
rect 378784 1005382 378836 1005388
rect 378796 998782 378824 1005382
rect 378784 998776 378836 998782
rect 378784 998718 378836 998724
rect 376760 998640 376812 998646
rect 376760 998582 376812 998588
rect 377588 996260 377640 996266
rect 377588 996202 377640 996208
rect 377600 995586 377628 996202
rect 380176 995586 380204 1006266
rect 402244 1006188 402296 1006194
rect 402244 1006130 402296 1006136
rect 382924 1006052 382976 1006058
rect 382924 1005994 382976 1006000
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 377588 995580 377640 995586
rect 377588 995522 377640 995528
rect 380164 995580 380216 995586
rect 380164 995522 380216 995528
rect 380912 995217 380940 1001166
rect 382280 998436 382332 998442
rect 382280 998378 382332 998384
rect 382094 997248 382150 997257
rect 382094 997183 382150 997192
rect 382108 996441 382136 997183
rect 382094 996432 382150 996441
rect 382094 996367 382150 996376
rect 382292 996305 382320 998378
rect 382278 996296 382334 996305
rect 382278 996231 382334 996240
rect 382740 995988 382792 995994
rect 382740 995930 382792 995936
rect 380898 995208 380954 995217
rect 380898 995143 380954 995152
rect 374826 994800 374882 994809
rect 374826 994735 374882 994744
rect 382752 994362 382780 995930
rect 382936 995489 382964 1005994
rect 383292 1000544 383344 1000550
rect 383292 1000486 383344 1000492
rect 383304 996033 383332 1000486
rect 383568 998776 383620 998782
rect 383620 998724 383700 998730
rect 383568 998718 383700 998724
rect 383580 998702 383700 998718
rect 383476 998640 383528 998646
rect 383476 998582 383528 998588
rect 383290 996024 383346 996033
rect 383290 995959 383346 995968
rect 383108 995852 383160 995858
rect 383108 995794 383160 995800
rect 382922 995480 382978 995489
rect 382922 995415 382978 995424
rect 383120 994537 383148 995794
rect 383488 995586 383516 998582
rect 383292 995580 383344 995586
rect 383292 995522 383344 995528
rect 383476 995580 383528 995586
rect 383476 995522 383528 995528
rect 383106 994528 383162 994537
rect 383304 994498 383332 995522
rect 383672 995330 383700 998702
rect 399944 997144 399996 997150
rect 399944 997086 399996 997092
rect 399956 996985 399984 997086
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 399850 996296 399906 996305
rect 399850 996231 399906 996240
rect 385038 995752 385094 995761
rect 388626 995752 388682 995761
rect 385094 995710 385342 995738
rect 385038 995687 385094 995696
rect 388682 995710 389022 995738
rect 388626 995687 388682 995696
rect 385604 995586 385986 995602
rect 385592 995580 385986 995586
rect 385644 995574 385986 995580
rect 385592 995522 385644 995528
rect 399864 995489 399892 996231
rect 387890 995480 387946 995489
rect 384316 995438 384698 995466
rect 387536 995438 387826 995466
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 387536 995178 387564 995438
rect 387890 995415 387946 995424
rect 388166 995480 388222 995489
rect 399850 995480 399906 995489
rect 388222 995438 388378 995466
rect 388812 995444 388864 995450
rect 388166 995415 388222 995424
rect 387524 995172 387576 995178
rect 387524 995114 387576 995120
rect 387904 995058 387932 995415
rect 388812 995386 388864 995392
rect 389100 995438 389666 995466
rect 389824 995444 389876 995450
rect 388824 995330 388852 995386
rect 389100 995330 389128 995438
rect 389824 995386 389876 995392
rect 388824 995302 389128 995330
rect 388442 995072 388498 995081
rect 387904 995030 388442 995058
rect 388442 995007 388498 995016
rect 389836 994498 389864 995386
rect 392136 994809 392164 995452
rect 392122 994800 392178 994809
rect 392122 994735 392178 994744
rect 383106 994463 383162 994472
rect 383292 994492 383344 994498
rect 383292 994434 383344 994440
rect 389824 994492 389876 994498
rect 389824 994434 389876 994440
rect 392688 994362 392716 995452
rect 393332 994634 393360 995452
rect 393976 994770 394004 995452
rect 395172 995042 395200 995452
rect 395160 995036 395212 995042
rect 395160 994978 395212 994984
rect 393964 994764 394016 994770
rect 393964 994706 394016 994712
rect 393320 994628 393372 994634
rect 393320 994570 393372 994576
rect 382740 994356 382792 994362
rect 382740 994298 382792 994304
rect 392676 994356 392728 994362
rect 392676 994298 392728 994304
rect 396368 994294 396396 995452
rect 397012 994906 397040 995452
rect 397656 995314 397684 995452
rect 398866 995438 398972 995466
rect 398944 995382 398972 995438
rect 399850 995415 399906 995424
rect 398932 995376 398984 995382
rect 398932 995318 398984 995324
rect 397644 995308 397696 995314
rect 397644 995250 397696 995256
rect 397000 994900 397052 994906
rect 397000 994842 397052 994848
rect 400876 994537 400904 1005994
rect 402256 996130 402284 1006130
rect 422680 1006097 422708 1006402
rect 431682 1006360 431738 1006369
rect 431682 1006295 431684 1006304
rect 431736 1006295 431738 1006304
rect 431684 1006266 431736 1006272
rect 429198 1006224 429254 1006233
rect 434640 1006194 434668 1007082
rect 505008 1007072 505060 1007078
rect 505006 1007040 505008 1007049
rect 505060 1007040 505062 1007049
rect 505006 1006975 505062 1006984
rect 510356 1006942 510384 1007150
rect 515588 1007072 515640 1007078
rect 515588 1007014 515640 1007020
rect 505376 1006936 505428 1006942
rect 505374 1006904 505376 1006913
rect 510344 1006936 510396 1006942
rect 505428 1006904 505430 1006913
rect 436744 1006868 436796 1006874
rect 510344 1006878 510396 1006884
rect 505374 1006839 505430 1006848
rect 510528 1006868 510580 1006874
rect 436744 1006810 436796 1006816
rect 510528 1006810 510580 1006816
rect 436756 1006466 436784 1006810
rect 451832 1006732 451884 1006738
rect 451832 1006674 451884 1006680
rect 436744 1006460 436796 1006466
rect 436744 1006402 436796 1006408
rect 448520 1006460 448572 1006466
rect 448520 1006402 448572 1006408
rect 429198 1006159 429200 1006168
rect 429252 1006159 429254 1006168
rect 434628 1006188 434680 1006194
rect 429200 1006130 429252 1006136
rect 434628 1006130 434680 1006136
rect 422666 1006088 422722 1006097
rect 422666 1006023 422722 1006032
rect 425518 1006088 425574 1006097
rect 430026 1006088 430082 1006097
rect 425518 1006023 425520 1006032
rect 425572 1006023 425574 1006032
rect 429200 1006052 429252 1006058
rect 425520 1005994 425572 1006000
rect 430026 1006023 430028 1006032
rect 429200 1005994 429252 1006000
rect 430080 1006023 430082 1006032
rect 430028 1005994 430080 1006000
rect 427544 1005712 427596 1005718
rect 427542 1005680 427544 1005689
rect 427596 1005680 427598 1005689
rect 427542 1005615 427598 1005624
rect 428372 1005576 428424 1005582
rect 428370 1005544 428372 1005553
rect 428424 1005544 428426 1005553
rect 428370 1005479 428426 1005488
rect 423496 1005440 423548 1005446
rect 423494 1005408 423496 1005417
rect 423548 1005408 423550 1005417
rect 423494 1005343 423550 1005352
rect 424324 1005304 424376 1005310
rect 424322 1005272 424324 1005281
rect 424376 1005272 424378 1005281
rect 424322 1005207 424378 1005216
rect 423494 1005000 423550 1005009
rect 422024 1004964 422076 1004970
rect 423494 1004935 423496 1004944
rect 422024 1004906 422076 1004912
rect 423548 1004935 423550 1004944
rect 423496 1004906 423548 1004912
rect 420828 1004828 420880 1004834
rect 420828 1004770 420880 1004776
rect 419448 1001972 419500 1001978
rect 419448 1001914 419500 1001920
rect 402244 996124 402296 996130
rect 402244 996066 402296 996072
rect 416134 995752 416190 995761
rect 416134 995687 416190 995696
rect 415398 995480 415454 995489
rect 415398 995415 415400 995424
rect 415452 995415 415454 995424
rect 415400 995386 415452 995392
rect 416148 995293 416176 995687
rect 416136 995287 416188 995293
rect 416136 995229 416188 995235
rect 419460 994702 419488 1001914
rect 419448 994696 419500 994702
rect 419448 994638 419500 994644
rect 420840 994566 420868 1004770
rect 422036 1003542 422064 1004906
rect 422666 1004864 422722 1004873
rect 422666 1004799 422668 1004808
rect 422720 1004799 422722 1004808
rect 422668 1004770 422720 1004776
rect 422208 1004624 422260 1004630
rect 424324 1004624 424376 1004630
rect 422208 1004566 422260 1004572
rect 424322 1004592 424324 1004601
rect 424376 1004592 424378 1004601
rect 422220 1003950 422248 1004566
rect 424322 1004527 424378 1004536
rect 425520 1004216 425572 1004222
rect 425518 1004184 425520 1004193
rect 425572 1004184 425574 1004193
rect 425518 1004119 425574 1004128
rect 425152 1004080 425204 1004086
rect 425150 1004048 425152 1004057
rect 425204 1004048 425206 1004057
rect 425150 1003983 425206 1003992
rect 422208 1003944 422260 1003950
rect 422208 1003886 422260 1003892
rect 422024 1003536 422076 1003542
rect 422024 1003478 422076 1003484
rect 423772 1003536 423824 1003542
rect 423772 1003478 423824 1003484
rect 423588 1002244 423640 1002250
rect 423588 1002186 423640 1002192
rect 421470 1002008 421526 1002017
rect 421470 1001943 421472 1001952
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 423600 1000958 423628 1002186
rect 423784 1001230 423812 1003478
rect 426346 1002552 426402 1002561
rect 426402 1002510 426572 1002538
rect 426346 1002487 426402 1002496
rect 426346 1002280 426402 1002289
rect 426346 1002215 426348 1002224
rect 426400 1002215 426402 1002224
rect 426348 1002186 426400 1002192
rect 425704 1001972 425756 1001978
rect 425704 1001914 425756 1001920
rect 423772 1001224 423824 1001230
rect 423772 1001166 423824 1001172
rect 423588 1000952 423640 1000958
rect 423588 1000894 423640 1000900
rect 425716 997762 425744 1001914
rect 426544 998714 426572 1002510
rect 427174 1002008 427230 1002017
rect 427174 1001943 427176 1001952
rect 427228 1001943 427230 1001952
rect 427176 1001914 427228 1001920
rect 426532 998708 426584 998714
rect 426532 998650 426584 998656
rect 429212 998442 429240 1005994
rect 440884 1005712 440936 1005718
rect 440884 1005654 440936 1005660
rect 433984 1004964 434036 1004970
rect 433984 1004906 434036 1004912
rect 430854 1004864 430910 1004873
rect 430854 1004799 430856 1004808
rect 430908 1004799 430910 1004808
rect 432050 1004864 432106 1004873
rect 432050 1004799 432052 1004808
rect 430856 1004770 430908 1004776
rect 432104 1004799 432106 1004808
rect 432052 1004770 432104 1004776
rect 430026 1004728 430082 1004737
rect 432878 1004728 432934 1004737
rect 430026 1004663 430028 1004672
rect 430080 1004663 430082 1004672
rect 431960 1004692 432012 1004698
rect 430028 1004634 430080 1004640
rect 432878 1004663 432880 1004672
rect 431960 1004634 432012 1004640
rect 432932 1004663 432934 1004672
rect 432880 1004634 432932 1004640
rect 429384 1000952 429436 1000958
rect 429384 1000894 429436 1000900
rect 429396 998578 429424 1000894
rect 429384 998572 429436 998578
rect 429384 998514 429436 998520
rect 429200 998436 429252 998442
rect 429200 998378 429252 998384
rect 425704 997756 425756 997762
rect 425704 997698 425756 997704
rect 431972 997150 432000 1004634
rect 433338 1002008 433394 1002017
rect 433338 1001943 433340 1001952
rect 433392 1001943 433394 1001952
rect 433340 1001914 433392 1001920
rect 433996 997626 434024 1004906
rect 436744 1004828 436796 1004834
rect 436744 1004770 436796 1004776
rect 435364 1001972 435416 1001978
rect 435364 1001914 435416 1001920
rect 433984 997620 434036 997626
rect 433984 997562 434036 997568
rect 431960 997144 432012 997150
rect 431960 997086 432012 997092
rect 420828 994560 420880 994566
rect 400862 994528 400918 994537
rect 420828 994502 420880 994508
rect 400862 994463 400918 994472
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 396356 994288 396408 994294
rect 396356 994230 396408 994236
rect 370504 985992 370556 985998
rect 370504 985934 370556 985940
rect 381188 983634 381216 994230
rect 435376 992934 435404 1001914
rect 429936 992928 429988 992934
rect 429936 992870 429988 992876
rect 435364 992928 435416 992934
rect 435364 992870 435416 992876
rect 414112 991500 414164 991506
rect 414112 991442 414164 991448
rect 397828 985992 397880 985998
rect 397828 985934 397880 985940
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 985934
rect 414124 983620 414152 991442
rect 429948 983634 429976 992870
rect 436756 985998 436784 1004770
rect 438124 1004692 438176 1004698
rect 438124 1004634 438176 1004640
rect 438136 986134 438164 1004634
rect 440896 998345 440924 1005654
rect 446404 1005576 446456 1005582
rect 446404 1005518 446456 1005524
rect 440882 998336 440938 998345
rect 440882 998271 440938 998280
rect 439688 997756 439740 997762
rect 439688 997698 439740 997704
rect 439700 996441 439728 997698
rect 439872 997620 439924 997626
rect 439872 997562 439924 997568
rect 439884 996985 439912 997562
rect 439870 996976 439926 996985
rect 439870 996911 439926 996920
rect 439686 996432 439742 996441
rect 439686 996367 439742 996376
rect 446416 995625 446444 1005518
rect 448532 1003338 448560 1006402
rect 451844 1004222 451872 1006674
rect 505376 1006664 505428 1006670
rect 505374 1006632 505376 1006641
rect 505428 1006632 505430 1006641
rect 469864 1006596 469916 1006602
rect 505374 1006567 505430 1006576
rect 469864 1006538 469916 1006544
rect 456800 1006324 456852 1006330
rect 456800 1006266 456852 1006272
rect 449164 1004216 449216 1004222
rect 449164 1004158 449216 1004164
rect 451832 1004216 451884 1004222
rect 451832 1004158 451884 1004164
rect 448520 1003332 448572 1003338
rect 448520 1003274 448572 1003280
rect 446402 995616 446458 995625
rect 446402 995551 446458 995560
rect 446128 994288 446180 994294
rect 449176 994265 449204 1004158
rect 456812 1004086 456840 1006266
rect 464344 1005440 464396 1005446
rect 464344 1005382 464396 1005388
rect 454868 1004080 454920 1004086
rect 454868 1004022 454920 1004028
rect 456800 1004080 456852 1004086
rect 456800 1004022 456852 1004028
rect 451648 1003332 451700 1003338
rect 451648 1003274 451700 1003280
rect 451660 995110 451688 1003274
rect 454880 995897 454908 1004022
rect 458824 1003944 458876 1003950
rect 458824 1003886 458876 1003892
rect 461584 1003944 461636 1003950
rect 461584 1003886 461636 1003892
rect 456800 1001224 456852 1001230
rect 456800 1001166 456852 1001172
rect 454866 995888 454922 995897
rect 454866 995823 454922 995832
rect 451648 995104 451700 995110
rect 451648 995046 451700 995052
rect 456812 994294 456840 1001166
rect 458836 994838 458864 1003886
rect 458824 994832 458876 994838
rect 458824 994774 458876 994780
rect 461596 994430 461624 1003886
rect 464356 994809 464384 1005382
rect 465724 1005304 465776 1005310
rect 465724 1005246 465776 1005252
rect 464342 994800 464398 994809
rect 464342 994735 464398 994744
rect 465736 994537 465764 1005246
rect 467564 1004216 467616 1004222
rect 467564 1004158 467616 1004164
rect 467576 998918 467604 1004158
rect 467564 998912 467616 998918
rect 467564 998854 467616 998860
rect 466460 998708 466512 998714
rect 466460 998650 466512 998656
rect 465722 994528 465778 994537
rect 465722 994463 465778 994472
rect 461584 994424 461636 994430
rect 461584 994366 461636 994372
rect 456800 994288 456852 994294
rect 446128 994230 446180 994236
rect 449162 994256 449218 994265
rect 438124 986128 438176 986134
rect 438124 986070 438176 986076
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 994230
rect 456800 994230 456852 994236
rect 449162 994191 449218 994200
rect 466472 994158 466500 998650
rect 469876 996169 469904 1006538
rect 510540 1006398 510568 1006810
rect 514208 1006664 514260 1006670
rect 514208 1006606 514260 1006612
rect 513564 1006460 513616 1006466
rect 513564 1006402 513616 1006408
rect 507860 1006392 507912 1006398
rect 507858 1006360 507860 1006369
rect 510528 1006392 510580 1006398
rect 507912 1006360 507914 1006369
rect 510528 1006334 510580 1006340
rect 507858 1006295 507914 1006304
rect 506204 1006256 506256 1006262
rect 506202 1006224 506204 1006233
rect 506256 1006224 506258 1006233
rect 471428 1006188 471480 1006194
rect 506202 1006159 506258 1006168
rect 471428 1006130 471480 1006136
rect 471244 1006052 471296 1006058
rect 471244 1005994 471296 1006000
rect 471256 996713 471284 1005994
rect 471242 996704 471298 996713
rect 471242 996639 471298 996648
rect 469862 996160 469918 996169
rect 469862 996095 469918 996104
rect 471440 995353 471468 1006130
rect 498842 1006088 498898 1006097
rect 496728 1006052 496780 1006058
rect 498842 1006023 498844 1006032
rect 496728 1005994 496780 1006000
rect 498896 1006023 498898 1006032
rect 500498 1006088 500554 1006097
rect 513576 1006058 513604 1006402
rect 514220 1006194 514248 1006606
rect 514208 1006188 514260 1006194
rect 514208 1006130 514260 1006136
rect 500498 1006023 500500 1006032
rect 498844 1005994 498896 1006000
rect 500552 1006023 500554 1006032
rect 513564 1006052 513616 1006058
rect 500500 1005994 500552 1006000
rect 513564 1005994 513616 1006000
rect 472624 998912 472676 998918
rect 472624 998854 472676 998860
rect 472440 998572 472492 998578
rect 472440 998514 472492 998520
rect 472256 998436 472308 998442
rect 472256 998378 472308 998384
rect 471426 995344 471482 995353
rect 471426 995279 471482 995288
rect 472268 995081 472296 998378
rect 472452 995466 472480 998514
rect 472636 995586 472664 998854
rect 488908 997348 488960 997354
rect 488908 997290 488960 997296
rect 488920 996985 488948 997290
rect 488906 996976 488962 996985
rect 488906 996911 488962 996920
rect 483754 995752 483810 995761
rect 485594 995752 485650 995761
rect 483810 995710 484150 995738
rect 485346 995710 485594 995738
rect 483754 995687 483810 995696
rect 485594 995687 485650 995696
rect 474738 995616 474794 995625
rect 473372 995586 473662 995602
rect 472624 995580 472676 995586
rect 472624 995522 472676 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 480718 995616 480774 995625
rect 474794 995574 474950 995602
rect 474738 995551 474794 995560
rect 481270 995616 481326 995625
rect 481114 995574 481270 995602
rect 480718 995551 480774 995560
rect 481270 995551 481326 995560
rect 473360 995522 473412 995528
rect 472452 995438 473032 995466
rect 473004 995330 473032 995438
rect 473924 995438 474306 995466
rect 476500 995438 476790 995466
rect 476960 995438 477342 995466
rect 473924 995330 473952 995438
rect 476500 995353 476528 995438
rect 473004 995302 473952 995330
rect 476486 995344 476542 995353
rect 476486 995279 476542 995288
rect 476960 995081 476988 995438
rect 472254 995072 472310 995081
rect 472254 995007 472310 995016
rect 476946 995072 477002 995081
rect 476946 995007 477002 995016
rect 474556 994968 474608 994974
rect 474556 994910 474608 994916
rect 474568 994294 474596 994910
rect 475384 994424 475436 994430
rect 475384 994366 475436 994372
rect 474556 994288 474608 994294
rect 474556 994230 474608 994236
rect 475396 994158 475424 994366
rect 477972 994265 478000 995452
rect 478616 994537 478644 995452
rect 480732 995081 480760 995551
rect 480718 995072 480774 995081
rect 480718 995007 480774 995016
rect 481652 994809 481680 995452
rect 482296 994838 482324 995452
rect 482940 994974 482968 995452
rect 485976 995110 486004 995452
rect 485964 995104 486016 995110
rect 485964 995046 486016 995052
rect 486620 994974 486648 995452
rect 482928 994968 482980 994974
rect 482928 994910 482980 994916
rect 486608 994968 486660 994974
rect 486608 994910 486660 994916
rect 482284 994832 482336 994838
rect 481638 994800 481694 994809
rect 482284 994774 482336 994780
rect 481638 994735 481694 994744
rect 478602 994528 478658 994537
rect 478602 994463 478658 994472
rect 487816 994430 487844 995452
rect 489920 994968 489972 994974
rect 489920 994910 489972 994916
rect 487804 994424 487856 994430
rect 487804 994366 487856 994372
rect 489932 994294 489960 994910
rect 496740 994430 496768 1005994
rect 509054 1005952 509110 1005961
rect 509054 1005887 509056 1005896
rect 509108 1005887 509110 1005896
rect 514024 1005916 514076 1005922
rect 509056 1005858 509108 1005864
rect 514024 1005858 514076 1005864
rect 498844 1005304 498896 1005310
rect 498842 1005272 498844 1005281
rect 498896 1005272 498898 1005281
rect 498842 1005207 498898 1005216
rect 499670 1005000 499726 1005009
rect 498108 1004964 498160 1004970
rect 499670 1004935 499672 1004944
rect 498108 1004906 498160 1004912
rect 499724 1004935 499726 1004944
rect 508226 1005000 508282 1005009
rect 508226 1004935 508228 1004944
rect 499672 1004906 499724 1004912
rect 508280 1004935 508282 1004944
rect 509882 1005000 509938 1005009
rect 509938 1004958 510108 1004986
rect 509882 1004935 509938 1004944
rect 508228 1004906 508280 1004912
rect 498120 1001230 498148 1004906
rect 501326 1004864 501382 1004873
rect 499304 1004828 499356 1004834
rect 501326 1004799 501328 1004808
rect 499304 1004770 499356 1004776
rect 501380 1004799 501382 1004808
rect 507030 1004864 507086 1004873
rect 507030 1004799 507032 1004808
rect 501328 1004770 501380 1004776
rect 507084 1004799 507086 1004808
rect 509884 1004828 509936 1004834
rect 507032 1004770 507084 1004776
rect 509884 1004770 509936 1004776
rect 498108 1001224 498160 1001230
rect 498108 1001166 498160 1001172
rect 499316 998442 499344 1004770
rect 503350 1004728 503406 1004737
rect 508226 1004728 508282 1004737
rect 503350 1004663 503352 1004672
rect 503404 1004663 503406 1004672
rect 507308 1004692 507360 1004698
rect 503352 1004634 503404 1004640
rect 508226 1004663 508228 1004672
rect 507308 1004634 507360 1004640
rect 508280 1004663 508282 1004672
rect 508228 1004634 508280 1004640
rect 499488 1004624 499540 1004630
rect 500500 1004624 500552 1004630
rect 499488 1004566 499540 1004572
rect 500498 1004592 500500 1004601
rect 500552 1004592 500554 1004601
rect 499500 1003950 499528 1004566
rect 500498 1004527 500554 1004536
rect 502524 1004080 502576 1004086
rect 502522 1004048 502524 1004057
rect 502576 1004048 502578 1004057
rect 502522 1003983 502578 1003992
rect 499488 1003944 499540 1003950
rect 499488 1003886 499540 1003892
rect 501694 1002280 501750 1002289
rect 501694 1002215 501696 1002224
rect 501748 1002215 501750 1002224
rect 504364 1002244 504416 1002250
rect 501696 1002186 501748 1002192
rect 504364 1002186 504416 1002192
rect 501694 1002008 501750 1002017
rect 500868 1001972 500920 1001978
rect 502522 1002008 502578 1002017
rect 501694 1001943 501696 1001952
rect 500868 1001914 500920 1001920
rect 501748 1001943 501750 1001952
rect 501880 1001972 501932 1001978
rect 501696 1001914 501748 1001920
rect 501880 1001914 501932 1001920
rect 502352 1001966 502522 1001994
rect 499304 998436 499356 998442
rect 499304 998378 499356 998384
rect 496728 994424 496780 994430
rect 496728 994366 496780 994372
rect 500880 994294 500908 1001914
rect 501892 994838 501920 1001914
rect 502352 997490 502380 1001966
rect 502522 1001943 502578 1001952
rect 503350 1002008 503406 1002017
rect 503350 1001943 503352 1001952
rect 503404 1001943 503406 1001952
rect 504178 1002008 504234 1002017
rect 504178 1001943 504180 1001952
rect 503352 1001914 503404 1001920
rect 504232 1001943 504234 1001952
rect 504180 1001914 504232 1001920
rect 504376 1001894 504404 1002186
rect 504546 1002144 504602 1002153
rect 504546 1002079 504548 1002088
rect 504600 1002079 504602 1002088
rect 507124 1002108 507176 1002114
rect 504548 1002050 504600 1002056
rect 507124 1002050 507176 1002056
rect 505744 1001972 505796 1001978
rect 505744 1001914 505796 1001920
rect 504376 1001866 504588 1001894
rect 504560 998073 504588 1001866
rect 504546 998064 504602 998073
rect 504546 997999 504602 998008
rect 502340 997484 502392 997490
rect 502340 997426 502392 997432
rect 505756 997082 505784 1001914
rect 505744 997076 505796 997082
rect 505744 997018 505796 997024
rect 506202 995888 506258 995897
rect 506202 995823 506204 995832
rect 506256 995823 506258 995832
rect 506204 995794 506256 995800
rect 507136 995110 507164 1002050
rect 507320 997762 507348 1004634
rect 507308 997756 507360 997762
rect 507308 997698 507360 997704
rect 509896 997626 509924 1004770
rect 510080 1004562 510108 1004958
rect 511264 1004964 511316 1004970
rect 511264 1004906 511316 1004912
rect 510620 1004692 510672 1004698
rect 510620 1004634 510672 1004640
rect 510068 1004556 510120 1004562
rect 510068 1004498 510120 1004504
rect 510342 1002008 510398 1002017
rect 510342 1001943 510344 1001952
rect 510396 1001943 510398 1001952
rect 510344 1001914 510396 1001920
rect 509884 997620 509936 997626
rect 509884 997562 509936 997568
rect 510632 997354 510660 1004634
rect 510620 997348 510672 997354
rect 510620 997290 510672 997296
rect 511276 996130 511304 1004906
rect 512644 1001972 512696 1001978
rect 512644 1001914 512696 1001920
rect 511264 996124 511316 996130
rect 511264 996066 511316 996072
rect 509056 995852 509108 995858
rect 509056 995794 509108 995800
rect 507124 995104 507176 995110
rect 509068 995081 509096 995794
rect 507124 995046 507176 995052
rect 509054 995072 509110 995081
rect 509054 995007 509110 995016
rect 511078 995072 511134 995081
rect 511078 995007 511134 995016
rect 501880 994832 501932 994838
rect 501880 994774 501932 994780
rect 489920 994288 489972 994294
rect 477958 994256 478014 994265
rect 489920 994230 489972 994236
rect 500868 994288 500920 994294
rect 500868 994230 500920 994236
rect 477958 994191 478014 994200
rect 466460 994152 466512 994158
rect 466460 994094 466512 994100
rect 475384 994152 475436 994158
rect 475384 994094 475436 994100
rect 478972 992928 479024 992934
rect 478972 992870 479024 992876
rect 462780 986128 462832 986134
rect 462780 986070 462832 986076
rect 429948 983606 430330 983634
rect 446140 983606 446522 983634
rect 462792 983620 462820 986070
rect 478984 983620 479012 992870
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 995007
rect 512656 991506 512684 1001914
rect 512644 991500 512696 991506
rect 512644 991442 512696 991448
rect 514036 985998 514064 1005858
rect 515404 1004556 515456 1004562
rect 515404 1004498 515456 1004504
rect 514668 1004080 514720 1004086
rect 514668 1004022 514720 1004028
rect 514680 998578 514708 1004022
rect 514668 998572 514720 998578
rect 514668 998514 514720 998520
rect 515416 986134 515444 1004498
rect 515600 998714 515628 1007014
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 516796 1001894 516824 1005246
rect 516796 1001866 517284 1001894
rect 515588 998708 515640 998714
rect 515588 998650 515640 998656
rect 516876 997756 516928 997762
rect 516876 997698 516928 997704
rect 516692 997484 516744 997490
rect 516692 997426 516744 997432
rect 516704 996441 516732 997426
rect 516888 996713 516916 997698
rect 517060 997620 517112 997626
rect 517060 997562 517112 997568
rect 517072 996985 517100 997562
rect 517058 996976 517114 996985
rect 517058 996911 517114 996920
rect 516874 996704 516930 996713
rect 516874 996639 516930 996648
rect 516690 996432 516746 996441
rect 516690 996367 516746 996376
rect 517256 993682 517284 1001866
rect 517520 998436 517572 998442
rect 517520 998378 517572 998384
rect 517532 995081 517560 998378
rect 517704 997076 517756 997082
rect 517704 997018 517756 997024
rect 517518 995072 517574 995081
rect 517518 995007 517574 995016
rect 517716 994537 517744 997018
rect 518176 994809 518204 1007150
rect 552294 1007040 552350 1007049
rect 552294 1006975 552296 1006984
rect 552348 1006975 552350 1006984
rect 568028 1007004 568080 1007010
rect 552296 1006946 552348 1006952
rect 568028 1006946 568080 1006952
rect 520924 1006868 520976 1006874
rect 520924 1006810 520976 1006816
rect 519544 1006460 519596 1006466
rect 519544 1006402 519596 1006408
rect 518348 1003944 518400 1003950
rect 518348 1003886 518400 1003892
rect 518162 994800 518218 994809
rect 518162 994735 518218 994744
rect 517702 994528 517758 994537
rect 517702 994463 517758 994472
rect 518360 994158 518388 1003886
rect 519556 996169 519584 1006402
rect 520372 1001224 520424 1001230
rect 520372 1001166 520424 1001172
rect 519542 996160 519598 996169
rect 519542 996095 519598 996104
rect 519820 994968 519872 994974
rect 519820 994910 519872 994916
rect 519832 994430 519860 994910
rect 519820 994424 519872 994430
rect 519820 994366 519872 994372
rect 518348 994152 518400 994158
rect 518348 994094 518400 994100
rect 520384 993818 520412 1001166
rect 520936 994265 520964 1006810
rect 557172 1006800 557224 1006806
rect 557170 1006768 557172 1006777
rect 565268 1006800 565320 1006806
rect 557224 1006768 557226 1006777
rect 565268 1006742 565320 1006748
rect 557170 1006703 557226 1006712
rect 553124 1006664 553176 1006670
rect 553122 1006632 553124 1006641
rect 562508 1006664 562560 1006670
rect 553176 1006632 553178 1006641
rect 562508 1006606 562560 1006612
rect 553122 1006567 553178 1006576
rect 551100 1006528 551152 1006534
rect 551098 1006496 551100 1006505
rect 556620 1006528 556672 1006534
rect 551152 1006496 551154 1006505
rect 556804 1006528 556856 1006534
rect 556620 1006470 556672 1006476
rect 556802 1006496 556804 1006505
rect 556856 1006496 556858 1006505
rect 551098 1006431 551154 1006440
rect 555424 1006392 555476 1006398
rect 555424 1006334 555476 1006340
rect 522304 1006324 522356 1006330
rect 522304 1006266 522356 1006272
rect 522316 995926 522344 1006266
rect 553952 1006256 554004 1006262
rect 553950 1006224 553952 1006233
rect 554004 1006224 554006 1006233
rect 522488 1006188 522540 1006194
rect 553950 1006159 554006 1006168
rect 522488 1006130 522540 1006136
rect 522304 995920 522356 995926
rect 522304 995862 522356 995868
rect 522500 995761 522528 1006130
rect 554318 1006088 554374 1006097
rect 554318 1006023 554320 1006032
rect 554372 1006023 554374 1006032
rect 554320 1005994 554372 1006000
rect 551466 1005136 551522 1005145
rect 551466 1005071 551468 1005080
rect 551520 1005071 551522 1005080
rect 551468 1005042 551520 1005048
rect 555148 1002448 555200 1002454
rect 555146 1002416 555148 1002425
rect 555200 1002416 555202 1002425
rect 555146 1002351 555202 1002360
rect 554318 1002280 554374 1002289
rect 551928 1002244 551980 1002250
rect 554318 1002215 554320 1002224
rect 551928 1002186 551980 1002192
rect 554372 1002215 554374 1002224
rect 554320 1002186 554372 1002192
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 523868 998708 523920 998714
rect 523868 998650 523920 998656
rect 522486 995752 522542 995761
rect 522486 995687 522542 995696
rect 523880 995489 523908 998650
rect 524052 998572 524104 998578
rect 524052 998514 524104 998520
rect 524064 997257 524092 998514
rect 549168 997824 549220 997830
rect 551468 997824 551520 997830
rect 549168 997766 549220 997772
rect 551466 997792 551468 997801
rect 551520 997792 551522 997801
rect 540888 997688 540940 997694
rect 540888 997630 540940 997636
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 540900 996985 540928 997630
rect 549180 997082 549208 997766
rect 551466 997727 551522 997736
rect 551940 997558 551968 1002186
rect 555146 1002008 555202 1002017
rect 554700 1001966 555146 1001994
rect 553122 998608 553178 998617
rect 553122 998543 553124 998552
rect 553176 998543 553178 998552
rect 553124 998514 553176 998520
rect 552294 998472 552350 998481
rect 552294 998407 552296 998416
rect 552348 998407 552350 998416
rect 552296 998378 552348 998384
rect 551928 997552 551980 997558
rect 551928 997494 551980 997500
rect 549168 997076 549220 997082
rect 549168 997018 549220 997024
rect 540886 996976 540942 996985
rect 540886 996911 540942 996920
rect 524050 996704 524106 996713
rect 524050 996639 524106 996648
rect 524064 995586 524092 996639
rect 549442 996432 549498 996441
rect 549442 996367 549444 996376
rect 549496 996367 549498 996376
rect 550640 996396 550692 996402
rect 549444 996338 549496 996344
rect 550640 996338 550692 996344
rect 540244 995852 540296 995858
rect 540244 995794 540296 995800
rect 526074 995752 526130 995761
rect 528558 995752 528614 995761
rect 526130 995710 526378 995738
rect 526074 995687 526130 995696
rect 529110 995752 529166 995761
rect 528614 995710 528770 995738
rect 528558 995687 528614 995696
rect 533526 995752 533582 995761
rect 529166 995710 529414 995738
rect 529110 995687 529166 995696
rect 536562 995752 536618 995761
rect 533582 995710 533738 995738
rect 533526 995687 533582 995696
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 525352 995586 525734 995602
rect 524052 995580 524104 995586
rect 524052 995522 524104 995528
rect 525340 995580 525734 995586
rect 525392 995574 525734 995580
rect 525340 995522 525392 995528
rect 523866 995480 523922 995489
rect 523866 995415 523922 995424
rect 524786 995480 524842 995489
rect 532698 995480 532754 995489
rect 524842 995438 525090 995466
rect 524786 995415 524842 995424
rect 528204 995110 528232 995452
rect 528192 995104 528244 995110
rect 530044 995081 530072 995452
rect 532148 995172 532200 995178
rect 532148 995114 532200 995120
rect 528192 995046 528244 995052
rect 530030 995072 530086 995081
rect 530030 995007 530086 995016
rect 530216 994968 530268 994974
rect 530216 994910 530268 994916
rect 523684 994424 523736 994430
rect 523684 994366 523736 994372
rect 520922 994256 520978 994265
rect 520922 994191 520978 994200
rect 523696 994158 523724 994366
rect 530228 994294 530256 994910
rect 530216 994288 530268 994294
rect 532160 994265 532188 995114
rect 532528 994537 532556 995452
rect 532754 995438 533094 995466
rect 532698 995415 532754 995424
rect 534368 994974 534396 995452
rect 534356 994968 534408 994974
rect 534356 994910 534408 994916
rect 532514 994528 532570 994537
rect 532514 994463 532570 994472
rect 530216 994230 530268 994236
rect 532146 994256 532202 994265
rect 532146 994191 532202 994200
rect 535564 994158 535592 995452
rect 537404 994809 537432 995452
rect 537680 995438 538062 995466
rect 537390 994800 537446 994809
rect 537390 994735 537446 994744
rect 537680 994294 537708 995438
rect 538126 995208 538182 995217
rect 538126 995143 538182 995152
rect 538310 995208 538366 995217
rect 538310 995143 538366 995152
rect 538140 994974 538168 995143
rect 538128 994968 538180 994974
rect 538128 994910 538180 994916
rect 538324 994430 538352 995143
rect 539244 994838 539272 995452
rect 540256 995178 540284 995794
rect 540244 995172 540296 995178
rect 540244 995114 540296 995120
rect 539232 994832 539284 994838
rect 539232 994774 539284 994780
rect 538312 994424 538364 994430
rect 538312 994366 538364 994372
rect 550652 994294 550680 996338
rect 554700 995586 554728 1001966
rect 555146 1001943 555202 1001952
rect 555436 997694 555464 1006334
rect 555976 1005440 556028 1005446
rect 555974 1005408 555976 1005417
rect 556028 1005408 556030 1005417
rect 555974 1005343 556030 1005352
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 555424 997688 555476 997694
rect 555424 997630 555476 997636
rect 554688 995580 554740 995586
rect 554688 995522 554740 995528
rect 556632 995110 556660 1006470
rect 556802 1006431 556858 1006440
rect 558828 1006392 558880 1006398
rect 558826 1006360 558828 1006369
rect 558880 1006360 558882 1006369
rect 558826 1006295 558882 1006304
rect 562520 1006194 562548 1006606
rect 564440 1006528 564492 1006534
rect 564440 1006470 564492 1006476
rect 562508 1006188 562560 1006194
rect 562508 1006130 562560 1006136
rect 564452 1005922 564480 1006470
rect 564440 1005916 564492 1005922
rect 564440 1005858 564492 1005864
rect 560850 1005000 560906 1005009
rect 560850 1004935 560852 1004944
rect 560904 1004935 560906 1004944
rect 560852 1004906 560904 1004912
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002552 558054 1002561
rect 557998 1002487 558000 1002496
rect 558052 1002487 558054 1002496
rect 558000 1002458 558052 1002464
rect 557540 1002448 557592 1002454
rect 557540 1002390 557592 1002396
rect 557552 997218 557580 1002390
rect 557998 1002280 558054 1002289
rect 557998 1002215 558000 1002224
rect 558052 1002215 558054 1002224
rect 558000 1002186 558052 1002192
rect 557540 997212 557592 997218
rect 557540 997154 557592 997160
rect 558196 996810 558224 1004770
rect 560850 1004728 560906 1004737
rect 559472 1004692 559524 1004698
rect 560850 1004663 560852 1004672
rect 559472 1004634 559524 1004640
rect 560904 1004663 560906 1004672
rect 565084 1004692 565136 1004698
rect 560852 1004634 560904 1004640
rect 565084 1004634 565136 1004640
rect 558826 1002416 558882 1002425
rect 558826 1002351 558828 1002360
rect 558880 1002351 558882 1002360
rect 558828 1002322 558880 1002328
rect 559484 1001894 559512 1004634
rect 560944 1002516 560996 1002522
rect 560944 1002458 560996 1002464
rect 560482 1002280 560538 1002289
rect 560300 1002244 560352 1002250
rect 560482 1002215 560484 1002224
rect 560300 1002186 560352 1002192
rect 560536 1002215 560538 1002224
rect 560484 1002186 560536 1002192
rect 559654 1002144 559710 1002153
rect 559654 1002079 559656 1002088
rect 559708 1002079 559710 1002088
rect 559656 1002050 559708 1002056
rect 560022 1002008 560078 1002017
rect 560022 1001943 560024 1001952
rect 560076 1001943 560078 1001952
rect 560024 1001914 560076 1001920
rect 559484 1001866 559604 1001894
rect 558184 996804 558236 996810
rect 558184 996746 558236 996752
rect 556620 995104 556672 995110
rect 556620 995046 556672 995052
rect 537668 994288 537720 994294
rect 537668 994230 537720 994236
rect 550640 994288 550692 994294
rect 550640 994230 550692 994236
rect 523684 994152 523736 994158
rect 523684 994094 523736 994100
rect 535552 994152 535604 994158
rect 535552 994094 535604 994100
rect 520372 993812 520424 993818
rect 520372 993754 520424 993760
rect 517244 993676 517296 993682
rect 517244 993618 517296 993624
rect 559576 991506 559604 1001866
rect 560312 995994 560340 1002186
rect 560300 995988 560352 995994
rect 560300 995930 560352 995936
rect 560956 992934 560984 1002458
rect 562508 1002380 562560 1002386
rect 562508 1002322 562560 1002328
rect 561678 1002144 561734 1002153
rect 561496 1002108 561548 1002114
rect 561678 1002079 561680 1002088
rect 561496 1002050 561548 1002056
rect 561732 1002079 561734 1002088
rect 561680 1002050 561732 1002056
rect 561508 1001994 561536 1002050
rect 561508 1001966 561720 1001994
rect 561692 995858 561720 1001966
rect 562324 1001972 562376 1001978
rect 562324 1001914 562376 1001920
rect 561680 995852 561732 995858
rect 561680 995794 561732 995800
rect 562140 995852 562192 995858
rect 562140 995794 562192 995800
rect 562152 995586 562180 995794
rect 562140 995580 562192 995586
rect 562140 995522 562192 995528
rect 560944 992928 560996 992934
rect 560944 992870 560996 992876
rect 543832 991500 543884 991506
rect 543832 991442 543884 991448
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 515404 986128 515456 986134
rect 515404 986070 515456 986076
rect 527640 986128 527692 986134
rect 527640 986070 527692 986076
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 986070
rect 543844 983620 543872 991442
rect 562336 990146 562364 1001914
rect 562520 993070 562548 1002322
rect 563060 1002244 563112 1002250
rect 563060 1002186 563112 1002192
rect 563072 996130 563100 1002186
rect 563704 1002108 563756 1002114
rect 563704 1002050 563756 1002056
rect 563060 996124 563112 996130
rect 563060 996066 563112 996072
rect 562508 993064 562560 993070
rect 562508 993006 562560 993012
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 563716 987426 563744 1002050
rect 563704 987420 563756 987426
rect 563704 987362 563756 987368
rect 565096 985998 565124 1004634
rect 565280 999122 565308 1006742
rect 567844 1005916 567896 1005922
rect 567844 1005858 567896 1005864
rect 566464 1004964 566516 1004970
rect 566464 1004906 566516 1004912
rect 565268 999116 565320 999122
rect 565268 999058 565320 999064
rect 565820 998572 565872 998578
rect 565820 998514 565872 998520
rect 565832 997354 565860 998514
rect 565820 997348 565872 997354
rect 565820 997290 565872 997296
rect 566476 986134 566504 1004906
rect 567856 994838 567884 1005858
rect 568040 998238 568068 1006946
rect 571984 1006324 572036 1006330
rect 571984 1006266 572036 1006272
rect 570604 1006188 570656 1006194
rect 570604 1006130 570656 1006136
rect 569224 1005100 569276 1005106
rect 569224 1005042 569276 1005048
rect 568212 999116 568264 999122
rect 568212 999058 568264 999064
rect 568028 998232 568080 998238
rect 568028 998174 568080 998180
rect 567844 994832 567896 994838
rect 567844 994774 567896 994780
rect 568224 994265 568252 999058
rect 568210 994256 568266 994265
rect 568210 994191 568266 994200
rect 569236 993954 569264 1005042
rect 570236 997348 570288 997354
rect 570236 997290 570288 997296
rect 570248 994809 570276 997290
rect 570616 995994 570644 1006130
rect 571996 997422 572024 1006266
rect 574744 1006052 574796 1006058
rect 574744 1005994 574796 1006000
rect 573364 1005440 573416 1005446
rect 573364 1005382 573416 1005388
rect 572720 998436 572772 998442
rect 572720 998378 572772 998384
rect 571984 997416 572036 997422
rect 571984 997358 572036 997364
rect 570788 997212 570840 997218
rect 570788 997154 570840 997160
rect 570604 995988 570656 995994
rect 570604 995930 570656 995936
rect 570800 994974 570828 997154
rect 572732 996946 572760 998378
rect 572904 998232 572956 998238
rect 572904 998174 572956 998180
rect 572720 996940 572772 996946
rect 572720 996882 572772 996888
rect 570788 994968 570840 994974
rect 570788 994910 570840 994916
rect 570234 994800 570290 994809
rect 570234 994735 570290 994744
rect 572916 994537 572944 998174
rect 573376 997694 573404 1005382
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 573364 997688 573416 997694
rect 573364 997630 573416 997636
rect 572902 994528 572958 994537
rect 572902 994463 572958 994472
rect 572720 994288 572772 994294
rect 572720 994230 572772 994236
rect 569224 993948 569276 993954
rect 569224 993890 569276 993896
rect 572732 989534 572760 994230
rect 574112 994090 574140 1001166
rect 574756 997286 574784 1005994
rect 591304 997960 591356 997966
rect 591304 997902 591356 997908
rect 625804 997960 625856 997966
rect 625804 997902 625856 997908
rect 590844 997824 590896 997830
rect 590844 997766 590896 997772
rect 590568 997416 590620 997422
rect 590568 997358 590620 997364
rect 574744 997280 574796 997286
rect 574744 997222 574796 997228
rect 590580 996985 590608 997358
rect 590856 997286 590884 997766
rect 591316 997558 591344 997902
rect 625620 997824 625672 997830
rect 625620 997766 625672 997772
rect 623688 997688 623740 997694
rect 623688 997630 623740 997636
rect 591304 997552 591356 997558
rect 591304 997494 591356 997500
rect 590844 997280 590896 997286
rect 590844 997222 590896 997228
rect 617156 997076 617208 997082
rect 617156 997018 617208 997024
rect 590566 996976 590622 996985
rect 590384 996940 590436 996946
rect 590566 996911 590622 996920
rect 590384 996882 590436 996888
rect 590396 996418 590424 996882
rect 590568 996736 590620 996742
rect 590566 996704 590568 996713
rect 590620 996704 590622 996713
rect 590566 996639 590622 996648
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 617168 995353 617196 997018
rect 623700 995586 623728 997630
rect 625632 996033 625660 997766
rect 625618 996024 625674 996033
rect 625618 995959 625674 995968
rect 625620 995852 625672 995858
rect 625620 995794 625672 995800
rect 623688 995580 623740 995586
rect 623688 995522 623740 995528
rect 617154 995344 617210 995353
rect 617154 995279 617210 995288
rect 590566 995072 590622 995081
rect 590566 995007 590622 995016
rect 590580 994566 590608 995007
rect 625632 994566 625660 995794
rect 625816 995761 625844 997902
rect 642088 995920 642140 995926
rect 642088 995862 642140 995868
rect 642100 995761 642128 995862
rect 625802 995752 625858 995761
rect 625802 995687 625858 995696
rect 627182 995752 627238 995761
rect 629758 995752 629814 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 630862 995752 630918 995761
rect 629814 995710 630016 995738
rect 629758 995687 629814 995696
rect 634542 995752 634598 995761
rect 630918 995710 631212 995738
rect 630862 995687 630918 995696
rect 637670 995752 637726 995761
rect 634598 995710 634892 995738
rect 637376 995710 637670 995738
rect 634542 995687 634598 995696
rect 637670 995687 637726 995696
rect 642086 995752 642142 995761
rect 642086 995687 642142 995696
rect 629574 995616 629630 995625
rect 626552 995586 626888 995602
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 629630 995574 629892 995602
rect 629574 995551 629630 995560
rect 626540 995522 626592 995528
rect 627932 995438 628176 995466
rect 590568 994560 590620 994566
rect 590568 994502 590620 994508
rect 625620 994560 625672 994566
rect 625620 994502 625672 994508
rect 627932 994265 627960 995438
rect 629864 995330 629892 995574
rect 630140 995438 630568 995466
rect 631520 995438 631856 995466
rect 634004 995438 634340 995466
rect 635200 995438 635536 995466
rect 635844 995438 636180 995466
rect 638572 995438 638908 995466
rect 630140 995330 630168 995438
rect 629864 995302 630168 995330
rect 631520 994537 631548 995438
rect 634004 994566 634032 995438
rect 635200 994809 635228 995438
rect 635844 995353 635872 995438
rect 635830 995344 635886 995353
rect 635830 995279 635886 995288
rect 635186 994800 635242 994809
rect 635186 994735 635242 994744
rect 633992 994560 634044 994566
rect 631506 994528 631562 994537
rect 633992 994502 634044 994508
rect 631506 994463 631562 994472
rect 627918 994256 627974 994265
rect 627918 994191 627974 994200
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 638880 992322 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640720 995438 641056 995466
rect 639064 994838 639092 995438
rect 639524 995110 639552 995438
rect 639512 995104 639564 995110
rect 639512 995046 639564 995052
rect 640720 994974 640748 995438
rect 660578 995072 660634 995081
rect 660578 995007 660580 995016
rect 660632 995007 660634 995016
rect 660580 994977 660632 994983
rect 640708 994968 640760 994974
rect 640708 994910 640760 994916
rect 639052 994832 639104 994838
rect 639052 994774 639104 994780
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993682 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660960 993818 660988 994502
rect 660948 993812 661000 993818
rect 660948 993754 661000 993760
rect 660764 993676 660816 993682
rect 660764 993618 660816 993624
rect 660304 993064 660356 993070
rect 660304 993006 660356 993012
rect 638868 992316 638920 992322
rect 638868 992258 638920 992264
rect 640800 992316 640852 992322
rect 640800 992258 640852 992264
rect 572720 989528 572772 989534
rect 572720 989470 572772 989476
rect 576308 989528 576360 989534
rect 576308 989470 576360 989476
rect 566464 986128 566516 986134
rect 566464 986070 566516 986076
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 989470
rect 608784 987420 608836 987426
rect 608784 987362 608836 987368
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608796 983620 608824 987362
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 624988 983620 625016 985934
rect 640812 983634 640840 992258
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 660316 937281 660344 993006
rect 668584 992928 668636 992934
rect 668584 992870 668636 992876
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660302 937272 660358 937281
rect 660302 937207 660358 937216
rect 661696 937038 661724 957743
rect 663064 948116 663116 948122
rect 663064 948058 663116 948064
rect 663076 941769 663104 948058
rect 663062 941760 663118 941769
rect 663062 941695 663118 941704
rect 665836 939865 665864 961862
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 668596 937553 668624 992870
rect 669964 990140 670016 990146
rect 669964 990082 670016 990088
rect 669976 938505 670004 990082
rect 672724 975724 672776 975730
rect 672724 975666 672776 975672
rect 672736 947345 672764 975666
rect 673366 966648 673422 966657
rect 673366 966583 673422 966592
rect 675114 966648 675170 966657
rect 675114 966583 675170 966592
rect 673182 960800 673238 960809
rect 673182 960735 673238 960744
rect 672998 952232 673054 952241
rect 672998 952167 673054 952176
rect 672722 947336 672778 947345
rect 672722 947271 672778 947280
rect 673012 943934 673040 952167
rect 673196 943934 673224 960735
rect 673012 943906 673132 943934
rect 673196 943906 673316 943934
rect 669962 938496 670018 938505
rect 669962 938431 670018 938440
rect 671802 938088 671858 938097
rect 671802 938023 671858 938032
rect 671618 937816 671674 937825
rect 671618 937751 671674 937760
rect 668582 937544 668638 937553
rect 668582 937479 668638 937488
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 670698 929520 670754 929529
rect 670698 929455 670754 929464
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 663064 921868 663116 921874
rect 663064 921810 663116 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 55862 892800 55918 892809
rect 55862 892735 55918 892744
rect 54482 892528 54538 892537
rect 54482 892463 54538 892472
rect 53286 892256 53342 892265
rect 53286 892191 53342 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62762 858664 62818 858673
rect 62762 858599 62818 858608
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799368 53158 799377
rect 53102 799303 53158 799312
rect 53104 793620 53156 793626
rect 53104 793562 53156 793568
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 669352 49018 669361
rect 48962 669287 49018 669296
rect 47872 634786 47992 634814
rect 47766 614136 47822 614145
rect 47766 614071 47822 614080
rect 47964 611726 47992 634786
rect 50356 626657 50384 714818
rect 51736 691393 51764 753510
rect 53116 730153 53144 793562
rect 54496 774353 54524 844562
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 55876 772857 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 62118 793591 62120 793600
rect 62172 793591 62174 793600
rect 62120 793562 62172 793568
rect 62776 788633 62804 858599
rect 652390 856352 652446 856361
rect 652390 856287 652446 856296
rect 652404 855642 652432 856287
rect 652392 855636 652444 855642
rect 652392 855578 652444 855584
rect 651838 843024 651894 843033
rect 651838 842959 651894 842968
rect 651852 841838 651880 842959
rect 651840 841832 651892 841838
rect 651840 841774 651892 841780
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 55862 772848 55918 772857
rect 55862 772783 55918 772792
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62776 743073 62804 780399
rect 652390 776656 652446 776665
rect 652390 776591 652446 776600
rect 652404 775606 652432 776591
rect 652392 775600 652444 775606
rect 652392 775542 652444 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 53102 730144 53158 730153
rect 53102 730079 53158 730088
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 51724 674892 51776 674898
rect 51724 674834 51776 674840
rect 51736 646649 51764 674834
rect 51722 646640 51778 646649
rect 51722 646575 51778 646584
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 652022 736808 652078 736817
rect 652022 736743 652078 736752
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 55876 643249 55904 701014
rect 62776 697921 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 651470 710288 651526 710297
rect 651470 710223 651526 710232
rect 651484 709374 651512 710223
rect 651472 709368 651524 709374
rect 651472 709310 651524 709316
rect 62762 697912 62818 697921
rect 62762 697847 62818 697856
rect 651472 696992 651524 696998
rect 651470 696960 651472 696969
rect 651524 696960 651526 696969
rect 651470 696895 651526 696904
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 651654 683632 651710 683641
rect 651654 683567 651710 683576
rect 651668 683194 651696 683567
rect 651656 683188 651708 683194
rect 651656 683130 651708 683136
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 651470 670440 651526 670449
rect 651470 670375 651526 670384
rect 651484 669390 651512 670375
rect 651472 669384 651524 669390
rect 651472 669326 651524 669332
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 651470 657112 651526 657121
rect 651470 657047 651526 657056
rect 651484 656946 651512 657047
rect 651472 656940 651524 656946
rect 651472 656882 651524 656888
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 50342 626648 50398 626657
rect 50342 626583 50398 626592
rect 50344 623824 50396 623830
rect 50344 623766 50396 623772
rect 47952 611720 48004 611726
rect 47952 611662 48004 611668
rect 50356 601361 50384 623766
rect 51736 601769 51764 636210
rect 651470 630592 651526 630601
rect 651470 630527 651526 630536
rect 651484 629338 651512 630527
rect 651472 629332 651524 629338
rect 651472 629274 651524 629280
rect 652036 627881 652064 736743
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 661684 815652 661736 815658
rect 661684 815594 661736 815600
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 652022 627872 652078 627881
rect 652022 627807 652078 627816
rect 660316 625297 660344 763166
rect 661696 673169 661724 815594
rect 663076 760481 663104 921810
rect 665824 909492 665876 909498
rect 665824 909434 665876 909440
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868737 664484 881826
rect 664442 868728 664498 868737
rect 664442 868663 664498 868672
rect 664444 855636 664496 855642
rect 664444 855578 664496 855584
rect 663062 760472 663118 760481
rect 663062 760407 663118 760416
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 661868 696992 661920 696998
rect 661868 696934 661920 696940
rect 661682 673160 661738 673169
rect 661682 673095 661738 673104
rect 661684 669384 661736 669390
rect 661684 669326 661736 669332
rect 661696 643793 661724 669326
rect 661682 643784 661738 643793
rect 661682 643719 661738 643728
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 50342 601352 50398 601361
rect 50342 601287 50398 601296
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 582448 47638 582457
rect 47582 582383 47638 582392
rect 45020 582346 45232 582374
rect 44822 556472 44878 556481
rect 44822 556407 44878 556416
rect 44822 556064 44878 556073
rect 44822 555999 44878 556008
rect 44836 555506 44864 555999
rect 45020 555665 45048 582346
rect 48976 557841 49004 597518
rect 51724 583772 51776 583778
rect 51724 583714 51776 583720
rect 48962 557832 49018 557841
rect 48962 557767 49018 557776
rect 51736 557569 51764 583714
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 51722 557560 51778 557569
rect 51722 557495 51778 557504
rect 45558 556880 45614 556889
rect 45558 556815 45614 556824
rect 45006 555656 45062 555665
rect 45006 555591 45062 555600
rect 44836 555478 44956 555506
rect 44362 555248 44418 555257
rect 44362 555183 44418 555192
rect 44178 548720 44234 548729
rect 44178 548655 44234 548664
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43640 379514 43668 547703
rect 43810 547088 43866 547097
rect 43810 547023 43866 547032
rect 43456 379486 43576 379514
rect 43640 379486 43760 379514
rect 42982 379400 43038 379409
rect 42982 379335 43038 379344
rect 42996 365809 43024 379335
rect 43350 371920 43406 371929
rect 43350 371855 43406 371864
rect 42982 365800 43038 365809
rect 42982 365735 43038 365744
rect 42536 356646 42840 356674
rect 42536 356606 42564 356646
rect 42168 356538 42196 356592
rect 42260 356578 42564 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 42430 356144 42486 356153
rect 42430 356079 42486 356088
rect 42444 355926 42472 356079
rect 42182 355898 42472 355926
rect 43364 355881 43392 371855
rect 43350 355872 43406 355881
rect 43350 355807 43406 355816
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 43548 355314 43576 379486
rect 43732 355586 43760 379486
rect 43824 355722 43852 547023
rect 44192 535265 44220 548655
rect 44178 535256 44234 535265
rect 44178 535191 44234 535200
rect 44376 428097 44404 555183
rect 44730 554432 44786 554441
rect 44730 554367 44786 554376
rect 44546 550760 44602 550769
rect 44546 550695 44602 550704
rect 44560 532817 44588 550695
rect 44546 532808 44602 532817
rect 44546 532743 44602 532752
rect 44362 428088 44418 428097
rect 44362 428023 44418 428032
rect 44454 427680 44510 427689
rect 44454 427615 44510 427624
rect 44270 426864 44326 426873
rect 44270 426799 44326 426808
rect 43994 419520 44050 419529
rect 43994 419455 44050 419464
rect 44008 355858 44036 419455
rect 44284 384033 44312 426799
rect 44468 384849 44496 427615
rect 44744 427281 44772 554367
rect 44928 428913 44956 555478
rect 45098 551576 45154 551585
rect 45098 551511 45154 551520
rect 45112 529689 45140 551511
rect 45282 549128 45338 549137
rect 45282 549063 45338 549072
rect 45296 534449 45324 549063
rect 45282 534440 45338 534449
rect 45282 534375 45338 534384
rect 45098 529680 45154 529689
rect 45098 529615 45154 529624
rect 45572 429729 45600 556815
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 45558 429720 45614 429729
rect 45558 429655 45614 429664
rect 45190 429312 45246 429321
rect 45190 429247 45246 429256
rect 44914 428904 44970 428913
rect 44914 428839 44970 428848
rect 45006 428496 45062 428505
rect 45006 428431 45062 428440
rect 44730 427272 44786 427281
rect 44730 427207 44786 427216
rect 44638 422512 44694 422521
rect 44638 422447 44694 422456
rect 44652 407153 44680 422447
rect 44822 420744 44878 420753
rect 44822 420679 44878 420688
rect 44638 407144 44694 407153
rect 44638 407079 44694 407088
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44454 384840 44510 384849
rect 44454 384775 44510 384784
rect 44270 384024 44326 384033
rect 44270 383959 44326 383968
rect 44454 379944 44510 379953
rect 44454 379879 44510 379888
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 44284 356697 44312 377431
rect 44468 359961 44496 379879
rect 44652 379514 44680 385183
rect 44836 379514 44864 420679
rect 45020 385665 45048 428431
rect 45204 386753 45232 429247
rect 45374 418296 45430 418305
rect 45374 418231 45430 418240
rect 45388 406881 45416 418231
rect 45374 406872 45430 406881
rect 45374 406807 45430 406816
rect 45190 386744 45246 386753
rect 45190 386679 45246 386688
rect 45190 386064 45246 386073
rect 45190 385999 45246 386008
rect 45006 385656 45062 385665
rect 45006 385591 45062 385600
rect 45204 385506 45232 385999
rect 45020 385478 45232 385506
rect 44652 379486 44772 379514
rect 44836 379486 44956 379514
rect 44744 360194 44772 379486
rect 44744 360166 44864 360194
rect 44454 359952 44510 359961
rect 44454 359887 44510 359896
rect 44270 356688 44326 356697
rect 44270 356623 44326 356632
rect 44008 355830 44312 355858
rect 44284 355722 44312 355830
rect 43824 355694 44220 355722
rect 44284 355706 44680 355722
rect 44284 355700 44692 355706
rect 44284 355694 44640 355700
rect 44192 355586 44220 355694
rect 44640 355642 44692 355648
rect 43732 355558 43944 355586
rect 44192 355558 44772 355586
rect 43916 355450 43944 355558
rect 43916 355422 44128 355450
rect 43548 355286 44036 355314
rect 44008 354634 44036 355286
rect 44100 354906 44128 355422
rect 44100 354890 44615 354906
rect 44100 354884 44627 354890
rect 44100 354878 44575 354884
rect 44575 354826 44627 354832
rect 44575 354680 44627 354686
rect 44008 354628 44575 354634
rect 44008 354622 44627 354628
rect 44008 354606 44615 354622
rect 44744 354498 44772 355558
rect 44836 354634 44864 360166
rect 44928 357434 44956 379486
rect 45020 360194 45048 385478
rect 45190 384432 45246 384441
rect 45190 384367 45246 384376
rect 45204 379514 45232 384367
rect 45374 383616 45430 383625
rect 45374 383551 45430 383560
rect 45204 379486 45324 379514
rect 45020 360166 45232 360194
rect 44928 357406 45048 357434
rect 45020 355842 45048 357406
rect 45008 355836 45060 355842
rect 45008 355778 45060 355784
rect 44836 354606 44956 354634
rect 44744 354482 44839 354498
rect 44744 354476 44851 354482
rect 44744 354470 44799 354476
rect 44799 354418 44851 354424
rect 44686 354340 44738 354346
rect 44686 354282 44738 354288
rect 43902 354240 43958 354249
rect 44698 354226 44726 354282
rect 43958 354198 44726 354226
rect 43902 354175 43958 354184
rect 44730 353832 44786 353841
rect 44928 353818 44956 354606
rect 45204 354090 45232 360166
rect 44786 353790 44956 353818
rect 45020 354062 45232 354090
rect 44730 353767 44786 353776
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 38290 346352 38346 346361
rect 38290 346287 38346 346296
rect 38304 345098 38332 346287
rect 28908 345092 28960 345098
rect 28908 345034 28960 345040
rect 38292 345092 38344 345098
rect 38292 345034 38344 345040
rect 28920 344321 28948 345034
rect 28906 344312 28962 344321
rect 28906 344247 28962 344256
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 45020 343369 45048 354062
rect 45006 343360 45062 343369
rect 45006 343295 45062 343304
rect 45296 341737 45324 379486
rect 45388 345014 45416 383551
rect 45558 380352 45614 380361
rect 45558 380287 45614 380296
rect 45572 357377 45600 380287
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 426456 46994 426465
rect 46938 426391 46994 426400
rect 46952 399809 46980 426391
rect 47122 423600 47178 423609
rect 47122 423535 47178 423544
rect 47136 400217 47164 423535
rect 47122 400208 47178 400217
rect 47122 400143 47178 400152
rect 46938 399800 46994 399809
rect 46938 399735 46994 399744
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 46938 380760 46994 380769
rect 46938 380695 46994 380704
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 46388 362976 46440 362982
rect 46388 362918 46440 362924
rect 45558 357368 45614 357377
rect 45558 357303 45614 357312
rect 45650 356688 45706 356697
rect 45480 356646 45650 356674
rect 45480 353274 45508 356646
rect 45650 356623 45706 356632
rect 45926 355872 45982 355881
rect 45652 355836 45704 355842
rect 45926 355807 45982 355816
rect 45652 355778 45704 355784
rect 45664 354074 45692 355778
rect 45652 354068 45704 354074
rect 45652 354010 45704 354016
rect 45940 353802 45968 355807
rect 45928 353796 45980 353802
rect 45928 353738 45980 353744
rect 45480 353258 45600 353274
rect 45480 353252 45612 353258
rect 45480 353246 45560 353252
rect 45560 353194 45612 353200
rect 45388 344986 45508 345014
rect 45282 341728 45338 341737
rect 45282 341663 45338 341672
rect 45282 341320 45338 341329
rect 45282 341255 45338 341264
rect 45296 340762 45324 341255
rect 45480 340921 45508 344986
rect 45466 340912 45522 340921
rect 45466 340847 45522 340856
rect 45296 340734 45508 340762
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37924 339516 37976 339522
rect 37924 339458 37976 339464
rect 34426 338600 34482 338609
rect 34426 338535 34482 338544
rect 34440 336161 34468 338535
rect 34426 336152 34482 336161
rect 34426 336087 34482 336096
rect 37936 328409 37964 339458
rect 43074 334656 43130 334665
rect 43074 334591 43130 334600
rect 43626 334656 43682 334665
rect 43626 334591 43682 334600
rect 44270 334656 44326 334665
rect 44270 334591 44326 334600
rect 42798 334384 42854 334393
rect 42798 334319 42854 334328
rect 37922 328400 37978 328409
rect 37922 328335 37978 328344
rect 41786 326768 41842 326777
rect 41786 326703 41842 326712
rect 41800 326264 41828 326703
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42472 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42444 321473 42472 323734
rect 42430 321464 42486 321473
rect 42430 321399 42486 321408
rect 42182 321354 42288 321382
rect 42260 321314 42288 321354
rect 42812 321314 42840 334319
rect 43088 325694 43116 334591
rect 42260 321286 42840 321314
rect 42904 325666 43116 325694
rect 42904 320770 42932 325666
rect 43442 323096 43498 323105
rect 43442 323031 43498 323040
rect 42536 320742 42932 320770
rect 42536 320739 42564 320742
rect 42182 320711 42564 320739
rect 42430 320104 42486 320113
rect 42182 320062 42430 320090
rect 42430 320039 42486 320048
rect 42182 319518 42472 319546
rect 42444 319433 42472 319518
rect 42430 319424 42486 319433
rect 42430 319359 42486 319368
rect 42246 317520 42302 317529
rect 42246 317455 42302 317464
rect 42260 317059 42288 317455
rect 42182 317031 42288 317059
rect 41786 316704 41842 316713
rect 41786 316639 41842 316648
rect 41800 316404 41828 316639
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42154 312352 42210 312361
rect 42154 312287 42210 312296
rect 42168 312052 42196 312287
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 42890 299704 42946 299713
rect 42890 299639 42946 299648
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 41326 296032 41382 296041
rect 41326 295967 41382 295976
rect 32402 294808 32458 294817
rect 32402 294743 32458 294752
rect 32416 284986 32444 294743
rect 41340 291394 41368 295967
rect 41800 292505 41828 296783
rect 41786 292496 41842 292505
rect 41786 292431 41842 292440
rect 41340 291366 41460 291394
rect 41432 290442 41460 291366
rect 41786 290456 41842 290465
rect 41432 290414 41786 290442
rect 41786 290391 41842 290400
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 285122 41368 290255
rect 41328 285116 41380 285122
rect 41328 285058 41380 285064
rect 41696 285116 41748 285122
rect 41748 285076 42380 285104
rect 41696 285058 41748 285064
rect 32404 284980 32456 284986
rect 32404 284922 32456 284928
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42288 284866
rect 42260 283059 42288 284838
rect 42182 283031 42288 283059
rect 42352 281874 42380 285076
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42430 278695 42486 278704
rect 42338 278488 42394 278497
rect 42338 278423 42394 278432
rect 42168 277953 42196 278188
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 42154 277944 42210 277953
rect 42154 277879 42210 277888
rect 41800 277508 41828 277879
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42062 273456 42118 273465
rect 42062 273391 42118 273400
rect 42076 273224 42104 273391
rect 42062 273048 42118 273057
rect 42062 272983 42118 272992
rect 42076 272544 42104 272983
rect 42352 272014 42380 278423
rect 42182 271986 42380 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 42430 270464 42486 270473
rect 42430 270399 42486 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 270399
rect 42182 269507 42472 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 35806 259992 35862 260001
rect 35806 259927 35862 259936
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35820 258369 35848 259927
rect 35806 258360 35862 258369
rect 35806 258295 35862 258304
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 42904 256873 42932 299639
rect 43258 298888 43314 298897
rect 43258 298823 43314 298832
rect 43074 295216 43130 295225
rect 43074 295151 43130 295160
rect 43088 276593 43116 295151
rect 43074 276584 43130 276593
rect 43074 276519 43130 276528
rect 42890 256864 42946 256873
rect 42890 256799 42946 256808
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42798 256456 42854 256465
rect 42798 256391 42854 256400
rect 35438 253464 35494 253473
rect 35438 253399 35494 253408
rect 35452 252618 35480 253399
rect 35622 253056 35678 253065
rect 35622 252991 35678 253000
rect 39028 253020 39080 253026
rect 35636 252754 35664 252991
rect 39028 252962 39080 252968
rect 41512 253020 41564 253026
rect 41512 252962 41564 252968
rect 35808 252884 35860 252890
rect 35808 252826 35860 252832
rect 35624 252748 35676 252754
rect 35624 252690 35676 252696
rect 35820 252657 35848 252826
rect 39040 252754 39068 252962
rect 40684 252884 40736 252890
rect 40684 252826 40736 252832
rect 39028 252748 39080 252754
rect 39028 252690 39080 252696
rect 35806 252648 35862 252657
rect 35440 252612 35492 252618
rect 35806 252583 35862 252592
rect 35440 252554 35492 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 36544 251252 36596 251258
rect 36544 251194 36596 251200
rect 36556 242894 36584 251194
rect 36544 242888 36596 242894
rect 40696 242865 40724 252826
rect 36544 242830 36596 242836
rect 40682 242856 40738 242865
rect 40682 242791 40738 242800
rect 41524 242706 41552 252962
rect 41696 252544 41748 252550
rect 41748 252492 42472 252498
rect 41696 252486 42472 252492
rect 41708 252470 42472 252486
rect 42444 248414 42472 252470
rect 42444 248386 42656 248414
rect 42260 242950 42472 242978
rect 41696 242888 41748 242894
rect 42260 242842 42288 242950
rect 41748 242836 42288 242842
rect 41696 242830 42288 242836
rect 41708 242814 42288 242830
rect 41524 242678 42288 242706
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42260 238754 42288 242678
rect 42260 238726 42380 238754
rect 42168 238513 42196 238649
rect 42154 238504 42210 238513
rect 42154 238439 42210 238448
rect 42352 238014 42380 238726
rect 42182 237986 42380 238014
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42246 235920 42302 235929
rect 42246 235855 42302 235864
rect 42260 234983 42288 235855
rect 42182 234955 42288 234983
rect 42246 234560 42302 234569
rect 42246 234495 42302 234504
rect 42260 234342 42288 234495
rect 42182 234314 42288 234342
rect 42246 234152 42302 234161
rect 42246 234087 42302 234096
rect 42260 233695 42288 234087
rect 42182 233667 42288 233695
rect 42154 233336 42210 233345
rect 42154 233271 42210 233280
rect 42168 233104 42196 233271
rect 42246 231704 42302 231713
rect 42246 231639 42302 231648
rect 42260 230670 42288 231639
rect 42182 230642 42288 230670
rect 42154 230208 42210 230217
rect 42154 230143 42210 230152
rect 42168 229976 42196 230143
rect 42246 229936 42302 229945
rect 42246 229871 42302 229880
rect 42260 229378 42288 229871
rect 42182 229350 42288 229378
rect 42444 228834 42472 242950
rect 42628 237425 42656 248386
rect 42614 237416 42670 237425
rect 42614 237351 42670 237360
rect 42182 228806 42472 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 40682 222864 40738 222873
rect 40682 222799 40738 222808
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214305 35572 217903
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 40696 213994 40724 222799
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 40684 213988 40736 213994
rect 40684 213930 40736 213936
rect 42812 213761 42840 256391
rect 43272 256057 43300 298823
rect 43456 257689 43484 323031
rect 43640 322833 43668 334591
rect 43626 322824 43682 322833
rect 43626 322759 43682 322768
rect 44284 320113 44312 334591
rect 44270 320104 44326 320113
rect 44270 320039 44326 320048
rect 44178 311536 44234 311545
rect 44178 311471 44234 311480
rect 44192 299305 44220 311471
rect 44362 311264 44418 311273
rect 44362 311199 44418 311208
rect 44376 300121 44404 311199
rect 44362 300112 44418 300121
rect 44362 300047 44418 300056
rect 44178 299296 44234 299305
rect 44178 299231 44234 299240
rect 45480 298489 45508 340734
rect 45834 340096 45890 340105
rect 45834 340031 45890 340040
rect 45650 339280 45706 339289
rect 45650 339215 45706 339224
rect 45664 312361 45692 339215
rect 45848 313721 45876 340031
rect 46018 338464 46074 338473
rect 46018 338399 46074 338408
rect 46032 319433 46060 338399
rect 46018 319424 46074 319433
rect 46018 319359 46074 319368
rect 45834 313712 45890 313721
rect 45834 313647 45890 313656
rect 45650 312352 45706 312361
rect 45650 312287 45706 312296
rect 46400 303113 46428 362918
rect 46952 356153 46980 380695
rect 47122 379128 47178 379137
rect 47122 379063 47178 379072
rect 47136 361593 47164 379063
rect 47122 361584 47178 361593
rect 47122 361519 47178 361528
rect 46938 356144 46994 356153
rect 46938 356079 46994 356088
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46386 303104 46442 303113
rect 46386 303039 46442 303048
rect 45466 298480 45522 298489
rect 45466 298415 45522 298424
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 44178 298072 44234 298081
rect 44178 298007 44234 298016
rect 43626 293992 43682 294001
rect 43626 293927 43682 293936
rect 43640 273057 43668 293927
rect 43994 293176 44050 293185
rect 43994 293111 44050 293120
rect 43810 291952 43866 291961
rect 43810 291887 43866 291896
rect 43824 277137 43852 291887
rect 44008 279857 44036 293111
rect 43994 279848 44050 279857
rect 43994 279783 44050 279792
rect 43810 277128 43866 277137
rect 43810 277063 43866 277072
rect 43626 273048 43682 273057
rect 43626 272983 43682 272992
rect 43442 257680 43498 257689
rect 43442 257615 43498 257624
rect 43258 256048 43314 256057
rect 43258 255983 43314 255992
rect 43626 255640 43682 255649
rect 43626 255575 43682 255584
rect 42982 254824 43038 254833
rect 42982 254759 43038 254768
rect 42798 213752 42854 213761
rect 42798 213687 42854 213696
rect 42996 212129 43024 254759
rect 43442 251152 43498 251161
rect 43442 251087 43498 251096
rect 43258 242856 43314 242865
rect 43258 242791 43314 242800
rect 43272 225729 43300 242791
rect 43456 226681 43484 251087
rect 43640 251002 43668 255575
rect 44192 255241 44220 298007
rect 45480 297378 45508 298114
rect 44836 297350 45508 297378
rect 44362 294400 44418 294409
rect 44362 294335 44418 294344
rect 44376 270473 44404 294335
rect 44638 293584 44694 293593
rect 44638 293519 44694 293528
rect 44652 273465 44680 293519
rect 44638 273456 44694 273465
rect 44638 273391 44694 273400
rect 44362 270464 44418 270473
rect 44362 270399 44418 270408
rect 44178 255232 44234 255241
rect 44178 255167 44234 255176
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43548 250974 43668 251002
rect 43548 229094 43576 250974
rect 43718 249112 43774 249121
rect 43718 249047 43774 249056
rect 43732 231713 43760 249047
rect 43718 231704 43774 231713
rect 43718 231639 43774 231648
rect 43548 229066 43668 229094
rect 43442 226672 43498 226681
rect 43442 226607 43498 226616
rect 43258 225720 43314 225729
rect 43258 225655 43314 225664
rect 43442 213344 43498 213353
rect 43442 213279 43498 213288
rect 42982 212120 43038 212129
rect 42982 212055 43038 212064
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35820 211206 35848 211375
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 41696 211200 41748 211206
rect 41696 211142 41748 211148
rect 41708 209001 41736 211142
rect 42798 209672 42854 209681
rect 42798 209607 42854 209616
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 41694 208992 41750 209001
rect 41694 208927 41750 208936
rect 35820 208418 35848 208927
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 207777 40080 208354
rect 40038 207768 40094 207777
rect 40038 207703 40094 207712
rect 35622 204096 35678 204105
rect 35622 204031 35678 204040
rect 35636 202201 35664 204031
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 35622 202192 35678 202201
rect 35622 202127 35678 202136
rect 37936 197849 37964 202846
rect 37922 197840 37978 197849
rect 37922 197775 37978 197784
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 41878 195800 41934 195809
rect 41878 195735 41934 195744
rect 41892 195432 41920 195735
rect 42614 195528 42670 195537
rect 42614 195463 42670 195472
rect 41970 195256 42026 195265
rect 41970 195191 42026 195200
rect 41984 194820 42012 195191
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42628 192953 42656 195463
rect 42168 192902 42288 192930
rect 42614 192944 42670 192953
rect 42614 192879 42670 192888
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41786 187232 41842 187241
rect 41786 187167 41842 187176
rect 41800 186796 41828 187167
rect 42338 186280 42394 186289
rect 42338 186215 42394 186224
rect 42168 186130 42196 186184
rect 42352 186130 42380 186215
rect 42168 186102 42380 186130
rect 41786 185872 41842 185881
rect 41786 185807 41842 185816
rect 41800 185605 41828 185807
rect 42430 184920 42486 184929
rect 42430 184855 42486 184864
rect 42444 183779 42472 184855
rect 42182 183751 42472 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42812 182491 42840 209607
rect 43258 208040 43314 208049
rect 43258 207975 43314 207984
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 183161 43300 207975
rect 43456 206281 43484 213279
rect 43640 212945 43668 229066
rect 43626 212936 43682 212945
rect 43626 212871 43682 212880
rect 44192 211313 44220 253943
rect 44638 251968 44694 251977
rect 44638 251903 44694 251912
rect 44652 251818 44680 251903
rect 44652 251790 44772 251818
rect 44546 248704 44602 248713
rect 44546 248639 44602 248648
rect 44362 248296 44418 248305
rect 44362 248231 44418 248240
rect 44376 235929 44404 248231
rect 44362 235920 44418 235929
rect 44362 235855 44418 235864
rect 44560 234342 44588 248639
rect 44744 238754 44772 251790
rect 44468 234314 44588 234342
rect 44652 238726 44772 238754
rect 44468 234161 44496 234314
rect 44454 234152 44510 234161
rect 44454 234087 44510 234096
rect 44652 233345 44680 238726
rect 44638 233336 44694 233345
rect 44638 233271 44694 233280
rect 44836 214985 44864 297350
rect 45006 297256 45062 297265
rect 45006 297191 45062 297200
rect 45020 254425 45048 297191
rect 45190 291680 45246 291689
rect 45190 291615 45246 291624
rect 45204 277953 45232 291615
rect 46202 290728 46258 290737
rect 46202 290663 46258 290672
rect 45190 277944 45246 277953
rect 45190 277879 45246 277888
rect 45006 254416 45062 254425
rect 45006 254351 45062 254360
rect 45558 250744 45614 250753
rect 45558 250679 45614 250688
rect 45572 229945 45600 250679
rect 45834 250336 45890 250345
rect 45834 250271 45890 250280
rect 45848 230217 45876 250271
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 234569 46060 249455
rect 46018 234560 46074 234569
rect 46018 234495 46074 234504
rect 45834 230208 45890 230217
rect 45834 230143 45890 230152
rect 45558 229936 45614 229945
rect 45558 229871 45614 229880
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 44178 211304 44234 211313
rect 44178 211239 44234 211248
rect 45006 210896 45062 210905
rect 45006 210831 45062 210840
rect 44178 210488 44234 210497
rect 44178 210423 44234 210432
rect 43626 206816 43682 206825
rect 43626 206751 43682 206760
rect 43442 206272 43498 206281
rect 43442 206207 43498 206216
rect 43442 202192 43498 202201
rect 43442 202127 43498 202136
rect 43258 183152 43314 183161
rect 43258 183087 43314 183096
rect 42182 182463 42840 182491
rect 43456 42838 43484 202127
rect 43640 193225 43668 206751
rect 43810 205592 43866 205601
rect 43810 205527 43866 205536
rect 43626 193216 43682 193225
rect 43626 193151 43682 193160
rect 43824 190505 43852 205527
rect 43994 205184 44050 205193
rect 43994 205119 44050 205128
rect 44008 191729 44036 205119
rect 43994 191720 44050 191729
rect 43994 191655 44050 191664
rect 43810 190496 43866 190505
rect 43810 190431 43866 190440
rect 44192 184929 44220 210423
rect 45020 209774 45048 210831
rect 45020 209746 45508 209774
rect 44362 208584 44418 208593
rect 44362 208519 44418 208528
rect 44376 189961 44404 208519
rect 44546 206000 44602 206009
rect 44546 205935 44602 205944
rect 44362 189952 44418 189961
rect 44362 189887 44418 189896
rect 44560 187649 44588 205935
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44546 187640 44602 187649
rect 44546 187575 44602 187584
rect 44178 184920 44234 184929
rect 44178 184855 44234 184864
rect 44836 74534 44864 204711
rect 45480 196654 45508 209746
rect 45468 196648 45520 196654
rect 45468 196590 45520 196596
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 290663
rect 46938 247072 46994 247081
rect 46938 247007 46994 247016
rect 46952 238513 46980 247007
rect 46938 238504 46994 238513
rect 46938 238439 46994 238448
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 47596 49026 47624 333095
rect 47780 300529 47808 389234
rect 48976 387025 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 49148 415472 49200 415478
rect 49148 415414 49200 415420
rect 48962 387016 49018 387025
rect 48962 386951 49018 386960
rect 49160 346361 49188 415414
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51724 375420 51776 375426
rect 51724 375362 51776 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 49146 346352 49202 346361
rect 49146 346287 49202 346296
rect 50344 336796 50396 336802
rect 50344 336738 50396 336744
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47780 53242 47808 247415
rect 47950 212528 48006 212537
rect 47950 212463 48006 212472
rect 47964 192409 47992 212463
rect 48596 196648 48648 196654
rect 48596 196590 48648 196596
rect 48608 194449 48636 196590
rect 48594 194440 48650 194449
rect 48594 194375 48650 194384
rect 47950 192400 48006 192409
rect 47950 192335 48006 192344
rect 47768 53236 47820 53242
rect 47768 53178 47820 53184
rect 48976 51882 49004 334047
rect 49146 289912 49202 289921
rect 49146 289847 49202 289856
rect 48964 51876 49016 51882
rect 48964 51818 49016 51824
rect 49160 51746 49188 289847
rect 50356 260001 50384 336738
rect 51736 301345 51764 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 660316 599593 660344 616830
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 652390 590744 652446 590753
rect 652390 590679 652392 590688
rect 652444 590679 652446 590688
rect 658924 590708 658976 590714
rect 652392 590650 652444 590656
rect 658924 590650 658976 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 652574 497720 652630 497729
rect 652574 497655 652630 497664
rect 652588 494766 652616 497655
rect 652576 494760 652628 494766
rect 652576 494702 652628 494708
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 658936 492017 658964 590650
rect 661880 581097 661908 696934
rect 663076 689353 663104 723114
rect 664456 716553 664484 855578
rect 665836 761569 665864 909434
rect 669226 879200 669282 879209
rect 669226 879135 669282 879144
rect 668766 877704 668822 877713
rect 668766 877639 668822 877648
rect 667846 866688 667902 866697
rect 667846 866623 667902 866632
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666466 778424 666522 778433
rect 666466 778359 666522 778368
rect 665822 761560 665878 761569
rect 665822 761495 665878 761504
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 663064 656940 663116 656946
rect 663064 656882 663116 656888
rect 661866 581088 661922 581097
rect 661866 581023 661922 581032
rect 659108 563100 659160 563106
rect 659108 563042 659160 563048
rect 659120 554033 659148 563042
rect 659106 554024 659162 554033
rect 659106 553959 659162 553968
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 658922 492008 658978 492017
rect 62120 491972 62172 491978
rect 658922 491943 658978 491952
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 53104 310548 53156 310554
rect 53104 310490 53156 310496
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 51722 289912 51778 289921
rect 51722 289847 51778 289856
rect 50342 259992 50398 260001
rect 50342 259927 50398 259936
rect 50526 247752 50582 247761
rect 50526 247687 50582 247696
rect 50342 246528 50398 246537
rect 50342 246463 50398 246472
rect 49514 208992 49570 209001
rect 49514 208927 49570 208936
rect 49330 206272 49386 206281
rect 49330 206207 49386 206216
rect 49344 190505 49372 206207
rect 49528 196489 49556 208927
rect 49514 196480 49570 196489
rect 49514 196415 49570 196424
rect 49330 190496 49386 190505
rect 49330 190431 49386 190440
rect 49148 51740 49200 51746
rect 49148 51682 49200 51688
rect 50356 50522 50384 246463
rect 50540 53378 50568 247687
rect 50710 203280 50766 203289
rect 50710 203215 50766 203224
rect 50528 53372 50580 53378
rect 50528 53314 50580 53320
rect 50724 52018 50752 203215
rect 50712 52012 50764 52018
rect 50712 51954 50764 51960
rect 50344 50516 50396 50522
rect 50344 50458 50396 50464
rect 51736 49162 51764 289847
rect 53116 217977 53144 310490
rect 55876 278769 55904 401610
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 652022 378176 652078 378185
rect 652022 378111 652078 378120
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 651654 364848 651710 364857
rect 651654 364783 651710 364792
rect 651668 364410 651696 364783
rect 651656 364404 651708 364410
rect 651656 364346 651708 364352
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 651470 351656 651526 351665
rect 651470 351591 651526 351600
rect 651484 350606 651512 351591
rect 651472 350600 651524 350606
rect 651472 350542 651524 350548
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 62776 267073 62804 350231
rect 651470 338328 651526 338337
rect 651470 338263 651526 338272
rect 651484 338162 651512 338263
rect 651472 338156 651524 338162
rect 651472 338098 651524 338104
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 651484 310554 651512 311743
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62946 285152 63002 285161
rect 62946 285087 63002 285096
rect 62762 267064 62818 267073
rect 62762 266999 62818 267008
rect 62764 228540 62816 228546
rect 62764 228482 62816 228488
rect 57704 227044 57756 227050
rect 57704 226986 57756 226992
rect 56508 222896 56560 222902
rect 56508 222838 56560 222844
rect 56324 218204 56376 218210
rect 56324 218146 56376 218152
rect 55956 218068 56008 218074
rect 55956 218010 56008 218016
rect 53102 217968 53158 217977
rect 53102 217903 53158 217912
rect 55968 217002 55996 218010
rect 55660 216974 55996 217002
rect 56336 217002 56364 218146
rect 56520 218074 56548 222838
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57716 217002 57744 226986
rect 61384 225616 61436 225622
rect 61384 225558 61436 225564
rect 60648 224528 60700 224534
rect 60648 224470 60700 224476
rect 59268 224256 59320 224262
rect 59268 224198 59320 224204
rect 58440 218068 58492 218074
rect 58440 218010 58492 218016
rect 58452 217002 58480 218010
rect 59280 217002 59308 224198
rect 60096 218748 60148 218754
rect 60096 218690 60148 218696
rect 60108 217002 60136 218690
rect 60660 217002 60688 224470
rect 61396 218074 61424 225558
rect 61752 221604 61804 221610
rect 61752 221546 61804 221552
rect 61384 218068 61436 218074
rect 61384 218010 61436 218016
rect 61764 217002 61792 221546
rect 62580 218884 62632 218890
rect 62580 218826 62632 218832
rect 62592 217002 62620 218826
rect 62776 218210 62804 228482
rect 62960 222873 62988 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 274666 65932 277780
rect 67008 274718 67036 277780
rect 66996 274712 67048 274718
rect 65904 274638 66300 274666
rect 66996 274654 67048 274660
rect 66272 268394 66300 274638
rect 68204 271318 68232 277780
rect 68192 271312 68244 271318
rect 68192 271254 68244 271260
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274990 71820 277780
rect 71780 274984 71832 274990
rect 71780 274926 71832 274932
rect 71044 274712 71096 274718
rect 71044 274654 71096 274660
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 66260 268388 66312 268394
rect 66260 268330 66312 268336
rect 71056 267034 71084 274654
rect 72988 271182 73016 277780
rect 74092 275194 74120 277780
rect 75302 277766 75868 277794
rect 74080 275188 74132 275194
rect 74080 275130 74132 275136
rect 73804 274984 73856 274990
rect 73804 274926 73856 274932
rect 72976 271176 73028 271182
rect 72976 271118 73028 271124
rect 73816 267170 73844 274926
rect 75840 269958 75868 277766
rect 76484 275602 76512 277780
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 77208 275188 77260 275194
rect 77208 275130 77260 275136
rect 77220 273970 77248 275130
rect 77208 273964 77260 273970
rect 77208 273906 77260 273912
rect 77680 272542 77708 277780
rect 78876 272950 78904 277780
rect 78864 272944 78916 272950
rect 78864 272886 78916 272892
rect 77668 272536 77720 272542
rect 77668 272478 77720 272484
rect 80072 270094 80100 277780
rect 81268 275738 81296 277780
rect 81256 275732 81308 275738
rect 81256 275674 81308 275680
rect 82372 274242 82400 277780
rect 83582 277766 84148 277794
rect 82360 274236 82412 274242
rect 82360 274178 82412 274184
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 84120 269686 84148 277766
rect 84764 274106 84792 277780
rect 85960 275466 85988 277780
rect 86868 275596 86920 275602
rect 86868 275538 86920 275544
rect 85948 275460 86000 275466
rect 85948 275402 86000 275408
rect 84752 274100 84804 274106
rect 84752 274042 84804 274048
rect 84108 269680 84160 269686
rect 84108 269622 84160 269628
rect 86880 268938 86908 275538
rect 87156 272678 87184 277780
rect 88352 276010 88380 277780
rect 89548 277394 89576 277780
rect 89548 277366 89668 277394
rect 88340 276004 88392 276010
rect 88340 275946 88392 275952
rect 89640 275890 89668 277366
rect 89640 275862 89760 275890
rect 88984 275732 89036 275738
rect 88984 275674 89036 275680
rect 87144 272672 87196 272678
rect 87144 272614 87196 272620
rect 86868 268932 86920 268938
rect 86868 268874 86920 268880
rect 88996 267714 89024 275674
rect 89732 271454 89760 275862
rect 90652 274718 90680 277780
rect 91862 277766 92428 277794
rect 90640 274712 90692 274718
rect 90640 274654 90692 274660
rect 89720 271448 89772 271454
rect 89720 271390 89772 271396
rect 92400 268530 92428 277766
rect 93044 271726 93072 277780
rect 94240 272814 94268 277780
rect 95436 275874 95464 277780
rect 95424 275868 95476 275874
rect 95424 275810 95476 275816
rect 96632 275602 96660 277780
rect 97750 277766 97948 277794
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 96620 275596 96672 275602
rect 96620 275538 96672 275544
rect 95884 274712 95936 274718
rect 95884 274654 95936 274660
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 93032 271720 93084 271726
rect 93032 271662 93084 271668
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 88984 267708 89036 267714
rect 88984 267650 89036 267656
rect 95896 267578 95924 274654
rect 97920 270230 97948 277766
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 99300 268666 99328 277766
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 95884 267572 95936 267578
rect 95884 267514 95936 267520
rect 100680 267306 100708 277766
rect 101324 274378 101352 277780
rect 101312 274372 101364 274378
rect 101312 274314 101364 274320
rect 102520 268802 102548 277780
rect 103716 275738 103744 277780
rect 104912 277394 104940 277780
rect 104912 277366 105032 277394
rect 104808 275868 104860 275874
rect 104808 275810 104860 275816
rect 103704 275732 103756 275738
rect 103704 275674 103756 275680
rect 104820 274650 104848 275810
rect 104808 274644 104860 274650
rect 104808 274586 104860 274592
rect 105004 273086 105032 277366
rect 106016 274786 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 274780 106056 274786
rect 106004 274722 106056 274728
rect 104992 273080 105044 273086
rect 104992 273022 105044 273028
rect 102508 268796 102560 268802
rect 102508 268738 102560 268744
rect 107580 267442 107608 277766
rect 108960 269074 108988 277766
rect 110248 270366 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 110420 274780 110472 274786
rect 110420 274722 110472 274728
rect 110432 271862 110460 274722
rect 110420 271856 110472 271862
rect 110420 271798 110472 271804
rect 111996 271590 112024 277780
rect 113192 275874 113220 277780
rect 113180 275868 113232 275874
rect 113180 275810 113232 275816
rect 114296 273222 114324 277780
rect 115506 277766 115888 277794
rect 114284 273216 114336 273222
rect 114284 273158 114336 273164
rect 111984 271584 112036 271590
rect 111984 271526 112036 271532
rect 115860 270502 115888 277766
rect 116688 270638 116716 277780
rect 117898 277766 118648 277794
rect 116676 270632 116728 270638
rect 116676 270574 116728 270580
rect 115848 270496 115900 270502
rect 115848 270438 115900 270444
rect 110236 270360 110288 270366
rect 110236 270302 110288 270308
rect 118620 269414 118648 277766
rect 119080 269550 119108 277780
rect 120290 277766 120948 277794
rect 120920 271726 120948 277766
rect 121380 274514 121408 277780
rect 122590 277766 122788 277794
rect 121368 274508 121420 274514
rect 121368 274450 121420 274456
rect 120724 271720 120776 271726
rect 120724 271662 120776 271668
rect 120908 271720 120960 271726
rect 120908 271662 120960 271668
rect 119804 269680 119856 269686
rect 119804 269622 119856 269628
rect 119068 269544 119120 269550
rect 119068 269486 119120 269492
rect 118608 269408 118660 269414
rect 118608 269350 118660 269356
rect 108948 269068 109000 269074
rect 108948 269010 109000 269016
rect 107568 267436 107620 267442
rect 107568 267378 107620 267384
rect 100668 267300 100720 267306
rect 100668 267242 100720 267248
rect 73804 267164 73856 267170
rect 73804 267106 73856 267112
rect 71044 267028 71096 267034
rect 71044 266970 71096 266976
rect 119816 266490 119844 269622
rect 120736 266762 120764 271662
rect 122760 268258 122788 277766
rect 123772 273834 123800 277780
rect 124982 277766 125548 277794
rect 126178 277766 126928 277794
rect 123760 273828 123812 273834
rect 123760 273770 123812 273776
rect 122748 268252 122800 268258
rect 122748 268194 122800 268200
rect 125520 267986 125548 277766
rect 126900 269550 126928 277766
rect 127360 272406 127388 277780
rect 127348 272400 127400 272406
rect 127348 272342 127400 272348
rect 128556 271046 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 128544 271040 128596 271046
rect 128544 270982 128596 270988
rect 130856 270910 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 270904 130896 270910
rect 130844 270846 130896 270852
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 125508 267980 125560 267986
rect 125508 267922 125560 267928
rect 132420 266898 132448 277766
rect 133800 268122 133828 277766
rect 134444 273698 134472 277780
rect 135640 275058 135668 277780
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136548 274916 136600 274922
rect 136548 274858 136600 274864
rect 134432 273692 134484 273698
rect 134432 273634 134484 273640
rect 136560 269793 136588 274858
rect 136546 269784 136602 269793
rect 136546 269719 136602 269728
rect 136836 269278 136864 277780
rect 137940 270774 137968 277780
rect 138664 272944 138716 272950
rect 138664 272886 138716 272892
rect 138480 271312 138532 271318
rect 138480 271254 138532 271260
rect 137928 270768 137980 270774
rect 137928 270710 137980 270716
rect 136824 269272 136876 269278
rect 136824 269214 136876 269220
rect 137284 268388 137336 268394
rect 137284 268330 137336 268336
rect 133788 268116 133840 268122
rect 133788 268058 133840 268064
rect 132408 266892 132460 266898
rect 132408 266834 132460 266840
rect 120724 266756 120776 266762
rect 120724 266698 120776 266704
rect 119804 266484 119856 266490
rect 119804 266426 119856 266432
rect 137296 264316 137324 268330
rect 138112 267028 138164 267034
rect 138112 266970 138164 266976
rect 138124 264316 138152 266970
rect 138492 264330 138520 271254
rect 138676 266626 138704 272886
rect 139136 272270 139164 277780
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 139124 272264 139176 272270
rect 139124 272206 139176 272212
rect 139768 269816 139820 269822
rect 139952 269816 140004 269822
rect 139768 269758 139820 269764
rect 139950 269784 139952 269793
rect 140004 269784 140006 269793
rect 138664 266620 138716 266626
rect 138664 266562 138716 266568
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 139950 269719 140006 269728
rect 140148 264330 140176 275266
rect 140332 274786 140360 277780
rect 141542 277766 141832 277794
rect 140320 274780 140372 274786
rect 140320 274722 140372 274728
rect 141804 272950 141832 277766
rect 142724 275330 142752 277780
rect 143356 276004 143408 276010
rect 143356 275946 143408 275952
rect 142712 275324 142764 275330
rect 142712 275266 142764 275272
rect 141792 272944 141844 272950
rect 141792 272886 141844 272892
rect 141608 272264 141660 272270
rect 141608 272206 141660 272212
rect 141424 267164 141476 267170
rect 141424 267106 141476 267112
rect 140148 264302 140622 264330
rect 141436 264316 141464 267106
rect 141620 267034 141648 272206
rect 142160 271176 142212 271182
rect 142160 271118 142212 271124
rect 141608 267028 141660 267034
rect 141608 266970 141660 266976
rect 142172 264330 142200 271118
rect 143368 269958 143396 275946
rect 143540 273964 143592 273970
rect 143540 273906 143592 273912
rect 142620 269952 142672 269958
rect 142620 269894 142672 269900
rect 143356 269952 143408 269958
rect 143356 269894 143408 269900
rect 142632 267734 142660 269894
rect 142632 267706 142752 267734
rect 142724 264330 142752 267706
rect 143552 264330 143580 273906
rect 143920 272270 143948 277780
rect 144644 274780 144696 274786
rect 144644 274722 144696 274728
rect 144656 273562 144684 274722
rect 145024 273970 145052 277780
rect 146220 274786 146248 277780
rect 147430 277766 147628 277794
rect 146760 275460 146812 275466
rect 146760 275402 146812 275408
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145564 274236 145616 274242
rect 145564 274178 145616 274184
rect 145012 273964 145064 273970
rect 145012 273906 145064 273912
rect 144644 273556 144696 273562
rect 144644 273498 144696 273504
rect 145104 272536 145156 272542
rect 145104 272478 145156 272484
rect 143908 272264 143960 272270
rect 143908 272206 143960 272212
rect 144736 268932 144788 268938
rect 144736 268874 144788 268880
rect 144552 267708 144604 267714
rect 144552 267650 144604 267656
rect 144564 267170 144592 267650
rect 144552 267164 144604 267170
rect 144552 267106 144604 267112
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 268874
rect 144920 267708 144972 267714
rect 144920 267650 144972 267656
rect 144932 266490 144960 267650
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 272478
rect 145576 266558 145604 274178
rect 146772 270094 146800 275402
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 146760 270088 146812 270094
rect 146760 270030 146812 270036
rect 145564 266552 145616 266558
rect 145564 266494 145616 266500
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 147600 268394 147628 277766
rect 148324 274100 148376 274106
rect 148324 274042 148376 274048
rect 147588 268388 147640 268394
rect 147588 268330 147640 268336
rect 147588 267980 147640 267986
rect 147588 267922 147640 267928
rect 147600 267170 147628 267922
rect 147404 267164 147456 267170
rect 147404 267106 147456 267112
rect 147588 267164 147640 267170
rect 147588 267106 147640 267112
rect 147416 267050 147444 267106
rect 147416 267022 147720 267050
rect 147220 266416 147272 266422
rect 147220 266358 147272 266364
rect 147232 264316 147260 266358
rect 147692 264330 147720 267022
rect 148336 266422 148364 274042
rect 148612 271182 148640 277780
rect 149808 274922 149836 277780
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 149888 274780 149940 274786
rect 149888 274722 149940 274728
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149900 267170 149928 274722
rect 151004 271318 151032 277780
rect 152004 272672 152056 272678
rect 152004 272614 152056 272620
rect 150992 271312 151044 271318
rect 150992 271254 151044 271260
rect 151084 270632 151136 270638
rect 151084 270574 151136 270580
rect 150532 267708 150584 267714
rect 150532 267650 150584 267656
rect 149060 267164 149112 267170
rect 149060 267106 149112 267112
rect 149888 267164 149940 267170
rect 149888 267106 149940 267112
rect 149072 266626 149100 267106
rect 149060 266620 149112 266626
rect 149060 266562 149112 266568
rect 148876 266552 148928 266558
rect 148876 266494 148928 266500
rect 148324 266416 148376 266422
rect 148324 266358 148376 266364
rect 147692 264302 148074 264330
rect 148888 264316 148916 266494
rect 149704 266416 149756 266422
rect 149704 266358 149756 266364
rect 149716 264316 149744 266358
rect 150544 264316 150572 267650
rect 151096 266490 151124 270574
rect 151360 270088 151412 270094
rect 151360 270030 151412 270036
rect 151084 266484 151136 266490
rect 151084 266426 151136 266432
rect 151372 264316 151400 270030
rect 152016 264330 152044 272614
rect 152200 272542 152228 277780
rect 152188 272536 152240 272542
rect 152188 272478 152240 272484
rect 153304 272134 153332 277780
rect 153292 272128 153344 272134
rect 153292 272070 153344 272076
rect 152648 271448 152700 271454
rect 152648 271390 152700 271396
rect 152660 264330 152688 271390
rect 153844 270088 153896 270094
rect 153844 270030 153896 270036
rect 152016 264302 152214 264330
rect 152660 264302 153042 264330
rect 153856 264316 153884 270030
rect 154500 269958 154528 277780
rect 155710 277766 155908 277794
rect 154488 269952 154540 269958
rect 154488 269894 154540 269900
rect 155880 268530 155908 277766
rect 156892 276010 156920 277780
rect 156880 276004 156932 276010
rect 156880 275946 156932 275952
rect 156604 275596 156656 275602
rect 156604 275538 156656 275544
rect 156052 272808 156104 272814
rect 156052 272750 156104 272756
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 155868 268524 155920 268530
rect 155868 268466 155920 268472
rect 154672 267572 154724 267578
rect 154672 267514 154724 267520
rect 154684 264316 154712 267514
rect 155512 264316 155540 268466
rect 156064 264330 156092 272750
rect 156616 266762 156644 275538
rect 157616 274644 157668 274650
rect 157616 274586 157668 274592
rect 156420 266756 156472 266762
rect 156420 266698 156472 266704
rect 156604 266756 156656 266762
rect 156604 266698 156656 266704
rect 156432 264602 156460 266698
rect 156432 264574 156736 264602
rect 156708 264330 156736 264574
rect 157628 264330 157656 274586
rect 158088 274106 158116 277780
rect 159298 277766 159956 277794
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 156064 264302 156354 264330
rect 156708 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159928 270094 159956 277766
rect 160100 275732 160152 275738
rect 160100 275674 160152 275680
rect 160112 274242 160140 275674
rect 160480 275466 160508 277780
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161584 274718 161612 277780
rect 162124 275188 162176 275194
rect 162124 275130 162176 275136
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 160928 274372 160980 274378
rect 160928 274314 160980 274320
rect 160100 274236 160152 274242
rect 160100 274178 160152 274184
rect 159916 270088 159968 270094
rect 159916 270030 159968 270036
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 159640 266756 159692 266762
rect 159640 266698 159692 266704
rect 159652 264316 159680 266698
rect 160480 264316 160508 268602
rect 160940 264330 160968 274314
rect 162136 267578 162164 275130
rect 162780 268666 162808 277780
rect 163976 275602 164004 277780
rect 163964 275596 164016 275602
rect 163964 275538 164016 275544
rect 163136 274712 163188 274718
rect 163136 274654 163188 274660
rect 163148 268802 163176 274654
rect 164240 274236 164292 274242
rect 164240 274178 164292 274184
rect 163320 273080 163372 273086
rect 163320 273022 163372 273028
rect 162952 268796 163004 268802
rect 162952 268738 163004 268744
rect 163136 268796 163188 268802
rect 163136 268738 163188 268744
rect 162768 268660 162820 268666
rect 162768 268602 162820 268608
rect 162124 267572 162176 267578
rect 162124 267514 162176 267520
rect 162124 267300 162176 267306
rect 162124 267242 162176 267248
rect 160940 264302 161322 264330
rect 162136 264316 162164 267242
rect 162964 264316 162992 268738
rect 163332 264330 163360 273022
rect 164252 264330 164280 274178
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 164988 264330 165016 271798
rect 165172 271454 165200 277780
rect 166382 277766 166948 277794
rect 165160 271448 165212 271454
rect 165160 271390 165212 271396
rect 166920 270230 166948 277766
rect 167564 273086 167592 277780
rect 167736 275460 167788 275466
rect 167736 275402 167788 275408
rect 167552 273080 167604 273086
rect 167552 273022 167604 273028
rect 166908 270224 166960 270230
rect 166908 270166 166960 270172
rect 166908 269408 166960 269414
rect 166908 269350 166960 269356
rect 166264 269068 166316 269074
rect 166264 269010 166316 269016
rect 163332 264302 163806 264330
rect 164252 264302 164634 264330
rect 164988 264302 165462 264330
rect 166276 264316 166304 269010
rect 166920 267306 166948 269350
rect 167748 267442 167776 275402
rect 168668 272678 168696 277780
rect 169878 277766 170168 277794
rect 169944 275868 169996 275874
rect 169944 275810 169996 275816
rect 169024 273216 169076 273222
rect 169024 273158 169076 273164
rect 168656 272672 168708 272678
rect 168656 272614 168708 272620
rect 168380 271584 168432 271590
rect 168380 271526 168432 271532
rect 167920 270360 167972 270366
rect 167920 270302 167972 270308
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 167736 267436 167788 267442
rect 167736 267378 167788 267384
rect 166908 267300 166960 267306
rect 166908 267242 166960 267248
rect 167104 264316 167132 267378
rect 167932 264316 167960 270302
rect 168392 264330 168420 271526
rect 169036 266762 169064 273158
rect 169576 267572 169628 267578
rect 169576 267514 169628 267520
rect 169024 266756 169076 266762
rect 169024 266698 169076 266704
rect 168392 264302 168774 264330
rect 169588 264316 169616 267514
rect 169956 264330 169984 275810
rect 170140 274718 170168 277766
rect 171060 275466 171088 277780
rect 172270 277766 172468 277794
rect 171048 275460 171100 275466
rect 171048 275402 171100 275408
rect 170128 274712 170180 274718
rect 170128 274654 170180 274660
rect 171784 272128 171836 272134
rect 171784 272070 171836 272076
rect 171232 270496 171284 270502
rect 171232 270438 171284 270444
rect 169956 264302 170430 264330
rect 171244 264316 171272 270438
rect 171796 267714 171824 272070
rect 172440 270502 172468 277766
rect 173072 274712 173124 274718
rect 173072 274654 173124 274660
rect 172428 270496 172480 270502
rect 172428 270438 172480 270444
rect 173084 270366 173112 274654
rect 173452 271590 173480 277780
rect 174662 277766 175136 277794
rect 173440 271584 173492 271590
rect 173440 271526 173492 271532
rect 173072 270360 173124 270366
rect 173072 270302 173124 270308
rect 173716 269680 173768 269686
rect 173716 269622 173768 269628
rect 171784 267708 171836 267714
rect 171784 267650 171836 267656
rect 172060 266756 172112 266762
rect 172060 266698 172112 266704
rect 172072 264316 172100 266698
rect 172888 266484 172940 266490
rect 172888 266426 172940 266432
rect 172900 264316 172928 266426
rect 173728 264316 173756 269622
rect 175108 267306 175136 277766
rect 175844 271862 175872 277780
rect 176752 274508 176804 274514
rect 176752 274450 176804 274456
rect 175832 271856 175884 271862
rect 175832 271798 175884 271804
rect 175280 271720 175332 271726
rect 175280 271662 175332 271668
rect 174544 267300 174596 267306
rect 174544 267242 174596 267248
rect 175096 267300 175148 267306
rect 175096 267242 175148 267248
rect 174556 264316 174584 267242
rect 175292 264330 175320 271662
rect 176200 268252 176252 268258
rect 176200 268194 176252 268200
rect 175292 264302 175398 264330
rect 176212 264316 176240 268194
rect 176764 264330 176792 274450
rect 176948 274242 176976 277780
rect 178144 275738 178172 277780
rect 178132 275732 178184 275738
rect 178132 275674 178184 275680
rect 176936 274236 176988 274242
rect 176936 274178 176988 274184
rect 177488 273828 177540 273834
rect 177488 273770 177540 273776
rect 177500 264330 177528 273770
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179340 268938 179368 277780
rect 180536 272814 180564 277780
rect 181732 275874 181760 277780
rect 181720 275868 181772 275874
rect 181720 275810 181772 275816
rect 182088 275052 182140 275058
rect 182088 274994 182140 275000
rect 180524 272808 180576 272814
rect 180524 272750 180576 272756
rect 179880 272400 179932 272406
rect 179880 272342 179932 272348
rect 179328 268932 179380 268938
rect 179328 268874 179380 268880
rect 179512 266620 179564 266626
rect 179512 266562 179564 266568
rect 179524 264316 179552 266562
rect 179892 264330 179920 272342
rect 181352 271040 181404 271046
rect 181352 270982 181404 270988
rect 181168 269816 181220 269822
rect 181168 269758 181220 269764
rect 179892 264302 180366 264330
rect 181180 264316 181208 269758
rect 181364 267734 181392 270982
rect 182100 269822 182128 274994
rect 182928 274514 182956 277780
rect 184138 277766 184796 277794
rect 183468 275324 183520 275330
rect 183468 275266 183520 275272
rect 182916 274508 182968 274514
rect 182916 274450 182968 274456
rect 182456 270904 182508 270910
rect 182456 270846 182508 270852
rect 182088 269816 182140 269822
rect 182088 269758 182140 269764
rect 182180 269272 182232 269278
rect 182180 269214 182232 269220
rect 181364 267706 181576 267734
rect 181548 264330 181576 267706
rect 182192 266422 182220 269214
rect 182180 266416 182232 266422
rect 182180 266358 182232 266364
rect 182468 264330 182496 270846
rect 183480 269550 183508 275266
rect 184204 273080 184256 273086
rect 184204 273022 184256 273028
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183652 268116 183704 268122
rect 183652 268058 183704 268064
rect 181548 264302 182022 264330
rect 182468 264302 182850 264330
rect 183664 264316 183692 268058
rect 184216 267034 184244 273022
rect 184768 269686 184796 277766
rect 185228 274718 185256 277780
rect 186424 275330 186452 277780
rect 186412 275324 186464 275330
rect 186412 275266 186464 275272
rect 185584 274916 185636 274922
rect 185584 274858 185636 274864
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 185032 273692 185084 273698
rect 185032 273634 185084 273640
rect 184756 269680 184808 269686
rect 184756 269622 184808 269628
rect 184020 267028 184072 267034
rect 184020 266970 184072 266976
rect 184204 267028 184256 267034
rect 184204 266970 184256 266976
rect 184032 266762 184060 266970
rect 184480 266892 184532 266898
rect 184480 266834 184532 266840
rect 184020 266756 184072 266762
rect 184020 266698 184072 266704
rect 184492 264316 184520 266834
rect 185044 264330 185072 273634
rect 185596 269074 185624 274858
rect 187148 274712 187200 274718
rect 187148 274654 187200 274660
rect 186964 269816 187016 269822
rect 186964 269758 187016 269764
rect 185584 269068 185636 269074
rect 185584 269010 185636 269016
rect 186136 266416 186188 266422
rect 186136 266358 186188 266364
rect 185044 264302 185334 264330
rect 186148 264316 186176 266358
rect 186976 264316 187004 269758
rect 187160 267578 187188 274654
rect 187620 273086 187648 277780
rect 188816 275330 188844 277780
rect 187792 275324 187844 275330
rect 187792 275266 187844 275272
rect 188804 275324 188856 275330
rect 188804 275266 188856 275272
rect 187804 274378 187832 275266
rect 187792 274372 187844 274378
rect 187792 274314 187844 274320
rect 187792 273556 187844 273562
rect 187792 273498 187844 273504
rect 187608 273080 187660 273086
rect 187608 273022 187660 273028
rect 187804 272898 187832 273498
rect 187712 272870 187832 272898
rect 189816 272944 189868 272950
rect 189816 272886 189868 272892
rect 187332 269816 187384 269822
rect 187332 269758 187384 269764
rect 187344 269550 187372 269758
rect 187332 269544 187384 269550
rect 187332 269486 187384 269492
rect 187148 267572 187200 267578
rect 187148 267514 187200 267520
rect 187712 265674 187740 272870
rect 187884 270768 187936 270774
rect 187884 270710 187936 270716
rect 187700 265668 187752 265674
rect 187700 265610 187752 265616
rect 187896 265554 187924 270710
rect 189448 266756 189500 266762
rect 189448 266698 189500 266704
rect 188252 265668 188304 265674
rect 188252 265610 188304 265616
rect 187804 265526 187924 265554
rect 187804 264316 187832 265526
rect 188264 264330 188292 265610
rect 188264 264302 188646 264330
rect 189460 264316 189488 266698
rect 189828 264330 189856 272886
rect 190012 271046 190040 277780
rect 191208 272950 191236 277780
rect 191196 272944 191248 272950
rect 191196 272886 191248 272892
rect 190736 272264 190788 272270
rect 190736 272206 190788 272212
rect 190000 271040 190052 271046
rect 190000 270982 190052 270988
rect 190748 264330 190776 272206
rect 192312 271726 192340 277780
rect 193508 273970 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 193864 276004 193916 276010
rect 193864 275946 193916 275952
rect 192484 273964 192536 273970
rect 192484 273906 192536 273912
rect 193496 273964 193548 273970
rect 193496 273906 193548 273912
rect 192300 271720 192352 271726
rect 192300 271662 192352 271668
rect 191932 269816 191984 269822
rect 191932 269758 191984 269764
rect 189828 264302 190302 264330
rect 190748 264302 191130 264330
rect 191944 264316 191972 269758
rect 192496 264330 192524 273906
rect 193588 268388 193640 268394
rect 193588 268330 193640 268336
rect 192496 264302 192786 264330
rect 193600 264316 193628 268330
rect 193876 267034 193904 275946
rect 194612 269822 194640 277366
rect 195900 274650 195928 277780
rect 197110 277766 197308 277794
rect 198306 277766 198688 277794
rect 195888 274644 195940 274650
rect 195888 274586 195940 274592
rect 195980 271312 196032 271318
rect 195980 271254 196032 271260
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 193864 267028 193916 267034
rect 193864 266970 193916 266976
rect 194428 264316 194456 267106
rect 194796 264330 194824 271118
rect 195992 264330 196020 271254
rect 196900 269068 196952 269074
rect 196900 269010 196952 269016
rect 194796 264302 195270 264330
rect 195992 264302 196098 264330
rect 196912 264316 196940 269010
rect 197280 268394 197308 277766
rect 197544 272536 197596 272542
rect 197544 272478 197596 272484
rect 197268 268388 197320 268394
rect 197268 268330 197320 268336
rect 197556 264330 197584 272478
rect 198660 269958 198688 277766
rect 199488 272542 199516 277780
rect 200592 277394 200620 277780
rect 200500 277366 200620 277394
rect 199660 274508 199712 274514
rect 199660 274450 199712 274456
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 198188 269952 198240 269958
rect 198188 269894 198240 269900
rect 198648 269952 198700 269958
rect 198648 269894 198700 269900
rect 198200 264330 198228 269894
rect 199384 267708 199436 267714
rect 199384 267650 199436 267656
rect 197556 264302 197754 264330
rect 198200 264302 198582 264330
rect 199396 264316 199424 267650
rect 199672 267170 199700 274450
rect 200500 270910 200528 277366
rect 201788 276010 201816 277780
rect 201776 276004 201828 276010
rect 201776 275946 201828 275952
rect 202144 275596 202196 275602
rect 202144 275538 202196 275544
rect 200672 274100 200724 274106
rect 200672 274042 200724 274048
rect 200488 270904 200540 270910
rect 200488 270846 200540 270852
rect 200212 268524 200264 268530
rect 200212 268466 200264 268472
rect 199660 267164 199712 267170
rect 199660 267106 199712 267112
rect 200224 264316 200252 268466
rect 200684 264330 200712 274042
rect 201868 267028 201920 267034
rect 201868 266970 201920 266976
rect 200684 264302 201066 264330
rect 201880 264316 201908 266970
rect 202156 266422 202184 275538
rect 202696 270088 202748 270094
rect 202696 270030 202748 270036
rect 202144 266416 202196 266422
rect 202144 266358 202196 266364
rect 202708 264316 202736 270030
rect 202984 268530 203012 277780
rect 203996 277766 204194 277794
rect 205390 277766 205588 277794
rect 203996 268802 204024 277766
rect 205560 270094 205588 277766
rect 206284 274644 206336 274650
rect 206284 274586 206336 274592
rect 205732 271448 205784 271454
rect 205732 271390 205784 271396
rect 205548 270088 205600 270094
rect 205548 270030 205600 270036
rect 203524 268796 203576 268802
rect 203524 268738 203576 268744
rect 203984 268796 204036 268802
rect 203984 268738 204036 268744
rect 202972 268524 203024 268530
rect 202972 268466 203024 268472
rect 203536 264316 203564 268738
rect 205180 268660 205232 268666
rect 205180 268602 205232 268608
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 205192 264316 205220 268602
rect 205744 264330 205772 271390
rect 206296 266762 206324 274586
rect 206572 274106 206600 277780
rect 207782 277766 208348 277794
rect 206560 274100 206612 274106
rect 206560 274042 206612 274048
rect 207664 271856 207716 271862
rect 207664 271798 207716 271804
rect 207388 270224 207440 270230
rect 207388 270166 207440 270172
rect 206284 266756 206336 266762
rect 206284 266698 206336 266704
rect 206836 266416 206888 266422
rect 206836 266358 206888 266364
rect 205744 264302 206034 264330
rect 206848 264316 206876 266358
rect 207400 264330 207428 270166
rect 207676 267714 207704 271798
rect 208320 269550 208348 277766
rect 208492 272672 208544 272678
rect 208492 272614 208544 272620
rect 208308 269544 208360 269550
rect 208308 269486 208360 269492
rect 207664 267708 207716 267714
rect 207664 267650 207716 267656
rect 207400 264302 207690 264330
rect 208504 264316 208532 272614
rect 208872 271182 208900 277780
rect 210068 274718 210096 277780
rect 210424 275460 210476 275466
rect 210424 275402 210476 275408
rect 210056 274712 210108 274718
rect 210056 274654 210108 274660
rect 208860 271176 208912 271182
rect 208860 271118 208912 271124
rect 209504 270496 209556 270502
rect 209504 270438 209556 270444
rect 209516 266898 209544 270438
rect 210148 270360 210200 270366
rect 210148 270302 210200 270308
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 209504 266892 209556 266898
rect 209504 266834 209556 266840
rect 209332 264316 209360 266834
rect 210160 264316 210188 270302
rect 210436 266422 210464 275402
rect 211264 273086 211292 277780
rect 211804 273216 211856 273222
rect 211804 273158 211856 273164
rect 211252 273080 211304 273086
rect 211252 273022 211304 273028
rect 211816 267442 211844 273158
rect 212460 270230 212488 277780
rect 213670 277766 213868 277794
rect 212632 271584 212684 271590
rect 212632 271526 212684 271532
rect 212448 270224 212500 270230
rect 212448 270166 212500 270172
rect 211804 267436 211856 267442
rect 211804 267378 211856 267384
rect 210976 266892 211028 266898
rect 210976 266834 211028 266840
rect 210424 266416 210476 266422
rect 210424 266358 210476 266364
rect 210988 264316 211016 266834
rect 211804 266416 211856 266422
rect 211804 266358 211856 266364
rect 211816 264316 211844 266358
rect 212644 264316 212672 271526
rect 213840 270366 213868 277766
rect 214656 274236 214708 274242
rect 214656 274178 214708 274184
rect 213828 270360 213880 270366
rect 213828 270302 213880 270308
rect 213828 269680 213880 269686
rect 213828 269622 213880 269628
rect 213460 267708 213512 267714
rect 213460 267650 213512 267656
rect 213472 264316 213500 267650
rect 213840 266626 213868 269622
rect 214288 267300 214340 267306
rect 214288 267242 214340 267248
rect 213828 266620 213880 266626
rect 213828 266562 213880 266568
rect 214300 264316 214328 267242
rect 214668 264330 214696 274178
rect 214852 271862 214880 277780
rect 214840 271856 214892 271862
rect 214840 271798 214892 271804
rect 215956 271318 215984 277780
rect 217166 277766 217456 277794
rect 216864 275732 216916 275738
rect 216864 275674 216916 275680
rect 215944 271312 215996 271318
rect 215944 271254 215996 271260
rect 216128 271040 216180 271046
rect 216128 270982 216180 270988
rect 215944 268932 215996 268938
rect 215944 268874 215996 268880
rect 214668 264302 215142 264330
rect 215956 264316 215984 268874
rect 216140 267714 216168 270982
rect 216876 267734 216904 275674
rect 217232 272808 217284 272814
rect 217232 272750 217284 272756
rect 216128 267708 216180 267714
rect 216128 267650 216180 267656
rect 216784 267706 216904 267734
rect 216784 264316 216812 267706
rect 217244 264330 217272 272750
rect 217428 272678 217456 277766
rect 218348 275466 218376 277780
rect 218888 275868 218940 275874
rect 218888 275810 218940 275816
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217416 272672 217468 272678
rect 217416 272614 217468 272620
rect 218428 267164 218480 267170
rect 218428 267106 218480 267112
rect 217244 264302 217626 264330
rect 218440 264316 218468 267106
rect 218900 264330 218928 275810
rect 219544 268666 219572 277780
rect 220556 277766 220754 277794
rect 220556 274242 220584 277766
rect 221936 275602 221964 277780
rect 223146 277766 223528 277794
rect 223500 276026 223528 277766
rect 222108 276004 222160 276010
rect 223500 275998 223620 276026
rect 222108 275946 222160 275952
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 220912 274372 220964 274378
rect 220912 274314 220964 274320
rect 220544 274236 220596 274242
rect 220544 274178 220596 274184
rect 220084 273080 220136 273086
rect 220084 273022 220136 273028
rect 219532 268660 219584 268666
rect 219532 268602 219584 268608
rect 220096 267306 220124 273022
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 220084 266620 220136 266626
rect 220084 266562 220136 266568
rect 218900 264302 219282 264330
rect 220096 264316 220124 266562
rect 220924 264316 220952 274314
rect 222120 271862 222148 275946
rect 222844 275324 222896 275330
rect 222844 275266 222896 275272
rect 221464 271856 221516 271862
rect 221464 271798 221516 271804
rect 222108 271856 222160 271862
rect 222108 271798 222160 271804
rect 221476 267170 221504 271798
rect 221740 267572 221792 267578
rect 221740 267514 221792 267520
rect 221464 267164 221516 267170
rect 221464 267106 221516 267112
rect 221752 264316 221780 267514
rect 222568 267436 222620 267442
rect 222568 267378 222620 267384
rect 222580 264316 222608 267378
rect 222856 266422 222884 275266
rect 223592 271454 223620 275998
rect 224236 275126 224264 277780
rect 225432 275330 225460 277780
rect 225420 275324 225472 275330
rect 225420 275266 225472 275272
rect 224224 275120 224276 275126
rect 224224 275062 224276 275068
rect 226156 275120 226208 275126
rect 226156 275062 226208 275068
rect 224868 272944 224920 272950
rect 224920 272892 225000 272898
rect 224868 272886 225000 272892
rect 224880 272870 225000 272886
rect 223580 271448 223632 271454
rect 223580 271390 223632 271396
rect 224224 270904 224276 270910
rect 224224 270846 224276 270852
rect 223396 267708 223448 267714
rect 223396 267650 223448 267656
rect 222844 266416 222896 266422
rect 222844 266358 222896 266364
rect 223408 264316 223436 267650
rect 224236 267442 224264 270846
rect 224224 267436 224276 267442
rect 224224 267378 224276 267384
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 224236 264316 224264 266358
rect 224972 264330 225000 272870
rect 225512 271720 225564 271726
rect 225512 271662 225564 271668
rect 225524 264330 225552 271662
rect 226168 271590 226196 275062
rect 226340 273964 226392 273970
rect 226340 273906 226392 273912
rect 226156 271584 226208 271590
rect 226156 271526 226208 271532
rect 226352 264330 226380 273906
rect 226628 269686 226656 277780
rect 227824 277394 227852 277780
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 227824 277366 227944 277394
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 227272 264330 227300 269758
rect 227916 268802 227944 277366
rect 228836 272814 228864 277766
rect 228824 272808 228876 272814
rect 228824 272750 228876 272756
rect 230400 269958 230428 277766
rect 231412 272542 231440 277780
rect 232530 277766 233188 277794
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 230020 269952 230072 269958
rect 230020 269894 230072 269900
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 227720 268796 227772 268802
rect 227720 268738 227772 268744
rect 227904 268796 227956 268802
rect 227904 268738 227956 268744
rect 227732 267034 227760 268738
rect 229192 268388 229244 268394
rect 229192 268330 229244 268336
rect 227720 267028 227772 267034
rect 227720 266970 227772 266976
rect 228364 266756 228416 266762
rect 228364 266698 228416 266704
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226352 264302 226734 264330
rect 227272 264302 227562 264330
rect 228376 264316 228404 266698
rect 229204 264316 229232 268330
rect 230032 264316 230060 269894
rect 230584 264330 230612 272478
rect 232136 271856 232188 271862
rect 232136 271798 232188 271804
rect 230756 269544 230808 269550
rect 230756 269486 230808 269492
rect 230768 266422 230796 269486
rect 231676 267436 231728 267442
rect 231676 267378 231728 267384
rect 230756 266416 230808 266422
rect 230756 266358 230808 266364
rect 230584 264302 230874 264330
rect 231688 264316 231716 267378
rect 232148 264330 232176 271798
rect 233160 270502 233188 277766
rect 233148 270496 233200 270502
rect 233148 270438 233200 270444
rect 233332 268524 233384 268530
rect 233332 268466 233384 268472
rect 232148 264302 232530 264330
rect 233344 264316 233372 268466
rect 233712 268394 233740 277780
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 268388 233752 268394
rect 233700 268330 233752 268336
rect 233896 267442 233924 275538
rect 234908 273970 234936 277780
rect 236104 275602 236132 277780
rect 237300 277394 237328 277780
rect 237208 277366 237328 277394
rect 236092 275596 236144 275602
rect 236092 275538 236144 275544
rect 235448 274100 235500 274106
rect 235448 274042 235500 274048
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 234988 270088 235040 270094
rect 234988 270030 235040 270036
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234160 267028 234212 267034
rect 234160 266970 234212 266976
rect 234172 264316 234200 266970
rect 235000 264316 235028 270030
rect 235460 264330 235488 274042
rect 237208 270638 237236 277366
rect 237380 275460 237432 275466
rect 237380 275402 237432 275408
rect 237392 274378 237420 275402
rect 238496 274718 238524 277780
rect 238484 274712 238536 274718
rect 238484 274654 238536 274660
rect 237840 274508 237892 274514
rect 237840 274450 237892 274456
rect 237380 274372 237432 274378
rect 237380 274314 237432 274320
rect 237472 271176 237524 271182
rect 237472 271118 237524 271124
rect 237196 270632 237248 270638
rect 237196 270574 237248 270580
rect 237288 270496 237340 270502
rect 237288 270438 237340 270444
rect 237300 267034 237328 270438
rect 237288 267028 237340 267034
rect 237288 266970 237340 266976
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237484 264316 237512 271118
rect 237852 264330 237880 274450
rect 239600 274106 239628 277780
rect 239772 274712 239824 274718
rect 239772 274654 239824 274660
rect 239588 274100 239640 274106
rect 239588 274042 239640 274048
rect 239784 270094 239812 274654
rect 240600 274236 240652 274242
rect 240600 274178 240652 274184
rect 240612 270994 240640 274178
rect 240796 271182 240824 277780
rect 242006 277766 242388 277794
rect 242360 272678 242388 277766
rect 242164 272672 242216 272678
rect 242164 272614 242216 272620
rect 242348 272672 242400 272678
rect 242348 272614 242400 272620
rect 242176 271402 242204 272614
rect 242176 271374 242296 271402
rect 242072 271312 242124 271318
rect 242072 271254 242124 271260
rect 240784 271176 240836 271182
rect 240784 271118 240836 271124
rect 240612 270966 240732 270994
rect 240508 270360 240560 270366
rect 240508 270302 240560 270308
rect 239956 270224 240008 270230
rect 239956 270166 240008 270172
rect 239772 270088 239824 270094
rect 239772 270030 239824 270036
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 237852 264302 238326 264330
rect 239140 264316 239168 267242
rect 239968 264316 239996 270166
rect 240520 264330 240548 270302
rect 240704 266762 240732 270966
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 240692 266756 240744 266762
rect 240692 266698 240744 266704
rect 240520 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271254
rect 242268 266422 242296 271374
rect 243188 271318 243216 277780
rect 244384 274718 244412 277780
rect 245108 275324 245160 275330
rect 245108 275266 245160 275272
rect 244372 274712 244424 274718
rect 244372 274654 244424 274660
rect 243728 274372 243780 274378
rect 243728 274314 243780 274320
rect 243176 271312 243228 271318
rect 243176 271254 243228 271260
rect 242256 266416 242308 266422
rect 242256 266358 242308 266364
rect 243268 266416 243320 266422
rect 243268 266358 243320 266364
rect 242084 264302 242466 264330
rect 243280 264316 243308 266358
rect 243740 264330 243768 274314
rect 244924 268660 244976 268666
rect 244924 268602 244976 268608
rect 243740 264302 244122 264330
rect 244936 264316 244964 268602
rect 245120 266626 245148 275266
rect 245580 268530 245608 277780
rect 246790 277766 246988 277794
rect 245568 268524 245620 268530
rect 245568 268466 245620 268472
rect 246580 267436 246632 267442
rect 246580 267378 246632 267384
rect 245752 266756 245804 266762
rect 245752 266698 245804 266704
rect 245108 266620 245160 266626
rect 245108 266562 245160 266568
rect 245764 264316 245792 266698
rect 246592 264316 246620 267378
rect 246960 267170 246988 277766
rect 247224 271584 247276 271590
rect 247224 271526 247276 271532
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 247236 265674 247264 271526
rect 247880 271454 247908 277780
rect 249090 277766 249656 277794
rect 249064 272808 249116 272814
rect 249064 272750 249116 272756
rect 247408 271448 247460 271454
rect 247408 271390 247460 271396
rect 247868 271448 247920 271454
rect 247868 271390 247920 271396
rect 247224 265668 247276 265674
rect 247224 265610 247276 265616
rect 247420 264316 247448 271390
rect 249076 266762 249104 272750
rect 249628 270502 249656 277766
rect 250272 275330 250300 277780
rect 250260 275324 250312 275330
rect 250260 275266 250312 275272
rect 251088 274712 251140 274718
rect 251088 274654 251140 274660
rect 249616 270496 249668 270502
rect 249616 270438 249668 270444
rect 251100 270230 251128 274654
rect 251088 270224 251140 270230
rect 251088 270166 251140 270172
rect 250904 270088 250956 270094
rect 250904 270030 250956 270036
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 249064 266756 249116 266762
rect 249064 266698 249116 266704
rect 249064 266620 249116 266626
rect 249064 266562 249116 266568
rect 247868 265668 247920 265674
rect 247868 265610 247920 265616
rect 247880 264330 247908 265610
rect 247880 264302 248262 264330
rect 249076 264316 249104 266562
rect 249904 264316 249932 269758
rect 250916 269686 250944 270030
rect 251468 269822 251496 277780
rect 252678 277766 252968 277794
rect 252940 272542 252968 277766
rect 252744 272536 252796 272542
rect 252744 272478 252796 272484
rect 252928 272536 252980 272542
rect 252928 272478 252980 272484
rect 252008 270360 252060 270366
rect 252008 270302 252060 270308
rect 251456 269816 251508 269822
rect 251456 269758 251508 269764
rect 250904 269680 250956 269686
rect 250904 269622 250956 269628
rect 250720 268796 250772 268802
rect 250720 268738 250772 268744
rect 250732 264316 250760 268738
rect 251548 266756 251600 266762
rect 251548 266698 251600 266704
rect 251560 264316 251588 266698
rect 252020 266422 252048 270302
rect 252376 269952 252428 269958
rect 252376 269894 252428 269900
rect 252008 266416 252060 266422
rect 252008 266358 252060 266364
rect 252388 264316 252416 269894
rect 252756 264330 252784 272478
rect 253664 270496 253716 270502
rect 253664 270438 253716 270444
rect 253676 267306 253704 270438
rect 253860 270230 253888 277780
rect 255070 277766 255268 277794
rect 253848 270224 253900 270230
rect 253848 270166 253900 270172
rect 255240 268394 255268 277766
rect 255504 275596 255556 275602
rect 255504 275538 255556 275544
rect 254860 268388 254912 268394
rect 254860 268330 254912 268336
rect 255228 268388 255280 268394
rect 255228 268330 255280 268336
rect 253664 267300 253716 267306
rect 253664 267242 253716 267248
rect 254032 267028 254084 267034
rect 254032 266970 254084 266976
rect 252756 264302 253230 264330
rect 254044 264316 254072 266970
rect 254872 264316 254900 268330
rect 255516 265674 255544 275538
rect 256160 273970 256188 277780
rect 257370 277766 258028 277794
rect 255688 273964 255740 273970
rect 255688 273906 255740 273912
rect 256148 273964 256200 273970
rect 256148 273906 256200 273912
rect 255504 265668 255556 265674
rect 255504 265610 255556 265616
rect 255700 264316 255728 273906
rect 258000 266898 258028 277766
rect 258552 277394 258580 277780
rect 258460 277366 258580 277394
rect 258460 269958 258488 277366
rect 258632 274100 258684 274106
rect 258632 274042 258684 274048
rect 258448 269952 258500 269958
rect 258448 269894 258500 269900
rect 258172 269680 258224 269686
rect 258172 269622 258224 269628
rect 257988 266892 258040 266898
rect 257988 266834 258040 266840
rect 257344 266416 257396 266422
rect 257344 266358 257396 266364
rect 256148 265668 256200 265674
rect 256148 265610 256200 265616
rect 256160 264330 256188 265610
rect 256160 264302 256542 264330
rect 257356 264316 257384 266358
rect 258184 264316 258212 269622
rect 258644 264330 258672 274042
rect 259552 272672 259604 272678
rect 259552 272614 259604 272620
rect 259564 265674 259592 272614
rect 259748 271590 259776 277780
rect 260944 275466 260972 277780
rect 260932 275460 260984 275466
rect 260932 275402 260984 275408
rect 259736 271584 259788 271590
rect 259736 271526 259788 271532
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 259828 271176 259880 271182
rect 259828 271118 259880 271124
rect 259552 265668 259604 265674
rect 259552 265610 259604 265616
rect 258644 264302 259026 264330
rect 259840 264316 259868 271118
rect 260380 265668 260432 265674
rect 260380 265610 260432 265616
rect 260392 264330 260420 265610
rect 261036 264330 261064 271254
rect 262140 271182 262168 277780
rect 263258 277766 263548 277794
rect 264454 277766 264928 277794
rect 265650 277766 266308 277794
rect 262128 271176 262180 271182
rect 262128 271118 262180 271124
rect 262312 270360 262364 270366
rect 262312 270302 262364 270308
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262324 264316 262352 270302
rect 263520 268530 263548 277766
rect 264336 271448 264388 271454
rect 264336 271390 264388 271396
rect 263140 268524 263192 268530
rect 263140 268466 263192 268472
rect 263508 268524 263560 268530
rect 263508 268466 263560 268472
rect 263152 264316 263180 268466
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263980 264316 264008 267106
rect 264348 264330 264376 271390
rect 264900 269278 264928 277766
rect 265072 270224 265124 270230
rect 265072 270166 265124 270172
rect 264888 269272 264940 269278
rect 264888 269214 264940 269220
rect 265084 266762 265112 270166
rect 266280 270094 266308 277766
rect 266636 275324 266688 275330
rect 266636 275266 266688 275272
rect 266268 270088 266320 270094
rect 266268 270030 266320 270036
rect 265624 267300 265676 267306
rect 265624 267242 265676 267248
rect 265072 266756 265124 266762
rect 265072 266698 265124 266704
rect 264348 264302 264822 264330
rect 265636 264316 265664 267242
rect 266648 264330 266676 275266
rect 266832 271318 266860 277780
rect 268028 272542 268056 277780
rect 267832 272536 267884 272542
rect 267832 272478 267884 272484
rect 268016 272536 268068 272542
rect 268016 272478 268068 272484
rect 266820 271312 266872 271318
rect 266820 271254 266872 271260
rect 267280 269816 267332 269822
rect 267280 269758 267332 269764
rect 266478 264302 266676 264330
rect 267292 264316 267320 269758
rect 267844 264330 267872 272478
rect 268384 271584 268436 271590
rect 268384 271526 268436 271532
rect 268396 266422 268424 271526
rect 269224 269822 269252 277780
rect 270420 274718 270448 277780
rect 270408 274712 270460 274718
rect 270408 274654 270460 274660
rect 271144 274712 271196 274718
rect 271144 274654 271196 274660
rect 270592 273964 270644 273970
rect 270592 273906 270644 273912
rect 269212 269816 269264 269822
rect 269212 269758 269264 269764
rect 269120 269272 269172 269278
rect 269120 269214 269172 269220
rect 268936 266756 268988 266762
rect 268936 266698 268988 266704
rect 268384 266416 268436 266422
rect 268384 266358 268436 266364
rect 267844 264302 268134 264330
rect 268948 264316 268976 266698
rect 269132 266558 269160 269214
rect 269764 268388 269816 268394
rect 269764 268330 269816 268336
rect 269120 266552 269172 266558
rect 269120 266494 269172 266500
rect 269776 264316 269804 268330
rect 270604 264316 270632 273906
rect 271156 266898 271184 274654
rect 271524 273970 271552 277780
rect 272734 277766 273116 277794
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 273088 269958 273116 277766
rect 273536 275460 273588 275466
rect 273536 275402 273588 275408
rect 272248 269952 272300 269958
rect 272248 269894 272300 269900
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 271420 267028 271472 267034
rect 271420 266970 271472 266976
rect 271144 266892 271196 266898
rect 271144 266834 271196 266840
rect 271432 264316 271460 266970
rect 272260 264316 272288 269894
rect 273076 266416 273128 266422
rect 273076 266358 273128 266364
rect 273088 264316 273116 266358
rect 273548 264330 273576 275402
rect 273916 275330 273944 277780
rect 273904 275324 273956 275330
rect 273904 275266 273956 275272
rect 275112 271454 275140 277780
rect 275100 271448 275152 271454
rect 275100 271390 275152 271396
rect 276308 271182 276336 277780
rect 277504 274990 277532 277780
rect 278700 277394 278728 277780
rect 278608 277366 278728 277394
rect 277492 274984 277544 274990
rect 277492 274926 277544 274932
rect 276664 271312 276716 271318
rect 276664 271254 276716 271260
rect 274640 271176 274692 271182
rect 274640 271118 274692 271124
rect 276296 271176 276348 271182
rect 276296 271118 276348 271124
rect 274652 264330 274680 271118
rect 275560 268524 275612 268530
rect 275560 268466 275612 268472
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 268466
rect 276676 267034 276704 271254
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276664 267028 276716 267034
rect 276664 266970 276716 266976
rect 276388 266552 276440 266558
rect 276388 266494 276440 266500
rect 276400 264316 276428 266494
rect 277228 264316 277256 270030
rect 278044 267028 278096 267034
rect 278044 266970 278096 266976
rect 278056 264316 278084 266970
rect 278608 266422 278636 277366
rect 279804 272542 279832 277780
rect 280804 273964 280856 273970
rect 280804 273906 280856 273912
rect 278780 272536 278832 272542
rect 278780 272478 278832 272484
rect 279792 272536 279844 272542
rect 279792 272478 279844 272484
rect 278596 266416 278648 266422
rect 278596 266358 278648 266364
rect 278792 264330 278820 272478
rect 279700 269816 279752 269822
rect 279700 269758 279752 269764
rect 278792 264302 278898 264330
rect 279712 264316 279740 269758
rect 280816 267734 280844 273906
rect 281000 273766 281028 277780
rect 282210 277766 282776 277794
rect 280988 273760 281040 273766
rect 280988 273702 281040 273708
rect 282184 269952 282236 269958
rect 282184 269894 282236 269900
rect 280816 267706 280936 267734
rect 280528 266892 280580 266898
rect 280528 266834 280580 266840
rect 280540 264316 280568 266834
rect 280908 264330 280936 267706
rect 280908 264302 281382 264330
rect 282196 264316 282224 269894
rect 282748 269142 282776 277766
rect 282920 275324 282972 275330
rect 282920 275266 282972 275272
rect 282736 269136 282788 269142
rect 282736 269078 282788 269084
rect 282932 264330 282960 275266
rect 283392 274854 283420 277780
rect 284588 275466 284616 277780
rect 284576 275460 284628 275466
rect 284576 275402 284628 275408
rect 284300 274984 284352 274990
rect 284300 274926 284352 274932
rect 283380 274848 283432 274854
rect 283380 274790 283432 274796
rect 283472 271448 283524 271454
rect 283472 271390 283524 271396
rect 283484 264330 283512 271390
rect 284312 265674 284340 274926
rect 285784 274718 285812 277780
rect 286888 277394 286916 277780
rect 286796 277366 286916 277394
rect 285772 274712 285824 274718
rect 285772 274654 285824 274660
rect 284484 271176 284536 271182
rect 284484 271118 284536 271124
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271118
rect 286796 269958 286824 277366
rect 286968 274712 287020 274718
rect 286968 274654 287020 274660
rect 286784 269952 286836 269958
rect 286784 269894 286836 269900
rect 286980 267034 287008 274654
rect 287520 273760 287572 273766
rect 287520 273702 287572 273708
rect 287152 272536 287204 272542
rect 287152 272478 287204 272484
rect 286968 267028 287020 267034
rect 286968 266970 287020 266976
rect 286324 266416 286376 266422
rect 286324 266358 286376 266364
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 286336 264316 286364 266358
rect 287164 264316 287192 272478
rect 287532 264330 287560 273702
rect 288084 272950 288112 277780
rect 289280 274922 289308 277780
rect 290096 275460 290148 275466
rect 290096 275402 290148 275408
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289084 274848 289136 274854
rect 289084 274790 289136 274796
rect 288072 272944 288124 272950
rect 288072 272886 288124 272892
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 287532 264302 288006 264330
rect 288820 264316 288848 269078
rect 289096 267734 289124 274790
rect 289096 267706 289216 267734
rect 289188 264330 289216 267706
rect 290108 264330 290136 275402
rect 290476 275262 290504 277780
rect 290464 275256 290516 275262
rect 290464 275198 290516 275204
rect 290464 272944 290516 272950
rect 290464 272886 290516 272892
rect 290476 266422 290504 272886
rect 291672 270502 291700 277780
rect 292868 274718 292896 277780
rect 293408 274916 293460 274922
rect 293408 274858 293460 274864
rect 292856 274712 292908 274718
rect 292856 274654 292908 274660
rect 291660 270496 291712 270502
rect 291660 270438 291712 270444
rect 292120 269952 292172 269958
rect 292120 269894 292172 269900
rect 291292 267028 291344 267034
rect 291292 266970 291344 266976
rect 290464 266416 290516 266422
rect 290464 266358 290516 266364
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 266970
rect 292132 264316 292160 269894
rect 292948 266416 293000 266422
rect 292948 266358 293000 266364
rect 292960 264316 292988 266358
rect 293420 264330 293448 274858
rect 293868 274712 293920 274718
rect 293868 274654 293920 274660
rect 293880 266422 293908 274654
rect 294064 269142 294092 277780
rect 294328 275256 294380 275262
rect 294328 275198 294380 275204
rect 294052 269136 294104 269142
rect 294052 269078 294104 269084
rect 293868 266416 293920 266422
rect 293868 266358 293920 266364
rect 294340 264330 294368 275198
rect 295168 274666 295196 277780
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 295168 274638 295380 274666
rect 296352 274654 296404 274660
rect 295352 269278 295380 274638
rect 297928 270502 297956 277766
rect 298756 274718 298784 277780
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298744 274712 298796 274718
rect 298744 274654 298796 274660
rect 295524 270496 295576 270502
rect 295524 270438 295576 270444
rect 297916 270496 297968 270502
rect 297916 270438 297968 270444
rect 295340 269272 295392 269278
rect 295340 269214 295392 269220
rect 295536 267734 295564 270438
rect 297916 269272 297968 269278
rect 297916 269214 297968 269220
rect 297088 269136 297140 269142
rect 297088 269078 297140 269084
rect 295444 267706 295564 267734
rect 293420 264302 293802 264330
rect 294340 264302 294630 264330
rect 295444 264316 295472 267706
rect 296260 266416 296312 266422
rect 296260 266358 296312 266364
rect 296272 264316 296300 266358
rect 297100 264316 297128 269078
rect 297928 264316 297956 269214
rect 298388 264330 298416 274654
rect 299952 270502 299980 277780
rect 301148 277394 301176 277780
rect 301056 277366 301176 277394
rect 302344 277394 302372 277780
rect 302344 277366 302464 277394
rect 300124 274712 300176 274718
rect 300124 274654 300176 274660
rect 299572 270496 299624 270502
rect 299572 270438 299624 270444
rect 299940 270496 299992 270502
rect 299940 270438 299992 270444
rect 298388 264302 298770 264330
rect 299584 264316 299612 270438
rect 300136 264330 300164 274654
rect 300860 270496 300912 270502
rect 300860 270438 300912 270444
rect 300872 264330 300900 270438
rect 301056 266422 301084 277366
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300136 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303448 270450 303476 277780
rect 304092 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 303448 270422 303660 270450
rect 303632 264330 303660 270422
rect 304092 264330 304120 277766
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 316052 277766 316526 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 267300 312872 267306
rect 312820 267242 312872 267248
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312360 266416 312412 266422
rect 312360 266358 312412 266364
rect 312372 264330 312400 266358
rect 312018 264302 312400 264330
rect 312832 264316 312860 267242
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313648 267436 313700 267442
rect 313648 267378 313700 267384
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313660 264316 313688 267378
rect 314488 264316 314516 269758
rect 314672 266422 314700 277766
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266416 314712 266422
rect 314660 266358 314712 266364
rect 315776 264330 315804 271254
rect 316052 267306 316080 277766
rect 317708 277394 317736 277780
rect 317708 277366 317828 277394
rect 316960 270292 317012 270298
rect 316960 270234 317012 270240
rect 316040 267300 316092 267306
rect 316040 267242 316092 267248
rect 316132 266892 316184 266898
rect 316132 266834 316184 266840
rect 315330 264302 315804 264330
rect 316144 264316 316172 266834
rect 316972 264316 317000 270234
rect 317800 267442 317828 277366
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317788 267436 317840 267442
rect 317788 267378 317840 267384
rect 317788 266416 317840 266422
rect 317788 266358 317840 266364
rect 317800 264316 317828 266358
rect 318628 264316 318656 271730
rect 318812 269822 318840 277780
rect 320008 271318 320036 277780
rect 320192 277766 321218 277794
rect 321572 277766 322414 277794
rect 323136 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318800 269816 318852 269822
rect 318800 269758 318852 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320192 266898 320220 277766
rect 321376 274712 321428 274718
rect 321376 274654 321428 274660
rect 320180 266892 320232 266898
rect 320180 266834 320232 266840
rect 320272 266756 320324 266762
rect 320272 266698 320324 266704
rect 320284 264316 320312 266698
rect 321388 264330 321416 274654
rect 321572 270298 321600 277766
rect 322572 272536 322624 272542
rect 322572 272478 322624 272484
rect 321560 270292 321612 270298
rect 321560 270234 321612 270240
rect 321928 269816 321980 269822
rect 321928 269758 321980 269764
rect 321126 264302 321416 264330
rect 321940 264316 321968 269758
rect 322584 264330 322612 272478
rect 323136 266422 323164 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 325516 271312 325568 271318
rect 325516 271254 325568 271260
rect 323584 269952 323636 269958
rect 323584 269894 323636 269900
rect 323124 266416 323176 266422
rect 323124 266358 323176 266364
rect 322584 264302 322782 264330
rect 323596 264316 323624 269894
rect 324412 267028 324464 267034
rect 324412 266970 324464 266976
rect 324424 264316 324452 266970
rect 325528 264330 325556 271254
rect 325712 269142 325740 277766
rect 326896 270088 326948 270094
rect 326896 270030 326948 270036
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326068 268252 326120 268258
rect 326068 268194 326120 268200
rect 325266 264302 325556 264330
rect 326080 264316 326108 268194
rect 326908 264316 326936 270030
rect 327092 266762 327120 277780
rect 328288 274718 328316 277780
rect 328472 277766 329498 277794
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 328092 271176 328144 271182
rect 328092 271118 328144 271124
rect 327080 266756 327132 266762
rect 327080 266698 327132 266704
rect 328104 264330 328132 271118
rect 328472 269822 328500 277766
rect 330680 272542 330708 277780
rect 331232 277766 331890 277794
rect 332612 277766 333086 277794
rect 331036 273964 331088 273970
rect 331036 273906 331088 273912
rect 330668 272536 330720 272542
rect 330668 272478 330720 272484
rect 328460 269816 328512 269822
rect 328460 269758 328512 269764
rect 329380 269816 329432 269822
rect 329380 269758 329432 269764
rect 328552 268524 328604 268530
rect 328552 268466 328604 268472
rect 327750 264302 328132 264330
rect 328564 264316 328592 268466
rect 329392 264316 329420 269758
rect 330208 266552 330260 266558
rect 330208 266494 330260 266500
rect 330220 264316 330248 266494
rect 331048 264316 331076 273906
rect 331232 269958 331260 277766
rect 331404 274712 331456 274718
rect 331404 274654 331456 274660
rect 331220 269952 331272 269958
rect 331220 269894 331272 269900
rect 331416 268258 331444 274654
rect 332612 270494 332640 277766
rect 333612 272672 333664 272678
rect 333612 272614 333664 272620
rect 332520 270466 332640 270494
rect 331404 268252 331456 268258
rect 331404 268194 331456 268200
rect 332520 267034 332548 270466
rect 332508 267028 332560 267034
rect 332508 266970 332560 266976
rect 331864 266892 331916 266898
rect 331864 266834 331916 266840
rect 331876 264316 331904 266834
rect 333624 266422 333652 272614
rect 334176 271318 334204 277780
rect 334348 275324 334400 275330
rect 334348 275266 334400 275272
rect 334164 271312 334216 271318
rect 334164 271254 334216 271260
rect 333888 269952 333940 269958
rect 333888 269894 333940 269900
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 333612 266416 333664 266422
rect 333612 266358 333664 266364
rect 332704 264316 332732 266358
rect 333900 264330 333928 269894
rect 334360 268530 334388 275266
rect 335372 274718 335400 277780
rect 335556 277766 336582 277794
rect 335360 274712 335412 274718
rect 335360 274654 335412 274660
rect 334808 271312 334860 271318
rect 334808 271254 334860 271260
rect 334348 268524 334400 268530
rect 334348 268466 334400 268472
rect 334348 267436 334400 267442
rect 334348 267378 334400 267384
rect 333546 264302 333928 264330
rect 334360 264316 334388 267378
rect 334820 266558 334848 271254
rect 335556 270094 335584 277766
rect 337764 271182 337792 277780
rect 338960 275330 338988 277780
rect 339512 277766 340170 277794
rect 338948 275324 339000 275330
rect 338948 275266 339000 275272
rect 338948 275188 339000 275194
rect 338948 275130 339000 275136
rect 338028 272536 338080 272542
rect 338028 272478 338080 272484
rect 337752 271176 337804 271182
rect 337752 271118 337804 271124
rect 335544 270088 335596 270094
rect 335544 270030 335596 270036
rect 336832 270088 336884 270094
rect 336832 270030 336884 270036
rect 335636 269408 335688 269414
rect 335636 269350 335688 269356
rect 335176 268388 335228 268394
rect 335176 268330 335228 268336
rect 334808 266552 334860 266558
rect 334808 266494 334860 266500
rect 335188 264316 335216 268330
rect 335648 266898 335676 269350
rect 336004 267164 336056 267170
rect 336004 267106 336056 267112
rect 335636 266892 335688 266898
rect 335636 266834 335688 266840
rect 336016 264316 336044 267106
rect 336844 264316 336872 270030
rect 338040 264330 338068 272478
rect 338960 264330 338988 275130
rect 339316 270292 339368 270298
rect 339316 270234 339368 270240
rect 337686 264302 338068 264330
rect 338514 264302 338988 264330
rect 339328 264316 339356 270234
rect 339512 269822 339540 277766
rect 340604 271448 340656 271454
rect 340604 271390 340656 271396
rect 339500 269816 339552 269822
rect 339500 269758 339552 269764
rect 340616 264330 340644 271390
rect 341352 271318 341380 277780
rect 341524 275460 341576 275466
rect 341524 275402 341576 275408
rect 341340 271312 341392 271318
rect 341340 271254 341392 271260
rect 341536 270298 341564 275402
rect 342456 273970 342484 277780
rect 343666 277766 343864 277794
rect 342904 274236 342956 274242
rect 342904 274178 342956 274184
rect 342444 273964 342496 273970
rect 342444 273906 342496 273912
rect 342168 271176 342220 271182
rect 342168 271118 342220 271124
rect 341524 270292 341576 270298
rect 341524 270234 341576 270240
rect 341800 269816 341852 269822
rect 341800 269758 341852 269764
rect 340972 266416 341024 266422
rect 340972 266358 341024 266364
rect 340170 264302 340644 264330
rect 340984 264316 341012 266358
rect 341812 264316 341840 269758
rect 342180 266422 342208 271118
rect 342916 267442 342944 274178
rect 343836 269414 343864 277766
rect 344848 272678 344876 277780
rect 345124 277766 346058 277794
rect 344836 272672 344888 272678
rect 344836 272614 344888 272620
rect 344652 271312 344704 271318
rect 344652 271254 344704 271260
rect 343824 269408 343876 269414
rect 343824 269350 343876 269356
rect 342904 267436 342956 267442
rect 342904 267378 342956 267384
rect 343456 267300 343508 267306
rect 343456 267242 343508 267248
rect 342628 266892 342680 266898
rect 342628 266834 342680 266840
rect 342168 266416 342220 266422
rect 342168 266358 342220 266364
rect 342640 264316 342668 266834
rect 343468 264316 343496 267242
rect 344664 264330 344692 271254
rect 345124 269958 345152 277766
rect 347240 274242 347268 277780
rect 347792 277766 348450 277794
rect 347228 274236 347280 274242
rect 347228 274178 347280 274184
rect 346124 274100 346176 274106
rect 346124 274042 346176 274048
rect 345112 269952 345164 269958
rect 345112 269894 345164 269900
rect 345940 268524 345992 268530
rect 345940 268466 345992 268472
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 344310 264302 344692 264330
rect 345124 264316 345152 266358
rect 345952 264316 345980 268466
rect 346136 266422 346164 274042
rect 347044 273284 347096 273290
rect 347044 273226 347096 273232
rect 347056 267170 347084 273226
rect 347596 269952 347648 269958
rect 347596 269894 347648 269900
rect 347044 267164 347096 267170
rect 347044 267106 347096 267112
rect 346768 266552 346820 266558
rect 346768 266494 346820 266500
rect 346124 266416 346176 266422
rect 346124 266358 346176 266364
rect 346780 264316 346808 266494
rect 347608 264316 347636 269894
rect 347792 268394 347820 277766
rect 349632 273290 349660 277780
rect 350552 277766 350750 277794
rect 349620 273284 349672 273290
rect 349620 273226 349672 273232
rect 350264 273284 350316 273290
rect 350264 273226 350316 273232
rect 348424 270360 348476 270366
rect 348424 270302 348476 270308
rect 347780 268388 347832 268394
rect 347780 268330 347832 268336
rect 348436 264316 348464 270302
rect 350080 268388 350132 268394
rect 350080 268330 350132 268336
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 268330
rect 350276 266422 350304 273226
rect 350552 270094 350580 277766
rect 350724 275596 350776 275602
rect 350724 275538 350776 275544
rect 350736 271318 350764 275538
rect 351932 272542 351960 277780
rect 353128 275330 353156 277780
rect 354324 275466 354352 277780
rect 355152 277766 355534 277794
rect 356164 277766 356730 277794
rect 357452 277766 357926 277794
rect 354312 275460 354364 275466
rect 354312 275402 354364 275408
rect 353116 275324 353168 275330
rect 353116 275266 353168 275272
rect 353944 275324 353996 275330
rect 353944 275266 353996 275272
rect 352932 272808 352984 272814
rect 352932 272750 352984 272756
rect 351920 272536 351972 272542
rect 351920 272478 351972 272484
rect 350724 271312 350776 271318
rect 350724 271254 350776 271260
rect 351828 271312 351880 271318
rect 351828 271254 351880 271260
rect 350540 270088 350592 270094
rect 350540 270030 350592 270036
rect 351644 269680 351696 269686
rect 351644 269622 351696 269628
rect 350908 267436 350960 267442
rect 350908 267378 350960 267384
rect 350264 266416 350316 266422
rect 350264 266358 350316 266364
rect 350920 264316 350948 267378
rect 351656 266558 351684 269622
rect 351644 266552 351696 266558
rect 351644 266494 351696 266500
rect 351840 265690 351868 271254
rect 351748 265662 351868 265690
rect 351748 264316 351776 265662
rect 352944 264330 352972 272750
rect 353956 267306 353984 275266
rect 355152 271454 355180 277766
rect 355140 271448 355192 271454
rect 355140 271390 355192 271396
rect 355324 271448 355376 271454
rect 355324 271390 355376 271396
rect 354220 270088 354272 270094
rect 354220 270030 354272 270036
rect 353944 267300 353996 267306
rect 353944 267242 353996 267248
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 352590 264302 352972 264330
rect 353404 264316 353432 266970
rect 354232 264316 354260 270030
rect 355336 267034 355364 271390
rect 356164 271182 356192 277766
rect 356336 275324 356388 275330
rect 356336 275266 356388 275272
rect 356348 273290 356376 275266
rect 356336 273284 356388 273290
rect 356336 273226 356388 273232
rect 356152 271176 356204 271182
rect 356152 271118 356204 271124
rect 356520 271108 356572 271114
rect 356520 271050 356572 271056
rect 355876 267164 355928 267170
rect 355876 267106 355928 267112
rect 355324 267028 355376 267034
rect 355324 266970 355376 266976
rect 355048 266756 355100 266762
rect 355048 266698 355100 266704
rect 355060 264316 355088 266698
rect 355888 264316 355916 267106
rect 356532 266898 356560 271050
rect 356704 270224 356756 270230
rect 356704 270166 356756 270172
rect 356520 266892 356572 266898
rect 356520 266834 356572 266840
rect 356716 264316 356744 270166
rect 357452 269822 357480 277766
rect 358636 272536 358688 272542
rect 358636 272478 358688 272484
rect 357440 269816 357492 269822
rect 357440 269758 357492 269764
rect 358360 266620 358412 266626
rect 358360 266562 358412 266568
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 357544 264316 357572 266358
rect 358372 264316 358400 266562
rect 358648 266422 358676 272478
rect 359016 271114 359044 277780
rect 360212 275466 360240 277780
rect 361408 275602 361436 277780
rect 361396 275596 361448 275602
rect 361396 275538 361448 275544
rect 361580 275596 361632 275602
rect 361580 275538 361632 275544
rect 360200 275460 360252 275466
rect 360200 275402 360252 275408
rect 360292 274712 360344 274718
rect 360292 274654 360344 274660
rect 360108 273964 360160 273970
rect 360108 273906 360160 273912
rect 359004 271108 359056 271114
rect 359004 271050 359056 271056
rect 359924 270496 359976 270502
rect 359924 270438 359976 270444
rect 359188 266892 359240 266898
rect 359188 266834 359240 266840
rect 358636 266416 358688 266422
rect 358636 266358 358688 266364
rect 359200 264316 359228 266834
rect 359936 266762 359964 270438
rect 359924 266756 359976 266762
rect 359924 266698 359976 266704
rect 360120 265690 360148 273906
rect 360304 268530 360332 274654
rect 361592 271674 361620 275538
rect 362604 274106 362632 277780
rect 363052 275460 363104 275466
rect 363052 275402 363104 275408
rect 362868 274508 362920 274514
rect 362868 274450 362920 274456
rect 362592 274100 362644 274106
rect 362592 274042 362644 274048
rect 361224 271646 361620 271674
rect 360292 268524 360344 268530
rect 360292 268466 360344 268472
rect 360752 268524 360804 268530
rect 360752 268466 360804 268472
rect 360764 267442 360792 268466
rect 360752 267436 360804 267442
rect 360752 267378 360804 267384
rect 360028 265662 360148 265690
rect 360028 264316 360056 265662
rect 361224 264330 361252 271646
rect 362224 271584 362276 271590
rect 362224 271526 362276 271532
rect 362236 266626 362264 271526
rect 362880 267734 362908 274450
rect 363064 270366 363092 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 365732 277766 366114 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 364156 271176 364208 271182
rect 364156 271118 364208 271124
rect 363052 270360 363104 270366
rect 363052 270302 363104 270308
rect 363052 268660 363104 268666
rect 363052 268602 363104 268608
rect 363064 267734 363092 268602
rect 362788 267706 362908 267734
rect 362972 267706 363092 267734
rect 362224 266620 362276 266626
rect 362224 266562 362276 266568
rect 362788 266490 362816 267706
rect 361672 266484 361724 266490
rect 361672 266426 361724 266432
rect 362776 266484 362828 266490
rect 362776 266426 362828 266432
rect 360870 264302 361252 264330
rect 361684 264316 361712 266426
rect 362972 266370 363000 267706
rect 363328 267436 363380 267442
rect 363328 267378 363380 267384
rect 362880 266342 363000 266370
rect 362880 264330 362908 266342
rect 362526 264302 362908 264330
rect 363340 264316 363368 267378
rect 364168 264316 364196 271118
rect 364352 269686 364380 277766
rect 365732 269958 365760 277766
rect 367296 275466 367324 277780
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 368492 275330 368520 277780
rect 369124 275460 369176 275466
rect 369124 275402 369176 275408
rect 368480 275324 368532 275330
rect 368480 275266 368532 275272
rect 367100 274712 367152 274718
rect 367100 274654 367152 274660
rect 366916 274236 366968 274242
rect 366916 274178 366968 274184
rect 365720 269952 365772 269958
rect 365720 269894 365772 269900
rect 364984 269816 365036 269822
rect 364984 269758 365036 269764
rect 364340 269680 364392 269686
rect 364340 269622 364392 269628
rect 364996 264316 365024 269758
rect 365812 267572 365864 267578
rect 365812 267514 365864 267520
rect 365824 264316 365852 267514
rect 366928 264330 366956 274178
rect 367112 268394 367140 274654
rect 368388 272672 368440 272678
rect 368388 272614 368440 272620
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 368204 267300 368256 267306
rect 368204 267242 368256 267248
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 366956 264330
rect 367480 264316 367508 266358
rect 368216 264330 368244 267242
rect 368400 266422 368428 272614
rect 369136 267170 369164 275402
rect 369688 274718 369716 277780
rect 369872 277766 370898 277794
rect 369676 274712 369728 274718
rect 369676 274654 369728 274660
rect 369400 270360 369452 270366
rect 369400 270302 369452 270308
rect 369124 267164 369176 267170
rect 369124 267106 369176 267112
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 369412 264330 369440 270302
rect 369872 268530 369900 277766
rect 370504 275732 370556 275738
rect 370504 275674 370556 275680
rect 369860 268524 369912 268530
rect 369860 268466 369912 268472
rect 370320 268524 370372 268530
rect 370320 268466 370372 268472
rect 370332 264330 370360 268466
rect 370516 267442 370544 275674
rect 372080 271318 372108 277780
rect 373000 277766 373290 277794
rect 373000 272814 373028 277766
rect 373172 272944 373224 272950
rect 373172 272886 373224 272892
rect 372988 272808 373040 272814
rect 372988 272750 373040 272756
rect 372528 271720 372580 271726
rect 372528 271662 372580 271668
rect 372068 271312 372120 271318
rect 372068 271254 372120 271260
rect 372344 269952 372396 269958
rect 372344 269894 372396 269900
rect 370780 267708 370832 267714
rect 370780 267650 370832 267656
rect 370504 267436 370556 267442
rect 370504 267378 370556 267384
rect 368216 264302 368322 264330
rect 369150 264302 369440 264330
rect 369978 264302 370360 264330
rect 370792 264316 370820 267650
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 371620 264316 371648 266358
rect 372356 264330 372384 269894
rect 372540 266422 372568 271662
rect 373184 267734 373212 272886
rect 374380 271454 374408 277780
rect 375392 277766 375590 277794
rect 375104 275324 375156 275330
rect 375104 275266 375156 275272
rect 374368 271448 374420 271454
rect 374368 271390 374420 271396
rect 374920 268388 374972 268394
rect 374920 268330 374972 268336
rect 373092 267706 373212 267734
rect 373092 266898 373120 267706
rect 373264 267436 373316 267442
rect 373264 267378 373316 267384
rect 373080 266892 373132 266898
rect 373080 266834 373132 266840
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267378
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 268330
rect 375116 266422 375144 275266
rect 375392 270094 375420 277766
rect 376772 270502 376800 277780
rect 377968 275466 377996 277780
rect 378152 277766 379178 277794
rect 377956 275460 378008 275466
rect 377956 275402 378008 275408
rect 377772 274100 377824 274106
rect 377772 274042 377824 274048
rect 376760 270496 376812 270502
rect 376760 270438 376812 270444
rect 377588 270496 377640 270502
rect 377588 270438 377640 270444
rect 375380 270088 375432 270094
rect 375380 270030 375432 270036
rect 376576 270088 376628 270094
rect 376576 270030 376628 270036
rect 375748 267164 375800 267170
rect 375748 267106 375800 267112
rect 375104 266416 375156 266422
rect 375104 266358 375156 266364
rect 375760 264316 375788 267106
rect 376588 264316 376616 270030
rect 377600 267578 377628 270438
rect 377588 267572 377640 267578
rect 377588 267514 377640 267520
rect 377784 264330 377812 274042
rect 378152 270230 378180 277766
rect 380360 272542 380388 277780
rect 381188 277766 381570 277794
rect 380716 272808 380768 272814
rect 380716 272750 380768 272756
rect 380348 272536 380400 272542
rect 380348 272478 380400 272484
rect 379428 271448 379480 271454
rect 379428 271390 379480 271396
rect 378140 270224 378192 270230
rect 378140 270166 378192 270172
rect 378232 267028 378284 267034
rect 378232 266970 378284 266976
rect 377430 264302 377812 264330
rect 378244 264316 378272 266970
rect 379440 264330 379468 271390
rect 380532 266552 380584 266558
rect 380532 266494 380584 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380544 264330 380572 266494
rect 380728 266422 380756 272750
rect 381188 271590 381216 277766
rect 382280 275460 382332 275466
rect 382280 275402 382332 275408
rect 381360 271856 381412 271862
rect 381360 271798 381412 271804
rect 381176 271584 381228 271590
rect 381176 271526 381228 271532
rect 381372 267714 381400 271798
rect 382292 270230 382320 275402
rect 382660 272950 382688 277780
rect 383856 273970 383884 277780
rect 385052 275602 385080 277780
rect 385040 275596 385092 275602
rect 385040 275538 385092 275544
rect 386052 274712 386104 274718
rect 386052 274654 386104 274660
rect 384948 274372 385000 274378
rect 384948 274314 385000 274320
rect 383844 273964 383896 273970
rect 383844 273906 383896 273912
rect 382648 272944 382700 272950
rect 382648 272886 382700 272892
rect 382924 272536 382976 272542
rect 382924 272478 382976 272484
rect 381544 270224 381596 270230
rect 381544 270166 381596 270172
rect 382280 270224 382332 270230
rect 382280 270166 382332 270172
rect 381360 267708 381412 267714
rect 381360 267650 381412 267656
rect 380716 266416 380768 266422
rect 380716 266358 380768 266364
rect 380544 264302 380742 264330
rect 381556 264316 381584 270166
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 382384 264316 382412 268874
rect 382936 266558 382964 272478
rect 384028 269680 384080 269686
rect 384028 269622 384080 269628
rect 383200 267572 383252 267578
rect 383200 267514 383252 267520
rect 382924 266552 382976 266558
rect 382924 266494 382976 266500
rect 383212 264316 383240 267514
rect 384040 264316 384068 269622
rect 384960 267734 384988 274314
rect 385500 273964 385552 273970
rect 385500 273906 385552 273912
rect 384868 267706 384988 267734
rect 384868 264316 384896 267706
rect 385512 267306 385540 273906
rect 386064 271182 386092 274654
rect 386248 274514 386276 277780
rect 386432 277766 387458 277794
rect 386236 274508 386288 274514
rect 386236 274450 386288 274456
rect 386052 271176 386104 271182
rect 386052 271118 386104 271124
rect 385684 270224 385736 270230
rect 385684 270166 385736 270172
rect 385500 267300 385552 267306
rect 385500 267242 385552 267248
rect 385696 264316 385724 270166
rect 386432 268666 386460 277766
rect 388640 275738 388668 277780
rect 389180 276004 389232 276010
rect 389180 275946 389232 275952
rect 388628 275732 388680 275738
rect 388628 275674 388680 275680
rect 388076 275596 388128 275602
rect 388076 275538 388128 275544
rect 387708 271312 387760 271318
rect 387708 271254 387760 271260
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386420 268660 386472 268666
rect 386420 268602 386472 268608
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271254
rect 388088 269686 388116 275538
rect 389192 274242 389220 275946
rect 389744 274718 389772 277780
rect 390572 277766 390954 277794
rect 391952 277766 392150 277794
rect 389732 274712 389784 274718
rect 389732 274654 389784 274660
rect 389180 274236 389232 274242
rect 389180 274178 389232 274184
rect 390284 274236 390336 274242
rect 390284 274178 390336 274184
rect 389088 271040 389140 271046
rect 389088 270982 389140 270988
rect 388076 269680 388128 269686
rect 388076 269622 388128 269628
rect 389100 267734 389128 270982
rect 389008 267706 389128 267734
rect 388168 266892 388220 266898
rect 388168 266834 388220 266840
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 266834
rect 389008 264316 389036 267706
rect 390296 264330 390324 274178
rect 390572 269822 390600 277766
rect 391756 272944 391808 272950
rect 391756 272886 391808 272892
rect 390560 269816 390612 269822
rect 390560 269758 390612 269764
rect 390468 269544 390520 269550
rect 390468 269486 390520 269492
rect 390480 267442 390508 269486
rect 390468 267436 390520 267442
rect 390468 267378 390520 267384
rect 390652 267436 390704 267442
rect 390652 267378 390704 267384
rect 389850 264302 390324 264330
rect 390664 264316 390692 267378
rect 391768 264330 391796 272886
rect 391952 270502 391980 277766
rect 393332 276010 393360 277780
rect 393792 277766 394542 277794
rect 393320 276004 393372 276010
rect 393320 275946 393372 275952
rect 393792 272678 393820 277766
rect 395724 273970 395752 277780
rect 396092 277766 396934 277794
rect 397472 277766 398038 277794
rect 395896 274508 395948 274514
rect 395896 274450 395948 274456
rect 395712 273964 395764 273970
rect 395712 273906 395764 273912
rect 393780 272672 393832 272678
rect 393780 272614 393832 272620
rect 393964 272672 394016 272678
rect 393964 272614 394016 272620
rect 391940 270496 391992 270502
rect 391940 270438 391992 270444
rect 392308 269816 392360 269822
rect 392308 269758 392360 269764
rect 391506 264302 391796 264330
rect 392320 264316 392348 269758
rect 393136 267708 393188 267714
rect 393136 267650 393188 267656
rect 393148 264316 393176 267650
rect 393976 267170 394004 272614
rect 394332 271584 394384 271590
rect 394332 271526 394384 271532
rect 393964 267164 394016 267170
rect 393964 267106 394016 267112
rect 394344 264330 394372 271526
rect 394700 269680 394752 269686
rect 394700 269622 394752 269628
rect 394712 267578 394740 269622
rect 394700 267572 394752 267578
rect 394700 267514 394752 267520
rect 394792 266552 394844 266558
rect 394792 266494 394844 266500
rect 393990 264302 394372 264330
rect 394804 264316 394832 266494
rect 395908 264330 395936 274450
rect 396092 270366 396120 277766
rect 396356 275868 396408 275874
rect 396356 275810 396408 275816
rect 396368 272814 396396 275810
rect 397276 273080 397328 273086
rect 397276 273022 397328 273028
rect 396356 272808 396408 272814
rect 396356 272750 396408 272756
rect 396264 270496 396316 270502
rect 396264 270438 396316 270444
rect 396080 270360 396132 270366
rect 396080 270302 396132 270308
rect 396276 266898 396304 270438
rect 397092 267300 397144 267306
rect 397092 267242 397144 267248
rect 396264 266892 396316 266898
rect 396264 266834 396316 266840
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 395646 264302 395936 264330
rect 396460 264316 396488 266358
rect 397104 264330 397132 267242
rect 397288 266422 397316 273022
rect 397472 268530 397500 277766
rect 399220 271862 399248 277780
rect 399208 271856 399260 271862
rect 399208 271798 399260 271804
rect 400416 271726 400444 277780
rect 401626 277766 401916 277794
rect 400588 275188 400640 275194
rect 400588 275130 400640 275136
rect 400404 271720 400456 271726
rect 400404 271662 400456 271668
rect 400128 270632 400180 270638
rect 400128 270574 400180 270580
rect 397644 268660 397696 268666
rect 397644 268602 397696 268608
rect 397460 268524 397512 268530
rect 397460 268466 397512 268472
rect 397656 266558 397684 268602
rect 399760 267572 399812 267578
rect 399760 267514 399812 267520
rect 398104 266756 398156 266762
rect 398104 266698 398156 266704
rect 397644 266552 397696 266558
rect 397644 266494 397696 266500
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 266698
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 267514
rect 400140 266422 400168 270574
rect 400600 268938 400628 275130
rect 401324 271720 401376 271726
rect 401324 271662 401376 271668
rect 400588 268932 400640 268938
rect 400588 268874 400640 268880
rect 400588 268524 400640 268530
rect 400588 268466 400640 268472
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 268466
rect 401336 264330 401364 271662
rect 401888 269958 401916 277766
rect 402440 277766 402822 277794
rect 402060 270360 402112 270366
rect 402060 270302 402112 270308
rect 401876 269952 401928 269958
rect 401876 269894 401928 269900
rect 401600 269544 401652 269550
rect 401600 269486 401652 269492
rect 401612 267442 401640 269486
rect 402072 267714 402100 270302
rect 402440 269414 402468 277766
rect 404004 275330 404032 277780
rect 404464 277766 405214 277794
rect 403992 275324 404044 275330
rect 403992 275266 404044 275272
rect 404268 274712 404320 274718
rect 404268 274654 404320 274660
rect 403992 272808 404044 272814
rect 403992 272750 404044 272756
rect 403072 270088 403124 270094
rect 403072 270030 403124 270036
rect 402428 269408 402480 269414
rect 402428 269350 402480 269356
rect 402060 267708 402112 267714
rect 402060 267650 402112 267656
rect 401600 267436 401652 267442
rect 401600 267378 401652 267384
rect 402244 266892 402296 266898
rect 402244 266834 402296 266840
rect 401336 264302 401442 264330
rect 402256 264316 402284 266834
rect 403084 264316 403112 270030
rect 404004 267734 404032 272750
rect 404280 269958 404308 274654
rect 404268 269952 404320 269958
rect 404268 269894 404320 269900
rect 404464 268394 404492 277766
rect 405004 273964 405056 273970
rect 405004 273906 405056 273912
rect 404452 268388 404504 268394
rect 404452 268330 404504 268336
rect 403912 267706 404032 267734
rect 403912 264316 403940 267706
rect 404728 267164 404780 267170
rect 404728 267106 404780 267112
rect 404740 264316 404768 267106
rect 405016 266898 405044 273906
rect 406304 272678 406332 277780
rect 407120 274848 407172 274854
rect 407120 274790 407172 274796
rect 406844 273828 406896 273834
rect 406844 273770 406896 273776
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 405556 267708 405608 267714
rect 405556 267650 405608 267656
rect 405004 266892 405056 266898
rect 405004 266834 405056 266840
rect 405568 264316 405596 267650
rect 406856 264330 406884 273770
rect 407132 271454 407160 274790
rect 407500 274718 407528 277780
rect 407488 274712 407540 274718
rect 407488 274654 407540 274660
rect 408696 274106 408724 277780
rect 409892 274718 409920 277780
rect 410064 275732 410116 275738
rect 410064 275674 410116 275680
rect 409144 274712 409196 274718
rect 409144 274654 409196 274660
rect 409880 274712 409932 274718
rect 409880 274654 409932 274660
rect 408684 274100 408736 274106
rect 408684 274042 408736 274048
rect 408408 272672 408460 272678
rect 408408 272614 408460 272620
rect 407120 271448 407172 271454
rect 407120 271390 407172 271396
rect 407212 268388 407264 268394
rect 407212 268330 407264 268336
rect 406410 264302 406884 264330
rect 407224 264316 407252 268330
rect 408420 264330 408448 272614
rect 409156 267034 409184 274654
rect 410076 272950 410104 275674
rect 411088 274854 411116 277780
rect 412284 275874 412312 277780
rect 413100 276004 413152 276010
rect 413100 275946 413152 275952
rect 412272 275868 412324 275874
rect 412272 275810 412324 275816
rect 411260 275324 411312 275330
rect 411260 275266 411312 275272
rect 411076 274848 411128 274854
rect 411076 274790 411128 274796
rect 410248 274644 410300 274650
rect 410248 274586 410300 274592
rect 410260 273834 410288 274586
rect 410248 273828 410300 273834
rect 410248 273770 410300 273776
rect 410064 272944 410116 272950
rect 410064 272886 410116 272892
rect 411272 271946 411300 275266
rect 413112 274514 413140 275946
rect 413100 274508 413152 274514
rect 413100 274450 413152 274456
rect 412456 272944 412508 272950
rect 412456 272886 412508 272892
rect 410904 271918 411300 271946
rect 409788 271448 409840 271454
rect 409788 271390 409840 271396
rect 409604 267436 409656 267442
rect 409604 267378 409656 267384
rect 409144 267028 409196 267034
rect 409144 266970 409196 266976
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408066 264302 408448 264330
rect 408880 264316 408908 266358
rect 409616 264330 409644 267378
rect 409800 266422 409828 271390
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410904 264330 410932 271918
rect 411904 271856 411956 271862
rect 411904 271798 411956 271804
rect 411916 266762 411944 271798
rect 412180 266892 412232 266898
rect 412180 266834 412232 266840
rect 411904 266756 411956 266762
rect 411904 266698 411956 266704
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 409616 264302 409722 264330
rect 410550 264302 410932 264330
rect 411364 264316 411392 266358
rect 412192 264316 412220 266834
rect 412468 266422 412496 272886
rect 413388 272542 413416 277780
rect 414584 275466 414612 277780
rect 414572 275460 414624 275466
rect 414572 275402 414624 275408
rect 415308 275460 415360 275466
rect 415308 275402 415360 275408
rect 413928 274100 413980 274106
rect 413928 274042 413980 274048
rect 413376 272536 413428 272542
rect 413376 272478 413428 272484
rect 413940 267734 413968 274042
rect 415124 272536 415176 272542
rect 415124 272478 415176 272484
rect 413848 267706 413968 267734
rect 413008 266756 413060 266762
rect 413008 266698 413060 266704
rect 412456 266416 412508 266422
rect 412456 266358 412508 266364
rect 413020 264316 413048 266698
rect 413848 264316 413876 267706
rect 415136 264330 415164 272478
rect 415320 271046 415348 275402
rect 415780 275194 415808 277780
rect 416792 277766 416990 277794
rect 416412 275868 416464 275874
rect 416412 275810 416464 275816
rect 415768 275188 415820 275194
rect 415768 275130 415820 275136
rect 415308 271040 415360 271046
rect 415308 270982 415360 270988
rect 416424 266422 416452 275810
rect 416596 270904 416648 270910
rect 416596 270846 416648 270852
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415164 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 270846
rect 416792 269686 416820 277766
rect 418172 275602 418200 277780
rect 418160 275596 418212 275602
rect 418160 275538 418212 275544
rect 418344 275596 418396 275602
rect 418344 275538 418396 275544
rect 418356 273086 418384 275538
rect 419368 274378 419396 277780
rect 419552 277766 420578 277794
rect 419356 274372 419408 274378
rect 419356 274314 419408 274320
rect 419172 273216 419224 273222
rect 419172 273158 419224 273164
rect 418344 273080 418396 273086
rect 418344 273022 418396 273028
rect 418068 270768 418120 270774
rect 418068 270710 418120 270716
rect 417148 269952 417200 269958
rect 417148 269894 417200 269900
rect 416780 269680 416832 269686
rect 416780 269622 416832 269628
rect 416346 264302 416636 264330
rect 417160 264316 417188 269894
rect 418080 267734 418108 270710
rect 418988 268932 419040 268938
rect 418988 268874 419040 268880
rect 417988 267706 418108 267734
rect 417988 264316 418016 267706
rect 419000 267578 419028 268874
rect 418988 267572 419040 267578
rect 418988 267514 419040 267520
rect 419184 264330 419212 273158
rect 419552 270230 419580 277766
rect 421668 271318 421696 277780
rect 422312 277766 422878 277794
rect 423692 277766 424074 277794
rect 421656 271312 421708 271318
rect 421656 271254 421708 271260
rect 422116 271312 422168 271318
rect 422116 271254 422168 271260
rect 419540 270224 419592 270230
rect 419540 270166 419592 270172
rect 419632 269408 419684 269414
rect 419632 269350 419684 269356
rect 418830 264302 419212 264330
rect 419644 264316 419672 269350
rect 420920 269272 420972 269278
rect 420920 269214 420972 269220
rect 420460 268252 420512 268258
rect 420460 268194 420512 268200
rect 420472 264316 420500 268194
rect 420932 267714 420960 269214
rect 420920 267708 420972 267714
rect 420920 267650 420972 267656
rect 422128 267034 422156 271254
rect 422312 269074 422340 277766
rect 423692 270502 423720 277766
rect 425256 275466 425284 277780
rect 425244 275460 425296 275466
rect 425244 275402 425296 275408
rect 425336 274780 425388 274786
rect 425336 274722 425388 274728
rect 424968 274372 425020 274378
rect 424968 274314 425020 274320
rect 423680 270496 423732 270502
rect 423680 270438 423732 270444
rect 424600 269680 424652 269686
rect 424600 269622 424652 269628
rect 422300 269068 422352 269074
rect 422300 269010 422352 269016
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422312 267306 422340 268738
rect 422300 267300 422352 267306
rect 422300 267242 422352 267248
rect 421288 267028 421340 267034
rect 421288 266970 421340 266976
rect 422116 267028 422168 267034
rect 422116 266970 422168 266976
rect 422300 267028 422352 267034
rect 422300 266970 422352 266976
rect 421300 264316 421328 266970
rect 422312 266914 422340 266970
rect 422220 266886 422340 266914
rect 422220 266506 422248 266886
rect 422944 266620 422996 266626
rect 422944 266562 422996 266568
rect 422220 266478 422294 266506
rect 422266 266234 422294 266478
rect 422128 266206 422294 266234
rect 422128 264316 422156 266206
rect 422956 264316 422984 266562
rect 423772 266416 423824 266422
rect 423772 266358 423824 266364
rect 423784 264316 423812 266358
rect 424612 264316 424640 269622
rect 424980 266422 425008 274314
rect 425348 271590 425376 274722
rect 426452 274242 426480 277780
rect 426636 277766 427662 277794
rect 426440 274236 426492 274242
rect 426440 274178 426492 274184
rect 426348 273080 426400 273086
rect 426348 273022 426400 273028
rect 425336 271584 425388 271590
rect 425336 271526 425388 271532
rect 426360 267734 426388 273022
rect 426636 269550 426664 277766
rect 428844 275738 428872 277780
rect 429396 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275732 428884 275738
rect 428832 275674 428884 275680
rect 429200 275460 429252 275466
rect 429200 275402 429252 275408
rect 427820 275188 427872 275194
rect 427820 275130 427872 275136
rect 427084 274508 427136 274514
rect 427084 274450 427136 274456
rect 426624 269544 426676 269550
rect 426624 269486 426676 269492
rect 426268 267706 426388 267734
rect 424968 266416 425020 266422
rect 424968 266358 425020 266364
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 267706
rect 427096 266422 427124 274450
rect 427832 271726 427860 275130
rect 428464 273828 428516 273834
rect 428464 273770 428516 273776
rect 427820 271720 427872 271726
rect 427820 271662 427872 271668
rect 428280 270224 428332 270230
rect 428280 270166 428332 270172
rect 427360 269544 427412 269550
rect 427360 269486 427412 269492
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427372 264330 427400 269486
rect 427912 267300 427964 267306
rect 427912 267242 427964 267248
rect 427110 264302 427400 264330
rect 427924 264316 427952 267242
rect 428292 266762 428320 270166
rect 428476 266898 428504 273770
rect 429212 272814 429240 275402
rect 429200 272808 429252 272814
rect 429200 272750 429252 272756
rect 429396 269822 429424 277766
rect 429568 270496 429620 270502
rect 429568 270438 429620 270444
rect 429384 269816 429436 269822
rect 429384 269758 429436 269764
rect 428464 266892 428516 266898
rect 428464 266834 428516 266840
rect 428280 266756 428332 266762
rect 428280 266698 428332 266704
rect 428740 266756 428792 266762
rect 428740 266698 428792 266704
rect 428752 264316 428780 266698
rect 429580 264316 429608 270438
rect 430592 270366 430620 277766
rect 432340 274786 432368 277780
rect 433352 277766 433550 277794
rect 433156 275732 433208 275738
rect 433156 275674 433208 275680
rect 432328 274780 432380 274786
rect 432328 274722 432380 274728
rect 431684 271176 431736 271182
rect 431684 271118 431736 271124
rect 430580 270360 430632 270366
rect 430580 270302 430632 270308
rect 430396 267572 430448 267578
rect 430396 267514 430448 267520
rect 430408 264316 430436 267514
rect 431696 264330 431724 271118
rect 431960 267844 432012 267850
rect 431960 267786 432012 267792
rect 431972 267170 432000 267786
rect 431960 267164 432012 267170
rect 431960 267106 432012 267112
rect 432328 267164 432380 267170
rect 432328 267106 432380 267112
rect 432340 264330 432368 267106
rect 433168 264330 433196 275674
rect 433352 268666 433380 277766
rect 434732 276010 434760 277780
rect 434720 276004 434772 276010
rect 434720 275946 434772 275952
rect 435928 275602 435956 277780
rect 436112 277766 437046 277794
rect 435916 275596 435968 275602
rect 435916 275538 435968 275544
rect 435548 274780 435600 274786
rect 435548 274722 435600 274728
rect 434628 272808 434680 272814
rect 434628 272750 434680 272756
rect 434444 269816 434496 269822
rect 434444 269758 434496 269764
rect 433340 268660 433392 268666
rect 433340 268602 433392 268608
rect 433708 266416 433760 266422
rect 433708 266358 433760 266364
rect 431250 264302 431724 264330
rect 432078 264302 432368 264330
rect 432906 264302 433196 264330
rect 433720 264316 433748 266358
rect 434456 264330 434484 269758
rect 434640 266422 434668 272750
rect 435364 271448 435416 271454
rect 435364 271390 435416 271396
rect 435376 267442 435404 271390
rect 435560 270638 435588 274722
rect 435548 270632 435600 270638
rect 435548 270574 435600 270580
rect 436112 268802 436140 277766
rect 437480 276004 437532 276010
rect 437480 275946 437532 275952
rect 437492 274650 437520 275946
rect 437480 274644 437532 274650
rect 437480 274586 437532 274592
rect 438228 271862 438256 277780
rect 439056 277766 439438 277794
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439056 274786 439084 277766
rect 439504 275596 439556 275602
rect 439504 275538 439556 275544
rect 439044 274780 439096 274786
rect 439044 274722 439096 274728
rect 438768 274236 438820 274242
rect 438768 274178 438820 274184
rect 438216 271856 438268 271862
rect 438216 271798 438268 271804
rect 437388 270632 437440 270638
rect 437388 270574 437440 270580
rect 436100 268796 436152 268802
rect 436100 268738 436152 268744
rect 436192 268116 436244 268122
rect 436192 268058 436244 268064
rect 435364 267436 435416 267442
rect 435364 267378 435416 267384
rect 435364 266892 435416 266898
rect 435364 266834 435416 266840
rect 434628 266416 434680 266422
rect 434628 266358 434680 266364
rect 434456 264302 434562 264330
rect 435376 264316 435404 266834
rect 436204 264316 436232 268058
rect 437400 264330 437428 270574
rect 438780 267734 438808 274178
rect 438688 267706 438808 267734
rect 437848 266416 437900 266422
rect 437848 266358 437900 266364
rect 437046 264302 437428 264330
rect 437860 264316 437888 266358
rect 438688 264316 438716 267706
rect 439516 266422 439544 275538
rect 439964 271040 440016 271046
rect 439964 270982 440016 270988
rect 439688 266892 439740 266898
rect 439688 266834 439740 266840
rect 439700 266490 439728 266834
rect 439688 266484 439740 266490
rect 439688 266426 439740 266432
rect 439504 266416 439556 266422
rect 439504 266358 439556 266364
rect 439976 264330 440004 270982
rect 440252 268938 440280 277766
rect 440884 274644 440936 274650
rect 440884 274586 440936 274592
rect 440240 268932 440292 268938
rect 440240 268874 440292 268880
rect 440332 267708 440384 267714
rect 440332 267650 440384 267656
rect 439530 264302 440004 264330
rect 440344 264316 440372 267650
rect 440896 267170 440924 274586
rect 441160 268932 441212 268938
rect 441160 268874 441212 268880
rect 440884 267164 440936 267170
rect 440884 267106 440936 267112
rect 441172 264316 441200 268874
rect 441632 268530 441660 277766
rect 443012 275194 443040 277780
rect 443000 275188 443052 275194
rect 443000 275130 443052 275136
rect 443368 275052 443420 275058
rect 443368 274994 443420 275000
rect 443380 271590 443408 274994
rect 444208 273970 444236 277780
rect 444392 277766 445326 277794
rect 444196 273964 444248 273970
rect 444196 273906 444248 273912
rect 443644 271856 443696 271862
rect 443644 271798 443696 271804
rect 443368 271584 443420 271590
rect 443368 271526 443420 271532
rect 441620 268524 441672 268530
rect 441620 268466 441672 268472
rect 442816 267980 442868 267986
rect 442816 267922 442868 267928
rect 441804 266892 441856 266898
rect 441804 266834 441856 266840
rect 441816 266626 441844 266834
rect 441804 266620 441856 266626
rect 441804 266562 441856 266568
rect 441988 266620 442040 266626
rect 441988 266562 442040 266568
rect 442000 264316 442028 266562
rect 442828 264316 442856 267922
rect 443656 266626 443684 271798
rect 444392 270094 444420 277766
rect 446508 275466 446536 277780
rect 447152 277766 447718 277794
rect 448532 277766 448914 277794
rect 446496 275460 446548 275466
rect 446496 275402 446548 275408
rect 445944 275188 445996 275194
rect 445944 275130 445996 275136
rect 445668 271584 445720 271590
rect 445668 271526 445720 271532
rect 444380 270088 444432 270094
rect 444380 270030 444432 270036
rect 443920 269068 443972 269074
rect 443920 269010 443972 269016
rect 443644 266620 443696 266626
rect 443644 266562 443696 266568
rect 443932 264330 443960 269010
rect 445680 266626 445708 271526
rect 445956 271318 445984 275130
rect 445944 271312 445996 271318
rect 445944 271254 445996 271260
rect 446956 270360 447008 270366
rect 446956 270302 447008 270308
rect 446128 268796 446180 268802
rect 446128 268738 446180 268744
rect 445944 267436 445996 267442
rect 445944 267378 445996 267384
rect 445956 267034 445984 267378
rect 445944 267028 445996 267034
rect 445944 266970 445996 266976
rect 444472 266620 444524 266626
rect 444472 266562 444524 266568
rect 445668 266620 445720 266626
rect 445668 266562 445720 266568
rect 445852 266620 445904 266626
rect 445852 266562 445904 266568
rect 443670 264302 443960 264330
rect 444484 264316 444512 266562
rect 445864 266506 445892 266562
rect 445680 266478 445892 266506
rect 445680 264330 445708 266478
rect 445326 264302 445708 264330
rect 446140 264316 446168 268738
rect 446968 264316 446996 270302
rect 447152 267850 447180 277766
rect 447600 272264 447652 272270
rect 447600 272206 447652 272212
rect 447140 267844 447192 267850
rect 447140 267786 447192 267792
rect 447612 266898 447640 272206
rect 447784 270088 447836 270094
rect 447784 270030 447836 270036
rect 447600 266892 447652 266898
rect 447600 266834 447652 266840
rect 447796 264316 447824 270030
rect 448532 269278 448560 277766
rect 450096 276010 450124 277780
rect 451306 277766 451504 277794
rect 450084 276004 450136 276010
rect 450084 275946 450136 275952
rect 449900 275460 449952 275466
rect 449900 275402 449952 275408
rect 449912 270094 449940 275402
rect 451188 273964 451240 273970
rect 451188 273906 451240 273912
rect 449900 270088 449952 270094
rect 449900 270030 449952 270036
rect 448520 269272 448572 269278
rect 448520 269214 448572 269220
rect 450728 269272 450780 269278
rect 450728 269214 450780 269220
rect 448612 268660 448664 268666
rect 448612 268602 448664 268608
rect 448624 264316 448652 268602
rect 450740 267442 450768 269214
rect 451200 267734 451228 273906
rect 451476 268394 451504 277766
rect 452488 272678 452516 277780
rect 453592 275058 453620 277780
rect 454512 277766 454802 277794
rect 453580 275052 453632 275058
rect 453580 274994 453632 275000
rect 453396 274916 453448 274922
rect 453396 274858 453448 274864
rect 453408 272950 453436 274858
rect 453396 272944 453448 272950
rect 453396 272886 453448 272892
rect 452476 272672 452528 272678
rect 452476 272614 452528 272620
rect 453856 272672 453908 272678
rect 453856 272614 453908 272620
rect 451740 272400 451792 272406
rect 451740 272342 451792 272348
rect 451464 268388 451516 268394
rect 451464 268330 451516 268336
rect 451108 267706 451228 267734
rect 450728 267436 450780 267442
rect 450728 267378 450780 267384
rect 450912 267436 450964 267442
rect 450912 267378 450964 267384
rect 449440 267300 449492 267306
rect 449440 267242 449492 267248
rect 449452 264316 449480 267242
rect 450268 267164 450320 267170
rect 450268 267106 450320 267112
rect 450280 264316 450308 267106
rect 450924 266626 450952 267378
rect 450912 266620 450964 266626
rect 450912 266562 450964 266568
rect 451108 264316 451136 267706
rect 451752 267034 451780 272342
rect 453304 271720 453356 271726
rect 453304 271662 453356 271668
rect 453316 267306 453344 271662
rect 453304 267300 453356 267306
rect 453304 267242 453356 267248
rect 451740 267028 451792 267034
rect 451740 266970 451792 266976
rect 452752 266892 452804 266898
rect 452752 266834 452804 266840
rect 451924 266620 451976 266626
rect 451924 266562 451976 266568
rect 451936 264316 451964 266562
rect 452764 264316 452792 266834
rect 453868 264330 453896 272614
rect 454512 271454 454540 277766
rect 455984 275330 456012 277780
rect 456800 276004 456852 276010
rect 456800 275946 456852 275952
rect 455972 275324 456024 275330
rect 455972 275266 456024 275272
rect 456156 275324 456208 275330
rect 456156 275266 456208 275272
rect 456168 271538 456196 275266
rect 456812 274106 456840 275946
rect 457180 274922 457208 277780
rect 457168 274916 457220 274922
rect 457168 274858 457220 274864
rect 456800 274100 456852 274106
rect 456800 274042 456852 274048
rect 458376 273834 458404 277780
rect 459376 274100 459428 274106
rect 459376 274042 459428 274048
rect 458364 273828 458416 273834
rect 458364 273770 458416 273776
rect 457444 273692 457496 273698
rect 457444 273634 457496 273640
rect 455892 271510 456196 271538
rect 454500 271448 454552 271454
rect 454500 271390 454552 271396
rect 454684 271448 454736 271454
rect 454684 271390 454736 271396
rect 454408 267028 454460 267034
rect 454408 266970 454460 266976
rect 453606 264302 453896 264330
rect 454420 264316 454448 266970
rect 454696 266626 454724 271390
rect 455236 267300 455288 267306
rect 455236 267242 455288 267248
rect 454684 266620 454736 266626
rect 454684 266562 454736 266568
rect 455248 264316 455276 267242
rect 455892 266898 455920 271510
rect 456064 268524 456116 268530
rect 456064 268466 456116 268472
rect 455880 266892 455932 266898
rect 455880 266834 455932 266840
rect 456076 264316 456104 268466
rect 457456 267578 457484 273634
rect 458088 272944 458140 272950
rect 458088 272886 458140 272892
rect 457720 270088 457772 270094
rect 457720 270030 457772 270036
rect 457444 267572 457496 267578
rect 457444 267514 457496 267520
rect 456892 266620 456944 266626
rect 456892 266562 456944 266568
rect 456904 264316 456932 266562
rect 457732 264316 457760 270030
rect 458100 266626 458128 272886
rect 459192 267572 459244 267578
rect 459192 267514 459244 267520
rect 458088 266620 458140 266626
rect 458088 266562 458140 266568
rect 458548 266620 458600 266626
rect 458548 266562 458600 266568
rect 458560 264316 458588 266562
rect 459204 264330 459232 267514
rect 459388 266626 459416 274042
rect 459572 270230 459600 277780
rect 460676 276010 460704 277780
rect 460664 276004 460716 276010
rect 460664 275946 460716 275952
rect 460848 276004 460900 276010
rect 460848 275946 460900 275952
rect 459560 270224 459612 270230
rect 459560 270166 459612 270172
rect 460860 267986 460888 275946
rect 461872 272542 461900 277780
rect 463068 275874 463096 277780
rect 463988 277766 464278 277794
rect 465092 277766 465474 277794
rect 463056 275868 463108 275874
rect 463056 275810 463108 275816
rect 462964 275052 463016 275058
rect 462964 274994 463016 275000
rect 462228 274780 462280 274786
rect 462228 274722 462280 274728
rect 461860 272536 461912 272542
rect 461860 272478 461912 272484
rect 461584 271312 461636 271318
rect 461584 271254 461636 271260
rect 460848 267980 460900 267986
rect 460848 267922 460900 267928
rect 459560 267028 459612 267034
rect 459560 266970 459612 266976
rect 460204 267028 460256 267034
rect 460204 266970 460256 266976
rect 459572 266626 459600 266970
rect 459376 266620 459428 266626
rect 459376 266562 459428 266568
rect 459560 266620 459612 266626
rect 459560 266562 459612 266568
rect 459204 264302 459402 264330
rect 460216 264316 460244 266970
rect 461032 266892 461084 266898
rect 461032 266834 461084 266840
rect 461044 264316 461072 266834
rect 461596 266626 461624 271254
rect 462240 270774 462268 274722
rect 462976 273222 463004 274994
rect 462964 273216 463016 273222
rect 462964 273158 463016 273164
rect 463516 272536 463568 272542
rect 463516 272478 463568 272484
rect 463148 272128 463200 272134
rect 463148 272070 463200 272076
rect 462228 270768 462280 270774
rect 462228 270710 462280 270716
rect 461860 270224 461912 270230
rect 461860 270166 461912 270172
rect 461584 266620 461636 266626
rect 461584 266562 461636 266568
rect 461872 264316 461900 270166
rect 463160 264330 463188 272070
rect 462714 264302 463188 264330
rect 463528 264316 463556 272478
rect 463988 270910 464016 277766
rect 463976 270904 464028 270910
rect 463976 270846 464028 270852
rect 464344 270904 464396 270910
rect 464344 270846 464396 270852
rect 464356 267578 464384 270846
rect 464804 270768 464856 270774
rect 464804 270710 464856 270716
rect 464344 267572 464396 267578
rect 464344 267514 464396 267520
rect 464816 264330 464844 270710
rect 465092 269958 465120 277766
rect 466656 274786 466684 277780
rect 467852 275058 467880 277780
rect 468312 277766 468970 277794
rect 469232 277766 470166 277794
rect 467840 275052 467892 275058
rect 467840 274994 467892 275000
rect 467748 274916 467800 274922
rect 467748 274858 467800 274864
rect 466644 274780 466696 274786
rect 466644 274722 466696 274728
rect 465724 273828 465776 273834
rect 465724 273770 465776 273776
rect 465080 269952 465132 269958
rect 465080 269894 465132 269900
rect 465172 267572 465224 267578
rect 465172 267514 465224 267520
rect 464370 264302 464844 264330
rect 465184 264316 465212 267514
rect 465736 266762 465764 273770
rect 467760 273254 467788 274858
rect 467668 273226 467788 273254
rect 466000 269952 466052 269958
rect 466000 269894 466052 269900
rect 465724 266756 465776 266762
rect 465724 266698 465776 266704
rect 466012 264316 466040 269894
rect 466828 268388 466880 268394
rect 466828 268330 466880 268336
rect 466840 264316 466868 268330
rect 467668 264316 467696 273226
rect 468312 269414 468340 277766
rect 469232 273254 469260 277766
rect 471152 275868 471204 275874
rect 471152 275810 471204 275816
rect 469232 273226 469444 273254
rect 469220 269816 469272 269822
rect 469220 269758 469272 269764
rect 469232 269414 469260 269758
rect 468300 269408 468352 269414
rect 468300 269350 468352 269356
rect 469220 269408 469272 269414
rect 469220 269350 469272 269356
rect 468758 269240 468814 269249
rect 468758 269175 468814 269184
rect 468772 264330 468800 269175
rect 469416 268258 469444 273226
rect 470048 272264 470100 272270
rect 470048 272206 470100 272212
rect 470060 271998 470088 272206
rect 470048 271992 470100 271998
rect 470048 271934 470100 271940
rect 471164 270638 471192 275810
rect 471348 275194 471376 277780
rect 471992 277766 472558 277794
rect 471336 275188 471388 275194
rect 471336 275130 471388 275136
rect 471428 272400 471480 272406
rect 471428 272342 471480 272348
rect 471440 272134 471468 272342
rect 471428 272128 471480 272134
rect 471428 272070 471480 272076
rect 471152 270632 471204 270638
rect 471152 270574 471204 270580
rect 470968 269816 471020 269822
rect 470968 269758 471020 269764
rect 469404 268252 469456 268258
rect 469404 268194 469456 268200
rect 470140 268252 470192 268258
rect 470140 268194 470192 268200
rect 470152 266898 470180 268194
rect 470140 266892 470192 266898
rect 470140 266834 470192 266840
rect 470140 266620 470192 266626
rect 470140 266562 470192 266568
rect 469312 266484 469364 266490
rect 469312 266426 469364 266432
rect 468510 264302 468800 264330
rect 469324 264316 469352 266426
rect 470152 264316 470180 266562
rect 470980 264316 471008 269758
rect 471992 269278 472020 277766
rect 473084 275052 473136 275058
rect 473084 274994 473136 275000
rect 471980 269272 472032 269278
rect 471980 269214 472032 269220
rect 471796 266892 471848 266898
rect 471796 266834 471848 266840
rect 471808 264316 471836 266834
rect 473096 264330 473124 274994
rect 473452 273216 473504 273222
rect 473452 273158 473504 273164
rect 472650 264302 473124 264330
rect 473464 264316 473492 273158
rect 473740 271998 473768 277780
rect 474936 274378 474964 277780
rect 476146 277766 476344 277794
rect 474924 274372 474976 274378
rect 474924 274314 474976 274320
rect 475568 273556 475620 273562
rect 475568 273498 475620 273504
rect 473728 271992 473780 271998
rect 473728 271934 473780 271940
rect 474740 270632 474792 270638
rect 474740 270574 474792 270580
rect 474280 269272 474332 269278
rect 474280 269214 474332 269220
rect 474292 264316 474320 269214
rect 474752 266490 474780 270574
rect 475384 269680 475436 269686
rect 475384 269622 475436 269628
rect 475396 269521 475424 269622
rect 475382 269512 475438 269521
rect 475382 269447 475438 269456
rect 475580 266898 475608 273498
rect 476028 269816 476080 269822
rect 475750 269784 475806 269793
rect 476028 269758 476080 269764
rect 475750 269719 475806 269728
rect 475764 269550 475792 269719
rect 475752 269544 475804 269550
rect 475752 269486 475804 269492
rect 476040 269249 476068 269758
rect 476316 269521 476344 277766
rect 477236 274514 477264 277780
rect 477224 274508 477276 274514
rect 477224 274450 477276 274456
rect 476580 274372 476632 274378
rect 476580 274314 476632 274320
rect 477684 274372 477736 274378
rect 477684 274314 477736 274320
rect 476302 269512 476358 269521
rect 476302 269447 476358 269456
rect 476026 269240 476082 269249
rect 476026 269175 476082 269184
rect 475568 266892 475620 266898
rect 475568 266834 475620 266840
rect 476592 266762 476620 274314
rect 477696 273562 477724 274314
rect 477684 273556 477736 273562
rect 477684 273498 477736 273504
rect 478432 273086 478460 277780
rect 478892 277766 479642 277794
rect 478420 273080 478472 273086
rect 478420 273022 478472 273028
rect 478696 271992 478748 271998
rect 478696 271934 478748 271940
rect 476764 269272 476816 269278
rect 476764 269214 476816 269220
rect 476580 266756 476632 266762
rect 476580 266698 476632 266704
rect 474740 266484 474792 266490
rect 474740 266426 474792 266432
rect 475936 266484 475988 266490
rect 475936 266426 475988 266432
rect 475108 266076 475160 266082
rect 475108 266018 475160 266024
rect 475120 264316 475148 266018
rect 475948 264316 475976 266426
rect 476776 264316 476804 269214
rect 477592 266892 477644 266898
rect 477592 266834 477644 266840
rect 477604 264316 477632 266834
rect 478708 264330 478736 271934
rect 478892 269793 478920 277766
rect 480824 272134 480852 277780
rect 482020 273834 482048 277780
rect 483216 277394 483244 277780
rect 483124 277366 483244 277394
rect 482008 273828 482060 273834
rect 482008 273770 482060 273776
rect 482468 273556 482520 273562
rect 482468 273498 482520 273504
rect 481364 273420 481416 273426
rect 481364 273362 481416 273368
rect 480812 272128 480864 272134
rect 480812 272070 480864 272076
rect 480258 270736 480314 270745
rect 480258 270671 480314 270680
rect 480272 270586 480300 270671
rect 480180 270558 480300 270586
rect 480180 270502 480208 270558
rect 480168 270496 480220 270502
rect 480168 270438 480220 270444
rect 480352 270496 480404 270502
rect 480352 270438 480404 270444
rect 478878 269784 478934 269793
rect 478878 269719 478934 269728
rect 480364 269498 480392 270438
rect 480180 269470 480392 269498
rect 480180 269414 480208 269470
rect 479064 269408 479116 269414
rect 479062 269376 479064 269385
rect 479248 269408 479300 269414
rect 479116 269376 479118 269385
rect 479248 269350 479300 269356
rect 480168 269408 480220 269414
rect 480352 269408 480404 269414
rect 480168 269350 480220 269356
rect 480350 269376 480352 269385
rect 480404 269376 480406 269385
rect 479062 269311 479118 269320
rect 478446 264302 478736 264330
rect 479260 264316 479288 269350
rect 480350 269311 480406 269320
rect 480076 265668 480128 265674
rect 480076 265610 480128 265616
rect 480088 264316 480116 265610
rect 481376 264330 481404 273362
rect 482284 270088 482336 270094
rect 482282 270056 482284 270065
rect 482336 270056 482338 270065
rect 482282 269991 482338 270000
rect 481732 266756 481784 266762
rect 481732 266698 481784 266704
rect 480930 264302 481404 264330
rect 481744 264316 481772 266698
rect 482480 264330 482508 273498
rect 483124 270745 483152 277366
rect 484320 273698 484348 277780
rect 484584 275188 484636 275194
rect 484584 275130 484636 275136
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483756 272128 483808 272134
rect 483756 272070 483808 272076
rect 483110 270736 483166 270745
rect 483110 270671 483166 270680
rect 482652 270088 482704 270094
rect 482652 270030 482704 270036
rect 482664 269822 482692 270030
rect 482652 269816 482704 269822
rect 482652 269758 482704 269764
rect 483768 264330 483796 272070
rect 484044 271238 484440 271266
rect 484044 271182 484072 271238
rect 484032 271176 484084 271182
rect 484032 271118 484084 271124
rect 484216 271176 484268 271182
rect 484216 271118 484268 271124
rect 484228 270774 484256 271118
rect 484412 270774 484440 271238
rect 484216 270768 484268 270774
rect 484216 270710 484268 270716
rect 484400 270768 484452 270774
rect 484400 270710 484452 270716
rect 484596 270065 484624 275130
rect 485044 273080 485096 273086
rect 485044 273022 485096 273028
rect 485056 272406 485084 273022
rect 485044 272400 485096 272406
rect 485044 272342 485096 272348
rect 485516 270774 485544 277780
rect 486712 274650 486740 277780
rect 487908 275738 487936 277780
rect 488736 277766 489118 277794
rect 489932 277766 490314 277794
rect 487896 275732 487948 275738
rect 487896 275674 487948 275680
rect 488080 275732 488132 275738
rect 488080 275674 488132 275680
rect 488092 275194 488120 275674
rect 488080 275188 488132 275194
rect 488080 275130 488132 275136
rect 488540 274712 488592 274718
rect 488540 274654 488592 274660
rect 486700 274644 486752 274650
rect 486700 274586 486752 274592
rect 487068 273692 487120 273698
rect 487068 273634 487120 273640
rect 485504 270768 485556 270774
rect 485504 270710 485556 270716
rect 485044 270496 485096 270502
rect 485044 270438 485096 270444
rect 486700 270496 486752 270502
rect 486700 270438 486752 270444
rect 484582 270056 484638 270065
rect 484582 269991 484638 270000
rect 485056 269686 485084 270438
rect 485044 269680 485096 269686
rect 485044 269622 485096 269628
rect 484306 269512 484362 269521
rect 484306 269447 484362 269456
rect 484320 267734 484348 269447
rect 482480 264302 482586 264330
rect 483414 264302 483796 264330
rect 484228 267706 484348 267734
rect 484228 264316 484256 267706
rect 484858 266792 484914 266801
rect 484858 266727 484860 266736
rect 484912 266727 484914 266736
rect 485044 266756 485096 266762
rect 484860 266698 484912 266704
rect 485044 266698 485096 266704
rect 485056 266490 485084 266698
rect 485044 266484 485096 266490
rect 485044 266426 485096 266432
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 485044 265940 485096 265946
rect 485044 265882 485096 265888
rect 485056 264316 485084 265882
rect 485884 264316 485912 266358
rect 486712 264316 486740 270438
rect 487080 266422 487108 273634
rect 488356 272400 488408 272406
rect 488356 272342 488408 272348
rect 487988 272264 488040 272270
rect 487988 272206 488040 272212
rect 487252 267028 487304 267034
rect 487252 266970 487304 266976
rect 487436 267028 487488 267034
rect 487436 266970 487488 266976
rect 487264 266490 487292 266970
rect 487448 266801 487476 266970
rect 487434 266792 487490 266801
rect 487434 266727 487490 266736
rect 487252 266484 487304 266490
rect 487252 266426 487304 266432
rect 487068 266416 487120 266422
rect 487068 266358 487120 266364
rect 488000 264330 488028 272206
rect 487554 264302 488028 264330
rect 488368 264316 488396 272342
rect 488552 268122 488580 274654
rect 488736 272814 488764 277766
rect 488724 272808 488776 272814
rect 488724 272750 488776 272756
rect 489368 270768 489420 270774
rect 489368 270710 489420 270716
rect 488540 268116 488592 268122
rect 488540 268058 488592 268064
rect 489184 267844 489236 267850
rect 489184 267786 489236 267792
rect 489196 264316 489224 267786
rect 489380 266898 489408 270710
rect 489932 269634 489960 277766
rect 491496 274514 491524 277780
rect 492232 277766 492614 277794
rect 492232 274718 492260 277766
rect 493796 275874 493824 277780
rect 493784 275868 493836 275874
rect 493784 275810 493836 275816
rect 493968 275868 494020 275874
rect 493968 275810 494020 275816
rect 492496 275188 492548 275194
rect 492496 275130 492548 275136
rect 492220 274712 492272 274718
rect 492220 274654 492272 274660
rect 491484 274508 491536 274514
rect 491484 274450 491536 274456
rect 492312 274508 492364 274514
rect 492312 274450 492364 274456
rect 491208 273828 491260 273834
rect 491208 273770 491260 273776
rect 489886 269606 489960 269634
rect 489886 269550 489914 269606
rect 489874 269544 489926 269550
rect 490012 269544 490064 269550
rect 489874 269486 489926 269492
rect 490010 269512 490012 269521
rect 490064 269512 490066 269521
rect 490010 269447 490066 269456
rect 489368 266892 489420 266898
rect 489368 266834 489420 266840
rect 490288 266348 490340 266354
rect 490288 266290 490340 266296
rect 490300 264330 490328 266290
rect 491220 264330 491248 273770
rect 492324 267734 492352 274450
rect 492508 273086 492536 275130
rect 493980 274802 494008 275810
rect 494992 275602 495020 277780
rect 494980 275596 495032 275602
rect 494980 275538 495032 275544
rect 493796 274774 494008 274802
rect 492496 273080 492548 273086
rect 492496 273022 492548 273028
rect 493600 273080 493652 273086
rect 493600 273022 493652 273028
rect 492048 267706 492352 267734
rect 493324 267708 493376 267714
rect 492048 264330 492076 267706
rect 493324 267650 493376 267656
rect 492496 267028 492548 267034
rect 492496 266970 492548 266976
rect 490038 264302 490328 264330
rect 490866 264302 491248 264330
rect 491694 264302 492076 264330
rect 492508 264316 492536 266970
rect 493336 266490 493364 267650
rect 493324 266484 493376 266490
rect 493324 266426 493376 266432
rect 493612 264330 493640 273022
rect 493796 271046 493824 274774
rect 494060 274712 494112 274718
rect 494060 274654 494112 274660
rect 493784 271040 493836 271046
rect 493784 270982 493836 270988
rect 494072 267918 494100 274654
rect 496188 274242 496216 277780
rect 497384 275874 497412 277780
rect 497372 275868 497424 275874
rect 497372 275810 497424 275816
rect 498200 275868 498252 275874
rect 498200 275810 498252 275816
rect 496820 275596 496872 275602
rect 496820 275538 496872 275544
rect 496360 274508 496412 274514
rect 496360 274450 496412 274456
rect 496636 274508 496688 274514
rect 496636 274450 496688 274456
rect 496372 274242 496400 274450
rect 496176 274236 496228 274242
rect 496176 274178 496228 274184
rect 496360 274236 496412 274242
rect 496360 274178 496412 274184
rect 496268 272808 496320 272814
rect 496268 272750 496320 272756
rect 494532 270558 494928 270586
rect 494242 270328 494298 270337
rect 494242 270263 494298 270272
rect 494060 267912 494112 267918
rect 494060 267854 494112 267860
rect 494256 267734 494284 270263
rect 494532 269550 494560 270558
rect 494900 270502 494928 270558
rect 494704 270496 494756 270502
rect 494704 270438 494756 270444
rect 494888 270496 494940 270502
rect 494888 270438 494940 270444
rect 494716 269550 494744 270438
rect 494520 269544 494572 269550
rect 494520 269486 494572 269492
rect 494704 269544 494756 269550
rect 494704 269486 494756 269492
rect 493350 264302 493640 264330
rect 494164 267706 494284 267734
rect 495624 267708 495676 267714
rect 494164 264316 494192 267706
rect 495624 267650 495676 267656
rect 495808 267708 495860 267714
rect 495808 267650 495860 267656
rect 495636 266898 495664 267650
rect 495440 266892 495492 266898
rect 495440 266834 495492 266840
rect 495624 266892 495676 266898
rect 495624 266834 495676 266840
rect 495452 266286 495480 266834
rect 495440 266280 495492 266286
rect 495440 266222 495492 266228
rect 494980 265804 495032 265810
rect 494980 265746 495032 265752
rect 494992 264316 495020 265746
rect 495820 264316 495848 267650
rect 496280 264330 496308 272750
rect 496452 267980 496504 267986
rect 496452 267922 496504 267928
rect 496464 267442 496492 267922
rect 496648 267714 496676 274450
rect 496832 273222 496860 275538
rect 496820 273216 496872 273222
rect 496820 273158 496872 273164
rect 498212 267986 498240 275810
rect 498580 274718 498608 277780
rect 499592 277766 499790 277794
rect 500512 277766 500894 277794
rect 498752 275732 498804 275738
rect 498752 275674 498804 275680
rect 498764 274786 498792 275674
rect 498752 274780 498804 274786
rect 498752 274722 498804 274728
rect 498568 274712 498620 274718
rect 498568 274654 498620 274660
rect 498752 274644 498804 274650
rect 498752 274586 498804 274592
rect 498764 274242 498792 274586
rect 498752 274236 498804 274242
rect 498752 274178 498804 274184
rect 499592 268938 499620 277766
rect 500512 271862 500540 277766
rect 502076 276010 502104 277780
rect 502352 277766 503286 277794
rect 502064 276004 502116 276010
rect 502064 275946 502116 275952
rect 501972 274236 502024 274242
rect 501972 274178 502024 274184
rect 500960 273216 501012 273222
rect 500960 273158 501012 273164
rect 500500 271856 500552 271862
rect 500500 271798 500552 271804
rect 500684 271856 500736 271862
rect 500684 271798 500736 271804
rect 500696 271046 500724 271798
rect 499948 271040 500000 271046
rect 499948 270982 500000 270988
rect 500684 271040 500736 271046
rect 500684 270982 500736 270988
rect 499580 268932 499632 268938
rect 499580 268874 499632 268880
rect 498200 267980 498252 267986
rect 498200 267922 498252 267928
rect 499120 267980 499172 267986
rect 499120 267922 499172 267928
rect 496636 267708 496688 267714
rect 496636 267650 496688 267656
rect 497464 267708 497516 267714
rect 497464 267650 497516 267656
rect 496452 267436 496504 267442
rect 496452 267378 496504 267384
rect 496820 267436 496872 267442
rect 496820 267378 496872 267384
rect 496832 266762 496860 267378
rect 496820 266756 496872 266762
rect 496820 266698 496872 266704
rect 497004 266756 497056 266762
rect 497004 266698 497056 266704
rect 497016 266422 497044 266698
rect 497004 266416 497056 266422
rect 497004 266358 497056 266364
rect 496280 264302 496662 264330
rect 497476 264316 497504 267650
rect 498568 266212 498620 266218
rect 498568 266154 498620 266160
rect 498580 264330 498608 266154
rect 498318 264302 498608 264330
rect 499132 264316 499160 267922
rect 499960 264316 499988 270982
rect 500776 268116 500828 268122
rect 500776 268058 500828 268064
rect 500224 267028 500276 267034
rect 500224 266970 500276 266976
rect 500236 266490 500264 266970
rect 500224 266484 500276 266490
rect 500224 266426 500276 266432
rect 500788 264316 500816 268058
rect 500972 266218 501000 273158
rect 500960 266212 501012 266218
rect 500960 266154 501012 266160
rect 501984 264330 502012 274178
rect 502352 269074 502380 277766
rect 504468 277394 504496 277780
rect 504468 277366 504588 277394
rect 504180 275868 504232 275874
rect 504180 275810 504232 275816
rect 504192 275466 504220 275810
rect 504180 275460 504232 275466
rect 504180 275402 504232 275408
rect 504364 275460 504416 275466
rect 504364 275402 504416 275408
rect 504376 275194 504404 275402
rect 504364 275188 504416 275194
rect 504364 275130 504416 275136
rect 504560 271590 504588 277366
rect 505664 275738 505692 277780
rect 505652 275732 505704 275738
rect 505652 275674 505704 275680
rect 506860 275194 506888 277780
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 507124 275732 507176 275738
rect 507124 275674 507176 275680
rect 505192 275188 505244 275194
rect 505192 275130 505244 275136
rect 506848 275188 506900 275194
rect 506848 275130 506900 275136
rect 504548 271584 504600 271590
rect 504548 271526 504600 271532
rect 504732 271584 504784 271590
rect 504732 271526 504784 271532
rect 504744 269906 504772 271526
rect 504914 270600 504970 270609
rect 504914 270535 504970 270544
rect 504928 270366 504956 270535
rect 504916 270360 504968 270366
rect 504916 270302 504968 270308
rect 505054 270360 505106 270366
rect 505054 270302 505106 270308
rect 505066 270178 505094 270302
rect 504560 269878 504772 269906
rect 504928 270150 505094 270178
rect 502616 269136 502668 269142
rect 502616 269078 502668 269084
rect 502340 269068 502392 269074
rect 502340 269010 502392 269016
rect 502432 267028 502484 267034
rect 502432 266970 502484 266976
rect 501630 264302 502012 264330
rect 502444 264316 502472 266970
rect 502628 266354 502656 269078
rect 503260 268932 503312 268938
rect 503260 268874 503312 268880
rect 502616 266348 502668 266354
rect 502616 266290 502668 266296
rect 503272 264316 503300 268874
rect 504560 264330 504588 269878
rect 504730 269784 504786 269793
rect 504730 269719 504786 269728
rect 504114 264302 504588 264330
rect 504744 264330 504772 269719
rect 504928 269550 504956 270150
rect 504916 269544 504968 269550
rect 504916 269486 504968 269492
rect 505054 269544 505106 269550
rect 505054 269486 505106 269492
rect 505066 269362 505094 269486
rect 505020 269334 505094 269362
rect 505020 269142 505048 269334
rect 505008 269136 505060 269142
rect 505008 269078 505060 269084
rect 505204 268802 505232 275130
rect 506112 269068 506164 269074
rect 506112 269010 506164 269016
rect 505192 268796 505244 268802
rect 505192 268738 505244 268744
rect 504914 267472 504970 267481
rect 504914 267407 504970 267416
rect 504928 267034 504956 267407
rect 504916 267028 504968 267034
rect 504916 266970 504968 266976
rect 506124 264330 506152 269010
rect 507136 267170 507164 275674
rect 507676 271040 507728 271046
rect 507676 270982 507728 270988
rect 507124 267164 507176 267170
rect 507124 267106 507176 267112
rect 507400 267164 507452 267170
rect 507400 267106 507452 267112
rect 506572 266892 506624 266898
rect 506572 266834 506624 266840
rect 504744 264302 504942 264330
rect 505770 264302 506152 264330
rect 506584 264316 506612 266834
rect 507412 264316 507440 267106
rect 507688 266898 507716 270982
rect 507872 270609 507900 277366
rect 509160 275874 509188 277780
rect 509344 277766 510370 277794
rect 509148 275868 509200 275874
rect 509148 275810 509200 275816
rect 508044 275188 508096 275194
rect 508044 275130 508096 275136
rect 508056 271862 508084 275130
rect 508044 271856 508096 271862
rect 508044 271798 508096 271804
rect 508964 271856 509016 271862
rect 508964 271798 509016 271804
rect 507858 270600 507914 270609
rect 507858 270535 507914 270544
rect 508228 268796 508280 268802
rect 508228 268738 508280 268744
rect 508042 267472 508098 267481
rect 507860 267436 507912 267442
rect 508042 267407 508044 267416
rect 507860 267378 507912 267384
rect 508096 267407 508098 267416
rect 508044 267378 508096 267384
rect 507872 266898 507900 267378
rect 507676 266892 507728 266898
rect 507676 266834 507728 266840
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 508240 264316 508268 268738
rect 508976 264330 509004 271798
rect 509344 268666 509372 277766
rect 510252 276004 510304 276010
rect 510252 275946 510304 275952
rect 509332 268660 509384 268666
rect 509332 268602 509384 268608
rect 509238 267064 509294 267073
rect 509238 266999 509240 267008
rect 509292 266999 509294 267008
rect 509240 266970 509292 266976
rect 510264 264330 510292 275946
rect 511552 271726 511580 277780
rect 512184 275868 512236 275874
rect 512184 275810 512236 275816
rect 511540 271720 511592 271726
rect 511540 271662 511592 271668
rect 511908 271720 511960 271726
rect 511908 271662 511960 271668
rect 510712 268660 510764 268666
rect 510712 268602 510764 268608
rect 508976 264302 509082 264330
rect 509910 264302 510292 264330
rect 510724 264316 510752 268602
rect 511920 267734 511948 271662
rect 512196 267734 512224 275810
rect 512748 275738 512776 277780
rect 512736 275732 512788 275738
rect 512736 275674 512788 275680
rect 512920 275732 512972 275738
rect 512920 275674 512972 275680
rect 512932 275330 512960 275674
rect 512920 275324 512972 275330
rect 512920 275266 512972 275272
rect 513194 274000 513250 274009
rect 513944 273970 513972 277780
rect 514114 274000 514170 274009
rect 513194 273935 513250 273944
rect 513932 273964 513984 273970
rect 512736 268524 512788 268530
rect 512736 268466 512788 268472
rect 512748 268410 512776 268466
rect 512380 268394 512776 268410
rect 512368 268388 512776 268394
rect 512420 268382 512776 268388
rect 512368 268330 512420 268336
rect 511552 267706 511948 267734
rect 512012 267706 512224 267734
rect 511552 264316 511580 267706
rect 511724 267300 511776 267306
rect 512012 267288 512040 267706
rect 511776 267260 512040 267288
rect 511724 267242 511776 267248
rect 512368 267096 512420 267102
rect 512368 267038 512420 267044
rect 512380 264316 512408 267038
rect 513208 264316 513236 273935
rect 514114 273935 514116 273944
rect 513932 273906 513984 273912
rect 514168 273935 514170 273944
rect 514116 273906 514168 273912
rect 515140 271454 515168 277780
rect 516244 275738 516272 277780
rect 516428 277766 517454 277794
rect 518360 277766 518650 277794
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 516428 272678 516456 277766
rect 516784 275732 516836 275738
rect 516784 275674 516836 275680
rect 516416 272672 516468 272678
rect 516416 272614 516468 272620
rect 516600 272672 516652 272678
rect 516600 272614 516652 272620
rect 516612 272490 516640 272614
rect 516060 272462 516640 272490
rect 515128 271448 515180 271454
rect 515128 271390 515180 271396
rect 514300 271312 514352 271318
rect 514298 271280 514300 271289
rect 514484 271312 514536 271318
rect 514352 271280 514354 271289
rect 514484 271254 514536 271260
rect 514298 271215 514354 271224
rect 514024 268796 514076 268802
rect 514024 268738 514076 268744
rect 513838 268424 513894 268433
rect 514036 268394 514064 268738
rect 513838 268359 513840 268368
rect 513892 268359 513894 268368
rect 514024 268388 514076 268394
rect 513840 268330 513892 268336
rect 514024 268330 514076 268336
rect 514496 264330 514524 271254
rect 514944 268660 514996 268666
rect 514944 268602 514996 268608
rect 514956 268433 514984 268602
rect 514942 268424 514998 268433
rect 514942 268359 514998 268368
rect 514666 267336 514722 267345
rect 514666 267271 514722 267280
rect 514680 267102 514708 267271
rect 514668 267096 514720 267102
rect 514668 267038 514720 267044
rect 514852 267096 514904 267102
rect 514852 267038 514904 267044
rect 514050 264302 514524 264330
rect 514864 264316 514892 267038
rect 516060 264330 516088 272462
rect 516796 267734 516824 275674
rect 517520 275460 517572 275466
rect 517520 275402 517572 275408
rect 517336 271448 517388 271454
rect 517336 271390 517388 271396
rect 516336 267706 516824 267734
rect 516336 267102 516364 267706
rect 517348 267102 517376 271390
rect 517532 268666 517560 275402
rect 518360 271289 518388 277766
rect 519832 275874 519860 277780
rect 519820 275868 519872 275874
rect 519820 275810 519872 275816
rect 520188 275732 520240 275738
rect 520188 275674 520240 275680
rect 519726 271688 519782 271697
rect 519726 271623 519782 271632
rect 518346 271280 518402 271289
rect 518346 271215 518402 271224
rect 519740 271182 519768 271623
rect 519728 271176 519780 271182
rect 519728 271118 519780 271124
rect 519912 271176 519964 271182
rect 519912 271118 519964 271124
rect 519924 270994 519952 271118
rect 520200 270994 520228 275674
rect 521028 275466 521056 277780
rect 521856 277766 522238 277794
rect 521016 275460 521068 275466
rect 521016 275402 521068 275408
rect 521200 275460 521252 275466
rect 521200 275402 521252 275408
rect 521212 274786 521240 275402
rect 521200 274780 521252 274786
rect 521200 274722 521252 274728
rect 521660 274780 521712 274786
rect 521660 274722 521712 274728
rect 521106 274000 521162 274009
rect 521106 273935 521162 273944
rect 519648 270966 519952 270994
rect 520016 270966 520228 270994
rect 519648 270910 519676 270966
rect 519636 270904 519688 270910
rect 519636 270846 519688 270852
rect 517520 268660 517572 268666
rect 517520 268602 517572 268608
rect 518440 268660 518492 268666
rect 518440 268602 518492 268608
rect 516324 267096 516376 267102
rect 516324 267038 516376 267044
rect 516508 267096 516560 267102
rect 516508 267038 516560 267044
rect 517336 267096 517388 267102
rect 517520 267096 517572 267102
rect 517336 267038 517388 267044
rect 517518 267064 517520 267073
rect 517572 267064 517574 267073
rect 515706 264302 516088 264330
rect 516520 264316 516548 267038
rect 517518 266999 517574 267008
rect 517334 266792 517390 266801
rect 517334 266727 517390 266736
rect 517348 264316 517376 266727
rect 518452 264330 518480 268602
rect 518898 267608 518954 267617
rect 518898 267543 518954 267552
rect 518912 267458 518940 267543
rect 518728 267430 518940 267458
rect 518728 267102 518756 267430
rect 518990 267336 519046 267345
rect 518990 267271 519046 267280
rect 519176 267300 519228 267306
rect 519004 267170 519032 267271
rect 519176 267242 519228 267248
rect 518992 267164 519044 267170
rect 518992 267106 519044 267112
rect 518716 267096 518768 267102
rect 519188 267073 519216 267242
rect 518716 267038 518768 267044
rect 519174 267064 519230 267073
rect 518992 267028 519044 267034
rect 519174 266999 519230 267008
rect 518992 266970 519044 266976
rect 518716 266960 518768 266966
rect 518716 266902 518768 266908
rect 518728 266801 518756 266902
rect 518714 266792 518770 266801
rect 518714 266727 518770 266736
rect 518190 264302 518480 264330
rect 519004 264316 519032 266970
rect 520016 264330 520044 270966
rect 520188 270904 520240 270910
rect 520188 270846 520240 270852
rect 520200 267034 520228 270846
rect 520188 267028 520240 267034
rect 520188 266970 520240 266976
rect 521120 264330 521148 273935
rect 521474 272504 521530 272513
rect 521474 272439 521530 272448
rect 519846 264302 520044 264330
rect 520674 264302 521148 264330
rect 521488 264316 521516 272439
rect 521672 267617 521700 274722
rect 521856 272950 521884 277766
rect 523420 275466 523448 277780
rect 524524 277394 524552 277780
rect 524432 277366 524552 277394
rect 523408 275460 523460 275466
rect 523408 275402 523460 275408
rect 524432 274394 524460 277366
rect 525522 275768 525578 275777
rect 525522 275703 525524 275712
rect 525576 275703 525578 275712
rect 525524 275674 525576 275680
rect 525524 275324 525576 275330
rect 525524 275266 525576 275272
rect 523512 274366 524460 274394
rect 523512 274106 523540 274366
rect 523868 274236 523920 274242
rect 523868 274178 523920 274184
rect 523500 274100 523552 274106
rect 523500 274042 523552 274048
rect 523880 273970 523908 274178
rect 524050 274000 524106 274009
rect 523868 273964 523920 273970
rect 524050 273935 524052 273944
rect 523868 273906 523920 273912
rect 524104 273935 524106 273944
rect 524052 273906 524104 273912
rect 521844 272944 521896 272950
rect 521844 272886 521896 272892
rect 524328 272672 524380 272678
rect 524328 272614 524380 272620
rect 523498 271416 523554 271425
rect 523498 271351 523554 271360
rect 523512 271182 523540 271351
rect 523868 271312 523920 271318
rect 523868 271254 523920 271260
rect 523500 271176 523552 271182
rect 523500 271118 523552 271124
rect 523880 270910 523908 271254
rect 524142 271144 524198 271153
rect 524142 271079 524198 271088
rect 523868 270904 523920 270910
rect 523868 270846 523920 270852
rect 523684 268524 523736 268530
rect 523684 268466 523736 268472
rect 523498 268288 523554 268297
rect 523696 268258 523724 268466
rect 523498 268223 523500 268232
rect 523552 268223 523554 268232
rect 523684 268252 523736 268258
rect 523500 268194 523552 268200
rect 523684 268194 523736 268200
rect 521658 267608 521714 267617
rect 521658 267543 521714 267552
rect 522670 267336 522726 267345
rect 522670 267271 522726 267280
rect 522684 264330 522712 267271
rect 523132 267028 523184 267034
rect 523132 266970 523184 266976
rect 522330 264302 522712 264330
rect 523144 264316 523172 266970
rect 524156 264330 524184 271079
rect 524340 267034 524368 272614
rect 525340 268524 525392 268530
rect 525340 268466 525392 268472
rect 524328 267028 524380 267034
rect 524328 266970 524380 266976
rect 524788 267028 524840 267034
rect 524788 266970 524840 266976
rect 523986 264302 524184 264330
rect 524800 264316 524828 266970
rect 525352 264330 525380 268466
rect 525536 267034 525564 275266
rect 525720 271425 525748 277780
rect 525892 275732 525944 275738
rect 525892 275674 525944 275680
rect 525904 271697 525932 275674
rect 526916 274786 526944 277780
rect 527560 277766 528126 277794
rect 527272 275732 527324 275738
rect 527272 275674 527324 275680
rect 527284 275330 527312 275674
rect 527088 275324 527140 275330
rect 527088 275266 527140 275272
rect 527272 275324 527324 275330
rect 527272 275266 527324 275272
rect 527100 274786 527128 275266
rect 526904 274780 526956 274786
rect 526904 274722 526956 274728
rect 527088 274780 527140 274786
rect 527088 274722 527140 274728
rect 525890 271688 525946 271697
rect 525890 271623 525946 271632
rect 525706 271416 525762 271425
rect 525706 271351 525762 271360
rect 526812 270904 526864 270910
rect 526812 270846 526864 270852
rect 525524 267028 525576 267034
rect 525524 266970 525576 266976
rect 526824 264330 526852 270846
rect 527178 268560 527234 268569
rect 527178 268495 527180 268504
rect 527232 268495 527234 268504
rect 527364 268524 527416 268530
rect 527180 268466 527232 268472
rect 527364 268466 527416 268472
rect 527376 267734 527404 268466
rect 527560 268297 527588 277766
rect 529308 277394 529336 277780
rect 529216 277366 529336 277394
rect 530136 277766 530518 277794
rect 527730 275768 527786 275777
rect 527730 275703 527732 275712
rect 527784 275703 527786 275712
rect 527732 275674 527784 275680
rect 528512 274408 528568 274417
rect 528512 274343 528514 274352
rect 528566 274343 528568 274352
rect 528652 274372 528704 274378
rect 528514 274314 528566 274320
rect 528652 274314 528704 274320
rect 528664 274258 528692 274314
rect 528526 274230 528692 274258
rect 528098 274136 528154 274145
rect 528526 274106 528554 274230
rect 528650 274136 528706 274145
rect 528098 274071 528154 274080
rect 528514 274100 528566 274106
rect 527914 272912 527970 272921
rect 527914 272847 527970 272856
rect 527928 272678 527956 272847
rect 527916 272672 527968 272678
rect 527916 272614 527968 272620
rect 527546 268288 527602 268297
rect 527546 268223 527602 268232
rect 527376 267706 527496 267734
rect 527272 267028 527324 267034
rect 527272 266970 527324 266976
rect 525352 264302 525642 264330
rect 526470 264302 526852 264330
rect 527284 264316 527312 266970
rect 527468 266801 527496 267706
rect 527454 266792 527510 266801
rect 527454 266727 527510 266736
rect 528112 264316 528140 274071
rect 528650 274071 528652 274080
rect 528514 274042 528566 274048
rect 528704 274071 528706 274080
rect 528652 274042 528704 274048
rect 528514 272944 528566 272950
rect 528652 272944 528704 272950
rect 528514 272886 528566 272892
rect 528650 272912 528652 272921
rect 528704 272912 528706 272921
rect 528526 272762 528554 272886
rect 528650 272847 528706 272856
rect 528526 272734 528784 272762
rect 528376 272672 528428 272678
rect 528376 272614 528428 272620
rect 528388 272513 528416 272614
rect 528560 272536 528612 272542
rect 528374 272504 528430 272513
rect 528374 272439 528430 272448
rect 528558 272504 528560 272513
rect 528756 272524 528784 272734
rect 529020 272536 529072 272542
rect 528612 272504 528614 272513
rect 528756 272496 529020 272524
rect 529020 272478 529072 272484
rect 528558 272439 528614 272448
rect 529216 270230 529244 277366
rect 530136 275466 530164 277766
rect 531608 277394 531636 277780
rect 531608 277366 531728 277394
rect 530124 275460 530176 275466
rect 530124 275402 530176 275408
rect 531320 275460 531372 275466
rect 531320 275402 531372 275408
rect 530766 274952 530822 274961
rect 531332 274922 531360 275402
rect 530766 274887 530822 274896
rect 531320 274916 531372 274922
rect 529846 271416 529902 271425
rect 529846 271351 529902 271360
rect 529204 270224 529256 270230
rect 529204 270166 529256 270172
rect 529664 270224 529716 270230
rect 529664 270166 529716 270172
rect 528926 268560 528982 268569
rect 528926 268495 528928 268504
rect 528980 268495 528982 268504
rect 528928 268466 528980 268472
rect 528558 268288 528614 268297
rect 528526 268258 528558 268274
rect 528514 268252 528558 268258
rect 528566 268223 528614 268232
rect 528514 268194 528566 268200
rect 528558 267608 528614 267617
rect 528558 267543 528614 267552
rect 528572 267458 528600 267543
rect 528526 267430 528600 267458
rect 528526 267306 528554 267430
rect 528650 267336 528706 267345
rect 528514 267300 528566 267306
rect 528650 267271 528652 267280
rect 528514 267242 528566 267248
rect 528704 267271 528706 267280
rect 528652 267242 528704 267248
rect 528466 267064 528522 267073
rect 528466 266999 528468 267008
rect 528520 266999 528522 267008
rect 528742 267064 528798 267073
rect 528742 266999 528744 267008
rect 528468 266970 528520 266976
rect 528796 266999 528798 267008
rect 528744 266970 528796 266976
rect 528742 266656 528798 266665
rect 528742 266591 528744 266600
rect 528796 266591 528798 266600
rect 528928 266620 528980 266626
rect 528744 266562 528796 266568
rect 528928 266562 528980 266568
rect 528940 264316 528968 266562
rect 529676 264330 529704 270166
rect 529860 266626 529888 271351
rect 530780 270230 530808 274887
rect 531320 274858 531372 274864
rect 531504 274916 531556 274922
rect 531504 274858 531556 274864
rect 530768 270224 530820 270230
rect 530768 270166 530820 270172
rect 530952 270224 531004 270230
rect 530952 270166 531004 270172
rect 529848 266620 529900 266626
rect 529848 266562 529900 266568
rect 530964 264330 530992 270166
rect 531320 269952 531372 269958
rect 531320 269894 531372 269900
rect 531332 269793 531360 269894
rect 531318 269784 531374 269793
rect 531318 269719 531374 269728
rect 531516 267578 531544 274858
rect 531700 272513 531728 277366
rect 532804 275330 532832 277780
rect 532792 275324 532844 275330
rect 532792 275266 532844 275272
rect 532976 275324 533028 275330
rect 532976 275266 533028 275272
rect 531686 272504 531742 272513
rect 531686 272439 531742 272448
rect 532988 270178 533016 275266
rect 534000 274922 534028 277780
rect 534736 277766 535210 277794
rect 535656 277766 536406 277794
rect 534170 274952 534226 274961
rect 533988 274916 534040 274922
rect 534170 274887 534172 274896
rect 533988 274858 534040 274864
rect 534224 274887 534226 274896
rect 534172 274858 534224 274864
rect 533710 272232 533766 272241
rect 533710 272167 533766 272176
rect 532804 270150 533016 270178
rect 532804 270065 532832 270150
rect 532790 270056 532846 270065
rect 532790 269991 532846 270000
rect 533066 270056 533122 270065
rect 533066 269991 533122 270000
rect 531688 269952 531740 269958
rect 531688 269894 531740 269900
rect 531504 267572 531556 267578
rect 531504 267514 531556 267520
rect 531700 264330 531728 269894
rect 531870 267608 531926 267617
rect 531870 267543 531872 267552
rect 531924 267543 531926 267552
rect 531872 267514 531924 267520
rect 532240 266620 532292 266626
rect 532240 266562 532292 266568
rect 529676 264302 529782 264330
rect 530610 264302 530992 264330
rect 531438 264302 531728 264330
rect 532252 264316 532280 266562
rect 533080 264316 533108 269991
rect 533724 264330 533752 272167
rect 534736 269793 534764 277766
rect 535274 275360 535330 275369
rect 535274 275295 535276 275304
rect 535328 275295 535330 275304
rect 535460 275324 535512 275330
rect 535276 275266 535328 275272
rect 535460 275266 535512 275272
rect 534722 269784 534778 269793
rect 534722 269719 534778 269728
rect 535472 269634 535500 275266
rect 534736 269606 535500 269634
rect 533724 264302 533922 264330
rect 534736 264316 534764 269606
rect 535656 268297 535684 277766
rect 537588 275466 537616 277780
rect 538784 277394 538812 277780
rect 538692 277366 538812 277394
rect 539612 277766 539902 277794
rect 538220 275596 538272 275602
rect 538220 275538 538272 275544
rect 537576 275460 537628 275466
rect 538232 275448 538260 275538
rect 538232 275420 538536 275448
rect 537576 275402 537628 275408
rect 537944 275324 537996 275330
rect 537944 275266 537996 275272
rect 537956 275210 537984 275266
rect 537220 275182 537984 275210
rect 537220 274922 537248 275182
rect 538218 275088 538274 275097
rect 538048 275058 538218 275074
rect 538036 275052 538218 275058
rect 538088 275046 538218 275052
rect 538218 275023 538274 275032
rect 538036 274994 538088 275000
rect 538508 274922 538536 275420
rect 537208 274916 537260 274922
rect 537208 274858 537260 274864
rect 537392 274916 537444 274922
rect 537392 274858 537444 274864
rect 538496 274916 538548 274922
rect 538496 274858 538548 274864
rect 536102 270600 536158 270609
rect 536102 270535 536158 270544
rect 536116 270230 536144 270535
rect 536104 270224 536156 270230
rect 536104 270166 536156 270172
rect 536288 270224 536340 270230
rect 536288 270166 536340 270172
rect 535642 268288 535698 268297
rect 535642 268223 535698 268232
rect 536300 267734 536328 270166
rect 536024 267706 536328 267734
rect 536024 264330 536052 267706
rect 536378 267064 536434 267073
rect 536378 266999 536434 267008
rect 535578 264302 536052 264330
rect 536392 264316 536420 266999
rect 537404 266665 537432 274858
rect 538218 274680 538274 274689
rect 538218 274615 538274 274624
rect 538232 274530 538260 274615
rect 537956 274502 538260 274530
rect 537956 274417 537984 274502
rect 537942 274408 537998 274417
rect 537942 274343 537998 274352
rect 538128 274372 538180 274378
rect 538128 274314 538180 274320
rect 538312 274372 538364 274378
rect 538312 274314 538364 274320
rect 538140 274145 538168 274314
rect 538324 274145 538352 274314
rect 538126 274136 538182 274145
rect 538126 274071 538182 274080
rect 538310 274136 538366 274145
rect 538310 274071 538366 274080
rect 538218 272776 538274 272785
rect 538218 272711 538274 272720
rect 538232 272626 538260 272711
rect 538140 272598 538260 272626
rect 538140 272542 538168 272598
rect 538128 272536 538180 272542
rect 538128 272478 538180 272484
rect 538312 272536 538364 272542
rect 538312 272478 538364 272484
rect 538324 272241 538352 272478
rect 538310 272232 538366 272241
rect 538310 272167 538366 272176
rect 538034 271416 538090 271425
rect 538034 271351 538090 271360
rect 538048 271266 538076 271351
rect 538048 271238 538214 271266
rect 538186 271182 538214 271238
rect 538036 271176 538088 271182
rect 538036 271118 538088 271124
rect 538174 271176 538226 271182
rect 538174 271118 538226 271124
rect 538048 270722 538076 271118
rect 538048 270694 538214 270722
rect 538186 270638 538214 270694
rect 538036 270632 538088 270638
rect 537850 270600 537906 270609
rect 537850 270535 537906 270544
rect 538034 270600 538036 270609
rect 538174 270632 538226 270638
rect 538088 270600 538090 270609
rect 538174 270574 538226 270580
rect 538034 270535 538090 270544
rect 537864 270314 537892 270535
rect 537864 270286 538214 270314
rect 538186 270230 538214 270286
rect 538036 270224 538088 270230
rect 538036 270166 538088 270172
rect 538174 270224 538226 270230
rect 538174 270166 538226 270172
rect 538048 269958 538076 270166
rect 538692 270094 538720 277366
rect 538862 275360 538918 275369
rect 538862 275295 538864 275304
rect 538916 275295 538918 275304
rect 538864 275266 538916 275272
rect 538862 273864 538918 273873
rect 538862 273799 538918 273808
rect 538680 270088 538732 270094
rect 538680 270030 538732 270036
rect 537852 269952 537904 269958
rect 537852 269894 537904 269900
rect 538036 269952 538088 269958
rect 538036 269894 538088 269900
rect 537864 269521 537892 269894
rect 538034 269784 538090 269793
rect 538034 269719 538090 269728
rect 537850 269512 537906 269521
rect 537850 269447 537906 269456
rect 537574 267608 537630 267617
rect 537574 267543 537630 267552
rect 537390 266656 537446 266665
rect 537390 266591 537446 266600
rect 537588 264330 537616 267543
rect 537234 264302 537616 264330
rect 538048 264316 538076 269719
rect 538402 269512 538458 269521
rect 538458 269470 538628 269498
rect 538402 269447 538458 269456
rect 538600 269414 538628 269470
rect 538588 269408 538640 269414
rect 538588 269350 538640 269356
rect 538220 269272 538272 269278
rect 538220 269214 538272 269220
rect 538232 269113 538260 269214
rect 538218 269104 538274 269113
rect 538218 269039 538274 269048
rect 538310 267608 538366 267617
rect 538174 267572 538226 267578
rect 538310 267543 538312 267552
rect 538174 267514 538226 267520
rect 538364 267543 538366 267552
rect 538312 267514 538364 267520
rect 538186 267458 538214 267514
rect 538186 267430 538260 267458
rect 538232 267345 538260 267430
rect 538218 267336 538274 267345
rect 538218 267271 538274 267280
rect 538876 267073 538904 273799
rect 539612 270609 539640 277766
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 541452 277766 542294 277794
rect 543200 277766 543490 277794
rect 544212 277766 544686 277794
rect 540992 275058 541020 277366
rect 540980 275052 541032 275058
rect 540980 274994 541032 275000
rect 540702 272504 540758 272513
rect 540702 272439 540758 272448
rect 539598 270600 539654 270609
rect 539598 270535 539654 270544
rect 539230 268016 539286 268025
rect 539230 267951 539286 267960
rect 538862 267064 538918 267073
rect 538862 266999 538918 267008
rect 539244 264330 539272 267951
rect 539690 267608 539746 267617
rect 539690 267543 539746 267552
rect 538890 264302 539272 264330
rect 539704 264316 539732 267543
rect 540428 267028 540480 267034
rect 540428 266970 540480 266976
rect 540242 266792 540298 266801
rect 540242 266727 540298 266736
rect 540256 266626 540284 266727
rect 540440 266626 540468 266970
rect 540244 266620 540296 266626
rect 540244 266562 540296 266568
rect 540428 266620 540480 266626
rect 540428 266562 540480 266568
rect 540716 264330 540744 272439
rect 541452 269822 541480 277766
rect 543004 275596 543056 275602
rect 543004 275538 543056 275544
rect 543016 275058 543044 275538
rect 543004 275052 543056 275058
rect 543004 274994 543056 275000
rect 543200 274689 543228 277766
rect 544212 275097 544240 277766
rect 545120 275596 545172 275602
rect 545120 275538 545172 275544
rect 544198 275088 544254 275097
rect 544198 275023 544254 275032
rect 544382 274952 544438 274961
rect 544382 274887 544438 274896
rect 543186 274680 543242 274689
rect 543186 274615 543242 274624
rect 543188 270360 543240 270366
rect 543188 270302 543240 270308
rect 543372 270360 543424 270366
rect 543372 270302 543424 270308
rect 543200 269958 543228 270302
rect 543188 269952 543240 269958
rect 543188 269894 543240 269900
rect 541440 269816 541492 269822
rect 541440 269758 541492 269764
rect 543004 269816 543056 269822
rect 543004 269758 543056 269764
rect 541438 269376 541494 269385
rect 541438 269311 541494 269320
rect 541452 269210 541480 269311
rect 541624 269272 541676 269278
rect 541624 269214 541676 269220
rect 541440 269204 541492 269210
rect 541440 269146 541492 269152
rect 540888 267028 540940 267034
rect 540888 266970 540940 266976
rect 540900 266801 540928 266970
rect 540886 266792 540942 266801
rect 540886 266727 540942 266736
rect 541636 264330 541664 269214
rect 542174 267064 542230 267073
rect 542174 266999 542230 267008
rect 540546 264302 540744 264330
rect 541374 264302 541664 264330
rect 542188 264316 542216 266999
rect 543016 264316 543044 269758
rect 543384 269414 543412 270302
rect 543372 269408 543424 269414
rect 543556 269408 543608 269414
rect 543372 269350 543424 269356
rect 543554 269376 543556 269385
rect 543608 269376 543610 269385
rect 543554 269311 543610 269320
rect 544396 269113 544424 274887
rect 545132 272785 545160 275538
rect 545868 274922 545896 277780
rect 546512 277766 547078 277794
rect 547892 277766 548182 277794
rect 546038 274952 546094 274961
rect 545856 274916 545908 274922
rect 546038 274887 546040 274896
rect 545856 274858 545908 274864
rect 546092 274887 546094 274896
rect 546040 274858 546092 274864
rect 545118 272776 545174 272785
rect 545118 272711 545174 272720
rect 546512 269550 546540 277766
rect 545856 269544 545908 269550
rect 545316 269504 545856 269532
rect 545316 269414 545344 269504
rect 545856 269486 545908 269492
rect 546500 269544 546552 269550
rect 546500 269486 546552 269492
rect 545304 269408 545356 269414
rect 545856 269408 545908 269414
rect 545304 269350 545356 269356
rect 545500 269368 545856 269396
rect 545500 269278 545528 269368
rect 545856 269350 545908 269356
rect 545488 269272 545540 269278
rect 545488 269214 545540 269220
rect 544382 269104 544438 269113
rect 544382 269039 544438 269048
rect 543692 268424 543748 268433
rect 543692 268359 543694 268368
rect 543746 268359 543748 268368
rect 543832 268388 543884 268394
rect 543694 268330 543746 268336
rect 543832 268330 543884 268336
rect 543844 268025 543872 268330
rect 543830 268016 543886 268025
rect 543830 267951 543886 267960
rect 544014 267880 544070 267889
rect 543706 267838 544014 267866
rect 543706 267714 543734 267838
rect 544014 267815 544070 267824
rect 543694 267708 543746 267714
rect 543694 267650 543746 267656
rect 543832 267708 543884 267714
rect 543832 267650 543884 267656
rect 543844 267345 543872 267650
rect 543830 267336 543886 267345
rect 543830 267271 543886 267280
rect 547892 266082 547920 277766
rect 549364 277394 549392 277780
rect 549272 277366 549392 277394
rect 549272 273254 549300 277366
rect 550560 274922 550588 277780
rect 550548 274916 550600 274922
rect 550548 274858 550600 274864
rect 549272 273226 549484 273254
rect 548708 269952 548760 269958
rect 548708 269894 548760 269900
rect 548892 269952 548944 269958
rect 548892 269894 548944 269900
rect 548720 269686 548748 269894
rect 548708 269680 548760 269686
rect 548708 269622 548760 269628
rect 548904 269414 548932 269894
rect 548892 269408 548944 269414
rect 548892 269350 548944 269356
rect 549260 269408 549312 269414
rect 549260 269350 549312 269356
rect 548800 268388 548852 268394
rect 548800 268330 548852 268336
rect 548812 268274 548840 268330
rect 548444 268258 548840 268274
rect 548432 268252 548840 268258
rect 548484 268246 548840 268252
rect 548432 268194 548484 268200
rect 549272 266762 549300 269350
rect 549456 268433 549484 273226
rect 551756 270774 551784 277780
rect 552492 277766 552966 277794
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552492 271998 552520 277766
rect 552664 275596 552716 275602
rect 552664 275538 552716 275544
rect 552848 275596 552900 275602
rect 552848 275538 552900 275544
rect 552676 275058 552704 275538
rect 552664 275052 552716 275058
rect 552664 274994 552716 275000
rect 552860 274922 552888 275538
rect 552848 274916 552900 274922
rect 552848 274858 552900 274864
rect 552480 271992 552532 271998
rect 552480 271934 552532 271940
rect 552664 271992 552716 271998
rect 552664 271934 552716 271940
rect 551744 270768 551796 270774
rect 551744 270710 551796 270716
rect 549442 268424 549498 268433
rect 549442 268359 549498 268368
rect 552676 267889 552704 271934
rect 553412 269550 553440 277766
rect 553400 269544 553452 269550
rect 553400 269486 553452 269492
rect 552662 267880 552718 267889
rect 552662 267815 552718 267824
rect 549260 266756 549312 266762
rect 549260 266698 549312 266704
rect 547880 266076 547932 266082
rect 547880 266018 547932 266024
rect 554792 265674 554820 277766
rect 556448 273426 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 273420 556488 273426
rect 556436 273362 556488 273368
rect 557552 269278 557580 277366
rect 558840 273562 558868 277780
rect 558828 273556 558880 273562
rect 558828 273498 558880 273504
rect 560036 272134 560064 277780
rect 560864 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 272128 560076 272134
rect 560024 272070 560076 272076
rect 560864 270502 560892 277766
rect 560852 270496 560904 270502
rect 560852 270438 560904 270444
rect 558920 269544 558972 269550
rect 558920 269486 558972 269492
rect 557540 269272 557592 269278
rect 557540 269214 557592 269220
rect 558932 266490 558960 269486
rect 558920 266484 558972 266490
rect 558920 266426 558972 266432
rect 561692 265946 561720 277766
rect 563532 273698 563560 277780
rect 564452 277766 564742 277794
rect 563520 273692 563572 273698
rect 563520 273634 563572 273640
rect 564452 269686 564480 277766
rect 565924 272270 565952 277780
rect 567120 272406 567148 277780
rect 567672 277766 568330 277794
rect 568592 277766 569526 277794
rect 567108 272400 567160 272406
rect 567108 272342 567160 272348
rect 565912 272264 565964 272270
rect 565912 272206 565964 272212
rect 564440 269680 564492 269686
rect 564440 269622 564492 269628
rect 567672 267850 567700 277766
rect 568592 269414 568620 277766
rect 570708 273834 570736 277780
rect 571812 274650 571840 277780
rect 572732 277766 573022 277794
rect 571800 274644 571852 274650
rect 571800 274586 571852 274592
rect 570696 273828 570748 273834
rect 570696 273770 570748 273776
rect 570604 273692 570656 273698
rect 570604 273634 570656 273640
rect 568580 269408 568632 269414
rect 568580 269350 568632 269356
rect 567660 267844 567712 267850
rect 567660 267786 567712 267792
rect 570616 267442 570644 273634
rect 572732 269550 572760 277766
rect 574204 273086 574232 277780
rect 574940 277766 575414 277794
rect 575860 277766 576610 277794
rect 574192 273080 574244 273086
rect 574192 273022 574244 273028
rect 574940 270337 574968 277766
rect 574926 270328 574982 270337
rect 574926 270263 574982 270272
rect 572720 269544 572772 269550
rect 572720 269486 572772 269492
rect 571984 267708 572036 267714
rect 571984 267650 572036 267656
rect 571996 267442 572024 267650
rect 570604 267436 570656 267442
rect 570604 267378 570656 267384
rect 571984 267436 572036 267442
rect 571984 267378 572036 267384
rect 572168 266892 572220 266898
rect 572168 266834 572220 266840
rect 572180 266626 572208 266834
rect 572168 266620 572220 266626
rect 572168 266562 572220 266568
rect 561680 265940 561732 265946
rect 561680 265882 561732 265888
rect 575860 265810 575888 277766
rect 577228 275460 577280 275466
rect 577228 275402 577280 275408
rect 577240 275194 577268 275402
rect 577044 275188 577096 275194
rect 577044 275130 577096 275136
rect 577228 275188 577280 275194
rect 577228 275130 577280 275136
rect 577056 274922 577084 275130
rect 577044 274916 577096 274922
rect 577044 274858 577096 274864
rect 577792 274514 577820 277780
rect 578896 275058 578924 277780
rect 578884 275052 578936 275058
rect 578884 274994 578936 275000
rect 577780 274508 577832 274514
rect 577780 274450 577832 274456
rect 578884 272400 578936 272406
rect 578884 272342 578936 272348
rect 578896 266762 578924 272342
rect 580092 271998 580120 277780
rect 581288 273222 581316 277780
rect 582484 277394 582512 277780
rect 582392 277366 582512 277394
rect 581276 273216 581328 273222
rect 581276 273158 581328 273164
rect 580264 273080 580316 273086
rect 580264 273022 580316 273028
rect 580080 271992 580132 271998
rect 580080 271934 580132 271940
rect 580276 267345 580304 273022
rect 582392 267986 582420 277366
rect 583680 274922 583708 277780
rect 583864 277766 584890 277794
rect 583668 274916 583720 274922
rect 583668 274858 583720 274864
rect 583864 268122 583892 277766
rect 585784 274508 585836 274514
rect 585784 274450 585836 274456
rect 583852 268116 583904 268122
rect 583852 268058 583904 268064
rect 582380 267980 582432 267986
rect 582380 267922 582432 267928
rect 585796 267714 585824 274450
rect 586072 274378 586100 277780
rect 586060 274372 586112 274378
rect 586060 274314 586112 274320
rect 587176 273834 587204 277780
rect 587912 277766 588386 277794
rect 589384 277766 589582 277794
rect 587164 273828 587216 273834
rect 587164 273770 587216 273776
rect 587912 268938 587940 277766
rect 589384 271590 589412 277766
rect 590764 275330 590792 277780
rect 591040 277766 591974 277794
rect 590752 275324 590804 275330
rect 590752 275266 590804 275272
rect 589372 271584 589424 271590
rect 589372 271526 589424 271532
rect 591040 269074 591068 277766
rect 591304 271584 591356 271590
rect 591304 271526 591356 271532
rect 591316 270774 591344 271526
rect 593156 271046 593184 277780
rect 594352 272406 594380 277780
rect 594812 277766 595470 277794
rect 594340 272400 594392 272406
rect 594340 272342 594392 272348
rect 593144 271040 593196 271046
rect 593144 270982 593196 270988
rect 591304 270768 591356 270774
rect 591304 270710 591356 270716
rect 591028 269068 591080 269074
rect 591028 269010 591080 269016
rect 587900 268932 587952 268938
rect 587900 268874 587952 268880
rect 594812 268394 594840 277766
rect 596652 271862 596680 277780
rect 597848 276010 597876 277780
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597836 276004 597888 276010
rect 597836 275946 597888 275952
rect 598952 274666 598980 277366
rect 599124 275460 599176 275466
rect 599124 275402 599176 275408
rect 599136 275194 599164 275402
rect 599124 275188 599176 275194
rect 599124 275130 599176 275136
rect 598860 274638 598980 274666
rect 596640 271856 596692 271862
rect 596640 271798 596692 271804
rect 598860 268802 598888 274638
rect 600240 271726 600268 277780
rect 601436 274378 601464 277780
rect 602172 277766 602554 277794
rect 601424 274372 601476 274378
rect 601424 274314 601476 274320
rect 602172 274242 602200 277766
rect 602160 274236 602212 274242
rect 602160 274178 602212 274184
rect 602344 274236 602396 274242
rect 602344 274178 602396 274184
rect 600228 271720 600280 271726
rect 600228 271662 600280 271668
rect 598848 268796 598900 268802
rect 598848 268738 598900 268744
rect 594800 268388 594852 268394
rect 594800 268330 594852 268336
rect 581276 267708 581328 267714
rect 581276 267650 581328 267656
rect 585784 267708 585836 267714
rect 585784 267650 585836 267656
rect 580262 267336 580318 267345
rect 580262 267271 580318 267280
rect 581288 267170 581316 267650
rect 602356 267442 602384 274178
rect 603736 271590 603764 277780
rect 604932 275874 604960 277780
rect 604920 275868 604972 275874
rect 604920 275810 604972 275816
rect 604460 274916 604512 274922
rect 604460 274858 604512 274864
rect 603724 271584 603776 271590
rect 603724 271526 603776 271532
rect 604472 271454 604500 274858
rect 606128 272814 606156 277780
rect 607324 274922 607352 277780
rect 607312 274916 607364 274922
rect 607312 274858 607364 274864
rect 608520 274242 608548 277780
rect 608704 277766 609730 277794
rect 608508 274236 608560 274242
rect 608508 274178 608560 274184
rect 606116 272808 606168 272814
rect 606116 272750 606168 272756
rect 607864 271584 607916 271590
rect 607864 271526 607916 271532
rect 604460 271448 604512 271454
rect 604460 271390 604512 271396
rect 602344 267436 602396 267442
rect 602344 267378 602396 267384
rect 581276 267164 581328 267170
rect 581276 267106 581328 267112
rect 581644 267164 581696 267170
rect 581644 267106 581696 267112
rect 581656 266898 581684 267106
rect 607876 267073 607904 271526
rect 608704 268666 608732 277766
rect 610820 271318 610848 277780
rect 612016 275738 612044 277780
rect 612004 275732 612056 275738
rect 612004 275674 612056 275680
rect 611360 275460 611412 275466
rect 611360 275402 611412 275408
rect 611372 272950 611400 275402
rect 613212 273970 613240 277780
rect 613200 273964 613252 273970
rect 613200 273906 613252 273912
rect 613384 273760 613436 273766
rect 613384 273702 613436 273708
rect 611360 272944 611412 272950
rect 611360 272886 611412 272892
rect 610808 271312 610860 271318
rect 610808 271254 610860 271260
rect 608692 268660 608744 268666
rect 608692 268602 608744 268608
rect 613396 267306 613424 273702
rect 614408 272678 614436 277780
rect 615604 273766 615632 277780
rect 616800 275466 616828 277780
rect 616788 275460 616840 275466
rect 616788 275402 616840 275408
rect 615592 273760 615644 273766
rect 615592 273702 615644 273708
rect 614396 272672 614448 272678
rect 614396 272614 614448 272620
rect 617996 271153 618024 277780
rect 619100 274786 619128 277780
rect 619744 277766 620310 277794
rect 619088 274780 619140 274786
rect 619088 274722 619140 274728
rect 619548 274712 619600 274718
rect 619548 274654 619600 274660
rect 619560 274106 619588 274654
rect 619548 274100 619600 274106
rect 619548 274042 619600 274048
rect 617982 271144 618038 271153
rect 617982 271079 618038 271088
rect 619744 268530 619772 277766
rect 621492 270910 621520 277780
rect 622412 277766 622702 277794
rect 621664 271312 621716 271318
rect 621664 271254 621716 271260
rect 621480 270904 621532 270910
rect 621480 270846 621532 270852
rect 619732 268524 619784 268530
rect 619732 268466 619784 268472
rect 621676 267578 621704 271254
rect 621664 267572 621716 267578
rect 621664 267514 621716 267520
rect 613384 267300 613436 267306
rect 613384 267242 613436 267248
rect 622412 267170 622440 277766
rect 623884 274718 623912 277780
rect 623872 274712 623924 274718
rect 623872 274654 623924 274660
rect 625080 271182 625108 277780
rect 626184 275466 626212 277780
rect 626644 277766 627394 277794
rect 627932 277766 628590 277794
rect 629312 277766 629786 277794
rect 630692 277766 630982 277794
rect 626172 275460 626224 275466
rect 626172 275402 626224 275408
rect 626448 275460 626500 275466
rect 626448 275402 626500 275408
rect 626460 272513 626488 275402
rect 626446 272504 626502 272513
rect 626446 272439 626502 272448
rect 625068 271176 625120 271182
rect 625068 271118 625120 271124
rect 626644 270230 626672 277766
rect 627932 270366 627960 277766
rect 627920 270360 627972 270366
rect 627920 270302 627972 270308
rect 626632 270224 626684 270230
rect 626632 270166 626684 270172
rect 622400 267164 622452 267170
rect 622400 267106 622452 267112
rect 607862 267064 607918 267073
rect 629312 267034 629340 277766
rect 630692 270065 630720 277766
rect 632164 272542 632192 277780
rect 633360 275194 633388 277780
rect 633636 277766 634478 277794
rect 633348 275188 633400 275194
rect 633348 275130 633400 275136
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 633636 270094 633664 277766
rect 635660 273873 635688 277780
rect 635646 273864 635702 273873
rect 635646 273799 635702 273808
rect 636856 271318 636884 277780
rect 637592 277766 638066 277794
rect 638972 277766 639262 277794
rect 636844 271312 636896 271318
rect 636844 271254 636896 271260
rect 633624 270088 633676 270094
rect 630678 270056 630734 270065
rect 633624 270030 633676 270036
rect 630678 269991 630734 270000
rect 637592 269793 637620 277766
rect 637578 269784 637634 269793
rect 637578 269719 637634 269728
rect 638972 268258 639000 277766
rect 640444 273086 640472 277780
rect 641640 275466 641668 277780
rect 641916 277766 642758 277794
rect 641628 275460 641680 275466
rect 641628 275402 641680 275408
rect 640432 273080 640484 273086
rect 640432 273022 640484 273028
rect 641916 269958 641944 277766
rect 643940 271590 643968 277780
rect 644492 277766 645150 277794
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 643928 271584 643980 271590
rect 643928 271526 643980 271532
rect 641904 269952 641956 269958
rect 641904 269894 641956 269900
rect 644492 269822 644520 277766
rect 644480 269816 644532 269822
rect 644480 269758 644532 269764
rect 638960 268252 639012 268258
rect 638960 268194 639012 268200
rect 607862 266999 607918 267008
rect 629300 267028 629352 267034
rect 629300 266970 629352 266976
rect 581644 266892 581696 266898
rect 581644 266834 581696 266840
rect 578884 266756 578936 266762
rect 578884 266698 578936 266704
rect 575848 265804 575900 265810
rect 575848 265746 575900 265752
rect 554780 265668 554832 265674
rect 554780 265610 554832 265616
rect 558184 265668 558236 265674
rect 558184 265610 558236 265616
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553490 255640 553546 255649
rect 553490 255575 553492 255584
rect 553544 255575 553546 255584
rect 555424 255604 555476 255610
rect 553492 255546 553544 255552
rect 555424 255546 555476 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 554136 251194 554188 251200
rect 553858 249112 553914 249121
rect 553858 249047 553914 249056
rect 553872 246362 553900 249047
rect 554410 246936 554466 246945
rect 554410 246871 554466 246880
rect 553860 246356 553912 246362
rect 553860 246298 553912 246304
rect 554424 245682 554452 246871
rect 554412 245676 554464 245682
rect 554412 245618 554464 245624
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 553950 242584 554006 242593
rect 553950 242519 554006 242528
rect 553964 241534 553992 242519
rect 553952 241528 554004 241534
rect 553952 241470 554004 241476
rect 553858 240408 553914 240417
rect 553858 240343 553914 240352
rect 553872 240174 553900 240343
rect 553860 240168 553912 240174
rect 553860 240110 553912 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 140792 231662 141174 231690
rect 141528 231662 141818 231690
rect 90364 230444 90416 230450
rect 90364 230386 90416 230392
rect 88248 230036 88300 230042
rect 88248 229978 88300 229984
rect 74448 229900 74500 229906
rect 74448 229842 74500 229848
rect 67548 229764 67600 229770
rect 67548 229706 67600 229712
rect 65984 228404 66036 228410
rect 65984 228346 66036 228352
rect 64788 225752 64840 225758
rect 64788 225694 64840 225700
rect 62946 222864 63002 222873
rect 62946 222799 63002 222808
rect 64604 221468 64656 221474
rect 64604 221410 64656 221416
rect 63408 220108 63460 220114
rect 63408 220050 63460 220056
rect 62764 218204 62816 218210
rect 62764 218146 62816 218152
rect 63420 217002 63448 220050
rect 64236 218068 64288 218074
rect 64236 218010 64288 218016
rect 64248 217002 64276 218010
rect 56336 216974 56488 217002
rect 57316 216974 57744 217002
rect 58144 216974 58480 217002
rect 58972 216974 59308 217002
rect 59800 216974 60136 217002
rect 60628 216974 60688 217002
rect 61456 216974 61792 217002
rect 62284 216974 62620 217002
rect 63112 216974 63448 217002
rect 63940 216974 64276 217002
rect 64616 217002 64644 221410
rect 64800 218074 64828 225694
rect 64788 218068 64840 218074
rect 64788 218010 64840 218016
rect 65996 217002 66024 228346
rect 66720 220244 66772 220250
rect 66720 220186 66772 220192
rect 66732 217002 66760 220186
rect 67560 217002 67588 229706
rect 73066 226944 73122 226953
rect 73066 226879 73122 226888
rect 69664 226160 69716 226166
rect 69664 226102 69716 226108
rect 68926 224224 68982 224233
rect 68926 224159 68982 224168
rect 68376 221740 68428 221746
rect 68376 221682 68428 221688
rect 68388 217002 68416 221682
rect 68940 217002 68968 224159
rect 69676 218754 69704 226102
rect 71688 221876 71740 221882
rect 71688 221818 71740 221824
rect 70030 220144 70086 220153
rect 70030 220079 70086 220088
rect 69664 218748 69716 218754
rect 69664 218690 69716 218696
rect 70044 217002 70072 220079
rect 70860 219020 70912 219026
rect 70860 218962 70912 218968
rect 70872 217002 70900 218962
rect 71700 217002 71728 221818
rect 72882 220416 72938 220425
rect 72882 220351 72938 220360
rect 72516 218068 72568 218074
rect 72516 218010 72568 218016
rect 72528 217002 72556 218010
rect 64616 216974 64768 217002
rect 65596 216974 66024 217002
rect 66424 216974 66760 217002
rect 67252 216974 67588 217002
rect 68080 216974 68416 217002
rect 68908 216974 68968 217002
rect 69736 216974 70072 217002
rect 70564 216974 70900 217002
rect 71392 216974 71728 217002
rect 72220 216974 72556 217002
rect 72896 217002 72924 220351
rect 73080 218074 73108 226879
rect 74460 219434 74488 229842
rect 82084 228676 82136 228682
rect 82084 228618 82136 228624
rect 79966 228304 80022 228313
rect 79966 228239 80022 228248
rect 75828 227180 75880 227186
rect 75828 227122 75880 227128
rect 74276 219406 74488 219434
rect 73068 218068 73120 218074
rect 73068 218010 73120 218016
rect 74276 217002 74304 219406
rect 75644 218340 75696 218346
rect 75644 218282 75696 218288
rect 75000 218068 75052 218074
rect 75000 218010 75052 218016
rect 75012 217002 75040 218010
rect 75656 217002 75684 218282
rect 75840 218074 75868 227122
rect 76472 223984 76524 223990
rect 76472 223926 76524 223932
rect 76484 218890 76512 223926
rect 78404 223168 78456 223174
rect 78404 223110 78456 223116
rect 76656 220380 76708 220386
rect 76656 220322 76708 220328
rect 76472 218884 76524 218890
rect 76472 218826 76524 218832
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76668 217002 76696 220322
rect 77208 218748 77260 218754
rect 77208 218690 77260 218696
rect 77220 217002 77248 218690
rect 78416 217002 78444 223110
rect 79784 218204 79836 218210
rect 79784 218146 79836 218152
rect 79140 218068 79192 218074
rect 79140 218010 79192 218016
rect 79152 217002 79180 218010
rect 79796 217002 79824 218146
rect 79980 218074 80008 228239
rect 81348 223440 81400 223446
rect 81348 223382 81400 223388
rect 80796 219428 80848 219434
rect 80796 219370 80848 219376
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80808 217002 80836 219370
rect 81360 217002 81388 223382
rect 82096 218210 82124 228618
rect 86684 227316 86736 227322
rect 86684 227258 86736 227264
rect 83464 226296 83516 226302
rect 83464 226238 83516 226244
rect 82544 224392 82596 224398
rect 82544 224334 82596 224340
rect 82084 218204 82136 218210
rect 82084 218146 82136 218152
rect 82556 217002 82584 224334
rect 83280 220516 83332 220522
rect 83280 220458 83332 220464
rect 83292 217002 83320 220458
rect 83476 218346 83504 226238
rect 85488 222760 85540 222766
rect 85488 222702 85540 222708
rect 85304 219156 85356 219162
rect 85304 219098 85356 219104
rect 83924 218884 83976 218890
rect 83924 218826 83976 218832
rect 83464 218340 83516 218346
rect 83464 218282 83516 218288
rect 83936 217002 83964 218826
rect 84936 218068 84988 218074
rect 84936 218010 84988 218016
rect 84948 217002 84976 218010
rect 72896 216974 73048 217002
rect 73876 216974 74304 217002
rect 74704 216974 75040 217002
rect 75532 216974 75684 217002
rect 76360 216974 76696 217002
rect 77188 216974 77248 217002
rect 78016 216974 78444 217002
rect 78844 216974 79180 217002
rect 79672 216974 79824 217002
rect 80500 216974 80836 217002
rect 81328 216974 81388 217002
rect 82156 216974 82584 217002
rect 82984 216974 83320 217002
rect 83812 216974 83964 217002
rect 84640 216974 84976 217002
rect 85316 217002 85344 219098
rect 85500 218074 85528 222702
rect 85488 218068 85540 218074
rect 85488 218010 85540 218016
rect 86696 217002 86724 227258
rect 88064 223576 88116 223582
rect 88064 223518 88116 223524
rect 87420 218068 87472 218074
rect 87420 218010 87472 218016
rect 87432 217002 87460 218010
rect 88076 217002 88104 223518
rect 88260 218074 88288 229978
rect 89628 227452 89680 227458
rect 89628 227394 89680 227400
rect 89168 222624 89220 222630
rect 89168 222566 89220 222572
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 89180 217002 89208 222566
rect 89640 217002 89668 227394
rect 90376 219434 90404 230386
rect 118424 230308 118476 230314
rect 118424 230250 118476 230256
rect 111064 230172 111116 230178
rect 111064 230114 111116 230120
rect 103610 229800 103666 229809
rect 103610 229735 103666 229744
rect 92480 229220 92532 229226
rect 92480 229162 92532 229168
rect 92492 225758 92520 229162
rect 102048 229084 102100 229090
rect 102048 229026 102100 229032
rect 97908 228948 97960 228954
rect 97908 228890 97960 228896
rect 96528 228676 96580 228682
rect 96528 228618 96580 228624
rect 93768 226024 93820 226030
rect 93768 225966 93820 225972
rect 92480 225752 92532 225758
rect 92480 225694 92532 225700
rect 92388 223032 92440 223038
rect 92388 222974 92440 222980
rect 91560 220652 91612 220658
rect 91560 220594 91612 220600
rect 90364 219428 90416 219434
rect 90364 219370 90416 219376
rect 90732 219428 90784 219434
rect 90732 219370 90784 219376
rect 90744 217002 90772 219370
rect 91572 217002 91600 220594
rect 92400 217002 92428 222974
rect 93780 219298 93808 225966
rect 94964 225888 95016 225894
rect 94964 225830 95016 225836
rect 93216 219292 93268 219298
rect 93216 219234 93268 219240
rect 93768 219292 93820 219298
rect 93768 219234 93820 219240
rect 93228 217002 93256 219234
rect 93768 218612 93820 218618
rect 93768 218554 93820 218560
rect 93780 217002 93808 218554
rect 94976 217002 95004 225830
rect 95700 222012 95752 222018
rect 95700 221954 95752 221960
rect 95712 217002 95740 221954
rect 96540 217002 96568 228618
rect 96712 223304 96764 223310
rect 96712 223246 96764 223252
rect 96724 223038 96752 223246
rect 96712 223032 96764 223038
rect 96712 222974 96764 222980
rect 97724 220788 97776 220794
rect 97724 220730 97776 220736
rect 97356 218068 97408 218074
rect 97356 218010 97408 218016
rect 97368 217002 97396 218010
rect 85316 216974 85468 217002
rect 86296 216974 86724 217002
rect 87124 216974 87460 217002
rect 87952 216974 88104 217002
rect 88780 216974 89208 217002
rect 89608 216974 89668 217002
rect 90436 216974 90772 217002
rect 91264 216974 91600 217002
rect 92092 216974 92428 217002
rect 92920 216974 93256 217002
rect 93748 216974 93808 217002
rect 94576 216974 95004 217002
rect 95404 216974 95740 217002
rect 96232 216974 96568 217002
rect 97060 216974 97396 217002
rect 97736 217002 97764 220730
rect 97920 218074 97948 228890
rect 100668 227588 100720 227594
rect 100668 227530 100720 227536
rect 98644 223032 98696 223038
rect 98644 222974 98696 222980
rect 98656 222630 98684 222974
rect 98644 222624 98696 222630
rect 98644 222566 98696 222572
rect 99104 222624 99156 222630
rect 99104 222566 99156 222572
rect 97908 218068 97960 218074
rect 97908 218010 97960 218016
rect 99116 217002 99144 222566
rect 100484 218476 100536 218482
rect 100484 218418 100536 218424
rect 99840 218068 99892 218074
rect 99840 218010 99892 218016
rect 99852 217002 99880 218010
rect 100496 217002 100524 218418
rect 100680 218074 100708 227530
rect 101862 221504 101918 221513
rect 101862 221439 101918 221448
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101496 218068 101548 218074
rect 101496 218010 101548 218016
rect 101508 217002 101536 218010
rect 97736 216974 97888 217002
rect 98716 216974 99144 217002
rect 99544 216974 99880 217002
rect 100372 216974 100524 217002
rect 101200 216974 101536 217002
rect 101876 217002 101904 221439
rect 102060 218074 102088 229026
rect 103244 225480 103296 225486
rect 103244 225422 103296 225428
rect 102048 218068 102100 218074
rect 102048 218010 102100 218016
rect 103256 217002 103284 225422
rect 103624 224534 103652 229735
rect 108488 228948 108540 228954
rect 108488 228890 108540 228896
rect 108120 228812 108172 228818
rect 108120 228754 108172 228760
rect 108132 228274 108160 228754
rect 108120 228268 108172 228274
rect 108120 228210 108172 228216
rect 108500 228138 108528 228890
rect 106188 228132 106240 228138
rect 106188 228074 106240 228080
rect 108488 228132 108540 228138
rect 108488 228074 108540 228080
rect 105728 225344 105780 225350
rect 105728 225286 105780 225292
rect 103612 224528 103664 224534
rect 103612 224470 103664 224476
rect 104808 224120 104860 224126
rect 104808 224062 104860 224068
rect 104624 222012 104676 222018
rect 104624 221954 104676 221960
rect 103980 218068 104032 218074
rect 103980 218010 104032 218016
rect 103992 217002 104020 218010
rect 104636 217002 104664 221954
rect 104820 218074 104848 224062
rect 104808 218068 104860 218074
rect 104808 218010 104860 218016
rect 105740 217002 105768 225286
rect 106200 217002 106228 228074
rect 109868 227724 109920 227730
rect 109868 227666 109920 227672
rect 106924 226908 106976 226914
rect 106924 226850 106976 226856
rect 106936 219434 106964 226850
rect 108304 225752 108356 225758
rect 108304 225694 108356 225700
rect 108316 225486 108344 225694
rect 108304 225480 108356 225486
rect 108304 225422 108356 225428
rect 108948 224528 109000 224534
rect 108948 224470 109000 224476
rect 108120 221060 108172 221066
rect 108120 221002 108172 221008
rect 107936 220924 107988 220930
rect 107936 220866 107988 220872
rect 107948 220658 107976 220866
rect 107936 220652 107988 220658
rect 107936 220594 107988 220600
rect 106924 219428 106976 219434
rect 106924 219370 106976 219376
rect 107292 218340 107344 218346
rect 107292 218282 107344 218288
rect 107304 217002 107332 218282
rect 108132 217002 108160 221002
rect 108304 219292 108356 219298
rect 108304 219234 108356 219240
rect 108316 218482 108344 219234
rect 108304 218476 108356 218482
rect 108304 218418 108356 218424
rect 108960 217002 108988 224470
rect 109880 217002 109908 227666
rect 111076 218074 111104 230114
rect 113088 228132 113140 228138
rect 113088 228074 113140 228080
rect 112904 222352 112956 222358
rect 112904 222294 112956 222300
rect 111432 219972 111484 219978
rect 111432 219914 111484 219920
rect 110328 218068 110380 218074
rect 110328 218010 110380 218016
rect 111064 218068 111116 218074
rect 111064 218010 111116 218016
rect 110340 217002 110368 218010
rect 111444 217002 111472 219914
rect 112916 218074 112944 222294
rect 112260 218068 112312 218074
rect 112260 218010 112312 218016
rect 112904 218068 112956 218074
rect 112904 218010 112956 218016
rect 112272 217002 112300 218010
rect 113100 217002 113128 228074
rect 117228 225344 117280 225350
rect 117228 225286 117280 225292
rect 116860 224936 116912 224942
rect 116860 224878 116912 224884
rect 115664 224664 115716 224670
rect 115664 224606 115716 224612
rect 114468 221332 114520 221338
rect 114468 221274 114520 221280
rect 113916 218204 113968 218210
rect 113916 218146 113968 218152
rect 113928 217002 113956 218146
rect 114480 217002 114508 221274
rect 115676 217002 115704 224606
rect 116872 224126 116900 224878
rect 116860 224120 116912 224126
rect 116860 224062 116912 224068
rect 117044 224120 117096 224126
rect 117044 224062 117096 224068
rect 116400 218068 116452 218074
rect 116400 218010 116452 218016
rect 116412 217002 116440 218010
rect 117056 217002 117084 224062
rect 117240 218074 117268 225286
rect 118436 224126 118464 230250
rect 140044 229628 140096 229634
rect 140044 229570 140096 229576
rect 131120 229492 131172 229498
rect 131120 229434 131172 229440
rect 122932 229356 122984 229362
rect 122932 229298 122984 229304
rect 122748 227996 122800 228002
rect 122748 227938 122800 227944
rect 121368 226772 121420 226778
rect 121368 226714 121420 226720
rect 119804 226636 119856 226642
rect 119804 226578 119856 226584
rect 118608 224800 118660 224806
rect 118608 224742 118660 224748
rect 118424 224120 118476 224126
rect 118424 224062 118476 224068
rect 117964 223304 118016 223310
rect 117964 223246 118016 223252
rect 118148 223304 118200 223310
rect 118148 223246 118200 223252
rect 117976 222494 118004 223246
rect 117964 222488 118016 222494
rect 117964 222430 118016 222436
rect 118160 222358 118188 223246
rect 118148 222352 118200 222358
rect 118148 222294 118200 222300
rect 117964 222148 118016 222154
rect 117964 222090 118016 222096
rect 118148 222148 118200 222154
rect 118148 222090 118200 222096
rect 117976 221202 118004 222090
rect 117964 221196 118016 221202
rect 117964 221138 118016 221144
rect 118160 221066 118188 222090
rect 118148 221060 118200 221066
rect 118148 221002 118200 221008
rect 118056 220924 118108 220930
rect 118056 220866 118108 220872
rect 117872 219428 117924 219434
rect 117872 219370 117924 219376
rect 117884 219162 117912 219370
rect 117872 219156 117924 219162
rect 117872 219098 117924 219104
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 118068 217002 118096 220866
rect 118620 217002 118648 224742
rect 119816 217002 119844 226578
rect 120540 218068 120592 218074
rect 120540 218010 120592 218016
rect 120552 217002 120580 218010
rect 121380 217002 121408 226714
rect 122288 224120 122340 224126
rect 122288 224062 122340 224068
rect 122300 217002 122328 224062
rect 122760 217002 122788 227938
rect 122944 224942 122972 229298
rect 125784 226908 125836 226914
rect 125784 226850 125836 226856
rect 125796 226506 125824 226850
rect 125784 226500 125836 226506
rect 125784 226442 125836 226448
rect 129648 226500 129700 226506
rect 129648 226442 129700 226448
rect 127440 225480 127492 225486
rect 127440 225422 127492 225428
rect 127452 225214 127480 225422
rect 127440 225208 127492 225214
rect 127440 225150 127492 225156
rect 128084 225208 128136 225214
rect 128084 225150 128136 225156
rect 126888 225072 126940 225078
rect 126888 225014 126940 225020
rect 122932 224936 122984 224942
rect 122932 224878 122984 224884
rect 126520 224936 126572 224942
rect 126520 224878 126572 224884
rect 126532 224398 126560 224878
rect 126520 224392 126572 224398
rect 126520 224334 126572 224340
rect 126704 224392 126756 224398
rect 126704 224334 126756 224340
rect 125140 223848 125192 223854
rect 125140 223790 125192 223796
rect 123482 222864 123538 222873
rect 123482 222799 123538 222808
rect 123496 219434 123524 222799
rect 124680 219836 124732 219842
rect 124680 219778 124732 219784
rect 123484 219428 123536 219434
rect 123484 219370 123536 219376
rect 123852 219156 123904 219162
rect 123852 219098 123904 219104
rect 123864 217002 123892 219098
rect 124692 217002 124720 219778
rect 101876 216974 102028 217002
rect 102856 216974 103284 217002
rect 103684 216974 104020 217002
rect 104512 216974 104664 217002
rect 105340 216974 105768 217002
rect 106168 216974 106228 217002
rect 106996 216974 107332 217002
rect 107824 216974 108160 217002
rect 108652 216974 108988 217002
rect 109480 216974 109908 217002
rect 110308 216974 110368 217002
rect 111136 216974 111472 217002
rect 111964 216974 112300 217002
rect 112792 216974 113128 217002
rect 113620 216974 113956 217002
rect 114448 216974 114508 217002
rect 115276 216974 115704 217002
rect 116104 216974 116440 217002
rect 116932 216974 117084 217002
rect 117760 216974 118096 217002
rect 118588 216974 118648 217002
rect 119416 216974 119844 217002
rect 120244 216974 120580 217002
rect 121072 216974 121408 217002
rect 121900 216974 122328 217002
rect 122728 216974 122788 217002
rect 123556 216974 123892 217002
rect 124384 216974 124720 217002
rect 125152 217002 125180 223790
rect 126336 218476 126388 218482
rect 126336 218418 126388 218424
rect 126348 217002 126376 218418
rect 125152 216974 125212 217002
rect 126040 216974 126376 217002
rect 126716 217002 126744 224334
rect 126900 218482 126928 225014
rect 127072 219156 127124 219162
rect 127072 219098 127124 219104
rect 127084 218482 127112 219098
rect 126888 218476 126940 218482
rect 126888 218418 126940 218424
rect 127072 218476 127124 218482
rect 127072 218418 127124 218424
rect 128096 217002 128124 225150
rect 128820 221060 128872 221066
rect 128820 221002 128872 221008
rect 128832 217002 128860 221002
rect 129660 217002 129688 226442
rect 131132 224398 131160 229434
rect 134614 228032 134670 228041
rect 134614 227967 134670 227976
rect 133788 227860 133840 227866
rect 133788 227802 133840 227808
rect 131120 224392 131172 224398
rect 131120 224334 131172 224340
rect 131304 224392 131356 224398
rect 131304 224334 131356 224340
rect 131316 224126 131344 224334
rect 131304 224120 131356 224126
rect 131304 224062 131356 224068
rect 131488 224120 131540 224126
rect 131488 224062 131540 224068
rect 131500 223854 131528 224062
rect 131488 223848 131540 223854
rect 131488 223790 131540 223796
rect 132224 223712 132276 223718
rect 132224 223654 132276 223660
rect 131028 219564 131080 219570
rect 131028 219506 131080 219512
rect 130476 219156 130528 219162
rect 130476 219098 130528 219104
rect 130488 217002 130516 219098
rect 131040 217002 131068 219506
rect 132236 217002 132264 223654
rect 133604 222352 133656 222358
rect 133604 222294 133656 222300
rect 132776 219428 132828 219434
rect 132776 219370 132828 219376
rect 132788 219026 132816 219370
rect 132776 219020 132828 219026
rect 132776 218962 132828 218968
rect 132960 219020 133012 219026
rect 132960 218962 133012 218968
rect 132972 217002 133000 218962
rect 133616 217002 133644 222294
rect 133800 219026 133828 227802
rect 133788 219020 133840 219026
rect 133788 218962 133840 218968
rect 134628 217002 134656 227967
rect 135260 227044 135312 227050
rect 135260 226986 135312 226992
rect 135444 227044 135496 227050
rect 135444 226986 135496 226992
rect 135272 226522 135300 226986
rect 135456 226642 135484 226986
rect 135444 226636 135496 226642
rect 135444 226578 135496 226584
rect 135628 226636 135680 226642
rect 135628 226578 135680 226584
rect 137560 226636 137612 226642
rect 137560 226578 137612 226584
rect 135640 226522 135668 226578
rect 137572 226522 137600 226578
rect 135272 226494 135668 226522
rect 137204 226506 137600 226522
rect 137192 226500 137600 226506
rect 137244 226494 137600 226500
rect 139306 226536 139362 226545
rect 139306 226471 139362 226480
rect 137192 226442 137244 226448
rect 136824 225616 136876 225622
rect 136824 225558 136876 225564
rect 137008 225616 137060 225622
rect 137008 225558 137060 225564
rect 136362 225312 136418 225321
rect 136362 225247 136418 225256
rect 134984 223848 135036 223854
rect 134984 223790 135036 223796
rect 126716 216974 126868 217002
rect 127696 216974 128124 217002
rect 128524 216974 128860 217002
rect 129352 216974 129688 217002
rect 130180 216974 130516 217002
rect 131008 216974 131068 217002
rect 131836 216974 132264 217002
rect 132664 216974 133000 217002
rect 133492 216974 133644 217002
rect 134320 216974 134656 217002
rect 134996 217002 135024 223790
rect 136376 217002 136404 225247
rect 136836 225162 136864 225558
rect 137020 225350 137048 225558
rect 137008 225344 137060 225350
rect 137008 225286 137060 225292
rect 136836 225134 137508 225162
rect 137480 225078 137508 225134
rect 137468 225072 137520 225078
rect 137468 225014 137520 225020
rect 137100 222896 137152 222902
rect 137100 222838 137152 222844
rect 137284 222896 137336 222902
rect 137284 222838 137336 222844
rect 137112 222358 137140 222838
rect 137296 222494 137324 222838
rect 137284 222488 137336 222494
rect 137284 222430 137336 222436
rect 137468 222488 137520 222494
rect 137468 222430 137520 222436
rect 136916 222352 136968 222358
rect 136916 222294 136968 222300
rect 137100 222352 137152 222358
rect 137480 222306 137508 222430
rect 137100 222294 137152 222300
rect 136928 222194 136956 222294
rect 137296 222278 137508 222306
rect 137296 222194 137324 222278
rect 136928 222166 137324 222194
rect 138570 221776 138626 221785
rect 138570 221711 138626 221720
rect 137284 221604 137336 221610
rect 137284 221546 137336 221552
rect 137468 221604 137520 221610
rect 137468 221546 137520 221552
rect 137296 221202 137324 221546
rect 137100 221196 137152 221202
rect 137100 221138 137152 221144
rect 137284 221196 137336 221202
rect 137284 221138 137336 221144
rect 137112 221082 137140 221138
rect 137480 221082 137508 221546
rect 138584 221474 138612 221711
rect 138572 221468 138624 221474
rect 138572 221410 138624 221416
rect 138756 221468 138808 221474
rect 138756 221410 138808 221416
rect 137112 221054 137508 221082
rect 137284 220788 137336 220794
rect 137284 220730 137336 220736
rect 137468 220788 137520 220794
rect 137468 220730 137520 220736
rect 137296 219706 137324 220730
rect 137284 219700 137336 219706
rect 137284 219642 137336 219648
rect 137480 219570 137508 220730
rect 137468 219564 137520 219570
rect 137468 219506 137520 219512
rect 137928 219564 137980 219570
rect 137928 219506 137980 219512
rect 137100 219020 137152 219026
rect 137100 218962 137152 218968
rect 137112 217002 137140 218962
rect 137940 217002 137968 219506
rect 138768 217002 138796 221410
rect 139320 217002 139348 226471
rect 140056 219434 140084 229570
rect 140792 228546 140820 231662
rect 140780 228540 140832 228546
rect 140780 228482 140832 228488
rect 140964 228540 141016 228546
rect 140964 228482 141016 228488
rect 140976 228274 141004 228482
rect 140964 228268 141016 228274
rect 140964 228210 141016 228216
rect 141148 228268 141200 228274
rect 141148 228210 141200 228216
rect 141160 228041 141188 228210
rect 141146 228032 141202 228041
rect 141146 227967 141202 227976
rect 141528 225078 141556 231662
rect 142158 227216 142214 227225
rect 142158 227151 142214 227160
rect 142172 226658 142200 227151
rect 142126 226630 142200 226658
rect 142126 226506 142154 226630
rect 142250 226536 142306 226545
rect 142114 226500 142166 226506
rect 142250 226471 142252 226480
rect 142114 226442 142166 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 142114 225344 142166 225350
rect 142252 225344 142304 225350
rect 142114 225286 142166 225292
rect 142250 225312 142252 225321
rect 142304 225312 142306 225321
rect 142126 225162 142154 225286
rect 142250 225247 142306 225256
rect 142448 225162 142476 231676
rect 143092 227225 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 145038 231662 145236 231690
rect 143078 227216 143134 227225
rect 143078 227151 143134 227160
rect 143552 226166 143580 231662
rect 143540 226160 143592 226166
rect 143540 226102 143592 226108
rect 142986 225584 143042 225593
rect 142986 225519 143042 225528
rect 142126 225134 142200 225162
rect 142448 225134 142660 225162
rect 141516 225072 141568 225078
rect 141516 225014 141568 225020
rect 141884 225072 141936 225078
rect 142172 225060 142200 225134
rect 142436 225072 142488 225078
rect 142172 225032 142436 225060
rect 141884 225014 141936 225020
rect 142436 225014 142488 225020
rect 141608 224256 141660 224262
rect 141608 224198 141660 224204
rect 141620 223990 141648 224198
rect 141424 223984 141476 223990
rect 141422 223952 141424 223961
rect 141608 223984 141660 223990
rect 141476 223952 141478 223961
rect 141608 223926 141660 223932
rect 141422 223887 141478 223896
rect 141054 220824 141110 220833
rect 141054 220759 141110 220768
rect 141068 220114 141096 220759
rect 141056 220108 141108 220114
rect 141056 220050 141108 220056
rect 141240 220108 141292 220114
rect 141240 220050 141292 220056
rect 140044 219428 140096 219434
rect 140044 219370 140096 219376
rect 140226 218648 140282 218657
rect 140226 218583 140228 218592
rect 140280 218583 140282 218592
rect 140412 218612 140464 218618
rect 140228 218554 140280 218560
rect 140412 218554 140464 218560
rect 140424 217002 140452 218554
rect 141252 217002 141280 220050
rect 141896 217002 141924 225014
rect 142068 224936 142120 224942
rect 142068 224878 142120 224884
rect 142080 224262 142108 224878
rect 142068 224256 142120 224262
rect 142068 224198 142120 224204
rect 142632 222358 142660 225134
rect 142620 222352 142672 222358
rect 142620 222294 142672 222300
rect 142804 221876 142856 221882
rect 142804 221818 142856 221824
rect 142816 221610 142844 221818
rect 142804 221604 142856 221610
rect 142804 221546 142856 221552
rect 142436 221468 142488 221474
rect 142436 221410 142488 221416
rect 142448 221241 142476 221410
rect 142434 221232 142490 221241
rect 142434 221167 142490 221176
rect 143000 219586 143028 225519
rect 143448 222284 143500 222290
rect 143448 222226 143500 222232
rect 143172 221876 143224 221882
rect 143172 221818 143224 221824
rect 143184 221474 143212 221818
rect 143172 221468 143224 221474
rect 143172 221410 143224 221416
rect 134996 216974 135148 217002
rect 135976 216974 136404 217002
rect 136804 216974 137140 217002
rect 137632 216974 137968 217002
rect 138460 216974 138796 217002
rect 139288 216974 139348 217002
rect 140116 216974 140452 217002
rect 140944 216974 141280 217002
rect 141772 216974 141924 217002
rect 142448 219558 143028 219586
rect 142448 217002 142476 219558
rect 142804 219428 142856 219434
rect 142804 219370 142856 219376
rect 142816 219026 142844 219370
rect 142804 219020 142856 219026
rect 142804 218962 142856 218968
rect 143172 219020 143224 219026
rect 143172 218962 143224 218968
rect 143184 218906 143212 218962
rect 142632 218878 143212 218906
rect 142632 218618 142660 218878
rect 142620 218612 142672 218618
rect 142620 218554 142672 218560
rect 143460 217002 143488 222226
rect 144012 221202 144040 231662
rect 144644 230580 144696 230586
rect 144644 230522 144696 230528
rect 144656 229770 144684 230522
rect 144644 229764 144696 229770
rect 144644 229706 144696 229712
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 222290 144868 229706
rect 145208 223990 145236 231662
rect 145668 229809 145696 231676
rect 146326 231662 146524 231690
rect 145654 229800 145710 229809
rect 145654 229735 145710 229744
rect 146298 229256 146354 229265
rect 146298 229191 146300 229200
rect 146352 229191 146354 229200
rect 146300 229162 146352 229168
rect 146496 229094 146524 231662
rect 146680 231662 146970 231690
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 148428 231662 148902 231690
rect 149072 231662 149546 231690
rect 146680 229094 146708 231662
rect 146944 229628 146996 229634
rect 146944 229570 146996 229576
rect 146956 229226 146984 229570
rect 146944 229220 146996 229226
rect 146944 229162 146996 229168
rect 146404 229066 146524 229094
rect 146588 229066 146708 229094
rect 145930 228032 145986 228041
rect 145930 227967 145986 227976
rect 145196 223984 145248 223990
rect 145380 223984 145432 223990
rect 145196 223926 145248 223932
rect 145378 223952 145380 223961
rect 145432 223952 145434 223961
rect 145378 223887 145434 223896
rect 145012 222352 145064 222358
rect 145012 222294 145064 222300
rect 144828 222284 144880 222290
rect 144828 222226 144880 222232
rect 145024 222170 145052 222294
rect 144656 222142 145052 222170
rect 144182 221232 144238 221241
rect 144000 221196 144052 221202
rect 144182 221167 144184 221176
rect 144000 221138 144052 221144
rect 144236 221167 144238 221176
rect 144184 221138 144236 221144
rect 143632 218884 143684 218890
rect 143632 218826 143684 218832
rect 143644 218657 143672 218826
rect 143630 218648 143686 218657
rect 143630 218583 143686 218592
rect 144656 217002 144684 222142
rect 145380 221468 145432 221474
rect 145380 221410 145432 221416
rect 145392 217002 145420 221410
rect 145944 217002 145972 227967
rect 146206 223952 146262 223961
rect 146206 223887 146262 223896
rect 146220 218890 146248 223887
rect 146404 220833 146432 229066
rect 146588 221785 146616 229066
rect 146944 226160 146996 226166
rect 146944 226102 146996 226108
rect 146956 225622 146984 226102
rect 146944 225616 146996 225622
rect 146944 225558 146996 225564
rect 147232 223990 147260 231662
rect 147968 229265 147996 231662
rect 147954 229256 148010 229265
rect 147954 229191 148010 229200
rect 147404 225616 147456 225622
rect 147402 225584 147404 225593
rect 147456 225584 147458 225593
rect 147402 225519 147458 225528
rect 147220 223984 147272 223990
rect 147680 223984 147732 223990
rect 147220 223926 147272 223932
rect 147678 223952 147680 223961
rect 147732 223952 147734 223961
rect 147678 223887 147734 223896
rect 147310 222184 147366 222193
rect 147310 222119 147366 222128
rect 146574 221776 146630 221785
rect 146574 221711 146630 221720
rect 147324 221610 147352 222119
rect 147494 221912 147550 221921
rect 147494 221847 147550 221856
rect 147508 221746 147536 221847
rect 147496 221740 147548 221746
rect 147496 221682 147548 221688
rect 147312 221604 147364 221610
rect 147312 221546 147364 221552
rect 148428 220833 148456 231662
rect 148784 229764 148836 229770
rect 148784 229706 148836 229712
rect 148796 229094 148824 229706
rect 148612 229066 148824 229094
rect 146390 220824 146446 220833
rect 146390 220759 146446 220768
rect 147218 220824 147274 220833
rect 147218 220759 147274 220768
rect 148414 220824 148470 220833
rect 148414 220759 148470 220768
rect 147232 220250 147260 220759
rect 147220 220244 147272 220250
rect 147220 220186 147272 220192
rect 147508 220114 147674 220130
rect 147508 220108 147686 220114
rect 147508 220102 147634 220108
rect 146208 218884 146260 218890
rect 146208 218826 146260 218832
rect 146714 217252 146766 217258
rect 146714 217194 146766 217200
rect 142448 216974 142600 217002
rect 143428 216974 143488 217002
rect 144256 216974 144684 217002
rect 145084 216974 145420 217002
rect 145912 216974 145972 217002
rect 146726 216988 146754 217194
rect 147508 217002 147536 220102
rect 147634 220050 147686 220056
rect 148612 218634 148640 229066
rect 149072 221921 149100 231662
rect 150176 228410 150204 231676
rect 150544 231662 150834 231690
rect 151004 231662 151478 231690
rect 151832 231662 152122 231690
rect 150544 230586 150572 231662
rect 150532 230580 150584 230586
rect 150532 230522 150584 230528
rect 151004 229094 151032 231662
rect 151358 229936 151414 229945
rect 151832 229922 151860 231662
rect 152188 230580 152240 230586
rect 152188 230522 152240 230528
rect 151358 229871 151414 229880
rect 151786 229894 151860 229922
rect 150820 229066 151032 229094
rect 150164 228404 150216 228410
rect 150164 228346 150216 228352
rect 150348 228404 150400 228410
rect 150348 228346 150400 228352
rect 150360 228041 150388 228346
rect 150346 228032 150402 228041
rect 150346 227967 150402 227976
rect 150346 226672 150402 226681
rect 150346 226607 150402 226616
rect 149058 221912 149114 221921
rect 149058 221847 149114 221856
rect 148784 221468 148836 221474
rect 148784 221410 148836 221416
rect 148520 218618 148640 218634
rect 148508 218612 148640 218618
rect 148560 218606 148640 218612
rect 148508 218554 148560 218560
rect 148796 217002 148824 221410
rect 149980 219292 150032 219298
rect 149980 219234 150032 219240
rect 150164 219292 150216 219298
rect 150164 219234 150216 219240
rect 149334 218784 149390 218793
rect 149334 218719 149336 218728
rect 149388 218719 149390 218728
rect 149520 218748 149572 218754
rect 149336 218690 149388 218696
rect 149520 218690 149572 218696
rect 149532 217002 149560 218690
rect 149992 218618 150020 219234
rect 149980 218612 150032 218618
rect 149980 218554 150032 218560
rect 150176 217002 150204 219234
rect 150360 218754 150388 226607
rect 150622 220824 150678 220833
rect 150622 220759 150678 220768
rect 150636 220386 150664 220759
rect 150624 220380 150676 220386
rect 150624 220322 150676 220328
rect 150820 220153 150848 229066
rect 151372 222494 151400 229871
rect 151786 229650 151814 229894
rect 151912 229764 151964 229770
rect 151912 229706 151964 229712
rect 151924 229650 151952 229706
rect 152200 229650 152228 230522
rect 152370 229936 152426 229945
rect 152370 229871 152426 229880
rect 152384 229770 152412 229871
rect 152372 229764 152424 229770
rect 152372 229706 152424 229712
rect 151786 229622 151860 229650
rect 151924 229622 152228 229650
rect 151832 229094 151860 229622
rect 151832 229066 152136 229094
rect 151818 227352 151874 227361
rect 151818 227287 151874 227296
rect 151832 227202 151860 227287
rect 151740 227186 151860 227202
rect 151728 227180 151860 227186
rect 151780 227174 151860 227180
rect 151728 227122 151780 227128
rect 151726 223816 151782 223825
rect 151726 223751 151782 223760
rect 151360 222488 151412 222494
rect 151360 222430 151412 222436
rect 150806 220144 150862 220153
rect 150806 220079 150862 220088
rect 150348 218748 150400 218754
rect 150348 218690 150400 218696
rect 151176 218612 151228 218618
rect 151176 218554 151228 218560
rect 151188 217002 151216 218554
rect 151740 217002 151768 223751
rect 152108 222193 152136 229066
rect 152280 227180 152332 227186
rect 152280 227122 152332 227128
rect 152292 226681 152320 227122
rect 152278 226672 152334 226681
rect 152278 226607 152334 226616
rect 152752 224369 152780 231676
rect 153396 229226 153424 231676
rect 153580 231662 154054 231690
rect 153384 229220 153436 229226
rect 153384 229162 153436 229168
rect 153580 229094 153608 231662
rect 153844 229220 153896 229226
rect 153844 229162 153896 229168
rect 153580 229066 153792 229094
rect 152922 226128 152978 226137
rect 152922 226063 152978 226072
rect 152738 224360 152794 224369
rect 152738 224295 152794 224304
rect 152280 223168 152332 223174
rect 152280 223110 152332 223116
rect 152464 223168 152516 223174
rect 152464 223110 152516 223116
rect 152292 222494 152320 223110
rect 152476 222902 152504 223110
rect 152464 222896 152516 222902
rect 152464 222838 152516 222844
rect 152280 222488 152332 222494
rect 152280 222430 152332 222436
rect 152094 222184 152150 222193
rect 152094 222119 152150 222128
rect 152648 220516 152700 220522
rect 152648 220458 152700 220464
rect 152660 219706 152688 220458
rect 152648 219700 152700 219706
rect 152648 219642 152700 219648
rect 152464 219020 152516 219026
rect 152464 218962 152516 218968
rect 152476 217258 152504 218962
rect 152464 217252 152516 217258
rect 152464 217194 152516 217200
rect 152936 217002 152964 226063
rect 153764 220561 153792 229066
rect 153856 224954 153884 229162
rect 154684 227361 154712 231676
rect 154670 227352 154726 227361
rect 154670 227287 154726 227296
rect 155328 226953 155356 231676
rect 155972 229906 156000 231676
rect 156156 231662 156630 231690
rect 155960 229900 156012 229906
rect 155960 229842 156012 229848
rect 155866 228032 155922 228041
rect 155866 227967 155922 227976
rect 155314 226944 155370 226953
rect 155314 226879 155370 226888
rect 154212 226296 154264 226302
rect 154264 226244 154804 226250
rect 154212 226238 154804 226244
rect 154224 226222 154804 226238
rect 154776 226166 154804 226222
rect 154764 226160 154816 226166
rect 154764 226102 154816 226108
rect 153856 224926 153976 224954
rect 153750 220552 153806 220561
rect 153750 220487 153806 220496
rect 153108 219700 153160 219706
rect 153108 219642 153160 219648
rect 153120 218618 153148 219642
rect 153948 218793 153976 224926
rect 154578 223986 154634 223995
rect 154578 223921 154634 223930
rect 154488 222896 154540 222902
rect 154488 222838 154540 222844
rect 153934 218784 153990 218793
rect 153934 218719 153990 218728
rect 153108 218612 153160 218618
rect 153108 218554 153160 218560
rect 153660 218612 153712 218618
rect 153660 218554 153712 218560
rect 153672 217002 153700 218554
rect 154500 217002 154528 222838
rect 155314 222456 155370 222465
rect 155314 222391 155370 222400
rect 155328 217002 155356 222391
rect 155880 217002 155908 227967
rect 156156 220833 156184 231662
rect 156604 229900 156656 229906
rect 156604 229842 156656 229848
rect 156616 229094 156644 229842
rect 156248 229066 156644 229094
rect 156248 224954 156276 229066
rect 156420 228540 156472 228546
rect 156420 228482 156472 228488
rect 156432 228426 156460 228482
rect 156432 228410 157012 228426
rect 156432 228404 157024 228410
rect 156432 228398 156972 228404
rect 156972 228346 157024 228352
rect 156512 227180 156564 227186
rect 156512 227122 156564 227128
rect 156524 227032 156552 227122
rect 156972 227044 157024 227050
rect 156524 227004 156972 227032
rect 156972 226986 157024 226992
rect 157260 224954 157288 231676
rect 157628 231662 157918 231690
rect 158272 231662 158562 231690
rect 158824 231662 159206 231690
rect 157430 228576 157486 228585
rect 157430 228511 157486 228520
rect 157444 228410 157472 228511
rect 157432 228404 157484 228410
rect 157432 228346 157484 228352
rect 157628 226250 157656 231662
rect 158272 230722 158300 231662
rect 158260 230716 158312 230722
rect 158260 230658 158312 230664
rect 157982 228984 158038 228993
rect 157982 228919 158038 228928
rect 157800 228404 157852 228410
rect 157800 228346 157852 228352
rect 157812 228041 157840 228346
rect 157798 228032 157854 228041
rect 157798 227967 157854 227976
rect 157444 226222 157656 226250
rect 157444 226166 157472 226222
rect 157432 226160 157484 226166
rect 157616 226160 157668 226166
rect 157432 226102 157484 226108
rect 157614 226128 157616 226137
rect 157668 226128 157670 226137
rect 157614 226063 157670 226072
rect 156248 224926 156368 224954
rect 156142 220824 156198 220833
rect 156142 220759 156198 220768
rect 156340 218754 156368 224926
rect 157076 224926 157288 224954
rect 156880 223984 156932 223990
rect 156880 223926 156932 223932
rect 156892 223825 156920 223926
rect 156878 223816 156934 223825
rect 156878 223751 156934 223760
rect 157076 222494 157104 224926
rect 157338 224496 157394 224505
rect 157338 224431 157394 224440
rect 157352 224346 157380 224431
rect 157306 224318 157380 224346
rect 157306 224262 157334 224318
rect 157294 224256 157346 224262
rect 157294 224198 157346 224204
rect 157432 224256 157484 224262
rect 157432 224198 157484 224204
rect 157444 224097 157472 224198
rect 157430 224088 157486 224097
rect 157430 224023 157486 224032
rect 157248 223440 157300 223446
rect 157246 223408 157248 223417
rect 157432 223440 157484 223446
rect 157300 223408 157302 223417
rect 157246 223343 157302 223352
rect 157430 223408 157432 223417
rect 157484 223408 157486 223417
rect 157430 223343 157486 223352
rect 157064 222488 157116 222494
rect 157248 222488 157300 222494
rect 157064 222430 157116 222436
rect 157246 222456 157248 222465
rect 157300 222456 157302 222465
rect 157246 222391 157302 222400
rect 157614 220416 157670 220425
rect 157614 220351 157616 220360
rect 157668 220351 157670 220360
rect 157800 220380 157852 220386
rect 157616 220322 157668 220328
rect 157800 220322 157852 220328
rect 156328 218748 156380 218754
rect 156328 218690 156380 218696
rect 156972 218748 157024 218754
rect 156972 218690 157024 218696
rect 156984 217002 157012 218690
rect 157812 217002 157840 220322
rect 157996 218346 158024 228919
rect 158824 228585 158852 231662
rect 158810 228576 158866 228585
rect 158810 228511 158866 228520
rect 159638 227488 159694 227497
rect 159638 227423 159640 227432
rect 159692 227423 159694 227432
rect 159640 227394 159692 227400
rect 159836 223446 159864 231676
rect 160480 228313 160508 231676
rect 161124 230450 161152 231676
rect 161112 230444 161164 230450
rect 161112 230386 161164 230392
rect 161296 230444 161348 230450
rect 161296 230386 161348 230392
rect 160466 228304 160522 228313
rect 160466 228239 160522 228248
rect 160008 227452 160060 227458
rect 160008 227394 160060 227400
rect 159824 223440 159876 223446
rect 158626 223408 158682 223417
rect 159824 223382 159876 223388
rect 158626 223343 158682 223352
rect 157984 218340 158036 218346
rect 157984 218282 158036 218288
rect 158640 217002 158668 223343
rect 159824 218204 159876 218210
rect 159824 218146 159876 218152
rect 159456 218068 159508 218074
rect 159456 218010 159508 218016
rect 159468 217002 159496 218010
rect 147508 216974 147568 217002
rect 148396 216974 148824 217002
rect 149224 216974 149560 217002
rect 150052 216974 150204 217002
rect 150880 216974 151216 217002
rect 151708 216974 151768 217002
rect 152536 216974 152964 217002
rect 153364 216974 153700 217002
rect 154192 216974 154528 217002
rect 155020 216974 155356 217002
rect 155848 216974 155908 217002
rect 156676 216974 157012 217002
rect 157504 216974 157840 217002
rect 158332 216974 158668 217002
rect 159160 216974 159496 217002
rect 159836 217002 159864 218146
rect 160020 218074 160048 227394
rect 161112 223440 161164 223446
rect 161112 223382 161164 223388
rect 160008 218068 160060 218074
rect 160008 218010 160060 218016
rect 161124 217002 161152 223382
rect 161308 219298 161336 230386
rect 161572 226024 161624 226030
rect 161572 225966 161624 225972
rect 161584 225593 161612 225966
rect 161570 225584 161626 225593
rect 161570 225519 161626 225528
rect 161768 224954 161796 231676
rect 162136 231662 162426 231690
rect 162964 231662 163070 231690
rect 161940 226296 161992 226302
rect 161940 226238 161992 226244
rect 161952 226030 161980 226238
rect 161940 226024 161992 226030
rect 161940 225966 161992 225972
rect 161584 224926 161796 224954
rect 161584 220425 161612 224926
rect 162136 222766 162164 231662
rect 162308 226296 162360 226302
rect 162308 226238 162360 226244
rect 162320 225078 162348 226238
rect 162308 225072 162360 225078
rect 162308 225014 162360 225020
rect 162768 225072 162820 225078
rect 162768 225014 162820 225020
rect 162308 223440 162360 223446
rect 162308 223382 162360 223388
rect 162320 222766 162348 223382
rect 162124 222760 162176 222766
rect 162124 222702 162176 222708
rect 162308 222760 162360 222766
rect 162308 222702 162360 222708
rect 161756 221740 161808 221746
rect 161756 221682 161808 221688
rect 161570 220416 161626 220425
rect 161570 220351 161626 220360
rect 161296 219292 161348 219298
rect 161296 219234 161348 219240
rect 161570 218376 161626 218385
rect 161570 218311 161572 218320
rect 161624 218311 161626 218320
rect 161572 218282 161624 218288
rect 161768 217002 161796 221682
rect 162308 219156 162360 219162
rect 162308 219098 162360 219104
rect 162320 218890 162348 219098
rect 162308 218884 162360 218890
rect 162308 218826 162360 218832
rect 162492 218884 162544 218890
rect 162492 218826 162544 218832
rect 161940 218748 161992 218754
rect 161940 218690 161992 218696
rect 161952 218346 161980 218690
rect 162308 218612 162360 218618
rect 162308 218554 162360 218560
rect 162320 218385 162348 218554
rect 162306 218376 162362 218385
rect 161940 218340 161992 218346
rect 162306 218311 162362 218320
rect 161940 218282 161992 218288
rect 162504 218210 162532 218826
rect 162492 218204 162544 218210
rect 162492 218146 162544 218152
rect 162780 217002 162808 225014
rect 162964 224505 162992 231662
rect 163700 229226 163728 231676
rect 163688 229220 163740 229226
rect 163688 229162 163740 229168
rect 163872 229220 163924 229226
rect 163872 229162 163924 229168
rect 163884 228993 163912 229162
rect 163870 228984 163926 228993
rect 163870 228919 163926 228928
rect 164344 227322 164372 231676
rect 164332 227316 164384 227322
rect 164332 227258 164384 227264
rect 162950 224496 163006 224505
rect 162950 224431 163006 224440
rect 163962 223952 164018 223961
rect 163962 223887 164018 223896
rect 163976 218618 164004 223887
rect 164988 223582 165016 231676
rect 165344 227316 165396 227322
rect 165344 227258 165396 227264
rect 164976 223576 165028 223582
rect 164976 223518 165028 223524
rect 164148 223440 164200 223446
rect 164148 223382 164200 223388
rect 163964 218612 164016 218618
rect 163964 218554 164016 218560
rect 163596 218204 163648 218210
rect 163596 218146 163648 218152
rect 163608 217002 163636 218146
rect 164160 217002 164188 223382
rect 165158 220280 165214 220289
rect 165158 220215 165214 220224
rect 165172 218346 165200 220215
rect 165160 218340 165212 218346
rect 165160 218282 165212 218288
rect 165356 217002 165384 227258
rect 165632 222873 165660 231676
rect 166080 230580 166132 230586
rect 166080 230522 166132 230528
rect 166092 223038 166120 230522
rect 166276 230042 166304 231676
rect 166460 231662 166934 231690
rect 167196 231662 167578 231690
rect 166264 230036 166316 230042
rect 166264 229978 166316 229984
rect 166460 227497 166488 231662
rect 166632 230036 166684 230042
rect 166632 229978 166684 229984
rect 166644 229226 166672 229978
rect 166632 229220 166684 229226
rect 166632 229162 166684 229168
rect 166630 228440 166686 228449
rect 166630 228375 166686 228384
rect 166446 227488 166502 227497
rect 166446 227423 166502 227432
rect 166644 225706 166672 228375
rect 166908 227452 166960 227458
rect 166908 227394 166960 227400
rect 166920 226386 166948 227394
rect 166920 226370 166994 226386
rect 166920 226364 167006 226370
rect 166920 226358 166954 226364
rect 166954 226306 167006 226312
rect 166816 226296 166868 226302
rect 166816 226238 166868 226244
rect 166828 225978 166856 226238
rect 166828 225950 166994 225978
rect 166966 225894 166994 225950
rect 166816 225888 166868 225894
rect 166814 225856 166816 225865
rect 166954 225888 167006 225894
rect 166868 225856 166870 225865
rect 166954 225830 167006 225836
rect 166814 225791 166870 225800
rect 166644 225678 166948 225706
rect 166722 225584 166778 225593
rect 166722 225519 166778 225528
rect 166736 225078 166764 225519
rect 166540 225072 166592 225078
rect 166538 225040 166540 225049
rect 166724 225072 166776 225078
rect 166592 225040 166594 225049
rect 166724 225014 166776 225020
rect 166538 224975 166594 224984
rect 166920 224954 166948 225678
rect 166736 224926 166948 224954
rect 166264 223576 166316 223582
rect 166264 223518 166316 223524
rect 166276 223310 166304 223518
rect 166446 223408 166502 223417
rect 166446 223343 166502 223352
rect 166264 223304 166316 223310
rect 166264 223246 166316 223252
rect 166460 223174 166488 223343
rect 166736 223258 166764 224926
rect 166644 223230 166764 223258
rect 166264 223168 166316 223174
rect 166262 223136 166264 223145
rect 166448 223168 166500 223174
rect 166316 223136 166318 223145
rect 166448 223110 166500 223116
rect 166262 223071 166318 223080
rect 166080 223032 166132 223038
rect 166080 222974 166132 222980
rect 165618 222864 165674 222873
rect 165618 222799 165674 222808
rect 166080 222624 166132 222630
rect 166078 222592 166080 222601
rect 166132 222592 166134 222601
rect 166078 222527 166134 222536
rect 165620 218612 165672 218618
rect 165620 218554 165672 218560
rect 165632 218074 165660 218554
rect 166644 218226 166672 223230
rect 166816 223032 166868 223038
rect 166816 222974 166868 222980
rect 166828 222698 166856 222974
rect 166816 222692 166868 222698
rect 166816 222634 166868 222640
rect 167000 222624 167052 222630
rect 166998 222592 167000 222601
rect 167052 222592 167054 222601
rect 166998 222527 167054 222536
rect 166814 222320 166870 222329
rect 167196 222306 167224 231662
rect 168208 230586 168236 231676
rect 168196 230580 168248 230586
rect 168196 230522 168248 230528
rect 167644 229220 167696 229226
rect 167644 229162 167696 229168
rect 166814 222255 166870 222264
rect 167104 222278 167224 222306
rect 166828 218618 166856 222255
rect 167104 222204 167132 222278
rect 167104 222176 167224 222204
rect 167196 220522 167224 222176
rect 167184 220516 167236 220522
rect 167184 220458 167236 220464
rect 167656 220289 167684 229162
rect 168852 227186 168880 231676
rect 169036 231662 169510 231690
rect 169864 231662 170154 231690
rect 170416 231662 170798 231690
rect 171152 231662 171442 231690
rect 168840 227180 168892 227186
rect 168840 227122 168892 227128
rect 169036 225078 169064 231662
rect 169484 227180 169536 227186
rect 169484 227122 169536 227128
rect 169024 225072 169076 225078
rect 169024 225014 169076 225020
rect 169208 225072 169260 225078
rect 169208 225014 169260 225020
rect 168104 223576 168156 223582
rect 168104 223518 168156 223524
rect 168288 223576 168340 223582
rect 168288 223518 168340 223524
rect 168116 223310 168144 223518
rect 168104 223304 168156 223310
rect 168104 223246 168156 223252
rect 168104 222760 168156 222766
rect 168104 222702 168156 222708
rect 168116 222329 168144 222702
rect 168102 222320 168158 222329
rect 168102 222255 168158 222264
rect 167642 220280 167698 220289
rect 167642 220215 167698 220224
rect 166816 218612 166868 218618
rect 166816 218554 166868 218560
rect 167000 218612 167052 218618
rect 167000 218554 167052 218560
rect 166552 218198 166672 218226
rect 166816 218204 166868 218210
rect 166552 218142 166580 218198
rect 166816 218146 166868 218152
rect 166080 218136 166132 218142
rect 166080 218078 166132 218084
rect 166540 218136 166592 218142
rect 166540 218078 166592 218084
rect 165620 218068 165672 218074
rect 165620 218010 165672 218016
rect 166092 217002 166120 218078
rect 166828 217002 166856 218146
rect 167012 218074 167040 218554
rect 168104 218204 168156 218210
rect 168104 218146 168156 218152
rect 167000 218068 167052 218074
rect 167000 218010 167052 218016
rect 167736 218068 167788 218074
rect 167736 218010 167788 218016
rect 167748 217002 167776 218010
rect 159836 216974 159988 217002
rect 160816 216974 161152 217002
rect 161644 216974 161796 217002
rect 162472 216974 162808 217002
rect 163300 216974 163636 217002
rect 164128 216974 164188 217002
rect 164956 216974 165384 217002
rect 165784 216974 166120 217002
rect 166612 216974 166856 217002
rect 167440 216974 167776 217002
rect 168116 217002 168144 218146
rect 168300 218074 168328 223518
rect 169220 219434 169248 225014
rect 169036 219406 169248 219434
rect 169036 219298 169064 219406
rect 169024 219292 169076 219298
rect 169024 219234 169076 219240
rect 169208 219292 169260 219298
rect 169208 219234 169260 219240
rect 169220 218618 169248 219234
rect 169208 218612 169260 218618
rect 169208 218554 169260 218560
rect 168288 218068 168340 218074
rect 168288 218010 168340 218016
rect 169496 217002 169524 227122
rect 169864 225865 169892 231662
rect 169850 225856 169906 225865
rect 169850 225791 169906 225800
rect 170416 223145 170444 231662
rect 171152 229094 171180 231662
rect 171152 229066 171456 229094
rect 171138 228984 171194 228993
rect 170968 228954 171138 228970
rect 170956 228948 171138 228954
rect 171008 228942 171138 228948
rect 171138 228919 171194 228928
rect 170956 228890 171008 228896
rect 171048 226024 171100 226030
rect 170862 225992 170918 226001
rect 171232 226024 171284 226030
rect 171048 225966 171100 225972
rect 171230 225992 171232 226001
rect 171284 225992 171286 226001
rect 170862 225927 170918 225936
rect 170876 225078 170904 225927
rect 171060 225842 171088 225966
rect 171230 225927 171286 225936
rect 171060 225814 171272 225842
rect 171244 225758 171272 225814
rect 171048 225752 171100 225758
rect 171046 225720 171048 225729
rect 171232 225752 171284 225758
rect 171100 225720 171102 225729
rect 171232 225694 171284 225700
rect 171046 225655 171102 225664
rect 170864 225072 170916 225078
rect 171048 225072 171100 225078
rect 170864 225014 170916 225020
rect 171046 225040 171048 225049
rect 171100 225040 171102 225049
rect 171046 224975 171102 224984
rect 170956 224256 171008 224262
rect 170954 224224 170956 224233
rect 171094 224256 171146 224262
rect 171008 224224 171010 224233
rect 171428 224233 171456 229066
rect 171600 228812 171652 228818
rect 171600 228754 171652 228760
rect 171612 228449 171640 228754
rect 172072 228682 172100 231676
rect 172242 228984 172298 228993
rect 172242 228919 172298 228928
rect 172426 228984 172482 228993
rect 172426 228919 172482 228928
rect 172256 228682 172284 228919
rect 172060 228676 172112 228682
rect 172060 228618 172112 228624
rect 172244 228676 172296 228682
rect 172244 228618 172296 228624
rect 171598 228440 171654 228449
rect 171598 228375 171654 228384
rect 171094 224198 171146 224204
rect 171414 224224 171470 224233
rect 170954 224159 171010 224168
rect 171106 224074 171134 224198
rect 171414 224159 171470 224168
rect 170968 224046 171134 224074
rect 170968 223961 170996 224046
rect 170954 223952 171010 223961
rect 170954 223887 171010 223896
rect 170402 223136 170458 223145
rect 170402 223071 170458 223080
rect 171140 222216 171192 222222
rect 171138 222184 171140 222193
rect 171192 222184 171194 222193
rect 171138 222119 171194 222128
rect 171324 222148 171376 222154
rect 171324 222090 171376 222096
rect 171336 222034 171364 222090
rect 171060 222018 171364 222034
rect 171048 222012 171364 222018
rect 171100 222006 171364 222012
rect 171048 221954 171100 221960
rect 170862 221912 170918 221921
rect 170862 221847 170918 221856
rect 171414 221912 171470 221921
rect 171414 221847 171416 221856
rect 170220 218612 170272 218618
rect 170220 218554 170272 218560
rect 170232 217002 170260 218554
rect 170876 218210 170904 221847
rect 171468 221847 171470 221856
rect 171416 221818 171468 221824
rect 171048 220516 171100 220522
rect 171048 220458 171100 220464
rect 170864 218204 170916 218210
rect 170864 218146 170916 218152
rect 171060 217002 171088 220458
rect 172440 219434 172468 228919
rect 172716 220658 172744 231676
rect 172992 231662 173374 231690
rect 173912 231662 174018 231690
rect 172992 222018 173020 231662
rect 173912 228954 173940 231662
rect 174082 228984 174138 228993
rect 173900 228948 173952 228954
rect 174082 228919 174084 228928
rect 173900 228890 173952 228896
rect 174136 228919 174138 228928
rect 174084 228890 174136 228896
rect 174266 228848 174322 228857
rect 174266 228783 174322 228792
rect 172980 222012 173032 222018
rect 172980 221954 173032 221960
rect 172704 220652 172756 220658
rect 172704 220594 172756 220600
rect 174280 219434 174308 228783
rect 174648 227594 174676 231676
rect 175292 229090 175320 231676
rect 175476 231662 175950 231690
rect 175280 229084 175332 229090
rect 175280 229026 175332 229032
rect 174636 227588 174688 227594
rect 174636 227530 174688 227536
rect 175004 227452 175056 227458
rect 175004 227394 175056 227400
rect 175016 222714 175044 227394
rect 175016 222686 175228 222714
rect 174820 222624 174872 222630
rect 174818 222592 174820 222601
rect 175004 222624 175056 222630
rect 174872 222592 174874 222601
rect 175004 222566 175056 222572
rect 174818 222527 174874 222536
rect 172348 219406 172468 219434
rect 174188 219406 174308 219434
rect 171876 218204 171928 218210
rect 171876 218146 171928 218152
rect 171888 217002 171916 218146
rect 168116 216974 168268 217002
rect 169096 216974 169524 217002
rect 169924 216974 170260 217002
rect 170752 216974 171088 217002
rect 171580 216974 171916 217002
rect 172348 217002 172376 219406
rect 174188 218482 174216 219406
rect 174176 218476 174228 218482
rect 174176 218418 174228 218424
rect 174360 218476 174412 218482
rect 174360 218418 174412 218424
rect 174372 218226 174400 218418
rect 174188 218198 174400 218226
rect 174188 218074 174216 218198
rect 173532 218068 173584 218074
rect 173532 218010 173584 218016
rect 174176 218068 174228 218074
rect 174176 218010 174228 218016
rect 174360 218068 174412 218074
rect 174360 218010 174412 218016
rect 173544 217002 173572 218010
rect 174372 217002 174400 218010
rect 175016 217002 175044 222566
rect 175200 218074 175228 222686
rect 175476 222601 175504 231662
rect 176580 229906 176608 231676
rect 176948 231662 177238 231690
rect 177408 231662 177882 231690
rect 178052 231662 178526 231690
rect 176568 229900 176620 229906
rect 176568 229842 176620 229848
rect 175648 229084 175700 229090
rect 175648 229026 175700 229032
rect 175660 228857 175688 229026
rect 175646 228848 175702 228857
rect 175646 228783 175702 228792
rect 176658 226128 176714 226137
rect 176658 226063 176714 226072
rect 176672 225978 176700 226063
rect 176626 225950 176700 225978
rect 176626 225894 176654 225950
rect 176292 225888 176344 225894
rect 175936 225836 176292 225842
rect 175936 225830 176344 225836
rect 176614 225888 176666 225894
rect 176614 225830 176666 225836
rect 176752 225888 176804 225894
rect 176752 225830 176804 225836
rect 175936 225814 176332 225830
rect 175936 225758 175964 225814
rect 175924 225752 175976 225758
rect 175924 225694 175976 225700
rect 176764 225321 176792 225830
rect 176948 225729 176976 231662
rect 176934 225720 176990 225729
rect 176934 225655 176990 225664
rect 176474 225312 176530 225321
rect 176474 225247 176530 225256
rect 176750 225312 176806 225321
rect 176750 225247 176806 225256
rect 175462 222592 175518 222601
rect 175462 222527 175518 222536
rect 176292 222012 176344 222018
rect 176292 221954 176344 221960
rect 176016 218204 176068 218210
rect 176016 218146 176068 218152
rect 175188 218068 175240 218074
rect 175188 218010 175240 218016
rect 176028 217002 176056 218146
rect 176304 218074 176332 221954
rect 176488 218210 176516 225247
rect 177408 222154 177436 231662
rect 177580 229900 177632 229906
rect 177580 229842 177632 229848
rect 177592 224954 177620 229842
rect 177592 224926 177896 224954
rect 177578 222184 177634 222193
rect 177396 222148 177448 222154
rect 177578 222119 177580 222128
rect 177396 222090 177448 222096
rect 177632 222119 177634 222128
rect 177580 222090 177632 222096
rect 177488 220652 177540 220658
rect 177488 220594 177540 220600
rect 177500 219978 177528 220594
rect 177488 219972 177540 219978
rect 177488 219914 177540 219920
rect 177672 219972 177724 219978
rect 177672 219914 177724 219920
rect 176476 218204 176528 218210
rect 176476 218146 176528 218152
rect 176292 218068 176344 218074
rect 176292 218010 176344 218016
rect 176568 218068 176620 218074
rect 176568 218010 176620 218016
rect 176580 217002 176608 218010
rect 177684 217002 177712 219914
rect 177868 218074 177896 224926
rect 178052 221513 178080 231662
rect 179156 229362 179184 231676
rect 179144 229356 179196 229362
rect 179144 229298 179196 229304
rect 179800 228682 179828 231676
rect 179984 231662 180458 231690
rect 180812 231662 181102 231690
rect 179788 228676 179840 228682
rect 179788 228618 179840 228624
rect 179328 227588 179380 227594
rect 179328 227530 179380 227536
rect 178038 221504 178094 221513
rect 178038 221439 178094 221448
rect 178314 221368 178370 221377
rect 178314 221303 178316 221312
rect 178368 221303 178370 221312
rect 178500 221332 178552 221338
rect 178316 221274 178368 221280
rect 178500 221274 178552 221280
rect 177856 218068 177908 218074
rect 177856 218010 177908 218016
rect 178512 217002 178540 221274
rect 179340 217002 179368 227530
rect 179984 222154 180012 231662
rect 180614 228984 180670 228993
rect 180614 228919 180670 228928
rect 179972 222148 180024 222154
rect 179972 222090 180024 222096
rect 180156 222148 180208 222154
rect 180156 222090 180208 222096
rect 180168 221338 180196 222090
rect 180156 221332 180208 221338
rect 180156 221274 180208 221280
rect 180156 218204 180208 218210
rect 180156 218146 180208 218152
rect 180168 217002 180196 218146
rect 172348 216974 172408 217002
rect 173236 216974 173572 217002
rect 174064 216974 174400 217002
rect 174892 216974 175044 217002
rect 175720 216974 176056 217002
rect 176548 216974 176608 217002
rect 177376 216974 177712 217002
rect 178204 216974 178540 217002
rect 179032 216974 179368 217002
rect 179860 216974 180196 217002
rect 180628 217002 180656 228919
rect 180812 226137 180840 231662
rect 181732 230042 181760 231676
rect 181720 230036 181772 230042
rect 181720 229978 181772 229984
rect 182088 229356 182140 229362
rect 182088 229298 182140 229304
rect 181720 229084 181772 229090
rect 181720 229026 181772 229032
rect 181260 228812 181312 228818
rect 181260 228754 181312 228760
rect 181272 228138 181300 228754
rect 181076 228132 181128 228138
rect 181076 228074 181128 228080
rect 181260 228132 181312 228138
rect 181260 228074 181312 228080
rect 181088 227882 181116 228074
rect 181732 228002 181760 229026
rect 181902 228984 181958 228993
rect 181902 228919 181904 228928
rect 181956 228919 181958 228928
rect 181904 228890 181956 228896
rect 181720 227996 181772 228002
rect 181720 227938 181772 227944
rect 181904 227996 181956 228002
rect 181904 227938 181956 227944
rect 181916 227882 181944 227938
rect 181088 227854 181944 227882
rect 180798 226128 180854 226137
rect 180798 226063 180854 226072
rect 181074 226128 181130 226137
rect 181074 226063 181130 226072
rect 181088 225894 181116 226063
rect 181076 225888 181128 225894
rect 181076 225830 181128 225836
rect 181628 225888 181680 225894
rect 181628 225830 181680 225836
rect 181444 225752 181496 225758
rect 181444 225694 181496 225700
rect 181456 225486 181484 225694
rect 181640 225486 181668 225830
rect 181444 225480 181496 225486
rect 181444 225422 181496 225428
rect 181628 225480 181680 225486
rect 181628 225422 181680 225428
rect 181260 224800 181312 224806
rect 181312 224748 181852 224754
rect 181260 224742 181852 224748
rect 181272 224726 181852 224742
rect 181824 224670 181852 224726
rect 181812 224664 181864 224670
rect 181812 224606 181864 224612
rect 181628 223032 181680 223038
rect 181628 222974 181680 222980
rect 181812 223032 181864 223038
rect 181812 222974 181864 222980
rect 181640 222766 181668 222974
rect 181628 222760 181680 222766
rect 181628 222702 181680 222708
rect 181260 222624 181312 222630
rect 181824 222578 181852 222974
rect 181312 222572 181852 222578
rect 181260 222566 181852 222572
rect 181272 222550 181852 222566
rect 181812 222148 181864 222154
rect 181812 222090 181864 222096
rect 181444 222012 181496 222018
rect 181444 221954 181496 221960
rect 181456 221338 181484 221954
rect 181444 221332 181496 221338
rect 181444 221274 181496 221280
rect 180984 219156 181036 219162
rect 180984 219098 181036 219104
rect 180996 218618 181024 219098
rect 180800 218612 180852 218618
rect 180800 218554 180852 218560
rect 180984 218612 181036 218618
rect 180984 218554 181036 218560
rect 180812 218074 180840 218554
rect 180800 218068 180852 218074
rect 180800 218010 180852 218016
rect 181824 217002 181852 222090
rect 182100 218074 182128 229298
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 182652 220658 182680 231662
rect 183284 225888 183336 225894
rect 183284 225830 183336 225836
rect 182640 220652 182692 220658
rect 182640 220594 182692 220600
rect 183296 219298 183324 225830
rect 183664 224534 183692 231676
rect 184308 230178 184336 231676
rect 184296 230172 184348 230178
rect 184296 230114 184348 230120
rect 184204 230036 184256 230042
rect 184204 229978 184256 229984
rect 183652 224528 183704 224534
rect 183652 224470 183704 224476
rect 184020 224528 184072 224534
rect 184020 224470 184072 224476
rect 183468 220652 183520 220658
rect 183468 220594 183520 220600
rect 182640 219292 182692 219298
rect 182640 219234 182692 219240
rect 183284 219292 183336 219298
rect 183284 219234 183336 219240
rect 182088 218068 182140 218074
rect 182088 218010 182140 218016
rect 182652 217002 182680 219234
rect 183480 217002 183508 220594
rect 183652 219292 183704 219298
rect 183652 219234 183704 219240
rect 183664 218482 183692 219234
rect 183652 218476 183704 218482
rect 183652 218418 183704 218424
rect 184032 217002 184060 224470
rect 184216 220658 184244 229978
rect 184952 228002 184980 231676
rect 185136 231662 185610 231690
rect 185780 231662 186254 231690
rect 184940 227996 184992 228002
rect 184940 227938 184992 227944
rect 184572 227724 184624 227730
rect 184572 227666 184624 227672
rect 184584 225758 184612 227666
rect 184572 225752 184624 225758
rect 184572 225694 184624 225700
rect 184846 225720 184902 225729
rect 184846 225655 184902 225664
rect 184204 220652 184256 220658
rect 184204 220594 184256 220600
rect 184388 220652 184440 220658
rect 184388 220594 184440 220600
rect 184400 219978 184428 220594
rect 184388 219972 184440 219978
rect 184388 219914 184440 219920
rect 184860 217002 184888 225655
rect 185136 221377 185164 231662
rect 185584 225480 185636 225486
rect 185584 225422 185636 225428
rect 185596 225185 185624 225422
rect 185582 225176 185638 225185
rect 185582 225111 185638 225120
rect 185780 223310 185808 231662
rect 186134 226128 186190 226137
rect 186134 226063 186190 226072
rect 186148 225978 186176 226063
rect 186412 226024 186464 226030
rect 186410 225992 186412 226001
rect 186596 226024 186648 226030
rect 186464 225992 186466 226001
rect 186148 225950 186314 225978
rect 186286 225894 186314 225950
rect 186596 225966 186648 225972
rect 186410 225927 186466 225936
rect 186136 225888 186188 225894
rect 186136 225830 186188 225836
rect 186274 225888 186326 225894
rect 186608 225842 186636 225966
rect 186274 225830 186326 225836
rect 186148 225457 186176 225830
rect 186424 225814 186636 225842
rect 186424 225729 186452 225814
rect 186410 225720 186466 225729
rect 186410 225655 186466 225664
rect 186134 225448 186190 225457
rect 186134 225383 186190 225392
rect 186884 224262 186912 231676
rect 187528 227730 187556 231676
rect 187896 231662 188186 231690
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 187056 225752 187108 225758
rect 187056 225694 187108 225700
rect 187068 225457 187096 225694
rect 187700 225480 187752 225486
rect 187054 225448 187110 225457
rect 187700 225422 187752 225428
rect 187054 225383 187110 225392
rect 187712 225214 187740 225422
rect 187700 225208 187752 225214
rect 187700 225150 187752 225156
rect 187056 224800 187108 224806
rect 187056 224742 187108 224748
rect 187516 224800 187568 224806
rect 187516 224742 187568 224748
rect 187068 224262 187096 224742
rect 186872 224256 186924 224262
rect 186872 224198 186924 224204
rect 187056 224256 187108 224262
rect 187056 224198 187108 224204
rect 185768 223304 185820 223310
rect 185768 223246 185820 223252
rect 186044 223304 186096 223310
rect 186044 223246 186096 223252
rect 185122 221368 185178 221377
rect 185122 221303 185178 221312
rect 186056 217002 186084 223246
rect 186780 218476 186832 218482
rect 186780 218418 186832 218424
rect 186792 217002 186820 218418
rect 187528 217002 187556 224742
rect 187896 220930 187924 231662
rect 188066 225992 188122 226001
rect 188066 225927 188122 225936
rect 188080 225214 188108 225927
rect 188068 225208 188120 225214
rect 188068 225150 188120 225156
rect 188816 224262 188844 231676
rect 189460 230314 189488 231676
rect 189448 230308 189500 230314
rect 189448 230250 189500 230256
rect 190104 226778 190132 231676
rect 190472 231662 190762 231690
rect 191406 231662 191604 231690
rect 190276 230036 190328 230042
rect 190276 229978 190328 229984
rect 190092 226772 190144 226778
rect 190092 226714 190144 226720
rect 188804 224256 188856 224262
rect 188804 224198 188856 224204
rect 188988 224256 189040 224262
rect 188988 224198 189040 224204
rect 187884 220924 187936 220930
rect 187884 220866 187936 220872
rect 188436 220924 188488 220930
rect 188436 220866 188488 220872
rect 188448 217002 188476 220866
rect 189000 217002 189028 224198
rect 190288 219434 190316 229978
rect 190472 229242 190500 231662
rect 190920 230308 190972 230314
rect 190920 230250 190972 230256
rect 190932 229770 190960 230250
rect 191288 230172 191340 230178
rect 191288 230114 191340 230120
rect 191300 229906 191328 230114
rect 191288 229900 191340 229906
rect 191288 229842 191340 229848
rect 190920 229764 190972 229770
rect 190920 229706 190972 229712
rect 190380 229214 190500 229242
rect 190380 228970 190408 229214
rect 190550 229120 190606 229129
rect 191380 229084 191432 229090
rect 190550 229055 190552 229064
rect 190604 229055 190606 229064
rect 190552 229026 190604 229032
rect 190932 229044 191380 229072
rect 190380 228942 190500 228970
rect 190472 226914 190500 228942
rect 190932 228818 190960 229044
rect 191380 229026 191432 229032
rect 190920 228812 190972 228818
rect 190920 228754 190972 228760
rect 190920 228268 190972 228274
rect 190920 228210 190972 228216
rect 190932 228002 190960 228210
rect 190920 227996 190972 228002
rect 190920 227938 190972 227944
rect 190460 226908 190512 226914
rect 190460 226850 190512 226856
rect 190552 225480 190604 225486
rect 190550 225448 190552 225457
rect 190736 225480 190788 225486
rect 190604 225448 190606 225457
rect 190736 225422 190788 225428
rect 190550 225383 190606 225392
rect 190748 224806 190776 225422
rect 191576 224954 191604 231662
rect 191748 227724 191800 227730
rect 191748 227666 191800 227672
rect 191392 224926 191604 224954
rect 190736 224800 190788 224806
rect 190736 224742 190788 224748
rect 191392 224670 191420 224926
rect 191380 224664 191432 224670
rect 191380 224606 191432 224612
rect 190920 219972 190972 219978
rect 190920 219914 190972 219920
rect 190196 219406 190316 219434
rect 190196 217002 190224 219406
rect 190932 217002 190960 219914
rect 191760 217002 191788 227666
rect 192036 222630 192064 231676
rect 192312 231662 192694 231690
rect 193338 231662 193536 231690
rect 192312 229129 192340 231662
rect 192298 229120 192354 229129
rect 192298 229055 192354 229064
rect 192208 228948 192260 228954
rect 192208 228890 192260 228896
rect 192220 223310 192248 228890
rect 192484 224664 192536 224670
rect 192484 224606 192536 224612
rect 192496 224126 192524 224606
rect 192484 224120 192536 224126
rect 192484 224062 192536 224068
rect 192668 224120 192720 224126
rect 192668 224062 192720 224068
rect 192208 223304 192260 223310
rect 192208 223246 192260 223252
rect 192484 223304 192536 223310
rect 192484 223246 192536 223252
rect 192024 222624 192076 222630
rect 192024 222566 192076 222572
rect 192496 218618 192524 223246
rect 192484 218612 192536 218618
rect 192484 218554 192536 218560
rect 192680 217002 192708 224062
rect 193508 219842 193536 231662
rect 193968 224398 193996 231676
rect 194612 229090 194640 231676
rect 194888 231662 195270 231690
rect 195532 231662 195914 231690
rect 194600 229084 194652 229090
rect 194600 229026 194652 229032
rect 194888 225457 194916 231662
rect 194874 225448 194930 225457
rect 194874 225383 194930 225392
rect 195532 225185 195560 231662
rect 195704 229084 195756 229090
rect 195704 229026 195756 229032
rect 195518 225176 195574 225185
rect 195518 225111 195574 225120
rect 195716 224954 195744 229026
rect 195888 226772 195940 226778
rect 195888 226714 195940 226720
rect 195900 225214 195928 226714
rect 195888 225208 195940 225214
rect 195888 225150 195940 225156
rect 195716 224926 195836 224954
rect 195808 224890 195836 224926
rect 195808 224862 195928 224890
rect 194324 224800 194376 224806
rect 194324 224742 194376 224748
rect 193956 224392 194008 224398
rect 193956 224334 194008 224340
rect 194140 224392 194192 224398
rect 194140 224334 194192 224340
rect 194152 224126 194180 224334
rect 194140 224120 194192 224126
rect 194140 224062 194192 224068
rect 193496 219836 193548 219842
rect 193496 219778 193548 219784
rect 193128 218612 193180 218618
rect 193128 218554 193180 218560
rect 193140 217002 193168 218554
rect 194336 217002 194364 224742
rect 194508 224664 194560 224670
rect 194508 224606 194560 224612
rect 195704 224664 195756 224670
rect 195704 224606 195756 224612
rect 194520 224126 194548 224606
rect 194508 224120 194560 224126
rect 194508 224062 194560 224068
rect 195244 221332 195296 221338
rect 195244 221274 195296 221280
rect 195428 221332 195480 221338
rect 195428 221274 195480 221280
rect 195256 221066 195284 221274
rect 195060 221060 195112 221066
rect 195060 221002 195112 221008
rect 195244 221060 195296 221066
rect 195244 221002 195296 221008
rect 194874 220824 194930 220833
rect 195072 220794 195100 221002
rect 195440 220930 195468 221274
rect 195428 220924 195480 220930
rect 195428 220866 195480 220872
rect 194874 220759 194876 220768
rect 194928 220759 194930 220768
rect 195060 220788 195112 220794
rect 194876 220730 194928 220736
rect 195060 220730 195112 220736
rect 194876 218068 194928 218074
rect 194876 218010 194928 218016
rect 194888 217002 194916 218010
rect 195716 217002 195744 224606
rect 195900 218074 195928 224862
rect 196544 224126 196572 231676
rect 196992 230308 197044 230314
rect 196992 230250 197044 230256
rect 196532 224120 196584 224126
rect 196532 224062 196584 224068
rect 196072 223304 196124 223310
rect 196072 223246 196124 223252
rect 196084 222766 196112 223246
rect 196072 222760 196124 222766
rect 196072 222702 196124 222708
rect 196070 220824 196126 220833
rect 196070 220759 196072 220768
rect 196124 220759 196126 220768
rect 196072 220730 196124 220736
rect 197004 219434 197032 230250
rect 197188 229498 197216 231676
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 198936 231662 199134 231690
rect 199304 231662 199778 231690
rect 197176 229492 197228 229498
rect 197176 229434 197228 229440
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197832 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 197832 220794 197860 229066
rect 198004 227996 198056 228002
rect 198004 227938 198056 227944
rect 197820 220788 197872 220794
rect 197820 220730 197872 220736
rect 197268 219836 197320 219842
rect 197268 219778 197320 219784
rect 196820 219406 197032 219434
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196820 217002 196848 219406
rect 197280 217002 197308 219778
rect 198016 219434 198044 227938
rect 198936 220930 198964 231662
rect 199304 226778 199332 231662
rect 200408 227866 200436 231676
rect 201052 228138 201080 231676
rect 201040 228132 201092 228138
rect 201040 228074 201092 228080
rect 201408 228132 201460 228138
rect 201408 228074 201460 228080
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 226908 200080 226914
rect 200028 226850 200080 226856
rect 199292 226772 199344 226778
rect 199292 226714 199344 226720
rect 199384 225208 199436 225214
rect 199384 225150 199436 225156
rect 198924 220924 198976 220930
rect 198924 220866 198976 220872
rect 198372 220788 198424 220794
rect 198372 220730 198424 220736
rect 198004 219428 198056 219434
rect 198004 219370 198056 219376
rect 198384 217002 198412 220730
rect 199396 219162 199424 225150
rect 199844 219428 199896 219434
rect 199844 219370 199896 219376
rect 199384 219156 199436 219162
rect 199384 219098 199436 219104
rect 198924 218068 198976 218074
rect 198924 218010 198976 218016
rect 198936 217002 198964 218010
rect 199856 217002 199884 219370
rect 200040 218074 200068 226850
rect 201224 224120 201276 224126
rect 201224 224062 201276 224068
rect 200028 218068 200080 218074
rect 200028 218010 200080 218016
rect 200856 218068 200908 218074
rect 200856 218010 200908 218016
rect 200868 217002 200896 218010
rect 180628 216974 180688 217002
rect 181516 216974 181852 217002
rect 182344 216974 182680 217002
rect 183172 216974 183508 217002
rect 184000 216974 184060 217002
rect 184828 216974 184888 217002
rect 185656 216974 186084 217002
rect 186484 216974 186820 217002
rect 187312 216974 187556 217002
rect 188140 216974 188476 217002
rect 188968 216974 189028 217002
rect 189796 216974 190224 217002
rect 190624 216974 190960 217002
rect 191452 216974 191788 217002
rect 192280 216974 192708 217002
rect 193108 216974 193168 217002
rect 193936 216974 194364 217002
rect 194764 216974 194916 217002
rect 195592 216974 195744 217002
rect 196420 216974 196848 217002
rect 197248 216974 197308 217002
rect 198076 216974 198412 217002
rect 198904 216974 198964 217002
rect 199732 216974 199884 217002
rect 200560 216974 200896 217002
rect 201236 217002 201264 224062
rect 201420 218074 201448 228074
rect 201696 223718 201724 231676
rect 202340 230178 202368 231676
rect 202328 230172 202380 230178
rect 202328 230114 202380 230120
rect 202984 225350 203012 231676
rect 203168 231662 203642 231690
rect 202972 225344 203024 225350
rect 202972 225286 203024 225292
rect 202602 225176 202658 225185
rect 202602 225111 202658 225120
rect 201684 223712 201736 223718
rect 201684 223654 201736 223660
rect 201408 218068 201460 218074
rect 201408 218010 201460 218016
rect 202616 217002 202644 225111
rect 203168 221354 203196 231662
rect 203892 229492 203944 229498
rect 203892 229434 203944 229440
rect 203708 222760 203760 222766
rect 203708 222702 203760 222708
rect 203522 222456 203578 222465
rect 203522 222391 203578 222400
rect 203536 222290 203564 222391
rect 203720 222358 203748 222702
rect 203708 222352 203760 222358
rect 203708 222294 203760 222300
rect 203524 222284 203576 222290
rect 203524 222226 203576 222232
rect 203076 221326 203196 221354
rect 203076 219570 203104 221326
rect 203248 221196 203300 221202
rect 203248 221138 203300 221144
rect 203260 220930 203288 221138
rect 203248 220924 203300 220930
rect 203248 220866 203300 220872
rect 203248 220244 203300 220250
rect 203248 220186 203300 220192
rect 203260 219570 203288 220186
rect 203064 219564 203116 219570
rect 203064 219506 203116 219512
rect 203248 219564 203300 219570
rect 203248 219506 203300 219512
rect 203904 218074 203932 229434
rect 204076 225616 204128 225622
rect 204076 225558 204128 225564
rect 204088 225350 204116 225558
rect 204076 225344 204128 225350
rect 204076 225286 204128 225292
rect 204272 223854 204300 231676
rect 204916 229094 204944 231676
rect 204548 229066 204944 229094
rect 205192 231662 205574 231690
rect 205836 231662 206218 231690
rect 206480 231662 206862 231690
rect 204548 228002 204576 229066
rect 204720 228540 204772 228546
rect 204720 228482 204772 228488
rect 204904 228540 204956 228546
rect 204904 228482 204956 228488
rect 204536 227996 204588 228002
rect 204536 227938 204588 227944
rect 204732 227866 204760 228482
rect 204916 228274 204944 228482
rect 204904 228268 204956 228274
rect 204904 228210 204956 228216
rect 204720 227860 204772 227866
rect 204720 227802 204772 227808
rect 205192 226506 205220 231662
rect 205364 230308 205416 230314
rect 205364 230250 205416 230256
rect 205376 229498 205404 230250
rect 205364 229492 205416 229498
rect 205364 229434 205416 229440
rect 205456 228132 205508 228138
rect 205456 228074 205508 228080
rect 205180 226500 205232 226506
rect 205180 226442 205232 226448
rect 204904 225616 204956 225622
rect 204904 225558 204956 225564
rect 204916 225214 204944 225558
rect 204904 225208 204956 225214
rect 205088 225208 205140 225214
rect 204904 225150 204956 225156
rect 205086 225176 205088 225185
rect 205140 225176 205142 225185
rect 205086 225111 205142 225120
rect 204732 224454 205128 224482
rect 204732 224126 204760 224454
rect 205100 224398 205128 224454
rect 204904 224392 204956 224398
rect 204904 224334 204956 224340
rect 205088 224392 205140 224398
rect 205088 224334 205140 224340
rect 204916 224126 204944 224334
rect 204720 224120 204772 224126
rect 204720 224062 204772 224068
rect 204904 224120 204956 224126
rect 204904 224062 204956 224068
rect 204260 223848 204312 223854
rect 204260 223790 204312 223796
rect 205272 223848 205324 223854
rect 205272 223790 205324 223796
rect 204076 223304 204128 223310
rect 204076 223246 204128 223252
rect 203340 218068 203392 218074
rect 203340 218010 203392 218016
rect 203892 218068 203944 218074
rect 203892 218010 203944 218016
rect 203352 217002 203380 218010
rect 204088 217002 204116 223246
rect 205088 222624 205140 222630
rect 205088 222566 205140 222572
rect 205100 222465 205128 222566
rect 205086 222456 205142 222465
rect 205086 222391 205142 222400
rect 204904 221604 204956 221610
rect 204904 221546 204956 221552
rect 205088 221604 205140 221610
rect 205088 221546 205140 221552
rect 204916 221066 204944 221546
rect 205100 221202 205128 221546
rect 205088 221196 205140 221202
rect 205088 221138 205140 221144
rect 204904 221060 204956 221066
rect 204904 221002 204956 221008
rect 205284 219434 205312 223790
rect 204720 219428 204772 219434
rect 204720 219370 204772 219376
rect 204916 219406 205312 219434
rect 204732 219162 204760 219370
rect 204720 219156 204772 219162
rect 204720 219098 204772 219104
rect 204916 219026 204944 219406
rect 204904 219020 204956 219026
rect 204904 218962 204956 218968
rect 204996 218068 205048 218074
rect 204996 218010 205048 218016
rect 205008 217002 205036 218010
rect 201236 216974 201388 217002
rect 202216 216974 202644 217002
rect 203044 216974 203380 217002
rect 203872 216974 204116 217002
rect 204700 216974 205036 217002
rect 205468 217002 205496 228074
rect 205836 219570 205864 231662
rect 206008 221196 206060 221202
rect 206008 221138 206060 221144
rect 205824 219564 205876 219570
rect 205824 219506 205876 219512
rect 206020 218074 206048 221138
rect 206480 220930 206508 231662
rect 207492 222358 207520 231676
rect 207768 231662 208150 231690
rect 207768 225350 207796 231662
rect 207756 225344 207808 225350
rect 207756 225286 207808 225292
rect 208124 225344 208176 225350
rect 208124 225286 208176 225292
rect 207480 222352 207532 222358
rect 207480 222294 207532 222300
rect 206468 220924 206520 220930
rect 206468 220866 206520 220872
rect 207480 219836 207532 219842
rect 207480 219778 207532 219784
rect 206652 219020 206704 219026
rect 206652 218962 206704 218968
rect 206008 218068 206060 218074
rect 206008 218010 206060 218016
rect 206664 217002 206692 218962
rect 207492 217002 207520 219778
rect 208136 217002 208164 225286
rect 208780 222630 208808 231676
rect 209424 224942 209452 231676
rect 210068 229634 210096 231676
rect 210056 229628 210108 229634
rect 210056 229570 210108 229576
rect 210240 229628 210292 229634
rect 210240 229570 210292 229576
rect 209412 224936 209464 224942
rect 209412 224878 209464 224884
rect 209688 224936 209740 224942
rect 209688 224878 209740 224884
rect 208768 222624 208820 222630
rect 208768 222566 208820 222572
rect 209504 222624 209556 222630
rect 209504 222566 209556 222572
rect 209136 218068 209188 218074
rect 209136 218010 209188 218016
rect 209148 217002 209176 218010
rect 205468 216974 205528 217002
rect 206356 216974 206692 217002
rect 207184 216974 207520 217002
rect 208012 216974 208164 217002
rect 208840 216974 209176 217002
rect 209516 217002 209544 222566
rect 209700 218074 209728 224878
rect 210252 222630 210280 229570
rect 210712 227866 210740 231676
rect 210700 227860 210752 227866
rect 210700 227802 210752 227808
rect 210240 222624 210292 222630
rect 210240 222566 210292 222572
rect 210884 222624 210936 222630
rect 210884 222566 210936 222572
rect 209688 218068 209740 218074
rect 209688 218010 209740 218016
rect 210896 217002 210924 222566
rect 211356 220250 211384 231676
rect 211632 231662 212014 231690
rect 211632 221066 211660 231662
rect 212644 229094 212672 231676
rect 212644 229066 212856 229094
rect 212632 228812 212684 228818
rect 212632 228754 212684 228760
rect 212644 228546 212672 228754
rect 212632 228540 212684 228546
rect 212632 228482 212684 228488
rect 212172 228404 212224 228410
rect 212172 228346 212224 228352
rect 212184 228002 212212 228346
rect 212172 227996 212224 228002
rect 212172 227938 212224 227944
rect 212356 226772 212408 226778
rect 212356 226714 212408 226720
rect 212172 222896 212224 222902
rect 212172 222838 212224 222844
rect 212184 222358 212212 222838
rect 212172 222352 212224 222358
rect 212172 222294 212224 222300
rect 211988 221468 212040 221474
rect 211988 221410 212040 221416
rect 212000 221066 212028 221410
rect 211620 221060 211672 221066
rect 211620 221002 211672 221008
rect 211988 221060 212040 221066
rect 211988 221002 212040 221008
rect 211344 220244 211396 220250
rect 211344 220186 211396 220192
rect 211620 220244 211672 220250
rect 211620 220186 211672 220192
rect 211632 217002 211660 220186
rect 212368 219434 212396 226714
rect 212828 223854 212856 229066
rect 213288 227050 213316 231676
rect 213946 231662 214144 231690
rect 213276 227044 213328 227050
rect 213276 226986 213328 226992
rect 213184 226500 213236 226506
rect 213184 226442 213236 226448
rect 212816 223848 212868 223854
rect 212816 223790 212868 223796
rect 212276 219406 212396 219434
rect 213000 219428 213052 219434
rect 212276 217002 212304 219406
rect 213000 219370 213052 219376
rect 213012 218346 213040 219370
rect 213196 218754 213224 226442
rect 213828 222760 213880 222766
rect 213828 222702 213880 222708
rect 213184 218748 213236 218754
rect 213184 218690 213236 218696
rect 213000 218340 213052 218346
rect 213000 218282 213052 218288
rect 213276 218340 213328 218346
rect 213276 218282 213328 218288
rect 213288 217002 213316 218282
rect 213840 217002 213868 222702
rect 214116 219706 214144 231662
rect 214300 231662 214590 231690
rect 214300 221066 214328 231662
rect 215220 230450 215248 231676
rect 215208 230444 215260 230450
rect 215208 230386 215260 230392
rect 215864 226166 215892 231676
rect 216232 231662 216522 231690
rect 215852 226160 215904 226166
rect 215852 226102 215904 226108
rect 215944 223848 215996 223854
rect 215944 223790 215996 223796
rect 214932 221604 214984 221610
rect 214932 221546 214984 221552
rect 214288 221060 214340 221066
rect 214288 221002 214340 221008
rect 214104 219700 214156 219706
rect 214104 219642 214156 219648
rect 214944 217002 214972 221546
rect 215956 218890 215984 223790
rect 216232 222358 216260 231662
rect 217152 229094 217180 231676
rect 217060 229066 217180 229094
rect 216496 226160 216548 226166
rect 216496 226102 216548 226108
rect 216220 222352 216272 222358
rect 216220 222294 216272 222300
rect 215944 218884 215996 218890
rect 215944 218826 215996 218832
rect 216312 218884 216364 218890
rect 216312 218826 216364 218832
rect 215760 218068 215812 218074
rect 215760 218010 215812 218016
rect 215772 217002 215800 218010
rect 216324 217002 216352 218826
rect 216508 218074 216536 226102
rect 217060 223990 217088 229066
rect 217796 226506 217824 231676
rect 218440 228002 218468 231676
rect 218624 231662 219098 231690
rect 218428 227996 218480 228002
rect 218428 227938 218480 227944
rect 217784 226500 217836 226506
rect 217784 226442 217836 226448
rect 217048 223984 217100 223990
rect 217048 223926 217100 223932
rect 217232 223984 217284 223990
rect 217232 223926 217284 223932
rect 217244 219434 217272 223926
rect 218624 220386 218652 231662
rect 219164 228812 219216 228818
rect 219164 228754 219216 228760
rect 218612 220380 218664 220386
rect 218612 220322 218664 220328
rect 217416 219700 217468 219706
rect 217416 219642 217468 219648
rect 217232 219428 217284 219434
rect 217232 219370 217284 219376
rect 216680 218340 216732 218346
rect 216680 218282 216732 218288
rect 216692 218074 216720 218282
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 216680 218068 216732 218074
rect 216680 218010 216732 218016
rect 217428 217002 217456 219642
rect 217968 219428 218020 219434
rect 217968 219370 218020 219376
rect 217980 217002 218008 219370
rect 219176 217002 219204 228754
rect 219728 222494 219756 231676
rect 220372 229226 220400 231676
rect 220360 229220 220412 229226
rect 220360 229162 220412 229168
rect 221016 226370 221044 231676
rect 221004 226364 221056 226370
rect 221004 226306 221056 226312
rect 221660 222902 221688 231676
rect 222016 226636 222068 226642
rect 222016 226578 222068 226584
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221648 222896 221700 222902
rect 221648 222838 221700 222844
rect 219716 222488 219768 222494
rect 219716 222430 219768 222436
rect 220084 222488 220136 222494
rect 220084 222430 220136 222436
rect 220096 219434 220124 222430
rect 220728 222352 220780 222358
rect 220728 222294 220780 222300
rect 220084 219428 220136 219434
rect 220084 219370 220136 219376
rect 219900 218748 219952 218754
rect 219900 218690 219952 218696
rect 219912 217002 219940 218690
rect 220740 217002 220768 222294
rect 221844 219434 221872 226442
rect 221660 219406 221872 219434
rect 221660 217002 221688 219406
rect 209516 216974 209668 217002
rect 210496 216974 210924 217002
rect 211324 216974 211660 217002
rect 212152 216974 212304 217002
rect 212980 216974 213316 217002
rect 213808 216974 213868 217002
rect 214636 216974 214972 217002
rect 215464 216974 215800 217002
rect 216292 216974 216352 217002
rect 217120 216974 217456 217002
rect 217948 216974 218008 217002
rect 218776 216974 219204 217002
rect 219604 216974 219940 217002
rect 220432 216974 220768 217002
rect 221260 216974 221688 217002
rect 222028 217002 222056 226578
rect 222304 223174 222332 231676
rect 222752 228404 222804 228410
rect 222752 228346 222804 228352
rect 222764 228002 222792 228346
rect 222752 227996 222804 228002
rect 222752 227938 222804 227944
rect 222476 226296 222528 226302
rect 222476 226238 222528 226244
rect 222488 225622 222516 226238
rect 222476 225616 222528 225622
rect 222476 225558 222528 225564
rect 222948 223854 222976 231676
rect 223396 230444 223448 230450
rect 223396 230386 223448 230392
rect 222936 223848 222988 223854
rect 222936 223790 222988 223796
rect 222292 223168 222344 223174
rect 222292 223110 222344 223116
rect 223408 219434 223436 230386
rect 223592 225078 223620 231676
rect 224040 228812 224092 228818
rect 224040 228754 224092 228760
rect 224052 228410 224080 228754
rect 224040 228404 224092 228410
rect 224040 228346 224092 228352
rect 224236 226114 224264 231676
rect 224052 226086 224264 226114
rect 224420 231662 224894 231690
rect 223580 225072 223632 225078
rect 223580 225014 223632 225020
rect 224052 223446 224080 226086
rect 224224 226024 224276 226030
rect 224224 225966 224276 225972
rect 224236 225622 224264 225966
rect 224224 225616 224276 225622
rect 224224 225558 224276 225564
rect 224040 223440 224092 223446
rect 224040 223382 224092 223388
rect 224224 223168 224276 223174
rect 224224 223110 224276 223116
rect 223316 219406 223436 219434
rect 224040 219428 224092 219434
rect 223316 217002 223344 219406
rect 224040 219370 224092 219376
rect 224052 218890 224080 219370
rect 224040 218884 224092 218890
rect 224040 218826 224092 218832
rect 224236 218346 224264 223110
rect 224420 221746 224448 231662
rect 225524 226302 225552 231676
rect 225696 228404 225748 228410
rect 225696 228346 225748 228352
rect 225512 226296 225564 226302
rect 225512 226238 225564 226244
rect 224684 225072 224736 225078
rect 224684 225014 224736 225020
rect 224408 221740 224460 221746
rect 224408 221682 224460 221688
rect 224224 218340 224276 218346
rect 224224 218282 224276 218288
rect 224696 218210 224724 225014
rect 225708 219434 225736 228346
rect 226168 228002 226196 231676
rect 226156 227996 226208 228002
rect 226156 227938 226208 227944
rect 226156 227860 226208 227866
rect 226156 227802 226208 227808
rect 225524 219406 225736 219434
rect 225524 218210 225552 219406
rect 225972 218884 226024 218890
rect 225972 218826 226024 218832
rect 224040 218204 224092 218210
rect 224040 218146 224092 218152
rect 224684 218204 224736 218210
rect 224684 218146 224736 218152
rect 224868 218204 224920 218210
rect 224868 218146 224920 218152
rect 225512 218204 225564 218210
rect 225512 218146 225564 218152
rect 225696 218204 225748 218210
rect 225696 218146 225748 218152
rect 224052 217002 224080 218146
rect 224880 217002 224908 218146
rect 225708 217002 225736 218146
rect 222028 216974 222088 217002
rect 222916 216974 223344 217002
rect 223744 216974 224080 217002
rect 224572 216974 224908 217002
rect 225400 216974 225736 217002
rect 225984 217002 226012 218826
rect 226168 218210 226196 227802
rect 226812 223582 226840 231676
rect 227456 227322 227484 231676
rect 227444 227316 227496 227322
rect 227444 227258 227496 227264
rect 226984 227044 227036 227050
rect 226984 226986 227036 226992
rect 226800 223576 226852 223582
rect 226800 223518 226852 223524
rect 226996 219298 227024 226986
rect 228100 223990 228128 231676
rect 228744 227186 228772 231676
rect 229296 231662 229402 231690
rect 229664 231662 230046 231690
rect 228732 227180 228784 227186
rect 228732 227122 228784 227128
rect 229054 227044 229106 227050
rect 229054 226986 229106 226992
rect 229066 226930 229094 226986
rect 229020 226902 229094 226930
rect 229020 226506 229048 226902
rect 229008 226500 229060 226506
rect 229008 226442 229060 226448
rect 228916 226296 228968 226302
rect 228916 226238 228968 226244
rect 228088 223984 228140 223990
rect 228088 223926 228140 223932
rect 227352 221060 227404 221066
rect 227352 221002 227404 221008
rect 226984 219292 227036 219298
rect 226984 219234 227036 219240
rect 226156 218204 226208 218210
rect 226156 218146 226208 218152
rect 227364 217002 227392 221002
rect 228180 218340 228232 218346
rect 228180 218282 228232 218288
rect 228192 217002 228220 218282
rect 228928 217002 228956 226238
rect 229296 220522 229324 231662
rect 229664 221882 229692 231662
rect 230676 229362 230704 231676
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230664 229356 230716 229362
rect 230664 229298 230716 229304
rect 229652 221876 229704 221882
rect 229652 221818 229704 221824
rect 230388 221740 230440 221746
rect 230388 221682 230440 221688
rect 229284 220516 229336 220522
rect 229284 220458 229336 220464
rect 229192 220380 229244 220386
rect 229192 220322 229244 220328
rect 229204 218346 229232 220322
rect 229192 218340 229244 218346
rect 229192 218282 229244 218288
rect 229836 218204 229888 218210
rect 229836 218146 229888 218152
rect 229848 217002 229876 218146
rect 230400 217002 230428 221682
rect 231136 218210 231164 229434
rect 231320 228818 231348 231676
rect 231308 228812 231360 228818
rect 231308 228754 231360 228760
rect 231964 227458 231992 231676
rect 232148 231662 232622 231690
rect 231952 227452 232004 227458
rect 231952 227394 232004 227400
rect 231584 223984 231636 223990
rect 231584 223926 231636 223932
rect 231124 218204 231176 218210
rect 231124 218146 231176 218152
rect 231596 217002 231624 223926
rect 232148 221474 232176 231662
rect 233252 227322 233280 231676
rect 233240 227316 233292 227322
rect 233240 227258 233292 227264
rect 232504 226500 232556 226506
rect 232504 226442 232556 226448
rect 232136 221468 232188 221474
rect 232136 221410 232188 221416
rect 232516 219434 232544 226442
rect 233896 226030 233924 231676
rect 234080 231662 234554 231690
rect 234816 231662 235198 231690
rect 233884 226024 233936 226030
rect 233884 225966 233936 225972
rect 233700 224528 233752 224534
rect 233700 224470 233752 224476
rect 233884 224528 233936 224534
rect 233884 224470 233936 224476
rect 233712 223854 233740 224470
rect 233896 224126 233924 224470
rect 233884 224120 233936 224126
rect 233884 224062 233936 224068
rect 233700 223848 233752 223854
rect 233700 223790 233752 223796
rect 233148 222896 233200 222902
rect 233148 222838 233200 222844
rect 232504 219428 232556 219434
rect 232504 219370 232556 219376
rect 232964 219428 233016 219434
rect 232964 219370 233016 219376
rect 232320 218204 232372 218210
rect 232320 218146 232372 218152
rect 232332 217002 232360 218146
rect 232976 217002 233004 219370
rect 233160 218210 233188 222838
rect 234080 220658 234108 231662
rect 234528 227316 234580 227322
rect 234528 227258 234580 227264
rect 234344 225616 234396 225622
rect 234344 225558 234396 225564
rect 234068 220652 234120 220658
rect 234068 220594 234120 220600
rect 233148 218204 233200 218210
rect 233148 218146 233200 218152
rect 233976 218204 234028 218210
rect 233976 218146 234028 218152
rect 233988 217002 234016 218146
rect 225984 216974 226228 217002
rect 227056 216974 227392 217002
rect 227884 216974 228220 217002
rect 228712 216974 228956 217002
rect 229540 216974 229876 217002
rect 230368 216974 230428 217002
rect 231196 216974 231624 217002
rect 232024 216974 232360 217002
rect 232852 216974 233004 217002
rect 233680 216974 234016 217002
rect 234356 217002 234384 225558
rect 234540 218210 234568 227258
rect 234816 223038 234844 231662
rect 235828 229770 235856 231676
rect 235816 229764 235868 229770
rect 235816 229706 235868 229712
rect 236472 227594 236500 231676
rect 236920 229764 236972 229770
rect 236920 229706 236972 229712
rect 236932 229094 236960 229706
rect 237116 229094 237144 231676
rect 237392 231662 237774 231690
rect 236932 229066 237052 229094
rect 237116 229066 237236 229094
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 235724 227180 235776 227186
rect 235724 227122 235776 227128
rect 234804 223032 234856 223038
rect 234804 222974 234856 222980
rect 235264 223032 235316 223038
rect 235264 222974 235316 222980
rect 235276 218482 235304 222974
rect 235264 218476 235316 218482
rect 235264 218418 235316 218424
rect 234528 218204 234580 218210
rect 234528 218146 234580 218152
rect 235736 217002 235764 227122
rect 237024 218210 237052 229066
rect 237208 228682 237236 229066
rect 237196 228676 237248 228682
rect 237196 228618 237248 228624
rect 237392 222018 237420 231662
rect 238404 223174 238432 231676
rect 239048 225894 239076 231676
rect 239404 228676 239456 228682
rect 239404 228618 239456 228624
rect 239036 225888 239088 225894
rect 239036 225830 239088 225836
rect 238668 223984 238720 223990
rect 238668 223926 238720 223932
rect 238392 223168 238444 223174
rect 238392 223110 238444 223116
rect 237380 222012 237432 222018
rect 237380 221954 237432 221960
rect 237288 221876 237340 221882
rect 237288 221818 237340 221824
rect 236460 218204 236512 218210
rect 236460 218146 236512 218152
rect 237012 218204 237064 218210
rect 237012 218146 237064 218152
rect 236472 217002 236500 218146
rect 237300 217002 237328 221818
rect 238116 219292 238168 219298
rect 238116 219234 238168 219240
rect 238128 217002 238156 219234
rect 238680 217002 238708 223926
rect 239416 219298 239444 228618
rect 239692 223854 239720 231676
rect 240152 231662 240350 231690
rect 239680 223848 239732 223854
rect 239680 223790 239732 223796
rect 240152 222154 240180 231662
rect 240980 229906 241008 231676
rect 240968 229900 241020 229906
rect 240968 229842 241020 229848
rect 241624 228954 241652 231676
rect 241612 228948 241664 228954
rect 241612 228890 241664 228896
rect 242268 225486 242296 231676
rect 242532 227792 242584 227798
rect 242532 227734 242584 227740
rect 242256 225480 242308 225486
rect 242256 225422 242308 225428
rect 240140 222148 240192 222154
rect 240140 222090 240192 222096
rect 241244 221468 241296 221474
rect 241244 221410 241296 221416
rect 240600 220516 240652 220522
rect 240600 220458 240652 220464
rect 239404 219292 239456 219298
rect 239404 219234 239456 219240
rect 239772 218476 239824 218482
rect 239772 218418 239824 218424
rect 239784 217002 239812 218418
rect 240612 217002 240640 220458
rect 241256 217002 241284 221410
rect 242256 218068 242308 218074
rect 242256 218010 242308 218016
rect 242268 217002 242296 218010
rect 234356 216974 234508 217002
rect 235336 216974 235764 217002
rect 236164 216974 236500 217002
rect 236992 216974 237328 217002
rect 237820 216974 238156 217002
rect 238648 216974 238708 217002
rect 239476 216974 239812 217002
rect 240304 216974 240640 217002
rect 241132 216974 241284 217002
rect 241960 216974 242296 217002
rect 242544 217002 242572 227734
rect 242912 225758 242940 231676
rect 243280 231662 243570 231690
rect 243832 231662 244214 231690
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 242900 225752 242952 225758
rect 242900 225694 242952 225700
rect 242716 223848 242768 223854
rect 242716 223790 242768 223796
rect 242728 218074 242756 223790
rect 243280 223038 243308 231662
rect 243544 226024 243596 226030
rect 243544 225966 243596 225972
rect 243268 223032 243320 223038
rect 243268 222974 243320 222980
rect 243556 218618 243584 225966
rect 243832 224262 243860 231662
rect 243820 224256 243872 224262
rect 243820 224198 243872 224204
rect 243912 222012 243964 222018
rect 243912 221954 243964 221960
rect 243544 218612 243596 218618
rect 243544 218554 243596 218560
rect 242716 218068 242768 218074
rect 242716 218010 242768 218016
rect 243924 217002 243952 221954
rect 244476 220114 244504 231662
rect 245120 221338 245148 231662
rect 246132 230042 246160 231676
rect 246120 230036 246172 230042
rect 246120 229978 246172 229984
rect 245660 229900 245712 229906
rect 245660 229842 245712 229848
rect 245672 227798 245700 229842
rect 246212 228812 246264 228818
rect 246212 228754 246264 228760
rect 245660 227792 245712 227798
rect 245660 227734 245712 227740
rect 245568 223168 245620 223174
rect 245568 223110 245620 223116
rect 245108 221332 245160 221338
rect 245108 221274 245160 221280
rect 244464 220108 244516 220114
rect 244464 220050 244516 220056
rect 244740 218068 244792 218074
rect 244740 218010 244792 218016
rect 244752 217002 244780 218010
rect 245580 217002 245608 223110
rect 246224 219162 246252 228754
rect 246776 224534 246804 231676
rect 247420 224806 247448 231676
rect 248064 227662 248092 231676
rect 248052 227656 248104 227662
rect 248052 227598 248104 227604
rect 248144 227452 248196 227458
rect 248144 227394 248196 227400
rect 247408 224800 247460 224806
rect 247408 224742 247460 224748
rect 246764 224528 246816 224534
rect 246764 224470 246816 224476
rect 247684 224528 247736 224534
rect 247684 224470 247736 224476
rect 246948 224256 247000 224262
rect 246948 224198 247000 224204
rect 246396 219428 246448 219434
rect 246396 219370 246448 219376
rect 246212 219156 246264 219162
rect 246212 219098 246264 219104
rect 246408 217002 246436 219370
rect 246960 217002 246988 224198
rect 247696 218074 247724 224470
rect 247684 218068 247736 218074
rect 247684 218010 247736 218016
rect 248156 217002 248184 227394
rect 248708 226030 248736 231676
rect 248892 231662 249366 231690
rect 249904 231662 250010 231690
rect 248696 226024 248748 226030
rect 248696 225966 248748 225972
rect 248892 224670 248920 231662
rect 249708 225888 249760 225894
rect 249708 225830 249760 225836
rect 248880 224664 248932 224670
rect 248880 224606 248932 224612
rect 249064 224664 249116 224670
rect 249064 224606 249116 224612
rect 249076 218210 249104 224606
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249524 218204 249576 218210
rect 249524 218146 249576 218152
rect 248880 218068 248932 218074
rect 248880 218010 248932 218016
rect 248892 217002 248920 218010
rect 249536 217002 249564 218146
rect 249720 218074 249748 225830
rect 249904 219978 249932 231662
rect 250640 229090 250668 231676
rect 251284 230178 251312 231676
rect 251272 230172 251324 230178
rect 251272 230114 251324 230120
rect 251732 230036 251784 230042
rect 251732 229978 251784 229984
rect 251744 229094 251772 229978
rect 251928 229094 251956 231676
rect 250628 229084 250680 229090
rect 251744 229066 251864 229094
rect 251928 229066 252048 229094
rect 250628 229026 250680 229032
rect 251088 228948 251140 228954
rect 251088 228890 251140 228896
rect 250904 223032 250956 223038
rect 250904 222974 250956 222980
rect 249892 219972 249944 219978
rect 249892 219914 249944 219920
rect 249708 218068 249760 218074
rect 249708 218010 249760 218016
rect 250536 218068 250588 218074
rect 250536 218010 250588 218016
rect 250548 217002 250576 218010
rect 242544 216974 242788 217002
rect 243616 216974 243952 217002
rect 244444 216974 244780 217002
rect 245272 216974 245608 217002
rect 246100 216974 246436 217002
rect 246928 216974 246988 217002
rect 247756 216974 248184 217002
rect 248584 216974 248920 217002
rect 249412 216974 249564 217002
rect 250240 216974 250576 217002
rect 250916 217002 250944 222974
rect 251100 218074 251128 228890
rect 251836 218210 251864 229066
rect 252020 226914 252048 229066
rect 252572 228274 252600 231676
rect 252756 231662 253230 231690
rect 252560 228268 252612 228274
rect 252560 228210 252612 228216
rect 252284 227588 252336 227594
rect 252284 227530 252336 227536
rect 252008 226908 252060 226914
rect 252008 226850 252060 226856
rect 251824 218204 251876 218210
rect 251824 218146 251876 218152
rect 251088 218068 251140 218074
rect 251088 218010 251140 218016
rect 252296 217002 252324 227530
rect 252756 220794 252784 231662
rect 253860 228818 253888 231676
rect 253848 228812 253900 228818
rect 253848 228754 253900 228760
rect 254504 225214 254532 231676
rect 254872 231662 255162 231690
rect 254492 225208 254544 225214
rect 254492 225150 254544 225156
rect 254872 223310 254900 231662
rect 255044 228812 255096 228818
rect 255044 228754 255096 228760
rect 254860 223304 254912 223310
rect 254860 223246 254912 223252
rect 252744 220788 252796 220794
rect 252744 220730 252796 220736
rect 253848 220652 253900 220658
rect 253848 220594 253900 220600
rect 253020 218612 253072 218618
rect 253020 218554 253072 218560
rect 253032 217002 253060 218554
rect 253860 217002 253888 220594
rect 254676 220108 254728 220114
rect 254676 220050 254728 220056
rect 254688 217002 254716 220050
rect 250916 216974 251068 217002
rect 251896 216974 252324 217002
rect 252724 216974 253060 217002
rect 253552 216974 253888 217002
rect 254380 216974 254716 217002
rect 255056 217002 255084 228754
rect 255792 224398 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 257080 228138 257108 231676
rect 257264 231662 257738 231690
rect 258092 231662 258382 231690
rect 257264 229094 257292 231662
rect 257264 229066 257384 229094
rect 257068 228132 257120 228138
rect 257068 228074 257120 228080
rect 255964 227792 256016 227798
rect 255964 227734 256016 227740
rect 255780 224392 255832 224398
rect 255780 224334 255832 224340
rect 255976 219026 256004 227734
rect 256332 222148 256384 222154
rect 256332 222090 256384 222096
rect 255964 219020 256016 219026
rect 255964 218962 256016 218968
rect 256344 217002 256372 222090
rect 257160 220788 257212 220794
rect 257160 220730 257212 220736
rect 257172 217002 257200 220730
rect 257356 219842 257384 229066
rect 257804 225752 257856 225758
rect 257804 225694 257856 225700
rect 257344 219836 257396 219842
rect 257344 219778 257396 219784
rect 257816 217002 257844 225694
rect 258092 221202 258120 231662
rect 259012 227798 259040 231676
rect 259276 229084 259328 229090
rect 259276 229026 259328 229032
rect 259000 227792 259052 227798
rect 259000 227734 259052 227740
rect 258080 221196 258132 221202
rect 258080 221138 258132 221144
rect 259092 219020 259144 219026
rect 259092 218962 259144 218968
rect 258816 218068 258868 218074
rect 258816 218010 258868 218016
rect 258828 217002 258856 218010
rect 255056 216974 255208 217002
rect 256036 216974 256372 217002
rect 256864 216974 257200 217002
rect 257692 216974 257844 217002
rect 258520 216974 258856 217002
rect 259104 217002 259132 218962
rect 259288 218074 259316 229026
rect 259656 224942 259684 231676
rect 259644 224936 259696 224942
rect 259644 224878 259696 224884
rect 260300 222630 260328 231676
rect 260944 225350 260972 231676
rect 261392 230308 261444 230314
rect 261392 230250 261444 230256
rect 261404 229094 261432 230250
rect 261588 229634 261616 231676
rect 261576 229628 261628 229634
rect 261576 229570 261628 229576
rect 261220 229066 261432 229094
rect 260932 225344 260984 225350
rect 260932 225286 260984 225292
rect 260564 223440 260616 223446
rect 260564 223382 260616 223388
rect 260288 222624 260340 222630
rect 260288 222566 260340 222572
rect 259276 218068 259328 218074
rect 259276 218010 259328 218016
rect 260576 217002 260604 223382
rect 261220 222154 261248 229066
rect 262232 226778 262260 231676
rect 262220 226772 262272 226778
rect 262220 226714 262272 226720
rect 262128 224392 262180 224398
rect 262128 224334 262180 224340
rect 261208 222148 261260 222154
rect 261208 222090 261260 222096
rect 261392 222148 261444 222154
rect 261392 222090 261444 222096
rect 261404 217002 261432 222090
rect 262140 217002 262168 224334
rect 262876 222766 262904 231676
rect 263060 231662 263534 231690
rect 263888 231662 264178 231690
rect 262864 222760 262916 222766
rect 262864 222702 262916 222708
rect 263060 220250 263088 231662
rect 263888 224670 263916 231662
rect 264808 226166 264836 231676
rect 265176 231662 265466 231690
rect 265728 231662 266110 231690
rect 264796 226160 264848 226166
rect 264796 226102 264848 226108
rect 264244 224936 264296 224942
rect 264244 224878 264296 224884
rect 263876 224664 263928 224670
rect 263876 224606 263928 224612
rect 263508 222760 263560 222766
rect 263508 222702 263560 222708
rect 263048 220244 263100 220250
rect 263048 220186 263100 220192
rect 263324 220244 263376 220250
rect 263324 220186 263376 220192
rect 262680 219156 262732 219162
rect 262680 219098 262732 219104
rect 262692 218618 262720 219098
rect 262680 218612 262732 218618
rect 262680 218554 262732 218560
rect 262956 218068 263008 218074
rect 262956 218010 263008 218016
rect 262968 217002 262996 218010
rect 259104 216974 259348 217002
rect 260176 216974 260604 217002
rect 261004 216974 261432 217002
rect 261832 216974 262168 217002
rect 262660 216974 262996 217002
rect 263336 217002 263364 220186
rect 263520 218074 263548 222702
rect 264256 218754 264284 224878
rect 264704 223304 264756 223310
rect 264704 223246 264756 223252
rect 264244 218748 264296 218754
rect 264244 218690 264296 218696
rect 263508 218068 263560 218074
rect 263508 218010 263560 218016
rect 264716 217002 264744 223246
rect 265176 219706 265204 231662
rect 265728 221610 265756 231662
rect 266740 226506 266768 231676
rect 267384 228546 267412 231676
rect 267372 228540 267424 228546
rect 267372 228482 267424 228488
rect 267556 228540 267608 228546
rect 267556 228482 267608 228488
rect 266728 226500 266780 226506
rect 266728 226442 266780 226448
rect 266268 226160 266320 226166
rect 267568 226114 267596 228482
rect 266268 226102 266320 226108
rect 265716 221604 265768 221610
rect 265716 221546 265768 221552
rect 265164 219700 265216 219706
rect 265164 219642 265216 219648
rect 266084 218748 266136 218754
rect 266084 218690 266136 218696
rect 265440 218068 265492 218074
rect 265440 218010 265492 218016
rect 265452 217002 265480 218010
rect 266096 217002 266124 218690
rect 266280 218074 266308 226102
rect 267384 226086 267596 226114
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 267096 218068 267148 218074
rect 267096 218010 267148 218016
rect 267108 217002 267136 218010
rect 263336 216974 263488 217002
rect 264316 216974 264744 217002
rect 265144 216974 265480 217002
rect 265972 216974 266124 217002
rect 266800 216974 267136 217002
rect 267384 217002 267412 226086
rect 267556 226024 267608 226030
rect 267556 225966 267608 225972
rect 267568 218074 267596 225966
rect 268028 222358 268056 231676
rect 268672 222494 268700 231676
rect 269316 224942 269344 231676
rect 269960 226642 269988 231676
rect 270316 227724 270368 227730
rect 270316 227666 270368 227672
rect 269948 226636 270000 226642
rect 269948 226578 270000 226584
rect 269304 224936 269356 224942
rect 269304 224878 269356 224884
rect 268844 223576 268896 223582
rect 268844 223518 268896 223524
rect 268660 222488 268712 222494
rect 268660 222430 268712 222436
rect 268016 222352 268068 222358
rect 268016 222294 268068 222300
rect 267740 221604 267792 221610
rect 267740 221546 267792 221552
rect 267752 218618 267780 221546
rect 267740 218612 267792 218618
rect 267740 218554 267792 218560
rect 267556 218068 267608 218074
rect 267556 218010 267608 218016
rect 268856 217002 268884 223518
rect 269580 218068 269632 218074
rect 269580 218010 269632 218016
rect 269592 217002 269620 218010
rect 270328 217002 270356 227666
rect 270604 225078 270632 231676
rect 271248 227050 271276 231676
rect 271892 230450 271920 231676
rect 271880 230444 271932 230450
rect 271880 230386 271932 230392
rect 272536 228002 272564 231676
rect 272720 231662 273194 231690
rect 272524 227996 272576 228002
rect 272524 227938 272576 227944
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 225072 270644 225078
rect 270592 225014 270644 225020
rect 271328 224664 271380 224670
rect 271328 224606 271380 224612
rect 271340 217002 271368 224606
rect 271800 217002 271828 226986
rect 272524 226908 272576 226914
rect 272524 226850 272576 226856
rect 272536 218482 272564 226850
rect 272720 221066 272748 231662
rect 273824 228410 273852 231676
rect 274008 231662 274482 231690
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274008 221610 274036 231662
rect 274180 230444 274232 230450
rect 274180 230386 274232 230392
rect 273996 221604 274048 221610
rect 273996 221546 274048 221552
rect 273720 221332 273772 221338
rect 273720 221274 273772 221280
rect 272708 221060 272760 221066
rect 272708 221002 272760 221008
rect 273076 219632 273128 219638
rect 273076 219574 273128 219580
rect 273088 219298 273116 219574
rect 273076 219292 273128 219298
rect 273076 219234 273128 219240
rect 272892 218612 272944 218618
rect 272892 218554 272944 218560
rect 272524 218476 272576 218482
rect 272524 218418 272576 218424
rect 272904 217002 272932 218554
rect 273732 217002 273760 221274
rect 274192 219434 274220 230386
rect 275112 226302 275140 231676
rect 275388 231662 275770 231690
rect 276124 231662 276414 231690
rect 275388 229094 275416 231662
rect 275296 229066 275416 229094
rect 275100 226296 275152 226302
rect 275100 226238 275152 226244
rect 275296 221898 275324 229066
rect 275652 225004 275704 225010
rect 275652 224946 275704 224952
rect 275204 221870 275324 221898
rect 275204 221746 275232 221870
rect 275192 221740 275244 221746
rect 275192 221682 275244 221688
rect 275376 221740 275428 221746
rect 275376 221682 275428 221688
rect 273916 219406 274220 219434
rect 273916 218074 273944 219406
rect 274548 218884 274600 218890
rect 274548 218826 274600 218832
rect 273904 218068 273956 218074
rect 273904 218010 273956 218016
rect 274560 217002 274588 218826
rect 275388 217002 275416 221682
rect 267384 216974 267628 217002
rect 268456 216974 268884 217002
rect 269284 216974 269620 217002
rect 270112 216974 270356 217002
rect 270940 216974 271368 217002
rect 271768 216974 271828 217002
rect 272596 216974 272932 217002
rect 273424 216974 273760 217002
rect 274252 216974 274588 217002
rect 275080 216974 275416 217002
rect 275664 217002 275692 224946
rect 276124 220386 276152 231662
rect 276848 230172 276900 230178
rect 276848 230114 276900 230120
rect 276860 225010 276888 230114
rect 277044 229498 277072 231676
rect 277032 229492 277084 229498
rect 277032 229434 277084 229440
rect 277124 228268 277176 228274
rect 277124 228210 277176 228216
rect 276848 225004 276900 225010
rect 276848 224946 276900 224952
rect 276112 220380 276164 220386
rect 276112 220322 276164 220328
rect 277136 217002 277164 228210
rect 277688 222902 277716 231676
rect 278332 227322 278360 231676
rect 278320 227316 278372 227322
rect 278320 227258 278372 227264
rect 278412 226296 278464 226302
rect 278412 226238 278464 226244
rect 277676 222896 277728 222902
rect 277676 222838 277728 222844
rect 278228 221604 278280 221610
rect 278228 221546 278280 221552
rect 277860 218068 277912 218074
rect 277860 218010 277912 218016
rect 277872 217002 277900 218010
rect 275664 216974 275908 217002
rect 276736 216974 277164 217002
rect 277564 216974 277900 217002
rect 278240 217002 278268 221546
rect 278424 218074 278452 226238
rect 278976 224126 279004 231676
rect 279252 231662 279634 231690
rect 278964 224120 279016 224126
rect 278964 224062 279016 224068
rect 279252 219638 279280 231662
rect 280264 227186 280292 231676
rect 280448 231662 280922 231690
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 280448 221882 280476 231662
rect 280804 227316 280856 227322
rect 280804 227258 280856 227264
rect 280436 221876 280488 221882
rect 280436 221818 280488 221824
rect 280068 219972 280120 219978
rect 280068 219914 280120 219920
rect 279240 219632 279292 219638
rect 279240 219574 279292 219580
rect 279516 218476 279568 218482
rect 279516 218418 279568 218424
rect 278412 218068 278464 218074
rect 278412 218010 278464 218016
rect 279528 217002 279556 218418
rect 280080 217002 280108 219914
rect 280816 218890 280844 227258
rect 281552 225622 281580 231676
rect 282196 229770 282224 231676
rect 282184 229764 282236 229770
rect 282184 229706 282236 229712
rect 282840 229094 282868 231676
rect 282472 229066 282868 229094
rect 283024 231662 283498 231690
rect 281540 225616 281592 225622
rect 281540 225558 281592 225564
rect 282472 223990 282500 229066
rect 282828 225004 282880 225010
rect 282828 224946 282880 224952
rect 282644 224800 282696 224806
rect 282644 224742 282696 224748
rect 282460 223984 282512 223990
rect 282460 223926 282512 223932
rect 281172 220380 281224 220386
rect 281172 220322 281224 220328
rect 280804 218884 280856 218890
rect 280804 218826 280856 218832
rect 280988 218884 281040 218890
rect 280988 218826 281040 218832
rect 281000 218482 281028 218826
rect 280988 218476 281040 218482
rect 280988 218418 281040 218424
rect 281184 217002 281212 220322
rect 282656 218074 282684 224742
rect 282000 218068 282052 218074
rect 282000 218010 282052 218016
rect 282644 218068 282696 218074
rect 282644 218010 282696 218016
rect 282012 217002 282040 218010
rect 282840 217002 282868 224946
rect 283024 220522 283052 231662
rect 284128 228682 284156 231676
rect 284116 228676 284168 228682
rect 284116 228618 284168 228624
rect 283932 228404 283984 228410
rect 283932 228346 283984 228352
rect 283012 220516 283064 220522
rect 283012 220458 283064 220464
rect 283656 218068 283708 218074
rect 283656 218010 283708 218016
rect 283668 217002 283696 218010
rect 278240 216974 278392 217002
rect 279220 216974 279556 217002
rect 280048 216974 280108 217002
rect 280876 216974 281212 217002
rect 281704 216974 282040 217002
rect 282532 216974 282868 217002
rect 283360 216974 283696 217002
rect 283944 217002 283972 228346
rect 284772 226914 284800 231676
rect 285048 231662 285430 231690
rect 285692 231662 286074 231690
rect 286336 231662 286718 231690
rect 284760 226908 284812 226914
rect 284760 226850 284812 226856
rect 285048 223854 285076 231662
rect 285312 229764 285364 229770
rect 285312 229706 285364 229712
rect 285324 225010 285352 229706
rect 285496 225616 285548 225622
rect 285496 225558 285548 225564
rect 285312 225004 285364 225010
rect 285312 224946 285364 224952
rect 285036 223848 285088 223854
rect 285036 223790 285088 223796
rect 284116 222896 284168 222902
rect 284116 222838 284168 222844
rect 284128 218074 284156 222838
rect 285508 219434 285536 225558
rect 285692 222018 285720 231662
rect 285680 222012 285732 222018
rect 285680 221954 285732 221960
rect 286336 221882 286364 231662
rect 287348 229906 287376 231676
rect 287624 231662 288006 231690
rect 287336 229900 287388 229906
rect 287336 229842 287388 229848
rect 286968 224120 287020 224126
rect 286968 224062 287020 224068
rect 285680 221876 285732 221882
rect 285680 221818 285732 221824
rect 286324 221876 286376 221882
rect 286324 221818 286376 221824
rect 285692 221474 285720 221818
rect 285680 221468 285732 221474
rect 285680 221410 285732 221416
rect 286048 221468 286100 221474
rect 286048 221410 286100 221416
rect 286060 219434 286088 221410
rect 285416 219406 285536 219434
rect 286048 219428 286100 219434
rect 284116 218068 284168 218074
rect 284116 218010 284168 218016
rect 285416 217002 285444 219406
rect 286048 219370 286100 219376
rect 286140 218476 286192 218482
rect 286140 218418 286192 218424
rect 286152 217002 286180 218418
rect 286980 217002 287008 224062
rect 287624 223174 287652 231662
rect 288072 228132 288124 228138
rect 288072 228074 288124 228080
rect 287612 223168 287664 223174
rect 287612 223110 287664 223116
rect 287796 218068 287848 218074
rect 287796 218010 287848 218016
rect 287808 217002 287836 218010
rect 283944 216974 284188 217002
rect 285016 216974 285444 217002
rect 285844 216974 286180 217002
rect 286672 216974 287008 217002
rect 287500 216974 287836 217002
rect 288084 217002 288112 228074
rect 288256 224936 288308 224942
rect 288256 224878 288308 224884
rect 288268 218074 288296 224878
rect 288636 224262 288664 231676
rect 289280 224534 289308 231676
rect 289268 224528 289320 224534
rect 289268 224470 289320 224476
rect 288624 224256 288676 224262
rect 288624 224198 288676 224204
rect 289544 224256 289596 224262
rect 289544 224198 289596 224204
rect 288256 218068 288308 218074
rect 288256 218010 288308 218016
rect 289556 217002 289584 224198
rect 289924 221474 289952 231676
rect 290568 225894 290596 231676
rect 291212 228954 291240 231676
rect 291200 228948 291252 228954
rect 291200 228890 291252 228896
rect 291856 227458 291884 231676
rect 292500 230042 292528 231676
rect 292488 230036 292540 230042
rect 292488 229978 292540 229984
rect 292396 228676 292448 228682
rect 292396 228618 292448 228624
rect 291844 227452 291896 227458
rect 291844 227394 291896 227400
rect 291844 226432 291896 226438
rect 291844 226374 291896 226380
rect 290556 225888 290608 225894
rect 290556 225830 290608 225836
rect 291108 223168 291160 223174
rect 291108 223110 291160 223116
rect 289912 221468 289964 221474
rect 289912 221410 289964 221416
rect 290280 221468 290332 221474
rect 290280 221410 290332 221416
rect 290292 217002 290320 221410
rect 291120 217002 291148 223110
rect 291660 219428 291712 219434
rect 291660 219370 291712 219376
rect 291672 217002 291700 219370
rect 291856 219162 291884 226374
rect 291844 219156 291896 219162
rect 291844 219098 291896 219104
rect 288084 216974 288328 217002
rect 289156 216974 289584 217002
rect 289984 216974 290320 217002
rect 290812 216974 291148 217002
rect 291640 216974 291700 217002
rect 292408 217002 292436 228618
rect 293144 227594 293172 231676
rect 293420 231662 293802 231690
rect 293132 227588 293184 227594
rect 293132 227530 293184 227536
rect 293420 220658 293448 231662
rect 293684 227452 293736 227458
rect 293684 227394 293736 227400
rect 293408 220652 293460 220658
rect 293408 220594 293460 220600
rect 293696 217002 293724 227394
rect 294432 223038 294460 231676
rect 295076 226438 295104 231676
rect 295720 228818 295748 231676
rect 295904 231662 296378 231690
rect 296824 231662 297022 231690
rect 295708 228812 295760 228818
rect 295708 228754 295760 228760
rect 295064 226432 295116 226438
rect 295064 226374 295116 226380
rect 295248 225888 295300 225894
rect 295248 225830 295300 225836
rect 294420 223032 294472 223038
rect 294420 222974 294472 222980
rect 293868 219836 293920 219842
rect 293868 219778 293920 219784
rect 293880 219026 293908 219778
rect 293868 219020 293920 219026
rect 293868 218962 293920 218968
rect 294420 219020 294472 219026
rect 294420 218962 294472 218968
rect 294432 217002 294460 218962
rect 295260 217002 295288 225830
rect 295904 220794 295932 231662
rect 296168 227180 296220 227186
rect 296168 227122 296220 227128
rect 295892 220788 295944 220794
rect 295892 220730 295944 220736
rect 296180 217002 296208 227122
rect 296628 220516 296680 220522
rect 296628 220458 296680 220464
rect 296640 217002 296668 220458
rect 296824 220114 296852 231662
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 296996 230036 297048 230042
rect 296996 229978 297048 229984
rect 297008 222766 297036 229978
rect 298296 229090 298324 231676
rect 298284 229084 298336 229090
rect 298284 229026 298336 229032
rect 297824 223576 297876 223582
rect 297824 223518 297876 223524
rect 296996 222760 297048 222766
rect 296996 222702 297048 222708
rect 296996 220652 297048 220658
rect 296996 220594 297048 220600
rect 296812 220108 296864 220114
rect 296812 220050 296864 220056
rect 297008 218618 297036 220594
rect 296996 218612 297048 218618
rect 296996 218554 297048 218560
rect 297836 217002 297864 223518
rect 298940 223446 298968 231676
rect 299204 227588 299256 227594
rect 299204 227530 299256 227536
rect 298928 223440 298980 223446
rect 298928 223382 298980 223388
rect 299216 218074 299244 227530
rect 299584 225758 299612 231676
rect 299952 231662 300242 231690
rect 299572 225752 299624 225758
rect 299572 225694 299624 225700
rect 299952 219842 299980 231662
rect 300124 229900 300176 229906
rect 300124 229842 300176 229848
rect 300136 223582 300164 229842
rect 300872 224398 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 302528 231662 302818 231690
rect 300860 224392 300912 224398
rect 300860 224334 300912 224340
rect 300124 223576 300176 223582
rect 300124 223518 300176 223524
rect 300308 223032 300360 223038
rect 300308 222974 300360 222980
rect 300124 220108 300176 220114
rect 300124 220050 300176 220056
rect 299940 219836 299992 219842
rect 299940 219778 299992 219784
rect 298560 218068 298612 218074
rect 298560 218010 298612 218016
rect 299204 218068 299256 218074
rect 299204 218010 299256 218016
rect 299388 218068 299440 218074
rect 299388 218010 299440 218016
rect 298572 217002 298600 218010
rect 299400 217002 299428 218010
rect 300136 217002 300164 220050
rect 300320 218074 300348 222974
rect 301056 220250 301084 231662
rect 301700 222154 301728 231662
rect 302528 230042 302556 231662
rect 302884 230308 302936 230314
rect 302884 230250 302936 230256
rect 302516 230036 302568 230042
rect 302516 229978 302568 229984
rect 301964 223440 302016 223446
rect 301964 223382 302016 223388
rect 301688 222148 301740 222154
rect 301688 222090 301740 222096
rect 301044 220244 301096 220250
rect 301044 220186 301096 220192
rect 300768 219020 300820 219026
rect 300768 218962 300820 218968
rect 300308 218068 300360 218074
rect 300308 218010 300360 218016
rect 300780 217002 300808 218962
rect 301976 217002 302004 223382
rect 302896 218754 302924 230250
rect 303448 226166 303476 231676
rect 303436 226160 303488 226166
rect 303436 226102 303488 226108
rect 304092 226030 304120 231676
rect 304080 226024 304132 226030
rect 304080 225966 304132 225972
rect 303436 224392 303488 224398
rect 303436 224334 303488 224340
rect 302884 218748 302936 218754
rect 302884 218690 302936 218696
rect 302700 218204 302752 218210
rect 302700 218146 302752 218152
rect 302712 217002 302740 218146
rect 303448 217002 303476 224334
rect 304736 223310 304764 231676
rect 305380 230314 305408 231676
rect 305368 230308 305420 230314
rect 305368 230250 305420 230256
rect 305644 230036 305696 230042
rect 305644 229978 305696 229984
rect 304908 225752 304960 225758
rect 304908 225694 304960 225700
rect 304724 223304 304776 223310
rect 304724 223246 304776 223252
rect 304724 221876 304776 221882
rect 304724 221818 304776 221824
rect 304736 218210 304764 221818
rect 304724 218204 304776 218210
rect 304724 218146 304776 218152
rect 304356 218068 304408 218074
rect 304356 218010 304408 218016
rect 304368 217002 304396 218010
rect 304920 217002 304948 225694
rect 305656 218074 305684 229978
rect 306024 223582 306052 231676
rect 306668 227730 306696 231676
rect 307312 228546 307340 231676
rect 307956 230450 307984 231676
rect 307944 230444 307996 230450
rect 307944 230386 307996 230392
rect 307852 230308 307904 230314
rect 307852 230250 307904 230256
rect 307300 228540 307352 228546
rect 307300 228482 307352 228488
rect 307668 228540 307720 228546
rect 307668 228482 307720 228488
rect 306656 227724 306708 227730
rect 306656 227666 306708 227672
rect 306012 223576 306064 223582
rect 306012 223518 306064 223524
rect 306104 223304 306156 223310
rect 306104 223246 306156 223252
rect 305644 218068 305696 218074
rect 305644 218010 305696 218016
rect 306116 217002 306144 223246
rect 306380 220788 306432 220794
rect 306380 220730 306432 220736
rect 306392 218482 306420 220730
rect 307484 218748 307536 218754
rect 307484 218690 307536 218696
rect 306380 218476 306432 218482
rect 306380 218418 306432 218424
rect 306840 218068 306892 218074
rect 306840 218010 306892 218016
rect 306852 217002 306880 218010
rect 307496 217002 307524 218690
rect 307680 218074 307708 228482
rect 307864 224262 307892 230250
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308588 226908 308640 226914
rect 308588 226850 308640 226856
rect 307852 224256 307904 224262
rect 307852 224198 307904 224204
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308600 217002 308628 226850
rect 308956 224256 309008 224262
rect 308956 224198 309008 224204
rect 292408 216974 292468 217002
rect 293296 216974 293724 217002
rect 294124 216974 294460 217002
rect 294952 216974 295288 217002
rect 295780 216974 296208 217002
rect 296608 216974 296668 217002
rect 297436 216974 297864 217002
rect 298264 216974 298600 217002
rect 299092 216974 299428 217002
rect 299920 216974 300164 217002
rect 300748 216974 300808 217002
rect 301576 216974 302004 217002
rect 302404 216974 302740 217002
rect 303232 216974 303476 217002
rect 304060 216974 304396 217002
rect 304888 216974 304948 217002
rect 305716 216974 306144 217002
rect 306544 216974 306880 217002
rect 307372 216974 307524 217002
rect 308200 216974 308628 217002
rect 308968 217002 308996 224198
rect 309244 221338 309272 231676
rect 309888 224670 309916 231676
rect 310546 231662 310744 231690
rect 309876 224664 309928 224670
rect 309876 224606 309928 224612
rect 310152 222012 310204 222018
rect 310152 221954 310204 221960
rect 309232 221332 309284 221338
rect 309232 221274 309284 221280
rect 310164 217002 310192 221954
rect 310716 220658 310744 231662
rect 310900 231662 311190 231690
rect 310900 221746 310928 231662
rect 311820 228274 311848 231676
rect 312096 231662 312478 231690
rect 311808 228268 311860 228274
rect 311808 228210 311860 228216
rect 312096 227322 312124 231662
rect 312544 230444 312596 230450
rect 312544 230386 312596 230392
rect 312084 227316 312136 227322
rect 312084 227258 312136 227264
rect 310888 221740 310940 221746
rect 310888 221682 310940 221688
rect 311532 221740 311584 221746
rect 311532 221682 311584 221688
rect 310704 220652 310756 220658
rect 310704 220594 310756 220600
rect 310980 218204 311032 218210
rect 310980 218146 311032 218152
rect 310992 217002 311020 218146
rect 311544 217002 311572 221682
rect 311716 220652 311768 220658
rect 311716 220594 311768 220600
rect 311728 219162 311756 220594
rect 311716 219156 311768 219162
rect 311716 219098 311768 219104
rect 312556 218890 312584 230386
rect 313108 230178 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230172 313148 230178
rect 313096 230114 313148 230120
rect 313096 226024 313148 226030
rect 313096 225966 313148 225972
rect 312544 218884 312596 218890
rect 312544 218826 312596 218832
rect 312636 218068 312688 218074
rect 312636 218010 312688 218016
rect 312648 217002 312676 218010
rect 308968 216974 309028 217002
rect 309856 216974 310192 217002
rect 310684 216974 311020 217002
rect 311512 216974 311572 217002
rect 312340 216974 312676 217002
rect 313108 217002 313136 225966
rect 313292 221610 313320 231662
rect 313280 221604 313332 221610
rect 313280 221546 313332 221552
rect 313936 219978 313964 231662
rect 315040 226302 315068 231676
rect 315684 230450 315712 231676
rect 315672 230444 315724 230450
rect 315672 230386 315724 230392
rect 315304 230172 315356 230178
rect 315304 230114 315356 230120
rect 315028 226296 315080 226302
rect 315028 226238 315080 226244
rect 314568 221604 314620 221610
rect 314568 221546 314620 221552
rect 313924 219972 313976 219978
rect 313924 219914 313976 219920
rect 314292 218884 314344 218890
rect 314292 218826 314344 218832
rect 314304 217002 314332 218826
rect 314580 218074 314608 221546
rect 315316 218210 315344 230114
rect 316328 224806 316356 231676
rect 316972 229094 317000 231676
rect 316696 229066 317000 229094
rect 317524 231662 317630 231690
rect 316316 224800 316368 224806
rect 316316 224742 316368 224748
rect 315856 224664 315908 224670
rect 315856 224606 315908 224612
rect 315672 219156 315724 219162
rect 315672 219098 315724 219104
rect 315304 218204 315356 218210
rect 315304 218146 315356 218152
rect 314568 218068 314620 218074
rect 314568 218010 314620 218016
rect 315120 218068 315172 218074
rect 315120 218010 315172 218016
rect 315132 217002 315160 218010
rect 315684 217002 315712 219098
rect 315868 218074 315896 224606
rect 316696 222902 316724 229066
rect 317328 226296 317380 226302
rect 317328 226238 317380 226244
rect 316684 222896 316736 222902
rect 316684 222838 316736 222844
rect 316868 222896 316920 222902
rect 316868 222838 316920 222844
rect 315856 218068 315908 218074
rect 315856 218010 315908 218016
rect 316880 217002 316908 222838
rect 317340 217002 317368 226238
rect 317524 220386 317552 231662
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 318064 228812 318116 228818
rect 318064 228754 318116 228760
rect 317512 220380 317564 220386
rect 317512 220322 317564 220328
rect 318076 219162 318104 228754
rect 318904 225622 318932 231676
rect 318892 225616 318944 225622
rect 318892 225558 318944 225564
rect 319548 224126 319576 231676
rect 319812 228948 319864 228954
rect 319812 228890 319864 228896
rect 319536 224120 319588 224126
rect 319536 224062 319588 224068
rect 318432 220244 318484 220250
rect 318432 220186 318484 220192
rect 318064 219156 318116 219162
rect 318064 219098 318116 219104
rect 318444 217002 318472 220186
rect 319260 218068 319312 218074
rect 319260 218010 319312 218016
rect 319272 217002 319300 218010
rect 319824 217002 319852 228890
rect 320192 228410 320220 231676
rect 320376 231662 320850 231690
rect 320180 228404 320232 228410
rect 320180 228346 320232 228352
rect 319996 224528 320048 224534
rect 319996 224470 320048 224476
rect 320008 218074 320036 224470
rect 320376 220794 320404 231662
rect 321480 228138 321508 231676
rect 321756 231662 322138 231690
rect 322400 231662 322782 231690
rect 321468 228132 321520 228138
rect 321468 228074 321520 228080
rect 321376 227724 321428 227730
rect 321376 227666 321428 227672
rect 320364 220788 320416 220794
rect 320364 220730 320416 220736
rect 320916 219156 320968 219162
rect 320916 219098 320968 219104
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 320928 217002 320956 219098
rect 313108 216974 313168 217002
rect 313996 216974 314332 217002
rect 314824 216974 315160 217002
rect 315652 216974 315712 217002
rect 316480 216974 316908 217002
rect 317308 216974 317368 217002
rect 318136 216974 318472 217002
rect 318964 216974 319300 217002
rect 319792 216974 319852 217002
rect 320620 216974 320956 217002
rect 321388 217002 321416 227666
rect 321756 221474 321784 231662
rect 322400 224942 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322664 225616 322716 225622
rect 322664 225558 322716 225564
rect 322388 224936 322440 224942
rect 322388 224878 322440 224884
rect 321744 221468 321796 221474
rect 321744 221410 321796 221416
rect 322676 217002 322704 225558
rect 323688 223174 323716 231662
rect 324044 229764 324096 229770
rect 324044 229706 324096 229712
rect 323676 223168 323728 223174
rect 323676 223110 323728 223116
rect 323400 220380 323452 220386
rect 323400 220322 323452 220328
rect 323412 217002 323440 220322
rect 324056 217002 324084 229706
rect 324700 219434 324728 231676
rect 325344 227458 325372 231676
rect 325332 227452 325384 227458
rect 325332 227394 325384 227400
rect 325608 226160 325660 226166
rect 325608 226102 325660 226108
rect 324688 219428 324740 219434
rect 324688 219370 324740 219376
rect 325424 219292 325476 219298
rect 325424 219234 325476 219240
rect 325056 218068 325108 218074
rect 325056 218010 325108 218016
rect 325068 217002 325096 218010
rect 321388 216974 321448 217002
rect 322276 216974 322704 217002
rect 323104 216974 323440 217002
rect 323932 216974 324084 217002
rect 324760 216974 325096 217002
rect 325436 217002 325464 219234
rect 325620 218074 325648 226102
rect 325988 225894 326016 231676
rect 326632 228682 326660 231676
rect 326620 228676 326672 228682
rect 326620 228618 326672 228624
rect 326804 228404 326856 228410
rect 326804 228346 326856 228352
rect 326344 227316 326396 227322
rect 326344 227258 326396 227264
rect 325976 225888 326028 225894
rect 325976 225830 326028 225836
rect 326356 219298 326384 227258
rect 326344 219292 326396 219298
rect 326344 219234 326396 219240
rect 325608 218068 325660 218074
rect 325608 218010 325660 218016
rect 326816 217002 326844 228346
rect 327276 220658 327304 231676
rect 327460 231662 327934 231690
rect 327264 220652 327316 220658
rect 327264 220594 327316 220600
rect 327460 220522 327488 231662
rect 328564 227594 328592 231676
rect 328552 227588 328604 227594
rect 328552 227530 328604 227536
rect 329208 227186 329236 231676
rect 329852 229906 329880 231676
rect 330036 231662 330510 231690
rect 329840 229900 329892 229906
rect 329840 229842 329892 229848
rect 329196 227180 329248 227186
rect 329196 227122 329248 227128
rect 329748 227180 329800 227186
rect 329748 227122 329800 227128
rect 329012 223576 329064 223582
rect 329012 223518 329064 223524
rect 328828 220788 328880 220794
rect 328828 220730 328880 220736
rect 327448 220516 327500 220522
rect 327448 220458 327500 220464
rect 328184 220516 328236 220522
rect 328184 220458 328236 220464
rect 327540 219292 327592 219298
rect 327540 219234 327592 219240
rect 327552 217002 327580 219234
rect 328196 217002 328224 220458
rect 328840 219026 328868 220730
rect 328828 219020 328880 219026
rect 328828 218962 328880 218968
rect 329024 218890 329052 223518
rect 329012 218884 329064 218890
rect 329012 218826 329064 218832
rect 329196 218068 329248 218074
rect 329196 218010 329248 218016
rect 329208 217002 329236 218010
rect 329760 217002 329788 227122
rect 330036 220114 330064 231662
rect 331140 223446 331168 231676
rect 331324 231662 331798 231690
rect 331968 231662 332442 231690
rect 331128 223440 331180 223446
rect 331128 223382 331180 223388
rect 330484 223168 330536 223174
rect 330484 223110 330536 223116
rect 330024 220108 330076 220114
rect 330024 220050 330076 220056
rect 330496 218074 330524 223110
rect 331324 223038 331352 231662
rect 331312 223032 331364 223038
rect 331312 222974 331364 222980
rect 331680 222148 331732 222154
rect 331680 222090 331732 222096
rect 330484 218068 330536 218074
rect 330484 218010 330536 218016
rect 330852 218068 330904 218074
rect 330852 218010 330904 218016
rect 330864 217002 330892 218010
rect 331692 217002 331720 222090
rect 331968 220794 331996 231662
rect 333072 224398 333100 231676
rect 333244 228676 333296 228682
rect 333244 228618 333296 228624
rect 333060 224392 333112 224398
rect 333060 224334 333112 224340
rect 331956 220788 332008 220794
rect 331956 220730 332008 220736
rect 332508 220108 332560 220114
rect 332508 220050 332560 220056
rect 332520 217002 332548 220050
rect 333256 219434 333284 228618
rect 333716 225758 333744 231676
rect 334084 231662 334374 231690
rect 333704 225752 333756 225758
rect 333704 225694 333756 225700
rect 333888 224392 333940 224398
rect 333888 224334 333940 224340
rect 333164 219406 333284 219434
rect 333164 218074 333192 219406
rect 333704 219020 333756 219026
rect 333704 218962 333756 218968
rect 333152 218068 333204 218074
rect 333152 218010 333204 218016
rect 333336 218068 333388 218074
rect 333336 218010 333388 218016
rect 333348 217002 333376 218010
rect 325436 216974 325588 217002
rect 326416 216974 326844 217002
rect 327244 216974 327580 217002
rect 328072 216974 328224 217002
rect 328900 216974 329236 217002
rect 329728 216974 329788 217002
rect 330556 216974 330892 217002
rect 331384 216974 331720 217002
rect 332212 216974 332548 217002
rect 333040 216974 333376 217002
rect 333716 217002 333744 218962
rect 333900 218074 333928 224334
rect 334084 221882 334112 231662
rect 335004 230042 335032 231676
rect 334992 230036 335044 230042
rect 334992 229978 335044 229984
rect 334256 229900 334308 229906
rect 334256 229842 334308 229848
rect 334268 226302 334296 229842
rect 335648 228546 335676 231676
rect 335636 228540 335688 228546
rect 335636 228482 335688 228488
rect 336292 227050 336320 231676
rect 336648 228540 336700 228546
rect 336648 228482 336700 228488
rect 336280 227044 336332 227050
rect 336280 226986 336332 226992
rect 336464 227044 336516 227050
rect 336464 226986 336516 226992
rect 334256 226296 334308 226302
rect 334256 226238 334308 226244
rect 335084 225752 335136 225758
rect 335084 225694 335136 225700
rect 334072 221876 334124 221882
rect 334072 221818 334124 221824
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 335096 217002 335124 225694
rect 336476 218074 336504 226986
rect 335820 218068 335872 218074
rect 335820 218010 335872 218016
rect 336464 218068 336516 218074
rect 336464 218010 336516 218016
rect 335832 217002 335860 218010
rect 336660 217002 336688 228482
rect 336936 223310 336964 231676
rect 337120 231662 337594 231690
rect 338132 231662 338238 231690
rect 338408 231662 338882 231690
rect 336924 223304 336976 223310
rect 336924 223246 336976 223252
rect 337120 218754 337148 231662
rect 337936 223032 337988 223038
rect 337936 222974 337988 222980
rect 337476 218884 337528 218890
rect 337476 218826 337528 218832
rect 337108 218748 337160 218754
rect 337108 218690 337160 218696
rect 337488 217002 337516 218826
rect 333716 216974 333868 217002
rect 334696 216974 335124 217002
rect 335524 216974 335860 217002
rect 336352 216974 336688 217002
rect 337180 216974 337516 217002
rect 337948 217002 337976 222974
rect 338132 222018 338160 231662
rect 338120 222012 338172 222018
rect 338120 221954 338172 221960
rect 338408 221746 338436 231662
rect 339512 224262 339540 231676
rect 340156 230178 340184 231676
rect 340144 230172 340196 230178
rect 340144 230114 340196 230120
rect 340604 227452 340656 227458
rect 340604 227394 340656 227400
rect 340144 225888 340196 225894
rect 340144 225830 340196 225836
rect 339500 224256 339552 224262
rect 339500 224198 339552 224204
rect 338396 221740 338448 221746
rect 338396 221682 338448 221688
rect 339132 221468 339184 221474
rect 339132 221410 339184 221416
rect 339144 217002 339172 221410
rect 340156 219162 340184 225830
rect 340616 219434 340644 227394
rect 340800 226030 340828 231676
rect 340788 226024 340840 226030
rect 340788 225966 340840 225972
rect 341444 224670 341472 231676
rect 341628 231662 342102 231690
rect 341432 224664 341484 224670
rect 341432 224606 341484 224612
rect 341628 221746 341656 231662
rect 341892 224256 341944 224262
rect 341892 224198 341944 224204
rect 341616 221740 341668 221746
rect 341616 221682 341668 221688
rect 341616 221604 341668 221610
rect 341616 221546 341668 221552
rect 340616 219406 340736 219434
rect 340144 219156 340196 219162
rect 340144 219098 340196 219104
rect 340512 218748 340564 218754
rect 340512 218690 340564 218696
rect 339960 218068 340012 218074
rect 339960 218010 340012 218016
rect 339972 217002 340000 218010
rect 340524 217002 340552 218690
rect 340708 218074 340736 219406
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341628 217002 341656 221546
rect 337948 216974 338008 217002
rect 338836 216974 339172 217002
rect 339664 216974 340000 217002
rect 340492 216974 340552 217002
rect 341320 216974 341656 217002
rect 341904 217002 341932 224198
rect 342732 223582 342760 231676
rect 343376 229094 343404 231676
rect 343192 229066 343404 229094
rect 343744 231662 344034 231690
rect 342720 223576 342772 223582
rect 342720 223518 342772 223524
rect 343192 222902 343220 229066
rect 343364 223304 343416 223310
rect 343364 223246 343416 223252
rect 343180 222896 343232 222902
rect 343180 222838 343232 222844
rect 343376 217002 343404 223246
rect 343744 220250 343772 231662
rect 344664 228818 344692 231676
rect 345308 229906 345336 231676
rect 345664 230104 345716 230110
rect 345664 230046 345716 230052
rect 345296 229900 345348 229906
rect 345296 229842 345348 229848
rect 344652 228812 344704 228818
rect 344652 228754 344704 228760
rect 344928 224664 344980 224670
rect 344928 224606 344980 224612
rect 343732 220244 343784 220250
rect 343732 220186 343784 220192
rect 344100 219292 344152 219298
rect 344100 219234 344152 219240
rect 344112 217002 344140 219234
rect 344940 217002 344968 224606
rect 345676 219434 345704 230046
rect 345952 228954 345980 231676
rect 345940 228948 345992 228954
rect 345940 228890 345992 228896
rect 346124 228812 346176 228818
rect 346124 228754 346176 228760
rect 345848 220244 345900 220250
rect 345848 220186 345900 220192
rect 345860 219434 345888 220186
rect 345572 219428 345704 219434
rect 345624 219406 345704 219428
rect 345768 219406 345888 219434
rect 345572 219370 345624 219376
rect 345768 217002 345796 219406
rect 341904 216974 342148 217002
rect 342976 216974 343404 217002
rect 343804 216974 344140 217002
rect 344632 216974 344968 217002
rect 345460 216974 345796 217002
rect 346136 217002 346164 228754
rect 346596 227730 346624 231676
rect 346584 227724 346636 227730
rect 346584 227666 346636 227672
rect 347044 225888 347096 225894
rect 347044 225830 347096 225836
rect 347056 219298 347084 225830
rect 347240 224534 347268 231676
rect 347884 226030 347912 231676
rect 348160 231662 348542 231690
rect 347872 226024 347924 226030
rect 347872 225966 347924 225972
rect 347228 224528 347280 224534
rect 347228 224470 347280 224476
rect 347504 222896 347556 222902
rect 347504 222838 347556 222844
rect 347044 219292 347096 219298
rect 347044 219234 347096 219240
rect 347516 217002 347544 222838
rect 348160 220386 348188 231662
rect 349172 226166 349200 231676
rect 349160 226160 349212 226166
rect 349160 226102 349212 226108
rect 349068 226024 349120 226030
rect 349068 225966 349120 225972
rect 348148 220380 348200 220386
rect 348148 220322 348200 220328
rect 348884 218204 348936 218210
rect 348884 218146 348936 218152
rect 348240 218068 348292 218074
rect 348240 218010 348292 218016
rect 348252 217002 348280 218010
rect 348896 217002 348924 218146
rect 349080 218074 349108 225966
rect 349816 225622 349844 231676
rect 350460 229770 350488 231676
rect 350448 229764 350500 229770
rect 350448 229706 350500 229712
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 349988 228948 350040 228954
rect 349988 228890 350040 228896
rect 349804 225616 349856 225622
rect 349804 225558 349856 225564
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 350000 217002 350028 228890
rect 350552 225026 350580 229570
rect 351104 228410 351132 231676
rect 351288 231662 351762 231690
rect 351288 229094 351316 231662
rect 351288 229066 351408 229094
rect 351092 228404 351144 228410
rect 351092 228346 351144 228352
rect 351184 225616 351236 225622
rect 351184 225558 351236 225564
rect 346136 216974 346288 217002
rect 347116 216974 347544 217002
rect 347944 216974 348280 217002
rect 348772 216974 348924 217002
rect 349600 216974 350028 217002
rect 350368 224998 350580 225026
rect 350368 217002 350396 224998
rect 351196 218210 351224 225558
rect 351380 220522 351408 229066
rect 352392 227322 352420 231676
rect 353036 230110 353064 231676
rect 353024 230104 353076 230110
rect 353024 230046 353076 230052
rect 352564 229900 352616 229906
rect 352564 229842 352616 229848
rect 352380 227316 352432 227322
rect 352380 227258 352432 227264
rect 351368 220516 351420 220522
rect 351368 220458 351420 220464
rect 352380 219428 352432 219434
rect 352380 219370 352432 219376
rect 351552 218612 351604 218618
rect 351552 218554 351604 218560
rect 351184 218204 351236 218210
rect 351184 218146 351236 218152
rect 351564 217002 351592 218554
rect 352392 217002 352420 219370
rect 352576 219026 352604 229842
rect 353680 227186 353708 231676
rect 353956 231662 354338 231690
rect 353668 227180 353720 227186
rect 353668 227122 353720 227128
rect 353956 222154 353984 231662
rect 354588 227180 354640 227186
rect 354588 227122 354640 227128
rect 353944 222148 353996 222154
rect 353944 222090 353996 222096
rect 353208 220380 353260 220386
rect 353208 220322 353260 220328
rect 352564 219020 352616 219026
rect 352564 218962 352616 218968
rect 353220 217002 353248 220322
rect 354404 219156 354456 219162
rect 354404 219098 354456 219104
rect 354036 218068 354088 218074
rect 354036 218010 354088 218016
rect 354048 217002 354076 218010
rect 350368 216974 350428 217002
rect 351256 216974 351592 217002
rect 352084 216974 352420 217002
rect 352912 216974 353248 217002
rect 353740 216974 354076 217002
rect 354416 217002 354444 219098
rect 354600 218074 354628 227122
rect 354968 223174 354996 231676
rect 355612 228682 355640 231676
rect 355600 228676 355652 228682
rect 355600 228618 355652 228624
rect 355324 228404 355376 228410
rect 355324 228346 355376 228352
rect 354956 223168 355008 223174
rect 354956 223110 355008 223116
rect 355336 218618 355364 228346
rect 355508 226908 355560 226914
rect 355508 226850 355560 226856
rect 355520 219162 355548 226850
rect 356256 224398 356284 231676
rect 356900 225758 356928 231676
rect 356888 225752 356940 225758
rect 356888 225694 356940 225700
rect 356244 224392 356296 224398
rect 356244 224334 356296 224340
rect 357348 224392 357400 224398
rect 357348 224334 357400 224340
rect 357164 223168 357216 223174
rect 357164 223110 357216 223116
rect 355508 219156 355560 219162
rect 355508 219098 355560 219104
rect 355692 219020 355744 219026
rect 355692 218962 355744 218968
rect 355324 218612 355376 218618
rect 355324 218554 355376 218560
rect 354588 218068 354640 218074
rect 354588 218010 354640 218016
rect 355704 217002 355732 218962
rect 356520 218068 356572 218074
rect 356520 218010 356572 218016
rect 356532 217002 356560 218010
rect 357176 217002 357204 223110
rect 357360 218074 357388 224334
rect 357544 220114 357572 231676
rect 358188 229906 358216 231676
rect 358176 229900 358228 229906
rect 358176 229842 358228 229848
rect 358084 229288 358136 229294
rect 358084 229230 358136 229236
rect 357532 220108 357584 220114
rect 357532 220050 357584 220056
rect 358096 218890 358124 229230
rect 358832 228546 358860 231676
rect 359200 231662 359490 231690
rect 358820 228540 358872 228546
rect 358820 228482 358872 228488
rect 359200 223038 359228 231662
rect 359464 227588 359516 227594
rect 359464 227530 359516 227536
rect 359188 223032 359240 223038
rect 359188 222974 359240 222980
rect 358728 219292 358780 219298
rect 358728 219234 358780 219240
rect 358084 218884 358136 218890
rect 358084 218826 358136 218832
rect 357348 218068 357400 218074
rect 357348 218010 357400 218016
rect 358176 218068 358228 218074
rect 358176 218010 358228 218016
rect 358188 217002 358216 218010
rect 358740 217002 358768 219234
rect 359476 218074 359504 227530
rect 360120 227050 360148 231676
rect 360764 229294 360792 231676
rect 360752 229288 360804 229294
rect 360752 229230 360804 229236
rect 360936 229288 360988 229294
rect 360936 229230 360988 229236
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359832 221740 359884 221746
rect 359832 221682 359884 221688
rect 359464 218068 359516 218074
rect 359464 218010 359516 218016
rect 359844 217002 359872 221682
rect 360660 220108 360712 220114
rect 360660 220050 360712 220056
rect 360672 217002 360700 220050
rect 360948 219434 360976 229230
rect 361408 227458 361436 231676
rect 361592 231662 362066 231690
rect 362236 231662 362710 231690
rect 361396 227452 361448 227458
rect 361396 227394 361448 227400
rect 361304 227316 361356 227322
rect 361304 227258 361356 227264
rect 360856 219406 360976 219434
rect 360856 218754 360884 219406
rect 360844 218748 360896 218754
rect 360844 218690 360896 218696
rect 361316 217002 361344 227258
rect 361592 221610 361620 231662
rect 362236 229094 362264 231662
rect 363340 229294 363368 231676
rect 363328 229288 363380 229294
rect 363328 229230 363380 229236
rect 362052 229066 362264 229094
rect 361580 221604 361632 221610
rect 361580 221546 361632 221552
rect 362052 221474 362080 229066
rect 362868 228404 362920 228410
rect 362868 228346 362920 228352
rect 362224 227316 362276 227322
rect 362224 227258 362276 227264
rect 362236 226914 362264 227258
rect 362224 226908 362276 226914
rect 362224 226850 362276 226856
rect 362040 221468 362092 221474
rect 362040 221410 362092 221416
rect 362316 221468 362368 221474
rect 362316 221410 362368 221416
rect 362328 217002 362356 221410
rect 362880 217002 362908 228346
rect 363984 223310 364012 231676
rect 364156 229900 364208 229906
rect 364156 229842 364208 229848
rect 363972 223304 364024 223310
rect 363972 223246 364024 223252
rect 364168 219434 364196 229842
rect 364628 224670 364656 231676
rect 364812 231662 365286 231690
rect 364616 224664 364668 224670
rect 364616 224606 364668 224612
rect 364812 224262 364840 231662
rect 365916 225894 365944 231676
rect 366192 231662 366574 231690
rect 366192 228818 366220 231662
rect 366180 228812 366232 228818
rect 366180 228754 366232 228760
rect 366916 228540 366968 228546
rect 366916 228482 366968 228488
rect 366272 227792 366324 227798
rect 366272 227734 366324 227740
rect 365904 225888 365956 225894
rect 365904 225830 365956 225836
rect 364800 224256 364852 224262
rect 364800 224198 364852 224204
rect 364984 224256 365036 224262
rect 364984 224198 365036 224204
rect 364076 219406 364196 219434
rect 364076 217002 364104 219406
rect 364996 219298 365024 224198
rect 364984 219292 365036 219298
rect 364984 219234 365036 219240
rect 366284 219162 366312 227734
rect 366272 219156 366324 219162
rect 366272 219098 366324 219104
rect 366732 218884 366784 218890
rect 366732 218826 366784 218832
rect 365628 218340 365680 218346
rect 365628 218282 365680 218288
rect 364800 218204 364852 218210
rect 364800 218146 364852 218152
rect 364812 217002 364840 218146
rect 365640 217002 365668 218282
rect 366456 218068 366508 218074
rect 366456 218010 366508 218016
rect 366468 217002 366496 218010
rect 354416 216974 354568 217002
rect 355396 216974 355732 217002
rect 356224 216974 356560 217002
rect 357052 216974 357204 217002
rect 357880 216974 358216 217002
rect 358708 216974 358768 217002
rect 359536 216974 359872 217002
rect 360364 216974 360700 217002
rect 361192 216974 361344 217002
rect 362020 216974 362356 217002
rect 362848 216974 362908 217002
rect 363676 216974 364104 217002
rect 364504 216974 364840 217002
rect 365332 216974 365668 217002
rect 366160 216974 366496 217002
rect 366744 217002 366772 218826
rect 366928 218074 366956 228482
rect 367204 226030 367232 231676
rect 367388 231662 367862 231690
rect 367192 226024 367244 226030
rect 367192 225966 367244 225972
rect 367388 220250 367416 231662
rect 367744 225888 367796 225894
rect 367744 225830 367796 225836
rect 367376 220244 367428 220250
rect 367376 220186 367428 220192
rect 367756 218210 367784 225830
rect 368492 222902 368520 231676
rect 369136 228954 369164 231676
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 369780 228682 369808 231676
rect 369768 228676 369820 228682
rect 369768 228618 369820 228624
rect 369124 227928 369176 227934
rect 369124 227870 369176 227876
rect 368480 222896 368532 222902
rect 368480 222838 368532 222844
rect 368112 220244 368164 220250
rect 368112 220186 368164 220192
rect 367744 218204 367796 218210
rect 367744 218146 367796 218152
rect 366916 218068 366968 218074
rect 366916 218010 366968 218016
rect 368124 217002 368152 220186
rect 369136 219026 369164 227870
rect 369768 227044 369820 227050
rect 369768 226986 369820 226992
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 369780 218210 369808 226986
rect 370424 225622 370452 231676
rect 371068 229770 371096 231676
rect 371436 231662 371726 231690
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 370964 229628 371016 229634
rect 370964 229570 371016 229576
rect 370412 225616 370464 225622
rect 370412 225558 370464 225564
rect 370504 223032 370556 223038
rect 370504 222974 370556 222980
rect 368940 218204 368992 218210
rect 368940 218146 368992 218152
rect 369768 218204 369820 218210
rect 369768 218146 369820 218152
rect 368952 217002 368980 218146
rect 370516 218074 370544 222974
rect 370976 219434 371004 229570
rect 371148 220516 371200 220522
rect 371148 220458 371200 220464
rect 370700 219406 371004 219434
rect 369768 218068 369820 218074
rect 369768 218010 369820 218016
rect 370504 218068 370556 218074
rect 370504 218010 370556 218016
rect 369780 217002 369808 218010
rect 370700 217002 370728 219406
rect 371160 217002 371188 220458
rect 371436 220386 371464 231662
rect 372356 227322 372384 231676
rect 373000 227798 373028 231676
rect 372988 227792 373040 227798
rect 372988 227734 373040 227740
rect 372344 227316 372396 227322
rect 372344 227258 372396 227264
rect 373264 227316 373316 227322
rect 373264 227258 373316 227264
rect 372344 225616 372396 225622
rect 372344 225558 372396 225564
rect 371424 220380 371476 220386
rect 371424 220322 371476 220328
rect 372356 217002 372384 225558
rect 373080 219156 373132 219162
rect 373080 219098 373132 219104
rect 373092 217002 373120 219098
rect 373276 218346 373304 227258
rect 373644 227186 373672 231676
rect 373816 228812 373868 228818
rect 373816 228754 373868 228760
rect 373632 227180 373684 227186
rect 373632 227122 373684 227128
rect 373828 219162 373856 228754
rect 374288 224398 374316 231676
rect 374932 227594 374960 231676
rect 375576 227934 375604 231676
rect 375564 227928 375616 227934
rect 375564 227870 375616 227876
rect 374920 227588 374972 227594
rect 374920 227530 374972 227536
rect 374276 224392 374328 224398
rect 374276 224334 374328 224340
rect 375288 224392 375340 224398
rect 375288 224334 375340 224340
rect 375104 222896 375156 222902
rect 375104 222838 375156 222844
rect 373816 219156 373868 219162
rect 373816 219098 373868 219104
rect 373724 219020 373776 219026
rect 373724 218962 373776 218968
rect 373264 218340 373316 218346
rect 373264 218282 373316 218288
rect 373736 217002 373764 218962
rect 374736 218068 374788 218074
rect 374736 218010 374788 218016
rect 374748 217002 374776 218010
rect 366744 216974 366988 217002
rect 367816 216974 368152 217002
rect 368644 216974 368980 217002
rect 369472 216974 369808 217002
rect 370300 216974 370728 217002
rect 371128 216974 371188 217002
rect 371956 216974 372384 217002
rect 372784 216974 373120 217002
rect 373612 216974 373764 217002
rect 374440 216974 374776 217002
rect 375116 217002 375144 222838
rect 375300 218074 375328 224334
rect 376220 223174 376248 231676
rect 376484 228676 376536 228682
rect 376484 228618 376536 228624
rect 376208 223168 376260 223174
rect 376208 223110 376260 223116
rect 375288 218068 375340 218074
rect 375288 218010 375340 218016
rect 376496 217002 376524 228618
rect 376864 221746 376892 231676
rect 377232 231662 377522 231690
rect 377232 227458 377260 231662
rect 377404 230444 377456 230450
rect 377404 230386 377456 230392
rect 377220 227452 377272 227458
rect 377220 227394 377272 227400
rect 376852 221740 376904 221746
rect 376852 221682 376904 221688
rect 377416 220114 377444 230386
rect 378152 224262 378180 231676
rect 378796 230450 378824 231676
rect 378784 230444 378836 230450
rect 378784 230386 378836 230392
rect 378968 229152 379020 229158
rect 378968 229094 379020 229100
rect 378140 224256 378192 224262
rect 378140 224198 378192 224204
rect 378048 221604 378100 221610
rect 378048 221546 378100 221552
rect 377404 220108 377456 220114
rect 377404 220050 377456 220056
rect 377220 218204 377272 218210
rect 377220 218146 377272 218152
rect 377232 217002 377260 218146
rect 378060 217002 378088 221546
rect 378980 219434 379008 229094
rect 379440 228410 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 379624 225894 379652 231662
rect 379612 225888 379664 225894
rect 379612 225830 379664 225836
rect 379336 225752 379388 225758
rect 379336 225694 379388 225700
rect 378704 219406 379008 219434
rect 378704 218890 378732 219406
rect 378692 218884 378744 218890
rect 378692 218826 378744 218832
rect 379152 218748 379204 218754
rect 379152 218690 379204 218696
rect 378876 218068 378928 218074
rect 378876 218010 378928 218016
rect 378888 217002 378916 218010
rect 375116 216974 375268 217002
rect 376096 216974 376524 217002
rect 376924 216974 377260 217002
rect 377752 216974 378088 217002
rect 378580 216974 378916 217002
rect 379164 217002 379192 218690
rect 379348 218074 379376 225694
rect 380268 221474 380296 231662
rect 380440 230036 380492 230042
rect 380440 229978 380492 229984
rect 380256 221468 380308 221474
rect 380256 221410 380308 221416
rect 380452 219434 380480 229978
rect 381372 229906 381400 231676
rect 381360 229900 381412 229906
rect 381360 229842 381412 229848
rect 382016 228546 382044 231676
rect 382476 231662 382674 231690
rect 382004 228540 382056 228546
rect 382004 228482 382056 228488
rect 381912 228404 381964 228410
rect 381912 228346 381964 228352
rect 380176 219406 380480 219434
rect 380176 219026 380204 219406
rect 380164 219020 380216 219026
rect 380164 218962 380216 218968
rect 380532 218476 380584 218482
rect 380532 218418 380584 218424
rect 379336 218068 379388 218074
rect 379336 218010 379388 218016
rect 380544 217002 380572 218418
rect 381924 218074 381952 228346
rect 382096 227180 382148 227186
rect 382096 227122 382148 227128
rect 381360 218068 381412 218074
rect 381360 218010 381412 218016
rect 381912 218068 381964 218074
rect 381912 218010 381964 218016
rect 381372 217002 381400 218010
rect 382108 217002 382136 227122
rect 382476 220250 382504 231662
rect 383304 227458 383332 231676
rect 383948 229158 383976 231676
rect 384304 229900 384356 229906
rect 384304 229842 384356 229848
rect 383936 229152 383988 229158
rect 383936 229094 383988 229100
rect 383292 227452 383344 227458
rect 383292 227394 383344 227400
rect 382832 227316 382884 227322
rect 382832 227258 382884 227264
rect 382464 220244 382516 220250
rect 382464 220186 382516 220192
rect 382844 218210 382872 227258
rect 383016 220244 383068 220250
rect 383016 220186 383068 220192
rect 382832 218204 382884 218210
rect 382832 218146 382884 218152
rect 383028 217002 383056 220186
rect 383568 219292 383620 219298
rect 383568 219234 383620 219240
rect 383580 217002 383608 219234
rect 384316 218482 384344 229842
rect 384592 223038 384620 231676
rect 384580 223032 384632 223038
rect 384580 222974 384632 222980
rect 385236 220522 385264 231676
rect 385880 227050 385908 231676
rect 386524 229770 386552 231676
rect 386512 229764 386564 229770
rect 386512 229706 386564 229712
rect 386972 229764 387024 229770
rect 386972 229706 387024 229712
rect 386984 229094 387012 229706
rect 387168 229094 387196 231676
rect 386984 229066 387104 229094
rect 387168 229066 387288 229094
rect 385868 227044 385920 227050
rect 385868 226986 385920 226992
rect 386328 227044 386380 227050
rect 386328 226986 386380 226992
rect 385224 220516 385276 220522
rect 385224 220458 385276 220464
rect 384672 219020 384724 219026
rect 384672 218962 384724 218968
rect 384304 218476 384356 218482
rect 384304 218418 384356 218424
rect 384684 217002 384712 218962
rect 386144 218884 386196 218890
rect 386144 218826 386196 218832
rect 385500 218068 385552 218074
rect 385500 218010 385552 218016
rect 385512 217002 385540 218010
rect 386156 217002 386184 218826
rect 386340 218074 386368 226986
rect 387076 219298 387104 229066
rect 387260 228818 387288 229066
rect 387248 228812 387300 228818
rect 387248 228754 387300 228760
rect 387812 224398 387840 231676
rect 388088 231662 388470 231690
rect 388088 225622 388116 231662
rect 389100 230042 389128 231676
rect 389088 230036 389140 230042
rect 389088 229978 389140 229984
rect 389744 228682 389772 231676
rect 390020 231662 390402 231690
rect 389732 228676 389784 228682
rect 389732 228618 389784 228624
rect 388076 225616 388128 225622
rect 388076 225558 388128 225564
rect 388444 225616 388496 225622
rect 388444 225558 388496 225564
rect 387800 224392 387852 224398
rect 387800 224334 387852 224340
rect 387708 223032 387760 223038
rect 387708 222974 387760 222980
rect 387064 219292 387116 219298
rect 387064 219234 387116 219240
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 387156 218068 387208 218074
rect 387156 218010 387208 218016
rect 387168 217002 387196 218010
rect 387720 217002 387748 222974
rect 388456 218074 388484 225558
rect 388904 224256 388956 224262
rect 388904 224198 388956 224204
rect 388444 218068 388496 218074
rect 388444 218010 388496 218016
rect 388916 217002 388944 224198
rect 390020 221610 390048 231662
rect 390284 228676 390336 228682
rect 390284 228618 390336 228624
rect 390008 221604 390060 221610
rect 390008 221546 390060 221552
rect 390296 218074 390324 228618
rect 391032 222902 391060 231676
rect 391676 227322 391704 231676
rect 392136 231662 392334 231690
rect 391848 228404 391900 228410
rect 391848 228346 391900 228352
rect 391664 227316 391716 227322
rect 391664 227258 391716 227264
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391296 221468 391348 221474
rect 391296 221410 391348 221416
rect 390468 220108 390520 220114
rect 390468 220050 390520 220056
rect 389640 218068 389692 218074
rect 389640 218010 389692 218016
rect 390284 218068 390336 218074
rect 390284 218010 390336 218016
rect 389652 217002 389680 218010
rect 390480 217002 390508 220050
rect 391308 217002 391336 221410
rect 391860 217002 391888 228346
rect 392136 218754 392164 231662
rect 392964 229094 392992 231676
rect 392872 229066 392992 229094
rect 392872 228546 392900 229066
rect 392860 228540 392912 228546
rect 392860 228482 392912 228488
rect 393044 228540 393096 228546
rect 393044 228482 393096 228488
rect 392124 218748 392176 218754
rect 392124 218690 392176 218696
rect 393056 217002 393084 228482
rect 393608 225758 393636 231676
rect 394252 229906 394280 231676
rect 394804 231662 394910 231690
rect 394240 229900 394292 229906
rect 394240 229842 394292 229848
rect 393964 227792 394016 227798
rect 393964 227734 394016 227740
rect 393596 225752 393648 225758
rect 393596 225694 393648 225700
rect 393976 219026 394004 227734
rect 394608 225752 394660 225758
rect 394608 225694 394660 225700
rect 393964 219020 394016 219026
rect 393964 218962 394016 218968
rect 394424 218204 394476 218210
rect 394424 218146 394476 218152
rect 393780 218068 393832 218074
rect 393780 218010 393832 218016
rect 393792 217002 393820 218010
rect 394436 217002 394464 218146
rect 394620 218074 394648 225694
rect 394804 220250 394832 231662
rect 395540 227798 395568 231676
rect 395528 227792 395580 227798
rect 395528 227734 395580 227740
rect 395988 227316 396040 227322
rect 395988 227258 396040 227264
rect 394792 220244 394844 220250
rect 394792 220186 394844 220192
rect 395804 218748 395856 218754
rect 395804 218690 395856 218696
rect 394608 218068 394660 218074
rect 394608 218010 394660 218016
rect 395436 218068 395488 218074
rect 395436 218010 395488 218016
rect 395448 217002 395476 218010
rect 379164 216974 379408 217002
rect 380236 216974 380572 217002
rect 381064 216974 381400 217002
rect 381892 216974 382136 217002
rect 382720 216974 383056 217002
rect 383548 216974 383608 217002
rect 384376 216974 384712 217002
rect 385204 216974 385540 217002
rect 386032 216974 386184 217002
rect 386860 216974 387196 217002
rect 387688 216974 387748 217002
rect 388516 216974 388944 217002
rect 389344 216974 389680 217002
rect 390172 216974 390508 217002
rect 391000 216974 391336 217002
rect 391828 216974 391888 217002
rect 392656 216974 393084 217002
rect 393484 216974 393820 217002
rect 394312 216974 394464 217002
rect 395140 216974 395476 217002
rect 395816 217002 395844 218690
rect 396000 218074 396028 227258
rect 396184 227186 396212 231676
rect 396828 229770 396856 231676
rect 396816 229764 396868 229770
rect 396816 229706 396868 229712
rect 397472 227798 397500 231676
rect 396724 227792 396776 227798
rect 396724 227734 396776 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396172 227180 396224 227186
rect 396172 227122 396224 227128
rect 396736 218890 396764 227734
rect 398116 223038 398144 231676
rect 398760 227050 398788 231676
rect 398748 227044 398800 227050
rect 398748 226986 398800 226992
rect 398748 226908 398800 226914
rect 398748 226850 398800 226856
rect 398104 223032 398156 223038
rect 398104 222974 398156 222980
rect 397184 222896 397236 222902
rect 397184 222838 397236 222844
rect 396724 218884 396776 218890
rect 396724 218826 396776 218832
rect 395988 218068 396040 218074
rect 395988 218010 396040 218016
rect 397196 217002 397224 222838
rect 397920 220244 397972 220250
rect 397920 220186 397972 220192
rect 397932 217002 397960 220186
rect 398760 217002 398788 226850
rect 399404 225622 399432 231676
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399392 225616 399444 225622
rect 399392 225558 399444 225564
rect 399576 218068 399628 218074
rect 399576 218010 399628 218016
rect 399588 217002 399616 218010
rect 395816 216974 395968 217002
rect 396796 216974 397224 217002
rect 397624 216974 397960 217002
rect 398452 216974 398788 217002
rect 399280 216974 399616 217002
rect 399864 217002 399892 229706
rect 400048 228682 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 401704 231662 401994 231690
rect 400036 228676 400088 228682
rect 400036 228618 400088 228624
rect 400036 228540 400088 228546
rect 400036 228482 400088 228488
rect 400048 218074 400076 228482
rect 400416 221474 400444 231662
rect 400968 224262 400996 231662
rect 401324 228812 401376 228818
rect 401324 228754 401376 228760
rect 400956 224256 401008 224262
rect 400956 224198 401008 224204
rect 400404 221468 400456 221474
rect 400404 221410 400456 221416
rect 400036 218068 400088 218074
rect 400036 218010 400088 218016
rect 401336 217002 401364 228754
rect 401704 220114 401732 231662
rect 402624 228410 402652 231676
rect 402612 228404 402664 228410
rect 402612 228346 402664 228352
rect 403268 227798 403296 231676
rect 403912 228274 403940 231676
rect 404268 230376 404320 230382
rect 404268 230318 404320 230324
rect 403900 228268 403952 228274
rect 403900 228210 403952 228216
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 404084 227792 404136 227798
rect 404084 227734 404136 227740
rect 401692 220108 401744 220114
rect 401692 220050 401744 220056
rect 402060 219020 402112 219026
rect 402060 218962 402112 218968
rect 402072 217002 402100 218962
rect 402256 218210 402284 227734
rect 402704 218884 402756 218890
rect 402704 218826 402756 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402716 217002 402744 218826
rect 403532 218068 403584 218074
rect 403532 218010 403584 218016
rect 403544 217002 403572 218010
rect 399864 216974 400108 217002
rect 400936 216974 401364 217002
rect 401764 216974 402100 217002
rect 402592 216974 402744 217002
rect 403420 216974 403572 217002
rect 404096 217002 404124 227734
rect 404280 218074 404308 230318
rect 404556 225758 404584 231676
rect 404740 231662 405214 231690
rect 404544 225752 404596 225758
rect 404544 225694 404596 225700
rect 404740 219434 404768 231662
rect 405372 221468 405424 221474
rect 405372 221410 405424 221416
rect 404556 219406 404768 219434
rect 404556 218754 404584 219406
rect 404544 218748 404596 218754
rect 404544 218690 404596 218696
rect 404268 218068 404320 218074
rect 404268 218010 404320 218016
rect 405384 217002 405412 221410
rect 405844 220250 405872 231676
rect 406488 227322 406516 231676
rect 407132 229094 407160 231676
rect 407132 229066 407252 229094
rect 406476 227316 406528 227322
rect 406476 227258 406528 227264
rect 407028 224936 407080 224942
rect 407028 224878 407080 224884
rect 405832 220244 405884 220250
rect 405832 220186 405884 220192
rect 406200 219564 406252 219570
rect 406200 219506 406252 219512
rect 406212 217002 406240 219506
rect 407040 217002 407068 224878
rect 407224 222902 407252 229066
rect 407776 228546 407804 231676
rect 408420 228818 408448 231676
rect 408696 231662 409078 231690
rect 408408 228812 408460 228818
rect 408408 228754 408460 228760
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 407764 227928 407816 227934
rect 407764 227870 407816 227876
rect 407212 222896 407264 222902
rect 407212 222838 407264 222844
rect 407580 219156 407632 219162
rect 407580 219098 407632 219104
rect 407592 217002 407620 219098
rect 407776 219026 407804 227870
rect 408696 226914 408724 231662
rect 408868 230240 408920 230246
rect 408868 230182 408920 230188
rect 408880 227798 408908 230182
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409604 228404 409656 228410
rect 409604 228346 409656 228352
rect 408868 227792 408920 227798
rect 408868 227734 408920 227740
rect 409144 227792 409196 227798
rect 409144 227734 409196 227740
rect 408684 226908 408736 226914
rect 408684 226850 408736 226856
rect 408408 222896 408460 222902
rect 408408 222838 408460 222844
rect 407764 219020 407816 219026
rect 407764 218962 407816 218968
rect 408420 217002 408448 222838
rect 409156 218890 409184 227734
rect 409144 218884 409196 218890
rect 409144 218826 409196 218832
rect 409616 217002 409644 228346
rect 410352 227798 410380 231676
rect 410996 230246 411024 231676
rect 410984 230240 411036 230246
rect 410984 230182 411036 230188
rect 410892 230036 410944 230042
rect 410892 229978 410944 229984
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410904 218074 410932 229978
rect 411076 228676 411128 228682
rect 411076 228618 411128 228624
rect 410340 218068 410392 218074
rect 410340 218010 410392 218016
rect 410892 218068 410944 218074
rect 410892 218010 410944 218016
rect 410352 217002 410380 218010
rect 411088 217002 411116 228618
rect 411640 227934 411668 231676
rect 412284 230382 412312 231676
rect 412744 231662 412942 231690
rect 412272 230376 412324 230382
rect 412272 230318 412324 230324
rect 412456 229764 412508 229770
rect 412456 229706 412508 229712
rect 411628 227928 411680 227934
rect 411628 227870 411680 227876
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411916 219162 411944 227734
rect 411904 219156 411956 219162
rect 411904 219098 411956 219104
rect 412468 218890 412496 229706
rect 412744 219570 412772 231662
rect 413572 227798 413600 231676
rect 413744 229084 413796 229090
rect 413744 229026 413796 229032
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219564 412784 219570
rect 412732 219506 412784 219512
rect 411996 218884 412048 218890
rect 411996 218826 412048 218832
rect 412456 218884 412508 218890
rect 412456 218826 412508 218832
rect 412008 217002 412036 218826
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 412560 217002 412588 218690
rect 413756 217002 413784 229026
rect 414216 221474 414244 231676
rect 414860 224942 414888 231676
rect 415504 228410 415532 231676
rect 416148 228682 416176 231676
rect 416136 228676 416188 228682
rect 416136 228618 416188 228624
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416596 227792 416648 227798
rect 416596 227734 416648 227740
rect 414848 224936 414900 224942
rect 414848 224878 414900 224884
rect 416412 224256 416464 224262
rect 416412 224198 416464 224204
rect 414204 221468 414256 221474
rect 414204 221410 414256 221416
rect 415124 221060 415176 221066
rect 415124 221002 415176 221008
rect 414480 220788 414532 220794
rect 414480 220730 414532 220736
rect 414492 217002 414520 220730
rect 415136 217002 415164 221002
rect 416424 219434 416452 224198
rect 416608 219434 416636 227734
rect 416792 222902 416820 231676
rect 417436 230042 417464 231676
rect 417712 231662 418094 231690
rect 418264 231662 418738 231690
rect 417424 230036 417476 230042
rect 417424 229978 417476 229984
rect 417712 229094 417740 231662
rect 417160 229066 417740 229094
rect 416780 222896 416832 222902
rect 416780 222838 416832 222844
rect 416424 219406 416544 219434
rect 416608 219406 416728 219434
rect 416136 218068 416188 218074
rect 416136 218010 416188 218016
rect 416148 217002 416176 218010
rect 404096 216974 404248 217002
rect 405076 216974 405412 217002
rect 405904 216974 406240 217002
rect 406732 216974 407068 217002
rect 407560 216974 407620 217002
rect 408388 216974 408448 217002
rect 409216 216974 409644 217002
rect 410044 216974 410380 217002
rect 410872 216974 411116 217002
rect 411700 216974 412036 217002
rect 412528 216974 412588 217002
rect 413356 216974 413784 217002
rect 414184 216974 414520 217002
rect 415012 216974 415164 217002
rect 415840 216974 416176 217002
rect 416516 217002 416544 219406
rect 416700 218074 416728 219406
rect 417160 218754 417188 229066
rect 418264 220794 418292 231662
rect 419368 229770 419396 231676
rect 419356 229764 419408 229770
rect 419356 229706 419408 229712
rect 419448 229288 419500 229294
rect 419448 229230 419500 229236
rect 418252 220788 418304 220794
rect 418252 220730 418304 220736
rect 417792 219428 417844 219434
rect 417792 219370 417844 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416688 218068 416740 218074
rect 416688 218010 416740 218016
rect 417804 217002 417832 219370
rect 419264 219156 419316 219162
rect 419264 219098 419316 219104
rect 418620 218068 418672 218074
rect 418620 218010 418672 218016
rect 418632 217002 418660 218010
rect 419276 217002 419304 219098
rect 419460 218074 419488 229230
rect 420012 229158 420040 231676
rect 420000 229152 420052 229158
rect 420000 229094 420052 229100
rect 420184 229152 420236 229158
rect 420184 229094 420236 229100
rect 420196 221066 420224 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420184 221060 420236 221066
rect 420184 221002 420236 221008
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420276 218068 420328 218074
rect 420276 218010 420328 218016
rect 420288 217002 420316 218010
rect 416516 216974 416668 217002
rect 417496 216974 417832 217002
rect 418324 216974 418660 217002
rect 419152 216974 419304 217002
rect 419980 216974 420316 217002
rect 420656 217002 420684 220798
rect 420840 218074 420868 222838
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 423784 231662 423890 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 224262 422248 229066
rect 422208 224256 422260 224262
rect 422208 224198 422260 224204
rect 421932 220108 421984 220114
rect 421932 220050 421984 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420828 218068 420880 218074
rect 420828 218010 420880 218016
rect 421944 217002 421972 220050
rect 422864 219434 422892 231662
rect 423588 224188 423640 224194
rect 423588 224130 423640 224136
rect 422680 219406 422892 219434
rect 422680 219162 422708 219406
rect 422668 219156 422720 219162
rect 422668 219098 422720 219104
rect 422760 218204 422812 218210
rect 422760 218146 422812 218152
rect 422772 217002 422800 218146
rect 423600 217002 423628 224130
rect 423784 220862 423812 231662
rect 424520 229294 424548 231676
rect 424508 229288 424560 229294
rect 424508 229230 424560 229236
rect 424324 229152 424376 229158
rect 424324 229094 424376 229100
rect 424336 224194 424364 229094
rect 424324 224188 424376 224194
rect 424324 224130 424376 224136
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 221944 425020 221950
rect 424968 221886 425020 221892
rect 423772 220856 423824 220862
rect 423772 220798 423824 220804
rect 424416 218068 424468 218074
rect 424416 218010 424468 218016
rect 424428 217002 424456 218010
rect 424980 217002 425008 221886
rect 425440 218210 425468 231662
rect 426452 224942 426480 231676
rect 426820 231662 427110 231690
rect 426440 224936 426492 224942
rect 426440 224878 426492 224884
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427924 231662 428398 231690
rect 428752 231662 429042 231690
rect 429212 231662 429686 231690
rect 429856 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 426992 224936 427044 224942
rect 426992 224878 427044 224884
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426808 218340 426860 218346
rect 426808 218282 426860 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 426072 218204 426124 218210
rect 426072 218146 426124 218152
rect 426084 217002 426112 218146
rect 426820 217002 426848 218282
rect 427004 218074 427032 224878
rect 427924 218210 427952 231662
rect 428752 219434 428780 231662
rect 429212 221950 429240 231662
rect 429200 221944 429252 221950
rect 429200 221886 429252 221892
rect 429856 219434 429884 231662
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 428476 219406 428780 219434
rect 429396 219406 429884 219434
rect 430212 219428 430264 219434
rect 427912 218204 427964 218210
rect 427912 218146 427964 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427728 218068 427780 218074
rect 427728 218010 427780 218016
rect 427740 217002 427768 218010
rect 428292 217002 428320 219370
rect 428476 218074 428504 219406
rect 429396 218346 429424 219406
rect 430212 219370 430264 219376
rect 429384 218340 429436 218346
rect 429384 218282 429436 218288
rect 428464 218068 428516 218074
rect 428464 218010 428516 218016
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217002 429148 218010
rect 430224 217002 430252 219370
rect 430684 218074 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220516 432288 220522
rect 432236 220458 432288 220464
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220458
rect 432708 219434 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 430960 219406 431264 219434
rect 431972 219406 432276 219434
rect 432696 219428 432748 219434
rect 430672 218068 430724 218074
rect 430672 218010 430724 218016
rect 430960 217002 430988 219406
rect 431972 218090 432000 219406
rect 432696 219370 432748 219376
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 431880 218062 432000 218090
rect 432696 218068 432748 218074
rect 431880 217002 431908 218062
rect 432696 218010 432748 218016
rect 432708 217002 432736 218010
rect 433260 217002 433288 218146
rect 420656 216974 420808 217002
rect 421636 216974 421972 217002
rect 422464 216974 422800 217002
rect 423292 216974 423628 217002
rect 424120 216974 424456 217002
rect 424948 216974 425008 217002
rect 425776 216974 426112 217002
rect 426604 216974 426848 217002
rect 427432 216974 427768 217002
rect 428260 216974 428320 217002
rect 429088 216974 429148 217002
rect 429916 216974 430252 217002
rect 430744 216974 430988 217002
rect 431572 216974 431908 217002
rect 432400 216974 432736 217002
rect 433228 216974 433288 217002
rect 433628 217002 433656 229066
rect 433812 218074 433840 229066
rect 434824 220522 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220516 434864 220522
rect 434812 220458 434864 220464
rect 435088 219428 435140 219434
rect 435088 219370 435140 219376
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 435100 217002 435128 219370
rect 435284 218210 435312 231662
rect 436100 229424 436152 229430
rect 436100 229366 436152 229372
rect 435916 218340 435968 218346
rect 435916 218282 435968 218288
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435928 217002 435956 218282
rect 436112 218226 436140 229366
rect 436296 218346 436324 231662
rect 436756 229430 436784 231676
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436744 229424 436796 229430
rect 436744 229366 436796 229372
rect 437032 219502 437060 231662
rect 437020 219496 437072 219502
rect 437020 219438 437072 219444
rect 437768 219434 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 437492 219406 437796 219434
rect 436284 218340 436336 218346
rect 436284 218282 436336 218288
rect 436112 218198 437060 218226
rect 436836 218068 436888 218074
rect 436836 218010 436888 218016
rect 436848 217002 436876 218010
rect 433628 216974 434056 217002
rect 434884 216974 435128 217002
rect 435712 216974 435956 217002
rect 436540 216974 436876 217002
rect 437032 217002 437060 218198
rect 437492 218074 437520 219406
rect 438964 218074 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438492 218068 438544 218074
rect 438492 218010 438544 218016
rect 438952 218068 439004 218074
rect 438952 218010 439004 218016
rect 438504 217002 438532 218010
rect 439332 217002 439360 230318
rect 440344 219434 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 440160 219406 440372 219434
rect 440160 217002 440188 219406
rect 440712 217002 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443210 231662 443408 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 441540 218062 441660 218090
rect 441540 217002 441568 218062
rect 437032 216974 437368 217002
rect 438196 216974 438532 217002
rect 439024 216974 439360 217002
rect 439852 216974 440188 217002
rect 440680 216974 440740 217002
rect 441508 216974 441568 217002
rect 442092 217002 442120 229094
rect 443380 217002 443408 231662
rect 443552 230444 443604 230450
rect 443552 230386 443604 230392
rect 442092 216974 442336 217002
rect 443164 216974 443408 217002
rect 443564 217002 443592 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 230110 444512 231676
rect 444668 231662 445142 231690
rect 444472 230104 444524 230110
rect 444472 230046 444524 230052
rect 444668 219434 444696 231662
rect 444840 230376 444892 230382
rect 444840 230318 444892 230324
rect 444852 229094 444880 230318
rect 445772 229094 445800 231676
rect 446416 230382 446444 231676
rect 446404 230376 446456 230382
rect 446404 230318 446456 230324
rect 447060 230246 447088 231676
rect 447244 231662 447718 231690
rect 447048 230240 447100 230246
rect 447048 230182 447100 230188
rect 444852 229066 445248 229094
rect 445772 229066 446076 229094
rect 444576 219406 444696 219434
rect 444576 217002 444604 219406
rect 445220 217002 445248 229066
rect 446048 217002 446076 229066
rect 447244 219434 447272 231662
rect 447600 230104 447652 230110
rect 447600 230046 447652 230052
rect 447152 219406 447272 219434
rect 447152 217870 447180 219406
rect 447140 217864 447192 217870
rect 447140 217806 447192 217812
rect 447612 217002 447640 230046
rect 448348 229094 448376 231676
rect 448992 229430 449020 231676
rect 449636 230382 449664 231676
rect 449164 230376 449216 230382
rect 449164 230318 449216 230324
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229424 449032 229430
rect 448980 229366 449032 229372
rect 448348 229066 448652 229094
rect 448624 217870 448652 229066
rect 447784 217864 447836 217870
rect 447784 217806 447836 217812
rect 448612 217864 448664 217870
rect 448612 217806 448664 217812
rect 443564 216974 443992 217002
rect 444576 216974 444820 217002
rect 445220 216974 445648 217002
rect 446048 216974 446476 217002
rect 447304 216974 447640 217002
rect 447796 217002 447824 217806
rect 449176 217002 449204 230318
rect 449900 230240 449952 230246
rect 449900 230182 449952 230188
rect 449912 229094 449940 230182
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 449912 229066 450216 229094
rect 449440 217864 449492 217870
rect 449440 217806 449492 217812
rect 447796 216974 448132 217002
rect 448960 216974 449204 217002
rect 449452 217002 449480 217806
rect 450188 217002 450216 229066
rect 450556 218414 450584 230318
rect 450924 229158 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451372 229424 451424 229430
rect 451372 229366 451424 229372
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 451384 224262 451412 229366
rect 451832 229288 451884 229294
rect 451832 229230 451884 229236
rect 451372 224256 451424 224262
rect 451372 224198 451424 224204
rect 450544 218408 450596 218414
rect 450544 218350 450596 218356
rect 451844 217002 451872 229230
rect 452016 224256 452068 224262
rect 452016 224198 452068 224204
rect 452028 219434 452056 224198
rect 452580 221474 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452568 221468 452620 221474
rect 452568 221410 452620 221416
rect 449452 216974 449788 217002
rect 450188 216974 450616 217002
rect 451444 216974 451872 217002
rect 451936 219406 452056 219434
rect 451936 217002 451964 219406
rect 452764 217002 452792 229094
rect 453316 218074 453344 230182
rect 453500 229362 453528 231676
rect 454144 230246 454172 231676
rect 454802 231662 455092 231690
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230240 454184 230246
rect 454132 230182 454184 230188
rect 453488 229356 453540 229362
rect 453488 229298 453540 229304
rect 453580 218408 453632 218414
rect 453580 218350 453632 218356
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 453592 217002 453620 218350
rect 454328 217002 454356 230318
rect 455064 218210 455092 231662
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455236 230240 455288 230246
rect 455236 230182 455288 230188
rect 455248 220794 455276 230182
rect 455788 229356 455840 229362
rect 455788 229298 455840 229304
rect 455800 229094 455828 229298
rect 456076 229094 456104 231676
rect 455800 229066 456012 229094
rect 456076 229066 456196 229094
rect 455236 220788 455288 220794
rect 455236 220730 455288 220736
rect 455052 218204 455104 218210
rect 455052 218146 455104 218152
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455432 217002 455460 218010
rect 455984 217002 456012 229066
rect 456168 224398 456196 229066
rect 456156 224392 456208 224398
rect 456156 224334 456208 224340
rect 456720 221610 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 457180 229094 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 457180 229066 457668 229094
rect 456708 221604 456760 221610
rect 456708 221546 456760 221552
rect 456708 221468 456760 221474
rect 456708 221410 456760 221416
rect 456720 219434 456748 221410
rect 456720 219406 456840 219434
rect 456812 217002 456840 219406
rect 457640 217002 457668 229066
rect 458008 223582 458036 231676
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 457996 223576 458048 223582
rect 457996 223518 458048 223524
rect 458548 220788 458600 220794
rect 458548 220730 458600 220736
rect 458560 217002 458588 220730
rect 459480 220250 459508 231662
rect 459652 224392 459704 224398
rect 459652 224334 459704 224340
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459664 217002 459692 224334
rect 459940 222902 459968 231676
rect 460584 224738 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224732 460624 224738
rect 460572 224674 460624 224680
rect 460204 223576 460256 223582
rect 460204 223518 460256 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 460216 219026 460244 223518
rect 461768 221604 461820 221610
rect 461768 221546 461820 221552
rect 460204 219020 460256 219026
rect 460204 218962 460256 218968
rect 461124 219020 461176 219026
rect 461124 218962 461176 218968
rect 460204 218204 460256 218210
rect 460204 218146 460256 218152
rect 460216 217002 460244 218146
rect 461136 217002 461164 218962
rect 461780 217002 461808 221546
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 229094 462544 231676
rect 462424 229066 462544 229094
rect 462424 224262 462452 229066
rect 462596 225820 462648 225826
rect 462596 225762 462648 225768
rect 462412 224256 462464 224262
rect 462412 224198 462464 224204
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462608 217002 462636 225762
rect 463160 225282 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225276 463200 225282
rect 463148 225218 463200 225224
rect 462964 224732 463016 224738
rect 462964 224674 463016 224680
rect 462976 218074 463004 224674
rect 462964 218068 463016 218074
rect 462964 218010 463016 218016
rect 463896 217002 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227594 465948 231662
rect 466104 231662 466394 231690
rect 465908 227588 465960 227594
rect 465908 227530 465960 227536
rect 466104 220862 466132 231662
rect 467024 230042 467052 231676
rect 467012 230036 467064 230042
rect 467012 229978 467064 229984
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467104 225276 467156 225282
rect 467104 225218 467156 225224
rect 466736 222896 466788 222902
rect 466736 222838 466788 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465172 220244 465224 220250
rect 465172 220186 465224 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464436 218068 464488 218074
rect 464436 218010 464488 218016
rect 451936 216974 452272 217002
rect 452764 216974 453100 217002
rect 453592 216974 453928 217002
rect 454328 216974 454756 217002
rect 455432 216974 455584 217002
rect 455984 216974 456412 217002
rect 456812 216974 457240 217002
rect 457640 216974 458068 217002
rect 458560 216974 458896 217002
rect 459664 216974 459724 217002
rect 460216 216974 460552 217002
rect 461136 216974 461380 217002
rect 461780 216974 462208 217002
rect 462608 216974 463036 217002
rect 463864 216974 463924 217002
rect 464448 217002 464476 218010
rect 465184 217002 465212 220186
rect 466000 218204 466052 218210
rect 466000 218146 466052 218152
rect 466012 217002 466040 218146
rect 466748 217002 466776 222838
rect 467116 218074 467144 225218
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230450 468340 231676
rect 468864 231662 468970 231690
rect 468300 230444 468352 230450
rect 468300 230386 468352 230392
rect 468864 229770 468892 231662
rect 469036 230444 469088 230450
rect 469036 230386 469088 230392
rect 468852 229764 468904 229770
rect 468852 229706 468904 229712
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468484 222148 468536 222154
rect 468484 222090 468536 222096
rect 467104 218068 467156 218074
rect 467104 218010 467156 218016
rect 467840 218068 467892 218074
rect 467840 218010 467892 218016
rect 467852 217002 467880 218010
rect 468496 217002 468524 222090
rect 469048 220250 469076 230386
rect 469600 229906 469628 231676
rect 469588 229900 469640 229906
rect 469588 229842 469640 229848
rect 469864 227588 469916 227594
rect 469864 227530 469916 227536
rect 469680 224256 469732 224262
rect 469680 224198 469732 224204
rect 469312 220720 469364 220726
rect 469312 220662 469364 220668
rect 469036 220244 469088 220250
rect 469036 220186 469088 220192
rect 469324 217002 469352 220662
rect 469692 217138 469720 224198
rect 469876 218550 469904 227530
rect 470244 224262 470272 231676
rect 470888 230246 470916 231676
rect 470876 230240 470928 230246
rect 470876 230182 470928 230188
rect 471532 227934 471560 231676
rect 471888 230240 471940 230246
rect 471888 230182 471940 230188
rect 471520 227928 471572 227934
rect 471520 227870 471572 227876
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230182
rect 472176 227050 472204 231676
rect 472834 231662 473308 231690
rect 472164 227044 472216 227050
rect 472164 226986 472216 226992
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471704 220856 471756 220862
rect 471704 220798 471756 220804
rect 469864 218544 469916 218550
rect 469864 218486 469916 218492
rect 470968 218544 471020 218550
rect 470968 218486 471020 218492
rect 469692 217110 470088 217138
rect 470060 217002 470088 217110
rect 470980 217002 471008 218486
rect 471716 218074 471744 220798
rect 473280 220386 473308 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474766 231662 475056 231690
rect 474004 230036 474056 230042
rect 474004 229978 474056 229984
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473452 222896 473504 222902
rect 473452 222838 473504 222844
rect 473268 220380 473320 220386
rect 473268 220322 473320 220328
rect 471980 219632 472032 219638
rect 471980 219574 472032 219580
rect 471704 218068 471756 218074
rect 471704 218010 471756 218016
rect 471992 217002 472020 219574
rect 472624 218068 472676 218074
rect 472624 218010 472676 218016
rect 472636 217002 472664 218010
rect 473464 217002 473492 222838
rect 474016 220794 474044 229978
rect 474476 229094 474504 231662
rect 474476 229066 474780 229094
rect 474752 222902 474780 229066
rect 475028 227798 475056 231662
rect 475396 230246 475424 231676
rect 475384 230240 475436 230246
rect 475384 230182 475436 230188
rect 475384 229764 475436 229770
rect 475384 229706 475436 229712
rect 475016 227792 475068 227798
rect 475016 227734 475068 227740
rect 474740 222896 474792 222902
rect 474740 222838 474792 222844
rect 475396 220794 475424 229706
rect 476040 229226 476068 231676
rect 476684 230382 476712 231676
rect 476672 230376 476724 230382
rect 476672 230318 476724 230324
rect 476856 229900 476908 229906
rect 476856 229842 476908 229848
rect 476028 229220 476080 229226
rect 476028 229162 476080 229168
rect 476672 225616 476724 225622
rect 476672 225558 476724 225564
rect 475752 223576 475804 223582
rect 475752 223518 475804 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475108 220788 475160 220794
rect 475108 220730 475160 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474280 220244 474332 220250
rect 474280 220186 474332 220192
rect 474292 217002 474320 220186
rect 475120 217002 475148 220730
rect 475764 219298 475792 223518
rect 476120 220788 476172 220794
rect 476120 220730 476172 220736
rect 475752 219292 475804 219298
rect 475752 219234 475804 219240
rect 476132 217002 476160 220730
rect 476684 217002 476712 225558
rect 476868 220794 476896 229842
rect 477328 225622 477356 231676
rect 477972 229634 478000 231676
rect 478340 231662 478630 231690
rect 477960 229628 478012 229634
rect 477960 229570 478012 229576
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 478340 223038 478368 231662
rect 479064 230240 479116 230246
rect 479064 230182 479116 230188
rect 478512 229628 478564 229634
rect 478512 229570 478564 229576
rect 478524 228154 478552 229570
rect 478696 229220 478748 229226
rect 478696 229162 478748 229168
rect 478708 228274 478736 229162
rect 478696 228268 478748 228274
rect 478696 228210 478748 228216
rect 478524 228126 478644 228154
rect 478328 223032 478380 223038
rect 478328 222974 478380 222980
rect 477592 222148 477644 222154
rect 477592 222090 477644 222096
rect 476856 220788 476908 220794
rect 476856 220730 476908 220736
rect 477604 217002 477632 222090
rect 478420 220788 478472 220794
rect 478420 220730 478472 220736
rect 478432 217002 478460 220730
rect 478616 220250 478644 228126
rect 479076 224398 479104 230182
rect 479260 229770 479288 231676
rect 479708 230376 479760 230382
rect 479708 230318 479760 230324
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 479720 228682 479748 230318
rect 479904 229294 479932 231676
rect 480548 230382 480576 231676
rect 480536 230376 480588 230382
rect 480536 230318 480588 230324
rect 479892 229288 479944 229294
rect 479892 229230 479944 229236
rect 479708 228676 479760 228682
rect 479708 228618 479760 228624
rect 479248 227928 479300 227934
rect 479248 227870 479300 227876
rect 479064 224392 479116 224398
rect 479064 224334 479116 224340
rect 478604 220244 478656 220250
rect 478604 220186 478656 220192
rect 479260 219434 479288 227870
rect 481192 227050 481220 231676
rect 481548 230376 481600 230382
rect 481548 230318 481600 230324
rect 480812 227044 480864 227050
rect 480812 226986 480864 226992
rect 481180 227044 481232 227050
rect 481180 226986 481232 226992
rect 479524 224256 479576 224262
rect 479524 224198 479576 224204
rect 479168 219406 479288 219434
rect 479168 217002 479196 219406
rect 479536 218346 479564 224198
rect 479524 218340 479576 218346
rect 479524 218282 479576 218288
rect 480352 218340 480404 218346
rect 480352 218282 480404 218288
rect 480364 217002 480392 218282
rect 480824 217002 480852 226986
rect 481560 220114 481588 230318
rect 481836 229906 481864 231676
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 482284 229288 482336 229294
rect 482284 229230 482336 229236
rect 482296 220386 482324 229230
rect 482480 228546 482508 231676
rect 483124 230382 483152 231676
rect 483112 230376 483164 230382
rect 483112 230318 483164 230324
rect 482468 228540 482520 228546
rect 482468 228482 482520 228488
rect 482836 227792 482888 227798
rect 482836 227734 482888 227740
rect 482848 222222 482876 227734
rect 483768 224262 483796 231676
rect 484426 231662 484808 231690
rect 484308 230376 484360 230382
rect 484308 230318 484360 230324
rect 483756 224256 483808 224262
rect 483756 224198 483808 224204
rect 482836 222216 482888 222222
rect 482836 222158 482888 222164
rect 481732 220380 481784 220386
rect 481732 220322 481784 220328
rect 482284 220380 482336 220386
rect 482284 220322 482336 220328
rect 481548 220108 481600 220114
rect 481548 220050 481600 220056
rect 481744 217002 481772 220322
rect 482560 219292 482612 219298
rect 482560 219234 482612 219240
rect 482572 217002 482600 219234
rect 482848 218074 482876 222158
rect 484320 221610 484348 230318
rect 484780 230042 484808 231662
rect 484768 230036 484820 230042
rect 484768 229978 484820 229984
rect 485056 227322 485084 231676
rect 485608 231662 485714 231690
rect 486358 231662 486648 231690
rect 485044 227316 485096 227322
rect 485044 227258 485096 227264
rect 485608 223038 485636 231662
rect 486620 224670 486648 231662
rect 486988 228410 487016 231676
rect 487160 229764 487212 229770
rect 487160 229706 487212 229712
rect 487172 228818 487200 229706
rect 487160 228812 487212 228818
rect 487160 228754 487212 228760
rect 487436 228676 487488 228682
rect 487436 228618 487488 228624
rect 486976 228404 487028 228410
rect 486976 228346 487028 228352
rect 487068 228268 487120 228274
rect 487068 228210 487120 228216
rect 486608 224664 486660 224670
rect 486608 224606 486660 224612
rect 485780 224392 485832 224398
rect 485780 224334 485832 224340
rect 485044 223032 485096 223038
rect 485044 222974 485096 222980
rect 485596 223032 485648 223038
rect 485596 222974 485648 222980
rect 484860 222896 484912 222902
rect 484860 222838 484912 222844
rect 484308 221604 484360 221610
rect 484308 221546 484360 221552
rect 484032 221468 484084 221474
rect 484032 221410 484084 221416
rect 482836 218068 482888 218074
rect 482836 218010 482888 218016
rect 484044 217002 484072 221410
rect 484872 219609 484900 222838
rect 484858 219600 484914 219609
rect 484858 219535 484914 219544
rect 484872 217002 484900 219535
rect 485056 218890 485084 222974
rect 485044 218884 485096 218890
rect 485044 218826 485096 218832
rect 485044 218068 485096 218074
rect 485044 218010 485096 218016
rect 464448 216974 464692 217002
rect 465184 216974 465520 217002
rect 466012 216974 466348 217002
rect 466748 216974 467176 217002
rect 467852 216974 468004 217002
rect 468496 216974 468832 217002
rect 469324 216974 469660 217002
rect 470060 216974 470488 217002
rect 470980 216974 471316 217002
rect 471992 216974 472144 217002
rect 472636 216974 472972 217002
rect 473464 216974 473800 217002
rect 474292 216974 474628 217002
rect 475120 216974 475456 217002
rect 476132 216974 476284 217002
rect 476684 216974 477112 217002
rect 477604 216974 477940 217002
rect 478432 216974 478768 217002
rect 479168 216974 479596 217002
rect 480364 216974 480424 217002
rect 480824 216974 481252 217002
rect 481744 216974 482080 217002
rect 482572 216974 482908 217002
rect 483736 216974 484072 217002
rect 484564 216974 484900 217002
rect 485056 217002 485084 218010
rect 485792 217002 485820 224334
rect 487080 220969 487108 228210
rect 487066 220960 487122 220969
rect 487066 220895 487122 220904
rect 487080 217002 487108 220895
rect 487448 219337 487476 228618
rect 487632 225758 487660 231676
rect 488276 230178 488304 231676
rect 488264 230172 488316 230178
rect 488264 230114 488316 230120
rect 488920 225894 488948 231676
rect 488908 225888 488960 225894
rect 488908 225830 488960 225836
rect 487620 225752 487672 225758
rect 487620 225694 487672 225700
rect 488540 225616 488592 225622
rect 488540 225558 488592 225564
rect 487434 219328 487490 219337
rect 487434 219263 487490 219272
rect 485056 216974 485392 217002
rect 485792 216974 486220 217002
rect 487048 216974 487108 217002
rect 487448 217002 487476 219263
rect 488552 217002 488580 225558
rect 489564 222902 489592 231676
rect 490208 230382 490236 231676
rect 490196 230376 490248 230382
rect 490196 230318 490248 230324
rect 490852 230042 490880 231676
rect 491208 230376 491260 230382
rect 491208 230318 491260 230324
rect 490840 230036 490892 230042
rect 490840 229978 490892 229984
rect 489920 229900 489972 229906
rect 489920 229842 489972 229848
rect 489932 229094 489960 229842
rect 489932 229066 490144 229094
rect 489920 228812 489972 228818
rect 489920 228754 489972 228760
rect 489552 222896 489604 222902
rect 489552 222838 489604 222844
rect 489184 220244 489236 220250
rect 489184 220186 489236 220192
rect 488906 217288 488962 217297
rect 488906 217223 488962 217232
rect 488920 217002 488948 217223
rect 487448 216974 487876 217002
rect 488552 216974 488948 217002
rect 489196 217002 489224 220186
rect 489932 218657 489960 228754
rect 490116 226370 490144 229066
rect 490104 226364 490156 226370
rect 490104 226306 490156 226312
rect 491220 220250 491248 230318
rect 491496 224534 491524 231676
rect 492154 231662 492628 231690
rect 491484 224528 491536 224534
rect 491484 224470 491536 224476
rect 492600 220386 492628 231662
rect 492784 230382 492812 231676
rect 493442 231662 494008 231690
rect 494086 231662 494376 231690
rect 492772 230376 492824 230382
rect 492772 230318 492824 230324
rect 493784 230376 493836 230382
rect 493980 230364 494008 231662
rect 493980 230336 494192 230364
rect 493784 230318 493836 230324
rect 491392 220380 491444 220386
rect 491392 220322 491444 220328
rect 492588 220380 492640 220386
rect 492588 220322 492640 220328
rect 491208 220244 491260 220250
rect 491208 220186 491260 220192
rect 490656 218884 490708 218890
rect 490656 218826 490708 218832
rect 489918 218648 489974 218657
rect 489918 218583 489974 218592
rect 490668 218113 490696 218826
rect 491206 218648 491262 218657
rect 491206 218583 491262 218592
rect 490654 218104 490710 218113
rect 490654 218039 490710 218048
rect 490668 217002 490696 218039
rect 491220 217002 491248 218583
rect 491404 218074 491432 220322
rect 492772 220108 492824 220114
rect 492772 220050 492824 220056
rect 491392 218068 491444 218074
rect 491392 218010 491444 218016
rect 492312 218068 492364 218074
rect 492312 218010 492364 218016
rect 492324 217002 492352 218010
rect 489196 216974 489532 217002
rect 490360 216974 490696 217002
rect 491188 216974 491248 217002
rect 492016 216974 492352 217002
rect 492784 217002 492812 220050
rect 493796 219978 493824 230318
rect 493968 230036 494020 230042
rect 493968 229978 494020 229984
rect 493980 228818 494008 229978
rect 493968 228812 494020 228818
rect 493968 228754 494020 228760
rect 493968 227044 494020 227050
rect 493968 226986 494020 226992
rect 493784 219972 493836 219978
rect 493784 219914 493836 219920
rect 493980 219502 494008 226986
rect 494164 225622 494192 230336
rect 494348 229770 494376 231662
rect 494716 230382 494744 231676
rect 494704 230376 494756 230382
rect 494704 230318 494756 230324
rect 494336 229764 494388 229770
rect 494336 229706 494388 229712
rect 495360 228682 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 228676 495400 228682
rect 495348 228618 495400 228624
rect 494704 228540 494756 228546
rect 494704 228482 494756 228488
rect 494152 225616 494204 225622
rect 494152 225558 494204 225564
rect 493968 219496 494020 219502
rect 493968 219438 494020 219444
rect 493980 217002 494008 219438
rect 494716 217705 494744 228482
rect 494888 226364 494940 226370
rect 494888 226306 494940 226312
rect 494900 219745 494928 226306
rect 496188 221746 496216 231662
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 496176 221740 496228 221746
rect 496176 221682 496228 221688
rect 495808 221604 495860 221610
rect 495808 221546 495860 221552
rect 494886 219736 494942 219745
rect 494886 219671 494942 219680
rect 494702 217696 494758 217705
rect 494702 217631 494758 217640
rect 494900 217002 494928 219671
rect 495162 217696 495218 217705
rect 495162 217631 495218 217640
rect 492784 216974 492844 217002
rect 493672 216974 494008 217002
rect 494500 216974 494928 217002
rect 495176 216753 495204 217631
rect 495820 217002 495848 221546
rect 496372 220522 496400 230318
rect 497292 227050 497320 231676
rect 497936 230314 497964 231676
rect 497924 230308 497976 230314
rect 497924 230250 497976 230256
rect 497464 229628 497516 229634
rect 497464 229570 497516 229576
rect 497280 227044 497332 227050
rect 497280 226986 497332 226992
rect 497280 224256 497332 224262
rect 497280 224198 497332 224204
rect 496360 220516 496412 220522
rect 496360 220458 496412 220464
rect 497292 219638 497320 224198
rect 497280 219632 497332 219638
rect 497280 219574 497332 219580
rect 497292 217002 497320 219574
rect 497476 218657 497504 229570
rect 498580 227186 498608 231676
rect 498844 227316 498896 227322
rect 498844 227258 498896 227264
rect 498568 227180 498620 227186
rect 498568 227122 498620 227128
rect 498200 223032 498252 223038
rect 498200 222974 498252 222980
rect 497462 218648 497518 218657
rect 497462 218583 497518 218592
rect 495820 216974 496156 217002
rect 496984 216974 497320 217002
rect 497476 217002 497504 218583
rect 498212 217870 498240 222974
rect 498200 217864 498252 217870
rect 498200 217806 498252 217812
rect 498856 217297 498884 227258
rect 499224 224398 499252 231676
rect 499868 230382 499896 231676
rect 500052 231662 500526 231690
rect 499856 230376 499908 230382
rect 499856 230318 499908 230324
rect 499580 230104 499632 230110
rect 499580 230046 499632 230052
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 499592 223582 499620 230046
rect 499580 223576 499632 223582
rect 499580 223518 499632 223524
rect 500052 221610 500080 231662
rect 501156 226030 501184 231676
rect 501328 230376 501380 230382
rect 501328 230318 501380 230324
rect 501340 227322 501368 230318
rect 501800 229294 501828 231676
rect 501788 229288 501840 229294
rect 501788 229230 501840 229236
rect 502444 228546 502472 231676
rect 503102 231662 503392 231690
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 501696 228404 501748 228410
rect 501696 228346 501748 228352
rect 501328 227316 501380 227322
rect 501328 227258 501380 227264
rect 501144 226024 501196 226030
rect 501144 225966 501196 225972
rect 501512 225752 501564 225758
rect 501512 225694 501564 225700
rect 500408 224664 500460 224670
rect 500408 224606 500460 224612
rect 500040 221604 500092 221610
rect 500040 221546 500092 221552
rect 500420 218385 500448 224606
rect 500406 218376 500462 218385
rect 500406 218311 500462 218320
rect 499120 217864 499172 217870
rect 499120 217806 499172 217812
rect 498842 217288 498898 217297
rect 498842 217223 498898 217232
rect 498856 217002 498884 217223
rect 497476 216974 497812 217002
rect 498640 216974 498884 217002
rect 499132 217002 499160 217806
rect 500420 217002 500448 218311
rect 501326 217560 501382 217569
rect 501326 217495 501382 217504
rect 501340 217025 501368 217495
rect 501326 217016 501382 217025
rect 499132 216974 499468 217002
rect 500296 216974 500448 217002
rect 501124 216974 501326 217002
rect 501524 217002 501552 225694
rect 501708 217569 501736 228346
rect 502984 225888 503036 225894
rect 502984 225830 503036 225836
rect 502996 217841 503024 225830
rect 503168 223576 503220 223582
rect 503168 223518 503220 223524
rect 503180 219201 503208 223518
rect 503364 223038 503392 231662
rect 503732 229634 503760 231676
rect 504390 231662 504680 231690
rect 504364 230240 504416 230246
rect 504364 230182 504416 230188
rect 503720 229628 503772 229634
rect 503720 229570 503772 229576
rect 503352 223032 503404 223038
rect 503352 222974 503404 222980
rect 503996 222896 504048 222902
rect 503996 222838 504048 222844
rect 503166 219192 503222 219201
rect 503166 219127 503222 219136
rect 502982 217832 503038 217841
rect 502982 217767 503038 217776
rect 501694 217560 501750 217569
rect 501694 217495 501750 217504
rect 503180 217002 503208 219127
rect 503626 217832 503682 217841
rect 503626 217767 503682 217776
rect 503640 217002 503668 217767
rect 501524 216974 501952 217002
rect 502780 216974 503208 217002
rect 503608 216974 503668 217002
rect 504008 217002 504036 222838
rect 504376 219842 504404 230182
rect 504652 222902 504680 231662
rect 505020 230382 505048 231676
rect 505678 231662 505968 231690
rect 505008 230376 505060 230382
rect 505008 230318 505060 230324
rect 505744 230376 505796 230382
rect 505744 230318 505796 230324
rect 504640 222896 504692 222902
rect 504640 222838 504692 222844
rect 505756 221882 505784 230318
rect 505940 230042 505968 231662
rect 505928 230036 505980 230042
rect 505928 229978 505980 229984
rect 505928 228812 505980 228818
rect 505928 228754 505980 228760
rect 505744 221876 505796 221882
rect 505744 221818 505796 221824
rect 505940 221241 505968 228754
rect 506308 228410 506336 231676
rect 506296 228404 506348 228410
rect 506296 228346 506348 228352
rect 506480 224528 506532 224534
rect 506480 224470 506532 224476
rect 505926 221232 505982 221241
rect 505926 221167 505982 221176
rect 505192 220108 505244 220114
rect 505192 220050 505244 220056
rect 504364 219836 504416 219842
rect 504364 219778 504416 219784
rect 505204 218929 505232 220050
rect 505190 218920 505246 218929
rect 505190 218855 505246 218864
rect 505204 218226 505232 218855
rect 505204 218198 505324 218226
rect 505100 218068 505152 218074
rect 505100 218010 505152 218016
rect 505112 217569 505140 218010
rect 505098 217560 505154 217569
rect 505098 217495 505154 217504
rect 505296 217002 505324 218198
rect 504008 216974 504436 217002
rect 505264 216974 505324 217002
rect 505940 217002 505968 221167
rect 506492 217002 506520 224470
rect 506952 223310 506980 231676
rect 507610 231662 507808 231690
rect 507124 229288 507176 229294
rect 507124 229230 507176 229236
rect 507136 228818 507164 229230
rect 507124 228812 507176 228818
rect 507124 228754 507176 228760
rect 506940 223304 506992 223310
rect 506940 223246 506992 223252
rect 507780 220386 507808 231662
rect 508240 224670 508268 231676
rect 508504 229628 508556 229634
rect 508504 229570 508556 229576
rect 508228 224664 508280 224670
rect 508228 224606 508280 224612
rect 508516 220658 508544 229570
rect 508884 225894 508912 231676
rect 509528 229498 509556 231676
rect 509884 229764 509936 229770
rect 509884 229706 509936 229712
rect 509516 229492 509568 229498
rect 509516 229434 509568 229440
rect 508872 225888 508924 225894
rect 508872 225830 508924 225836
rect 509700 225616 509752 225622
rect 509700 225558 509752 225564
rect 508504 220652 508556 220658
rect 508504 220594 508556 220600
rect 507400 220380 507452 220386
rect 507400 220322 507452 220328
rect 507768 220380 507820 220386
rect 507768 220322 507820 220328
rect 507412 219201 507440 220322
rect 508228 219972 508280 219978
rect 508228 219914 508280 219920
rect 507214 219192 507270 219201
rect 507214 219127 507216 219136
rect 507268 219127 507270 219136
rect 507398 219192 507454 219201
rect 507398 219127 507454 219136
rect 507216 219098 507268 219104
rect 507412 217002 507440 219127
rect 508240 217841 508268 219914
rect 509238 219192 509294 219201
rect 509238 219127 509294 219136
rect 509514 219192 509570 219201
rect 509514 219127 509516 219136
rect 509252 219042 509280 219127
rect 509568 219127 509570 219136
rect 509516 219098 509568 219104
rect 509252 219014 509556 219042
rect 509528 218958 509556 219014
rect 509516 218952 509568 218958
rect 509238 218920 509294 218929
rect 509516 218894 509568 218900
rect 509238 218855 509294 218864
rect 509252 218686 509280 218855
rect 509240 218680 509292 218686
rect 509240 218622 509292 218628
rect 508042 217832 508098 217841
rect 508042 217767 508044 217776
rect 508096 217767 508098 217776
rect 508226 217832 508282 217841
rect 508226 217767 508282 217776
rect 509330 217832 509386 217841
rect 509330 217767 509386 217776
rect 509514 217832 509570 217841
rect 509514 217767 509516 217776
rect 508044 217738 508096 217744
rect 508240 217002 508268 217767
rect 509344 217682 509372 217767
rect 509568 217767 509570 217776
rect 509516 217738 509568 217744
rect 509344 217654 509464 217682
rect 509436 217598 509464 217654
rect 509424 217592 509476 217598
rect 509424 217534 509476 217540
rect 509712 217002 509740 225558
rect 509896 218210 509924 229706
rect 510172 225622 510200 231676
rect 510620 229900 510672 229906
rect 510620 229842 510672 229848
rect 510632 227798 510660 229842
rect 510620 227792 510672 227798
rect 510620 227734 510672 227740
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510816 224534 510844 231676
rect 511460 230246 511488 231676
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 511448 228676 511500 228682
rect 511448 228618 511500 228624
rect 510804 224528 510856 224534
rect 510804 224470 510856 224476
rect 510988 220244 511040 220250
rect 510988 220186 511040 220192
rect 509884 218204 509936 218210
rect 509884 218146 509936 218152
rect 510528 218204 510580 218210
rect 510528 218146 510580 218152
rect 510540 217002 510568 218146
rect 505940 216974 506092 217002
rect 506492 216974 506920 217002
rect 507412 216974 507748 217002
rect 508240 216974 508576 217002
rect 509404 216974 509740 217002
rect 510232 216974 510568 217002
rect 511000 217002 511028 220186
rect 511460 217002 511488 228618
rect 512104 228274 512132 231676
rect 512762 231662 513144 231690
rect 513116 229094 513144 231662
rect 513392 229906 513420 231676
rect 513380 229900 513432 229906
rect 513380 229842 513432 229848
rect 513116 229066 513236 229094
rect 512092 228268 512144 228274
rect 512092 228210 512144 228216
rect 513012 227792 513064 227798
rect 513012 227734 513064 227740
rect 513024 219230 513052 227734
rect 513208 224262 513236 229066
rect 514036 227050 514064 231676
rect 513840 227044 513892 227050
rect 513840 226986 513892 226992
rect 514024 227044 514076 227050
rect 514024 226986 514076 226992
rect 513196 224256 513248 224262
rect 513196 224198 513248 224204
rect 513564 221740 513616 221746
rect 513564 221682 513616 221688
rect 513576 220862 513604 221682
rect 513564 220856 513616 220862
rect 513564 220798 513616 220804
rect 513012 219224 513064 219230
rect 513012 219166 513064 219172
rect 513024 217002 513052 219166
rect 513576 217002 513604 220798
rect 513852 219434 513880 226986
rect 514680 226166 514708 231676
rect 515324 229634 515352 231676
rect 515772 230036 515824 230042
rect 515772 229978 515824 229984
rect 515312 229628 515364 229634
rect 515312 229570 515364 229576
rect 514668 226160 514720 226166
rect 514668 226102 514720 226108
rect 515784 224806 515812 229978
rect 515968 227458 515996 231676
rect 516612 230382 516640 231676
rect 516600 230376 516652 230382
rect 516600 230318 516652 230324
rect 516784 230240 516836 230246
rect 516784 230182 516836 230188
rect 515956 227452 516008 227458
rect 515956 227394 516008 227400
rect 516048 227180 516100 227186
rect 516048 227122 516100 227128
rect 515772 224800 515824 224806
rect 515772 224742 515824 224748
rect 516060 220998 516088 227122
rect 516416 224392 516468 224398
rect 516416 224334 516468 224340
rect 516048 220992 516100 220998
rect 516048 220934 516100 220940
rect 515220 220516 515272 220522
rect 515220 220458 515272 220464
rect 515232 219842 515260 220458
rect 515220 219836 515272 219842
rect 515220 219778 515272 219784
rect 513852 219406 513972 219434
rect 511000 216974 511060 217002
rect 511460 216974 511888 217002
rect 512716 216974 513052 217002
rect 513544 216974 513604 217002
rect 513944 217002 513972 219406
rect 515232 217002 515260 219778
rect 516060 217002 516088 220934
rect 513944 216974 514372 217002
rect 515200 216974 515260 217002
rect 516028 216974 516088 217002
rect 516428 217002 516456 224334
rect 516796 223446 516824 230182
rect 517256 230042 517284 231676
rect 517428 230376 517480 230382
rect 517428 230318 517480 230324
rect 517244 230036 517296 230042
rect 517244 229978 517296 229984
rect 516784 223440 516836 223446
rect 516784 223382 516836 223388
rect 517440 219774 517468 230318
rect 517900 228954 517928 231676
rect 518164 229492 518216 229498
rect 518164 229434 518216 229440
rect 517888 228948 517940 228954
rect 517888 228890 517940 228896
rect 517796 227316 517848 227322
rect 517796 227258 517848 227264
rect 517612 222012 517664 222018
rect 517612 221954 517664 221960
rect 517624 221610 517652 221954
rect 517612 221604 517664 221610
rect 517612 221546 517664 221552
rect 517808 221513 517836 227258
rect 518176 221610 518204 229434
rect 518544 227594 518572 231676
rect 519188 229498 519216 231676
rect 519176 229492 519228 229498
rect 519176 229434 519228 229440
rect 519832 229090 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 521120 230246 521148 231676
rect 521568 230376 521620 230382
rect 521568 230318 521620 230324
rect 521108 230240 521160 230246
rect 521108 230182 521160 230188
rect 519820 229084 519872 229090
rect 519820 229026 519872 229032
rect 519728 228812 519780 228818
rect 519728 228754 519780 228760
rect 518532 227588 518584 227594
rect 518532 227530 518584 227536
rect 519360 225752 519412 225758
rect 519360 225694 519412 225700
rect 518532 222012 518584 222018
rect 518532 221954 518584 221960
rect 518164 221604 518216 221610
rect 518164 221546 518216 221552
rect 517794 221504 517850 221513
rect 517794 221439 517850 221448
rect 517978 221504 518034 221513
rect 517978 221439 518034 221448
rect 517428 219768 517480 219774
rect 517428 219710 517480 219716
rect 517992 219434 518020 221439
rect 517992 219406 518112 219434
rect 518084 217002 518112 219406
rect 518544 217002 518572 221954
rect 519176 219224 519228 219230
rect 518990 219192 519046 219201
rect 518990 219127 519046 219136
rect 519174 219192 519176 219201
rect 519228 219192 519230 219201
rect 519174 219127 519230 219136
rect 518716 218952 518768 218958
rect 518852 218920 518908 218929
rect 518768 218900 518852 218906
rect 518716 218894 518852 218900
rect 518728 218878 518852 218894
rect 518852 218855 518908 218864
rect 518714 218784 518770 218793
rect 518714 218719 518770 218728
rect 518728 218550 518756 218719
rect 518854 218680 518906 218686
rect 518852 218648 518854 218657
rect 518906 218648 518908 218657
rect 518852 218583 518908 218592
rect 518716 218544 518768 218550
rect 518716 218486 518768 218492
rect 519004 218498 519032 219127
rect 519004 218470 519124 218498
rect 519096 218414 519124 218470
rect 519084 218408 519136 218414
rect 519084 218350 519136 218356
rect 519176 217592 519228 217598
rect 519176 217534 519228 217540
rect 519188 217297 519216 217534
rect 518990 217288 519046 217297
rect 518990 217223 519046 217232
rect 519174 217288 519230 217297
rect 519174 217223 519230 217232
rect 519004 217138 519032 217223
rect 519004 217122 519124 217138
rect 519004 217116 519136 217122
rect 519004 217110 519084 217116
rect 519084 217058 519136 217064
rect 519372 217002 519400 225694
rect 519740 221785 519768 228754
rect 520924 228540 520976 228546
rect 520924 228482 520976 228488
rect 519726 221776 519782 221785
rect 519726 221711 519782 221720
rect 516428 216974 516856 217002
rect 517684 216974 518112 217002
rect 518512 216974 518572 217002
rect 519340 216974 519400 217002
rect 519740 217002 519768 221711
rect 520936 217002 520964 228482
rect 521580 220114 521608 230318
rect 521764 227322 521792 231676
rect 522422 231662 522712 231690
rect 522304 230036 522356 230042
rect 522304 229978 522356 229984
rect 521752 227316 521804 227322
rect 521752 227258 521804 227264
rect 521936 223032 521988 223038
rect 521936 222974 521988 222980
rect 521568 220108 521620 220114
rect 521568 220050 521620 220056
rect 521948 217002 521976 222974
rect 522316 222194 522344 229978
rect 522684 223174 522712 231662
rect 523052 230042 523080 231676
rect 523040 230036 523092 230042
rect 523040 229978 523092 229984
rect 522672 223168 522724 223174
rect 522672 223110 522724 223116
rect 523696 223038 523724 231676
rect 524340 226030 524368 231676
rect 524998 231662 525288 231690
rect 525064 229900 525116 229906
rect 525064 229842 525116 229848
rect 524328 226024 524380 226030
rect 524328 225966 524380 225972
rect 523684 223032 523736 223038
rect 523684 222974 523736 222980
rect 523776 222896 523828 222902
rect 523776 222838 523828 222844
rect 522316 222166 522896 222194
rect 522868 220658 522896 222166
rect 522672 220652 522724 220658
rect 522672 220594 522724 220600
rect 522856 220652 522908 220658
rect 522856 220594 522908 220600
rect 522684 219978 522712 220594
rect 522672 219972 522724 219978
rect 522672 219914 522724 219920
rect 522684 217002 522712 219914
rect 523788 217802 523816 222838
rect 523960 221876 524012 221882
rect 523960 221818 524012 221824
rect 523776 217796 523828 217802
rect 523776 217738 523828 217744
rect 523788 217002 523816 217738
rect 519740 216974 520168 217002
rect 520936 216988 520996 217002
rect 520936 216974 521010 216988
rect 521824 216974 521976 217002
rect 522652 216974 522712 217002
rect 523480 216974 523816 217002
rect 523972 217002 524000 221818
rect 525076 221338 525104 229842
rect 525260 229770 525288 231662
rect 525248 229764 525300 229770
rect 525248 229706 525300 229712
rect 525248 224800 525300 224806
rect 525248 224742 525300 224748
rect 525064 221332 525116 221338
rect 525064 221274 525116 221280
rect 525260 218074 525288 224742
rect 525628 224398 525656 231676
rect 526076 229628 526128 229634
rect 526076 229570 526128 229576
rect 526088 224806 526116 229570
rect 526272 228818 526300 231676
rect 526916 230450 526944 231676
rect 526904 230444 526956 230450
rect 526904 230386 526956 230392
rect 526260 228812 526312 228818
rect 526260 228754 526312 228760
rect 526536 228404 526588 228410
rect 526536 228346 526588 228352
rect 526076 224800 526128 224806
rect 526076 224742 526128 224748
rect 525616 224392 525668 224398
rect 525616 224334 525668 224340
rect 526352 223304 526404 223310
rect 526352 223246 526404 223252
rect 525248 218068 525300 218074
rect 525248 218010 525300 218016
rect 525260 217002 525288 218010
rect 525938 217252 525990 217258
rect 525938 217194 525990 217200
rect 523972 216974 524308 217002
rect 525136 216974 525288 217002
rect 525950 216988 525978 217194
rect 526364 217002 526392 223246
rect 526548 217258 526576 228346
rect 527560 225758 527588 231676
rect 527824 229492 527876 229498
rect 527824 229434 527876 229440
rect 527548 225752 527600 225758
rect 527548 225694 527600 225700
rect 527836 221746 527864 229434
rect 528204 228682 528232 231676
rect 528848 229906 528876 231676
rect 529506 231662 529888 231690
rect 528836 229900 528888 229906
rect 528836 229842 528888 229848
rect 528928 229764 528980 229770
rect 528928 229706 528980 229712
rect 528192 228676 528244 228682
rect 528192 228618 528244 228624
rect 528940 227730 528968 229706
rect 528928 227724 528980 227730
rect 528928 227666 528980 227672
rect 528928 225888 528980 225894
rect 528928 225830 528980 225836
rect 528008 224664 528060 224670
rect 528008 224606 528060 224612
rect 527824 221740 527876 221746
rect 527824 221682 527876 221688
rect 527272 220380 527324 220386
rect 527272 220322 527324 220328
rect 527284 218686 527312 220322
rect 527272 218680 527324 218686
rect 527272 218622 527324 218628
rect 526536 217252 526588 217258
rect 526536 217194 526588 217200
rect 527284 217002 527312 218622
rect 528020 217002 528048 224606
rect 528652 218816 528704 218822
rect 528572 218764 528652 218770
rect 528572 218758 528704 218764
rect 528572 218742 528692 218758
rect 528572 218657 528600 218742
rect 528558 218648 528614 218657
rect 528558 218583 528614 218592
rect 528742 218648 528798 218657
rect 528742 218583 528798 218592
rect 528756 218498 528784 218583
rect 528572 218470 528784 218498
rect 528572 218414 528600 218470
rect 528560 218408 528612 218414
rect 528560 218350 528612 218356
rect 528650 217832 528706 217841
rect 528650 217767 528706 217776
rect 528664 217598 528692 217767
rect 528284 217592 528336 217598
rect 528284 217534 528336 217540
rect 528652 217592 528704 217598
rect 528652 217534 528704 217540
rect 528296 217297 528324 217534
rect 528282 217288 528338 217297
rect 528282 217223 528338 217232
rect 528466 217288 528522 217297
rect 528466 217223 528522 217232
rect 528480 217122 528508 217223
rect 528468 217116 528520 217122
rect 528468 217058 528520 217064
rect 528940 217002 528968 225830
rect 529860 221882 529888 231662
rect 530136 225894 530164 231676
rect 530308 230240 530360 230246
rect 530308 230182 530360 230188
rect 530124 225888 530176 225894
rect 530124 225830 530176 225836
rect 530320 223310 530348 230182
rect 530780 229634 530808 231676
rect 530768 229628 530820 229634
rect 530768 229570 530820 229576
rect 531424 228546 531452 231676
rect 531412 228540 531464 228546
rect 531412 228482 531464 228488
rect 530584 225616 530636 225622
rect 530584 225558 530636 225564
rect 530308 223304 530360 223310
rect 530308 223246 530360 223252
rect 529848 221876 529900 221882
rect 529848 221818 529900 221824
rect 530032 221604 530084 221610
rect 530032 221546 530084 221552
rect 530044 220386 530072 221546
rect 530596 221134 530624 225558
rect 532068 224534 532096 231676
rect 532712 230314 532740 231676
rect 533370 231662 533752 231690
rect 532700 230308 532752 230314
rect 532700 230250 532752 230256
rect 533528 230172 533580 230178
rect 533528 230114 533580 230120
rect 533540 229906 533568 230114
rect 533528 229900 533580 229906
rect 533528 229842 533580 229848
rect 533528 228268 533580 228274
rect 533528 228210 533580 228216
rect 531780 224528 531832 224534
rect 531780 224470 531832 224476
rect 532056 224528 532108 224534
rect 532056 224470 532108 224476
rect 530584 221128 530636 221134
rect 530584 221070 530636 221076
rect 530032 220380 530084 220386
rect 530032 220322 530084 220328
rect 529110 217832 529166 217841
rect 529110 217767 529112 217776
rect 529164 217767 529166 217776
rect 529112 217738 529164 217744
rect 530044 217002 530072 220322
rect 530596 217002 530624 221070
rect 531792 217002 531820 224470
rect 532148 223440 532200 223446
rect 532148 223382 532200 223388
rect 532160 219026 532188 223382
rect 532884 220652 532936 220658
rect 532884 220594 532936 220600
rect 533344 220652 533396 220658
rect 533344 220594 533396 220600
rect 532698 220416 532754 220425
rect 532896 220386 532924 220594
rect 532698 220351 532700 220360
rect 532752 220351 532754 220360
rect 532884 220380 532936 220386
rect 532700 220322 532752 220328
rect 532884 220322 532936 220328
rect 533356 219978 533384 220594
rect 533344 219972 533396 219978
rect 533344 219914 533396 219920
rect 532148 219020 532200 219026
rect 532148 218962 532200 218968
rect 532608 219020 532660 219026
rect 532608 218962 532660 218968
rect 531964 218952 532016 218958
rect 531964 218894 532016 218900
rect 531976 218482 532004 218894
rect 531964 218476 532016 218482
rect 531964 218418 532016 218424
rect 532620 217002 532648 218962
rect 533344 218340 533396 218346
rect 533344 218282 533396 218288
rect 533356 218074 533384 218282
rect 533344 218068 533396 218074
rect 533344 218010 533396 218016
rect 533540 217002 533568 228210
rect 533724 222902 533752 231662
rect 534000 227186 534028 231676
rect 534644 229906 534672 231676
rect 534816 230036 534868 230042
rect 534816 229978 534868 229984
rect 534632 229900 534684 229906
rect 534632 229842 534684 229848
rect 533988 227180 534040 227186
rect 533988 227122 534040 227128
rect 534448 224256 534500 224262
rect 534448 224198 534500 224204
rect 533712 222896 533764 222902
rect 533712 222838 533764 222844
rect 534170 220416 534226 220425
rect 534034 220380 534086 220386
rect 534170 220351 534172 220360
rect 534034 220322 534086 220328
rect 534224 220351 534226 220360
rect 534172 220322 534224 220328
rect 534046 220266 534074 220322
rect 534046 220238 534120 220266
rect 534092 219978 534120 220238
rect 534080 219972 534132 219978
rect 534080 219914 534132 219920
rect 534264 218816 534316 218822
rect 534264 218758 534316 218764
rect 534276 218657 534304 218758
rect 534078 218648 534134 218657
rect 534078 218583 534134 218592
rect 534262 218648 534318 218657
rect 534262 218583 534318 218592
rect 534092 218498 534120 218583
rect 534092 218470 534212 218498
rect 534184 218346 534212 218470
rect 534172 218340 534224 218346
rect 534172 218282 534224 218288
rect 534264 217592 534316 217598
rect 534264 217534 534316 217540
rect 534276 217297 534304 217534
rect 534078 217288 534134 217297
rect 534078 217223 534134 217232
rect 534262 217288 534318 217297
rect 534262 217223 534318 217232
rect 533712 217116 533764 217122
rect 533712 217058 533764 217064
rect 533724 217002 533752 217058
rect 526364 216974 526792 217002
rect 527284 216974 527620 217002
rect 528020 216988 528448 217002
rect 528020 216974 528462 216988
rect 528940 216974 529276 217002
rect 530044 216974 530104 217002
rect 530596 216974 530932 217002
rect 531760 216974 531820 217002
rect 532588 216974 532648 217002
rect 533416 216974 533752 217002
rect 501326 216951 501382 216960
rect 495162 216744 495218 216753
rect 520982 216730 521010 216974
rect 528434 216866 528462 216974
rect 528434 216852 528600 216866
rect 528448 216850 528600 216852
rect 528448 216844 528612 216850
rect 528448 216838 528560 216844
rect 528560 216786 528612 216792
rect 495218 216702 495328 216730
rect 520982 216716 521332 216730
rect 520996 216714 521332 216716
rect 520996 216708 521344 216714
rect 520996 216702 521292 216708
rect 495162 216679 495218 216688
rect 521292 216650 521344 216656
rect 534092 216578 534120 217223
rect 534460 217002 534488 224198
rect 534828 221610 534856 229978
rect 535288 224262 535316 231676
rect 535460 226160 535512 226166
rect 535460 226102 535512 226108
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 534816 221604 534868 221610
rect 534816 221546 534868 221552
rect 535092 221332 535144 221338
rect 535092 221274 535144 221280
rect 535104 217002 535132 221274
rect 535472 219366 535500 226102
rect 535932 225622 535960 231676
rect 536576 229770 536604 231676
rect 536564 229764 536616 229770
rect 536564 229706 536616 229712
rect 537220 227050 537248 231676
rect 537484 230444 537536 230450
rect 537484 230386 537536 230392
rect 536104 227044 536156 227050
rect 536104 226986 536156 226992
rect 537208 227044 537260 227050
rect 537208 226986 537260 226992
rect 535920 225616 535972 225622
rect 535920 225558 535972 225564
rect 536116 224954 536144 226986
rect 536024 224926 536144 224954
rect 535460 219360 535512 219366
rect 535460 219302 535512 219308
rect 536024 217258 536052 224926
rect 537116 224800 537168 224806
rect 537116 224742 537168 224748
rect 536380 219360 536432 219366
rect 536380 219302 536432 219308
rect 536012 217252 536064 217258
rect 536012 217194 536064 217200
rect 536024 217002 536052 217194
rect 534244 216974 534488 217002
rect 535072 216974 535132 217002
rect 535900 216974 536052 217002
rect 536392 217002 536420 219302
rect 537128 219162 537156 224742
rect 537300 219972 537352 219978
rect 537300 219914 537352 219920
rect 537312 219366 537340 219914
rect 537496 219910 537524 230386
rect 537864 228410 537892 231676
rect 538508 230042 538536 231676
rect 538692 231662 539166 231690
rect 538496 230036 538548 230042
rect 538496 229978 538548 229984
rect 537852 228404 537904 228410
rect 537852 228346 537904 228352
rect 538496 227452 538548 227458
rect 538496 227394 538548 227400
rect 537484 219904 537536 219910
rect 537484 219846 537536 219852
rect 537300 219360 537352 219366
rect 537300 219302 537352 219308
rect 537116 219156 537168 219162
rect 537116 219098 537168 219104
rect 537128 217002 537156 219098
rect 537852 218884 537904 218890
rect 537852 218826 537904 218832
rect 537864 218074 537892 218826
rect 537852 218068 537904 218074
rect 537852 218010 537904 218016
rect 538508 217462 538536 227394
rect 538692 221474 538720 231662
rect 547144 230308 547196 230314
rect 547144 230250 547196 230256
rect 543924 230172 543976 230178
rect 543924 230114 543976 230120
rect 540244 229628 540296 229634
rect 540244 229570 540296 229576
rect 540060 228948 540112 228954
rect 540060 228890 540112 228896
rect 540072 221474 540100 228890
rect 538680 221468 538732 221474
rect 538680 221410 538732 221416
rect 540060 221468 540112 221474
rect 540060 221410 540112 221416
rect 540256 219774 540284 229570
rect 543188 229084 543240 229090
rect 543188 229026 543240 229032
rect 541624 227588 541676 227594
rect 541624 227530 541676 227536
rect 540888 221468 540940 221474
rect 540888 221410 540940 221416
rect 539048 219768 539100 219774
rect 539048 219710 539100 219716
rect 540244 219768 540296 219774
rect 540244 219710 540296 219716
rect 538864 219020 538916 219026
rect 538864 218962 538916 218968
rect 538876 218618 538904 218962
rect 538864 218612 538916 218618
rect 538864 218554 538916 218560
rect 538496 217456 538548 217462
rect 538496 217398 538548 217404
rect 538508 217002 538536 217398
rect 536392 216974 536728 217002
rect 537128 216974 537556 217002
rect 538384 216974 538536 217002
rect 539060 217002 539088 219710
rect 539692 219360 539744 219366
rect 539692 219302 539744 219308
rect 539232 219156 539284 219162
rect 539232 219098 539284 219104
rect 539244 218346 539272 219098
rect 539232 218340 539284 218346
rect 539232 218282 539284 218288
rect 539704 217002 539732 219302
rect 540900 217002 540928 221410
rect 539060 216974 539212 217002
rect 539704 216988 540040 217002
rect 539704 216974 540054 216988
rect 540868 216974 540928 217002
rect 541636 217002 541664 227530
rect 542452 221740 542504 221746
rect 542452 221682 542504 221688
rect 542464 219026 542492 221682
rect 542452 219020 542504 219026
rect 542452 218962 542504 218968
rect 542464 217002 542492 218962
rect 543200 217870 543228 229026
rect 543936 223446 543964 230114
rect 545764 227316 545816 227322
rect 545764 227258 545816 227264
rect 543924 223440 543976 223446
rect 543924 223382 543976 223388
rect 544936 223304 544988 223310
rect 544936 223246 544988 223252
rect 543556 221332 543608 221338
rect 543556 221274 543608 221280
rect 543372 220108 543424 220114
rect 543372 220050 543424 220056
rect 543384 219366 543412 220050
rect 543568 219994 543596 221274
rect 543922 220280 543978 220289
rect 543922 220215 543978 220224
rect 543568 219966 543780 219994
rect 543752 219910 543780 219966
rect 543740 219904 543792 219910
rect 543740 219846 543792 219852
rect 543372 219360 543424 219366
rect 543372 219302 543424 219308
rect 543740 219156 543792 219162
rect 543740 219098 543792 219104
rect 543752 218090 543780 219098
rect 543936 218890 543964 220215
rect 544948 220017 544976 223246
rect 544934 220008 544990 220017
rect 544934 219943 544990 219952
rect 544292 219360 544344 219366
rect 544292 219302 544344 219308
rect 543924 218884 543976 218890
rect 543924 218826 543976 218832
rect 544108 218884 544160 218890
rect 544108 218826 544160 218832
rect 544120 218226 544148 218826
rect 543936 218210 544148 218226
rect 543924 218204 544148 218210
rect 543976 218198 544148 218204
rect 543924 218146 543976 218152
rect 543706 218074 543780 218090
rect 544108 218136 544160 218142
rect 544108 218078 544160 218084
rect 543694 218068 543780 218074
rect 543746 218062 543780 218068
rect 543694 218010 543746 218016
rect 543832 218000 543884 218006
rect 543832 217942 543884 217948
rect 543188 217864 543240 217870
rect 543188 217806 543240 217812
rect 543200 217410 543228 217806
rect 543844 217598 543872 217942
rect 544120 217734 544148 218078
rect 544108 217728 544160 217734
rect 544108 217670 544160 217676
rect 543464 217592 543516 217598
rect 543464 217534 543516 217540
rect 543832 217592 543884 217598
rect 543832 217534 543884 217540
rect 543108 217382 543228 217410
rect 543108 217002 543136 217382
rect 543476 217297 543504 217534
rect 543462 217288 543518 217297
rect 543462 217223 543518 217232
rect 543646 217288 543702 217297
rect 543646 217223 543702 217232
rect 541636 216974 541696 217002
rect 542464 216974 542524 217002
rect 543108 216974 543352 217002
rect 534080 216572 534132 216578
rect 534080 216514 534132 216520
rect 540026 216458 540054 216974
rect 543660 216578 543688 217223
rect 544304 217002 544332 219302
rect 544180 216974 544332 217002
rect 544948 217002 544976 219943
rect 545776 217598 545804 227258
rect 546776 223168 546828 223174
rect 546776 223110 546828 223116
rect 546788 222194 546816 223110
rect 546788 222166 546908 222194
rect 546316 219292 546368 219298
rect 546316 219234 546368 219240
rect 546328 218482 546356 219234
rect 546880 219144 546908 222166
rect 547156 222154 547184 230250
rect 555436 230178 555464 255546
rect 556804 251252 556856 251258
rect 556804 251194 556856 251200
rect 555424 230172 555476 230178
rect 555424 230114 555476 230120
rect 555240 229900 555292 229906
rect 555240 229842 555292 229848
rect 551192 228812 551244 228818
rect 551192 228754 551244 228760
rect 549904 227724 549956 227730
rect 549904 227666 549956 227672
rect 547880 226024 547932 226030
rect 547880 225966 547932 225972
rect 547144 222148 547196 222154
rect 547144 222090 547196 222096
rect 547420 221604 547472 221610
rect 547420 221546 547472 221552
rect 547142 220280 547198 220289
rect 547142 220215 547198 220224
rect 546788 219116 546908 219144
rect 546592 219020 546644 219026
rect 546592 218962 546644 218968
rect 546604 218482 546632 218962
rect 546316 218476 546368 218482
rect 546316 218418 546368 218424
rect 546592 218476 546644 218482
rect 546592 218418 546644 218424
rect 545764 217592 545816 217598
rect 545764 217534 545816 217540
rect 545776 217002 545804 217534
rect 546788 217002 546816 219116
rect 546960 219020 547012 219026
rect 546960 218962 547012 218968
rect 546972 218754 547000 218962
rect 547156 218754 547184 220215
rect 546960 218748 547012 218754
rect 546960 218690 547012 218696
rect 547144 218748 547196 218754
rect 547144 218690 547196 218696
rect 544948 216974 545008 217002
rect 545776 216974 545836 217002
rect 546664 216974 546816 217002
rect 547432 217002 547460 221546
rect 547892 221270 547920 225966
rect 548156 223032 548208 223038
rect 548156 222974 548208 222980
rect 547880 221264 547932 221270
rect 547880 221206 547932 221212
rect 548168 217002 548196 222974
rect 549076 221264 549128 221270
rect 549076 221206 549128 221212
rect 548338 220688 548394 220697
rect 548338 220623 548394 220632
rect 548352 220114 548380 220623
rect 548340 220108 548392 220114
rect 548340 220050 548392 220056
rect 548524 220040 548576 220046
rect 548524 219982 548576 219988
rect 548536 219774 548564 219982
rect 548524 219768 548576 219774
rect 548524 219710 548576 219716
rect 548892 217864 548944 217870
rect 548628 217812 548892 217818
rect 548628 217806 548944 217812
rect 548628 217790 548932 217806
rect 548628 217002 548656 217790
rect 547432 216974 547828 217002
rect 548168 216974 548656 217002
rect 549088 217002 549116 221206
rect 549916 219774 549944 227666
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 550652 221270 550680 224334
rect 550640 221264 550692 221270
rect 550640 221206 550692 221212
rect 549904 219768 549956 219774
rect 549904 219710 549956 219716
rect 549916 217002 549944 219710
rect 550652 217002 550680 221206
rect 551204 217002 551232 228754
rect 553676 228676 553728 228682
rect 553676 228618 553728 228624
rect 553308 225752 553360 225758
rect 553308 225694 553360 225700
rect 553320 224954 553348 225694
rect 553228 224926 553348 224954
rect 553688 224954 553716 228618
rect 553688 224926 554452 224954
rect 553228 221746 553256 224926
rect 553216 221740 553268 221746
rect 553044 221700 553216 221728
rect 552664 221604 552716 221610
rect 552664 221546 552716 221552
rect 552386 220688 552442 220697
rect 552386 220623 552442 220632
rect 552400 217002 552428 220623
rect 552676 218754 552704 221546
rect 552846 220280 552902 220289
rect 552846 220215 552902 220224
rect 552860 219026 552888 220215
rect 552848 219020 552900 219026
rect 552848 218962 552900 218968
rect 553044 218872 553072 221700
rect 553216 221682 553268 221688
rect 553676 221604 553728 221610
rect 553676 221546 553728 221552
rect 553860 221604 553912 221610
rect 553860 221546 553912 221552
rect 553688 220425 553716 221546
rect 553674 220416 553730 220425
rect 553674 220351 553730 220360
rect 553872 220046 553900 221546
rect 554042 220688 554098 220697
rect 554042 220623 554098 220632
rect 554056 220046 554084 220623
rect 553860 220040 553912 220046
rect 553352 220008 553408 220017
rect 553860 219982 553912 219988
rect 554044 220040 554096 220046
rect 554044 219982 554096 219988
rect 553352 219943 553408 219952
rect 553366 219774 553394 219943
rect 553216 219768 553268 219774
rect 553216 219710 553268 219716
rect 553354 219768 553406 219774
rect 553354 219710 553406 219716
rect 553228 218872 553256 219710
rect 553492 219292 553544 219298
rect 553492 219234 553544 219240
rect 553504 219026 553532 219234
rect 553952 219224 554004 219230
rect 553952 219166 554004 219172
rect 553492 219020 553544 219026
rect 553492 218962 553544 218968
rect 553768 218884 553820 218890
rect 553044 218844 553164 218872
rect 553228 218844 553302 218872
rect 552664 218748 552716 218754
rect 552664 218690 552716 218696
rect 553136 217002 553164 218844
rect 553274 218754 553302 218844
rect 553964 218872 553992 219166
rect 554228 219020 554280 219026
rect 554228 218962 554280 218968
rect 553820 218844 553992 218872
rect 553768 218826 553820 218832
rect 553262 218748 553314 218754
rect 553262 218690 553314 218696
rect 554240 218498 554268 218962
rect 554056 218470 554268 218498
rect 554056 218385 554084 218470
rect 554042 218376 554098 218385
rect 554042 218311 554098 218320
rect 554226 218376 554282 218385
rect 554226 218311 554282 218320
rect 554240 218142 554268 218311
rect 554228 218136 554280 218142
rect 554228 218078 554280 218084
rect 554424 217002 554452 224926
rect 554872 223440 554924 223446
rect 554872 223382 554924 223388
rect 554594 220280 554650 220289
rect 554594 220215 554650 220224
rect 549088 216974 549148 217002
rect 549916 216974 549976 217002
rect 550652 216974 550804 217002
rect 551204 216974 551632 217002
rect 552400 216974 552460 217002
rect 553136 216974 553288 217002
rect 554116 216974 554452 217002
rect 547800 216578 547828 216974
rect 554608 216578 554636 220215
rect 554884 217002 554912 223382
rect 555252 222426 555280 229842
rect 556160 225888 556212 225894
rect 556160 225830 556212 225836
rect 555240 222420 555292 222426
rect 555240 222362 555292 222368
rect 555700 221876 555752 221882
rect 555700 221818 555752 221824
rect 555712 218006 555740 221818
rect 555700 218000 555752 218006
rect 555700 217942 555752 217948
rect 555712 217002 555740 217942
rect 556172 217002 556200 225830
rect 556816 225758 556844 251194
rect 558196 236094 558224 265610
rect 645872 261526 645900 277766
rect 647252 265674 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 265668 647292 265674
rect 647240 265610 647292 265616
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 565084 259480 565136 259486
rect 565084 259422 565136 259428
rect 560944 256760 560996 256766
rect 560944 256702 560996 256708
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 559564 230036 559616 230042
rect 559564 229978 559616 229984
rect 558184 228540 558236 228546
rect 558184 228482 558236 228488
rect 556804 225752 556856 225758
rect 556804 225694 556856 225700
rect 558196 222154 558224 228482
rect 558920 224528 558972 224534
rect 558920 224470 558972 224476
rect 558000 222148 558052 222154
rect 558000 222090 558052 222096
rect 558184 222148 558236 222154
rect 558184 222090 558236 222096
rect 558012 221610 558040 222090
rect 557080 221604 557132 221610
rect 557080 221546 557132 221552
rect 558000 221604 558052 221610
rect 558000 221546 558052 221552
rect 557092 217002 557120 221546
rect 558196 217002 558224 222090
rect 558932 217002 558960 224470
rect 559576 221882 559604 229978
rect 560956 227594 560984 256702
rect 563704 252612 563756 252618
rect 563704 252554 563756 252560
rect 562324 229764 562376 229770
rect 562324 229706 562376 229712
rect 560944 227588 560996 227594
rect 560944 227530 560996 227536
rect 561496 227180 561548 227186
rect 561496 227122 561548 227128
rect 560668 222896 560720 222902
rect 560668 222838 560720 222844
rect 559564 221876 559616 221882
rect 559564 221818 559616 221824
rect 559840 221604 559892 221610
rect 559840 221546 559892 221552
rect 559852 217002 559880 221546
rect 560680 217002 560708 222838
rect 561508 217002 561536 227122
rect 562140 222420 562192 222426
rect 562140 222362 562192 222368
rect 562152 217002 562180 222362
rect 562336 222057 562364 229706
rect 563716 223650 563744 252554
rect 564716 225616 564768 225622
rect 564716 225558 564768 225564
rect 563980 224256 564032 224262
rect 563980 224198 564032 224204
rect 563704 223644 563756 223650
rect 563704 223586 563756 223592
rect 562968 222896 563020 222902
rect 562968 222838 563020 222844
rect 562980 222442 563008 222838
rect 563992 222698 564020 224198
rect 563980 222692 564032 222698
rect 563980 222634 564032 222640
rect 562980 222414 563192 222442
rect 562874 222320 562930 222329
rect 562874 222255 562930 222264
rect 562888 222154 562916 222255
rect 562876 222148 562928 222154
rect 562876 222090 562928 222096
rect 562322 222048 562378 222057
rect 562322 221983 562378 221992
rect 562690 222048 562746 222057
rect 562690 221983 562692 221992
rect 562744 221983 562746 221992
rect 562692 221954 562744 221960
rect 563164 221762 563192 222414
rect 563334 222320 563390 222329
rect 563334 222255 563390 222264
rect 563348 222194 563376 222255
rect 563348 222166 563744 222194
rect 563518 222048 563574 222057
rect 563518 221983 563520 221992
rect 563572 221983 563574 221992
rect 563520 221954 563572 221960
rect 563336 221876 563388 221882
rect 563336 221818 563388 221824
rect 563348 221762 563376 221818
rect 563164 221734 563376 221762
rect 563716 221610 563744 222166
rect 563152 221604 563204 221610
rect 563152 221546 563204 221552
rect 563704 221604 563756 221610
rect 563704 221546 563756 221552
rect 563164 220674 563192 221546
rect 563992 220814 564020 222634
rect 564728 220814 564756 225558
rect 565096 222426 565124 259422
rect 566188 228404 566240 228410
rect 566188 228346 566240 228352
rect 565360 227044 565412 227050
rect 565360 226986 565412 226992
rect 565084 222420 565136 222426
rect 565084 222362 565136 222368
rect 564898 222320 564954 222329
rect 564898 222255 564954 222264
rect 564912 222154 564940 222255
rect 565372 222154 565400 226986
rect 564900 222148 564952 222154
rect 564900 222090 564952 222096
rect 565360 222148 565412 222154
rect 565360 222090 565412 222096
rect 565082 222048 565138 222057
rect 565082 221983 565138 221992
rect 563992 220786 564388 220814
rect 564728 220786 565032 220814
rect 563426 220688 563482 220697
rect 563164 220646 563426 220674
rect 563426 220623 563482 220632
rect 563242 220552 563298 220561
rect 563298 220510 563468 220538
rect 563242 220487 563298 220496
rect 562876 220040 562928 220046
rect 562876 219982 562928 219988
rect 563244 220040 563296 220046
rect 563244 219982 563296 219988
rect 562888 219722 562916 219982
rect 562888 219694 563100 219722
rect 563072 219638 563100 219694
rect 562876 219632 562928 219638
rect 562876 219574 562928 219580
rect 563060 219632 563112 219638
rect 563060 219574 563112 219580
rect 562888 219366 562916 219574
rect 563256 219366 563284 219982
rect 563440 219366 563468 220510
rect 563794 220416 563850 220425
rect 563794 220351 563850 220360
rect 563610 220144 563666 220153
rect 563610 220079 563666 220088
rect 562508 219360 562560 219366
rect 562508 219302 562560 219308
rect 562876 219360 562928 219366
rect 562876 219302 562928 219308
rect 563244 219360 563296 219366
rect 563244 219302 563296 219308
rect 563428 219360 563480 219366
rect 563428 219302 563480 219308
rect 554884 216988 554944 217002
rect 554884 216974 554958 216988
rect 555712 216974 555772 217002
rect 556172 216974 556600 217002
rect 557092 216974 557488 217002
rect 558196 216974 558256 217002
rect 558932 216974 559084 217002
rect 559852 216974 559912 217002
rect 560680 216974 560740 217002
rect 561508 216974 561568 217002
rect 562152 216974 562396 217002
rect 554930 216594 554958 216974
rect 554930 216580 555096 216594
rect 554944 216578 555096 216580
rect 543648 216572 543700 216578
rect 543648 216514 543700 216520
rect 547788 216572 547840 216578
rect 547788 216514 547840 216520
rect 554596 216572 554648 216578
rect 554944 216572 555108 216578
rect 554944 216566 555056 216572
rect 554596 216514 554648 216520
rect 555056 216514 555108 216520
rect 540150 216472 540206 216481
rect 540026 216444 540150 216458
rect 540040 216430 540150 216444
rect 540150 216407 540206 216416
rect 557078 216472 557134 216481
rect 557460 216458 557488 216974
rect 557722 216472 557778 216481
rect 557460 216430 557722 216458
rect 557078 216407 557080 216416
rect 557132 216407 557134 216416
rect 557722 216407 557778 216416
rect 558550 216472 558606 216481
rect 562520 216442 562548 219302
rect 563624 219230 563652 220079
rect 563612 219224 563664 219230
rect 563612 219166 563664 219172
rect 563808 219042 563836 220351
rect 564070 219906 564126 219915
rect 564070 219841 564126 219850
rect 562704 219014 563836 219042
rect 562704 216578 562732 219014
rect 564084 218906 564112 219841
rect 562888 218890 564112 218906
rect 562876 218884 564112 218890
rect 562928 218878 564112 218884
rect 562876 218826 562928 218832
rect 563198 218476 563250 218482
rect 563250 218436 563376 218464
rect 563198 218418 563250 218424
rect 563348 216578 563376 218436
rect 563612 218272 563664 218278
rect 563612 218214 563664 218220
rect 563624 218006 563652 218214
rect 563612 218000 563664 218006
rect 563612 217942 563664 217948
rect 563796 218000 563848 218006
rect 563796 217942 563848 217948
rect 563808 217598 563836 217942
rect 563796 217592 563848 217598
rect 563796 217534 563848 217540
rect 564360 217274 564388 220786
rect 564622 220144 564678 220153
rect 564678 220102 564848 220130
rect 564622 220079 564678 220088
rect 564820 218278 564848 220102
rect 564532 218272 564584 218278
rect 564532 218214 564584 218220
rect 564808 218272 564860 218278
rect 564808 218214 564860 218220
rect 564544 217598 564572 218214
rect 564532 217592 564584 217598
rect 564532 217534 564584 217540
rect 563624 217246 564388 217274
rect 562692 216572 562744 216578
rect 562692 216514 562744 216520
rect 563336 216572 563388 216578
rect 563336 216514 563388 216520
rect 563624 216458 563652 217246
rect 565004 217138 565032 220786
rect 564452 217110 565032 217138
rect 564452 217002 564480 217110
rect 565096 217002 565124 221983
rect 564052 216974 564480 217002
rect 564880 216974 565124 217002
rect 565372 217002 565400 222090
rect 566200 217002 566228 228346
rect 567660 227588 567712 227594
rect 567660 227530 567712 227536
rect 567672 224954 567700 227530
rect 568592 224954 568620 260850
rect 570616 234598 570644 261462
rect 632704 246356 632756 246362
rect 632704 246298 632756 246304
rect 598204 245676 598256 245682
rect 598204 245618 598256 245624
rect 587164 242208 587216 242214
rect 587164 242150 587216 242156
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 571340 230172 571392 230178
rect 571340 230114 571392 230120
rect 571352 229094 571380 230114
rect 571352 229066 571472 229094
rect 570696 225752 570748 225758
rect 570696 225694 570748 225700
rect 567672 224926 567792 224954
rect 568592 224926 569448 224954
rect 567198 222320 567254 222329
rect 567198 222255 567254 222264
rect 567212 217002 567240 222255
rect 567764 217002 567792 224926
rect 568672 222420 568724 222426
rect 568672 222362 568724 222368
rect 568684 217002 568712 222362
rect 569420 217002 569448 224926
rect 570328 223032 570380 223038
rect 570328 222974 570380 222980
rect 570144 222420 570196 222426
rect 570144 222362 570196 222368
rect 570156 219230 570184 222362
rect 570144 219224 570196 219230
rect 570144 219166 570196 219172
rect 570340 218754 570368 222974
rect 570510 222592 570566 222601
rect 570510 222527 570566 222536
rect 570524 219774 570552 222527
rect 570512 219768 570564 219774
rect 570512 219710 570564 219716
rect 570328 218748 570380 218754
rect 570328 218690 570380 218696
rect 570708 217002 570736 225694
rect 571248 223644 571300 223650
rect 571248 223586 571300 223592
rect 571062 222048 571118 222057
rect 571062 221983 571118 221992
rect 570878 219906 570934 219915
rect 570878 219841 570934 219850
rect 570892 218414 570920 219841
rect 571076 219722 571104 221983
rect 570984 219694 571104 219722
rect 570984 218770 571012 219694
rect 571260 219042 571288 223586
rect 571444 222902 571472 229066
rect 575388 223032 575440 223038
rect 575388 222974 575440 222980
rect 571432 222896 571484 222902
rect 571432 222838 571484 222844
rect 571892 222896 571944 222902
rect 571892 222838 571944 222844
rect 571432 219156 571484 219162
rect 571432 219098 571484 219104
rect 571260 219014 571380 219042
rect 570984 218742 571288 218770
rect 570880 218408 570932 218414
rect 570880 218350 570932 218356
rect 571064 218408 571116 218414
rect 571064 218350 571116 218356
rect 565372 216974 565708 217002
rect 566200 216974 566536 217002
rect 567212 216974 567364 217002
rect 567764 216974 568192 217002
rect 568684 216974 569020 217002
rect 569420 216974 569848 217002
rect 570676 216974 570736 217002
rect 558550 216407 558552 216416
rect 557080 216378 557132 216384
rect 558604 216407 558606 216416
rect 562508 216436 562560 216442
rect 558552 216378 558604 216384
rect 563224 216430 563652 216458
rect 571076 216442 571104 218350
rect 571260 216442 571288 218742
rect 571352 217002 571380 219014
rect 571444 218770 571472 219098
rect 571904 219042 571932 222838
rect 574652 222692 574704 222698
rect 574652 222634 574704 222640
rect 572260 222556 572312 222562
rect 572260 222498 572312 222504
rect 572076 220040 572128 220046
rect 572076 219982 572128 219988
rect 572088 219212 572116 219982
rect 572272 219416 572300 222498
rect 574468 222420 574520 222426
rect 574468 222362 574520 222368
rect 572442 222320 572498 222329
rect 572442 222255 572498 222264
rect 572456 221082 572484 222255
rect 572456 221054 572576 221082
rect 572548 220674 572576 221054
rect 572456 220646 572576 220674
rect 572824 220646 574232 220674
rect 572456 219722 572484 220646
rect 572626 220552 572682 220561
rect 572626 220487 572682 220496
rect 572640 220114 572668 220487
rect 572824 220289 572852 220646
rect 572810 220280 572866 220289
rect 572810 220215 572866 220224
rect 573454 220280 573510 220289
rect 573454 220215 573510 220224
rect 573914 220280 573970 220289
rect 573914 220215 573970 220224
rect 572628 220108 572680 220114
rect 572628 220050 572680 220056
rect 573270 220008 573326 220017
rect 572640 219966 573270 219994
rect 572640 219910 572668 219966
rect 573270 219943 573326 219952
rect 572628 219904 572680 219910
rect 572628 219846 572680 219852
rect 572812 219904 572864 219910
rect 572812 219846 572864 219852
rect 572824 219722 572852 219846
rect 572456 219694 572852 219722
rect 572272 219388 572576 219416
rect 572548 219348 572576 219388
rect 573468 219366 573496 220215
rect 573180 219360 573232 219366
rect 572548 219320 572668 219348
rect 572352 219224 572404 219230
rect 572088 219184 572352 219212
rect 572352 219166 572404 219172
rect 572352 219088 572404 219094
rect 571904 219014 572116 219042
rect 572640 219076 572668 219320
rect 573180 219302 573232 219308
rect 573456 219360 573508 219366
rect 573456 219302 573508 219308
rect 572996 219088 573048 219094
rect 572640 219048 572996 219076
rect 572352 219030 572404 219036
rect 572996 219030 573048 219036
rect 571800 218952 571852 218958
rect 571800 218894 571852 218900
rect 571812 218770 571840 218894
rect 571444 218742 571840 218770
rect 572088 218634 572116 219014
rect 571444 218606 572116 218634
rect 571444 217138 571472 218606
rect 572364 218385 572392 219030
rect 573192 218958 573220 219302
rect 573928 219178 573956 220215
rect 573928 219150 574048 219178
rect 572536 218952 572588 218958
rect 572536 218894 572588 218900
rect 573180 218952 573232 218958
rect 573180 218894 573232 218900
rect 572548 218618 572576 218894
rect 572536 218612 572588 218618
rect 572536 218554 572588 218560
rect 574020 218498 574048 219150
rect 573088 218476 573140 218482
rect 573088 218418 573140 218424
rect 573928 218470 574048 218498
rect 572350 218376 572406 218385
rect 572350 218311 572406 218320
rect 571800 218272 571852 218278
rect 571852 218220 572576 218226
rect 571800 218214 572576 218220
rect 571812 218198 572576 218214
rect 572548 218113 572576 218198
rect 572904 218136 572956 218142
rect 572534 218104 572590 218113
rect 572904 218078 572956 218084
rect 572534 218039 572590 218048
rect 572916 217841 572944 218078
rect 573100 217988 573128 218418
rect 573928 218346 573956 218470
rect 573732 218340 573784 218346
rect 573732 218282 573784 218288
rect 573916 218340 573968 218346
rect 573916 218282 573968 218288
rect 573744 218054 573772 218282
rect 573744 218026 574140 218054
rect 573272 218000 573324 218006
rect 573100 217960 573272 217988
rect 573272 217942 573324 217948
rect 571890 217832 571946 217841
rect 571890 217767 571946 217776
rect 572166 217832 572222 217841
rect 572166 217767 572222 217776
rect 572902 217832 572958 217841
rect 572902 217767 572958 217776
rect 571904 217682 571932 217767
rect 572180 217682 572208 217767
rect 571904 217654 572024 217682
rect 572180 217654 572852 217682
rect 571996 217138 572024 217654
rect 572824 217598 572852 217654
rect 572260 217592 572312 217598
rect 572260 217534 572312 217540
rect 572812 217592 572864 217598
rect 572812 217534 572864 217540
rect 572272 217274 572300 217534
rect 572272 217246 573312 217274
rect 571444 217110 571932 217138
rect 571996 217110 573220 217138
rect 571904 217002 571932 217110
rect 571352 216974 571504 217002
rect 571904 216974 572332 217002
rect 572996 216980 573048 216986
rect 572996 216922 573048 216928
rect 573008 216594 573036 216922
rect 573192 216730 573220 217110
rect 573284 216832 573312 217246
rect 573456 216844 573508 216850
rect 573284 216804 573456 216832
rect 573456 216786 573508 216792
rect 573192 216702 573956 216730
rect 573008 216566 573864 216594
rect 571064 216436 571116 216442
rect 562508 216378 562560 216384
rect 571064 216378 571116 216384
rect 571248 216436 571300 216442
rect 571248 216378 571300 216384
rect 573836 213364 573864 216566
rect 573928 213500 573956 216702
rect 574112 215830 574140 218026
rect 574204 215914 574232 220646
rect 574204 215886 574324 215914
rect 574100 215824 574152 215830
rect 574100 215766 574152 215772
rect 574296 215150 574324 215886
rect 574284 215144 574336 215150
rect 574284 215086 574336 215092
rect 574480 214742 574508 222362
rect 574664 218482 574692 222634
rect 574834 222592 574890 222601
rect 574834 222527 574890 222536
rect 574848 219774 574876 222527
rect 575202 220688 575258 220697
rect 575202 220623 575258 220632
rect 574836 219768 574888 219774
rect 574836 219710 574888 219716
rect 574836 219360 574888 219366
rect 574836 219302 574888 219308
rect 574652 218476 574704 218482
rect 574652 218418 574704 218424
rect 574652 218000 574704 218006
rect 574652 217942 574704 217948
rect 574664 216374 574692 217942
rect 574652 216368 574704 216374
rect 574652 216310 574704 216316
rect 574652 215960 574704 215966
rect 574652 215902 574704 215908
rect 574468 214736 574520 214742
rect 574468 214678 574520 214684
rect 574664 214606 574692 215902
rect 574848 215014 574876 219302
rect 575020 218952 575072 218958
rect 575020 218894 575072 218900
rect 575032 218210 575060 218894
rect 575020 218204 575072 218210
rect 575020 218146 575072 218152
rect 575020 216708 575072 216714
rect 575020 216650 575072 216656
rect 574836 215008 574888 215014
rect 574836 214950 574888 214956
rect 574652 214600 574704 214606
rect 574652 214542 574704 214548
rect 575032 213654 575060 216650
rect 575216 215354 575244 220623
rect 575400 218754 575428 222974
rect 576030 222048 576086 222057
rect 576030 221983 576086 221992
rect 575388 218748 575440 218754
rect 575388 218690 575440 218696
rect 575664 218476 575716 218482
rect 575664 218418 575716 218424
rect 575676 217598 575704 218418
rect 575388 217592 575440 217598
rect 575388 217534 575440 217540
rect 575664 217592 575716 217598
rect 575664 217534 575716 217540
rect 575400 215490 575428 217534
rect 575572 216980 575624 216986
rect 575572 216922 575624 216928
rect 575388 215484 575440 215490
rect 575388 215426 575440 215432
rect 575204 215348 575256 215354
rect 575204 215290 575256 215296
rect 575020 213648 575072 213654
rect 575020 213590 575072 213596
rect 574100 213512 574152 213518
rect 573928 213472 574100 213500
rect 574100 213454 574152 213460
rect 574100 213376 574152 213382
rect 573836 213336 574100 213364
rect 574100 213318 574152 213324
rect 575584 213246 575612 216922
rect 576044 214878 576072 221983
rect 577320 218000 577372 218006
rect 577320 217942 577372 217948
rect 577332 216986 577360 217942
rect 577320 216980 577372 216986
rect 577320 216922 577372 216928
rect 576400 215348 576452 215354
rect 576400 215290 576452 215296
rect 576032 214872 576084 214878
rect 576032 214814 576084 214820
rect 576412 213790 576440 215290
rect 576400 213784 576452 213790
rect 576400 213726 576452 213732
rect 575572 213240 575624 213246
rect 575572 213182 575624 213188
rect 577516 99346 577544 240110
rect 587176 238746 587204 242150
rect 587164 238740 587216 238746
rect 587164 238682 587216 238688
rect 598216 235278 598244 245618
rect 623044 244316 623096 244322
rect 623044 244258 623096 244264
rect 598204 235272 598256 235278
rect 598204 235214 598256 235220
rect 593972 222284 594024 222290
rect 593972 222226 594024 222232
rect 596640 222284 596692 222290
rect 596640 222226 596692 222232
rect 591946 222048 592002 222057
rect 591946 221983 591948 221992
rect 592000 221983 592002 221992
rect 592132 222012 592184 222018
rect 591948 221954 592000 221960
rect 592132 221954 592184 221960
rect 592144 220862 592172 221954
rect 592132 220856 592184 220862
rect 592132 220798 592184 220804
rect 592316 220788 592368 220794
rect 592316 220730 592368 220736
rect 578238 220416 578294 220425
rect 578238 220351 578294 220360
rect 592038 220416 592094 220425
rect 592038 220351 592094 220360
rect 578252 218346 578280 220351
rect 582746 220280 582802 220289
rect 591854 220280 591910 220289
rect 582746 220215 582748 220224
rect 582800 220215 582802 220224
rect 582932 220244 582984 220250
rect 582748 220186 582800 220192
rect 582932 220186 582984 220192
rect 591672 220244 591724 220250
rect 592052 220266 592080 220351
rect 591910 220238 592080 220266
rect 591854 220215 591910 220224
rect 591672 220186 591724 220192
rect 582010 220008 582066 220017
rect 582562 220008 582618 220017
rect 582066 219966 582562 219994
rect 582010 219943 582066 219952
rect 582562 219943 582618 219952
rect 582196 219904 582248 219910
rect 582196 219846 582248 219852
rect 582380 219904 582432 219910
rect 582380 219846 582432 219852
rect 582208 219366 582236 219846
rect 582392 219366 582420 219846
rect 582196 219360 582248 219366
rect 582196 219302 582248 219308
rect 582380 219360 582432 219366
rect 582380 219302 582432 219308
rect 582944 219230 582972 220186
rect 591684 219230 591712 220186
rect 592038 220008 592094 220017
rect 592038 219943 592040 219952
rect 592092 219943 592094 219952
rect 592040 219914 592092 219920
rect 591856 219904 591908 219910
rect 591856 219846 591908 219852
rect 591868 219366 591896 219846
rect 592328 219366 592356 220730
rect 592500 220244 592552 220250
rect 592500 220186 592552 220192
rect 591856 219360 591908 219366
rect 591856 219302 591908 219308
rect 592316 219360 592368 219366
rect 592316 219302 592368 219308
rect 592512 219230 592540 220186
rect 582932 219224 582984 219230
rect 582932 219166 582984 219172
rect 591672 219224 591724 219230
rect 591672 219166 591724 219172
rect 592500 219224 592552 219230
rect 592500 219166 592552 219172
rect 584404 218612 584456 218618
rect 584404 218554 584456 218560
rect 582104 218476 582156 218482
rect 582104 218418 582156 218424
rect 582748 218476 582800 218482
rect 582748 218418 582800 218424
rect 577688 218340 577740 218346
rect 577688 218282 577740 218288
rect 578240 218340 578292 218346
rect 578240 218282 578292 218288
rect 577700 218074 577728 218282
rect 582116 218113 582144 218418
rect 582564 218340 582616 218346
rect 582564 218282 582616 218288
rect 582576 218113 582604 218282
rect 582102 218104 582158 218113
rect 577688 218068 577740 218074
rect 582102 218039 582158 218048
rect 582562 218104 582618 218113
rect 582562 218039 582618 218048
rect 577688 218010 577740 218016
rect 582760 217841 582788 218418
rect 582562 217832 582618 217841
rect 582562 217767 582618 217776
rect 582746 217832 582802 217841
rect 582746 217767 582802 217776
rect 582576 216238 582604 217767
rect 584416 216714 584444 218554
rect 592132 218340 592184 218346
rect 592132 218282 592184 218288
rect 592144 217734 592172 218282
rect 592132 217728 592184 217734
rect 592132 217670 592184 217676
rect 592316 217728 592368 217734
rect 592316 217670 592368 217676
rect 591946 217560 592002 217569
rect 592002 217518 592172 217546
rect 591946 217495 592002 217504
rect 592144 217054 592172 217518
rect 592132 217048 592184 217054
rect 592132 216990 592184 216996
rect 591948 216980 592000 216986
rect 591948 216922 592000 216928
rect 591960 216866 591988 216922
rect 592328 216866 592356 217670
rect 591960 216838 592356 216866
rect 590106 216744 590162 216753
rect 584404 216708 584456 216714
rect 590106 216679 590162 216688
rect 584404 216650 584456 216656
rect 582564 216232 582616 216238
rect 582564 216174 582616 216180
rect 590120 215626 590148 216679
rect 590108 215620 590160 215626
rect 590108 215562 590160 215568
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578516 211656
rect 578568 211647 578570 211656
rect 578516 211618 578568 211624
rect 578896 208350 578924 213959
rect 580448 211676 580500 211682
rect 580448 211618 580500 211624
rect 579252 209840 579304 209846
rect 579250 209808 579252 209817
rect 579304 209808 579306 209817
rect 579250 209743 579306 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 580460 207670 580488 211618
rect 593984 210202 594012 222226
rect 596652 220998 596680 222226
rect 596824 222148 596876 222154
rect 596824 222090 596876 222096
rect 600412 222148 600464 222154
rect 600412 222090 600464 222096
rect 596640 220992 596692 220998
rect 596640 220934 596692 220940
rect 596836 220930 596864 222090
rect 599306 222048 599362 222057
rect 599124 222012 599176 222018
rect 599306 221983 599308 221992
rect 599124 221954 599176 221960
rect 599360 221983 599362 221992
rect 599308 221954 599360 221960
rect 597926 221232 597982 221241
rect 597926 221167 597982 221176
rect 596824 220924 596876 220930
rect 596824 220866 596876 220872
rect 597468 218748 597520 218754
rect 597468 218690 597520 218696
rect 594260 217790 594656 217818
rect 594260 217734 594288 217790
rect 594248 217728 594300 217734
rect 594248 217670 594300 217676
rect 594432 217728 594484 217734
rect 594432 217670 594484 217676
rect 594444 217462 594472 217670
rect 594628 217546 594656 217790
rect 596362 217560 596418 217569
rect 594628 217518 594840 217546
rect 594432 217456 594484 217462
rect 594432 217398 594484 217404
rect 594616 217456 594668 217462
rect 594616 217398 594668 217404
rect 594628 217190 594656 217398
rect 594812 217190 594840 217518
rect 596362 217495 596418 217504
rect 594616 217184 594668 217190
rect 594616 217126 594668 217132
rect 594800 217184 594852 217190
rect 594800 217126 594852 217132
rect 595168 217048 595220 217054
rect 595168 216990 595220 216996
rect 594798 213208 594854 213217
rect 594798 213143 594854 213152
rect 594812 210202 594840 213143
rect 595180 210202 595208 216990
rect 595720 215620 595772 215626
rect 595720 215562 595772 215568
rect 595732 210202 595760 215562
rect 596376 210202 596404 217495
rect 596822 217288 596878 217297
rect 596822 217223 596878 217232
rect 596640 217116 596692 217122
rect 596640 217058 596692 217064
rect 596652 216850 596680 217058
rect 596640 216844 596692 216850
rect 596640 216786 596692 216792
rect 596836 210202 596864 217223
rect 597480 217025 597508 218690
rect 597744 218340 597796 218346
rect 597744 218282 597796 218288
rect 597466 217016 597522 217025
rect 597466 216951 597522 216960
rect 597756 216714 597784 218282
rect 597744 216708 597796 216714
rect 597744 216650 597796 216656
rect 597560 216232 597612 216238
rect 597560 216174 597612 216180
rect 597572 210202 597600 216174
rect 597940 215294 597968 221167
rect 597848 215266 597968 215294
rect 599136 215294 599164 221954
rect 599306 220416 599362 220425
rect 599306 220351 599362 220360
rect 599136 215266 599256 215294
rect 597848 210202 597876 215266
rect 598480 213784 598532 213790
rect 598480 213726 598532 213732
rect 598492 210202 598520 213726
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597848 210174 598276 210202
rect 598492 210174 598828 210202
rect 599228 210118 599256 215266
rect 599320 210202 599348 220351
rect 600424 210202 600452 222090
rect 600596 222012 600648 222018
rect 600596 221954 600648 221960
rect 600608 210202 600636 221954
rect 609980 221876 610032 221882
rect 609980 221818 610032 221824
rect 608968 221740 609020 221746
rect 608968 221682 609020 221688
rect 608784 221604 608836 221610
rect 608784 221546 608836 221552
rect 606024 221468 606076 221474
rect 606024 221410 606076 221416
rect 603448 221128 603500 221134
rect 603448 221070 603500 221076
rect 601344 220918 601740 220946
rect 601344 220522 601372 220918
rect 601712 220794 601740 220918
rect 601516 220788 601568 220794
rect 601516 220730 601568 220736
rect 601700 220788 601752 220794
rect 601700 220730 601752 220736
rect 601332 220516 601384 220522
rect 601528 220504 601556 220730
rect 601976 220516 602028 220522
rect 601528 220476 601976 220504
rect 601332 220458 601384 220464
rect 601976 220458 602028 220464
rect 601516 220244 601568 220250
rect 601516 220186 601568 220192
rect 601700 220244 601752 220250
rect 601700 220186 601752 220192
rect 601528 219230 601556 220186
rect 601712 219230 601740 220186
rect 601516 219224 601568 219230
rect 601516 219166 601568 219172
rect 601700 219224 601752 219230
rect 601700 219166 601752 219172
rect 601424 218408 601476 218414
rect 601422 218376 601424 218385
rect 601476 218376 601478 218385
rect 601422 218311 601478 218320
rect 601606 218376 601662 218385
rect 601606 218311 601662 218320
rect 601422 218104 601478 218113
rect 601620 218090 601648 218311
rect 601478 218062 601648 218090
rect 601422 218039 601478 218048
rect 601160 217926 601740 217954
rect 600962 217016 601018 217025
rect 601160 216986 601188 217926
rect 601516 217864 601568 217870
rect 601516 217806 601568 217812
rect 601332 217728 601384 217734
rect 601332 217670 601384 217676
rect 600962 216951 601018 216960
rect 601148 216980 601200 216986
rect 600976 216730 601004 216951
rect 601148 216922 601200 216928
rect 601344 216889 601372 217670
rect 601528 217410 601556 217806
rect 601712 217734 601740 217926
rect 601976 217864 602028 217870
rect 601976 217806 602028 217812
rect 601700 217728 601752 217734
rect 601700 217670 601752 217676
rect 601654 217592 601706 217598
rect 601652 217560 601654 217569
rect 601792 217592 601844 217598
rect 601706 217560 601708 217569
rect 601792 217534 601844 217540
rect 601652 217495 601708 217504
rect 601804 217410 601832 217534
rect 601988 217410 602016 217806
rect 603262 217560 603318 217569
rect 603262 217495 603318 217504
rect 601528 217382 601832 217410
rect 601896 217382 602016 217410
rect 601516 217320 601568 217326
rect 601516 217262 601568 217268
rect 601700 217320 601752 217326
rect 601896 217308 601924 217382
rect 601752 217280 601924 217308
rect 601700 217262 601752 217268
rect 601528 217161 601556 217262
rect 601976 217252 602028 217258
rect 601976 217194 602028 217200
rect 601514 217152 601570 217161
rect 601514 217087 601570 217096
rect 601790 217152 601846 217161
rect 601790 217087 601792 217096
rect 601844 217087 601846 217096
rect 601792 217058 601844 217064
rect 601988 217002 602016 217194
rect 603276 217122 603304 217495
rect 603080 217116 603132 217122
rect 603080 217058 603132 217064
rect 603264 217116 603316 217122
rect 603264 217058 603316 217064
rect 601516 216980 601568 216986
rect 601712 216974 602016 217002
rect 601712 216968 601740 216974
rect 601516 216922 601568 216928
rect 601666 216940 601740 216968
rect 601330 216880 601386 216889
rect 601330 216815 601386 216824
rect 601528 216730 601556 216922
rect 600976 216702 601556 216730
rect 601666 216714 601694 216940
rect 601790 216880 601846 216889
rect 601790 216815 601846 216824
rect 601804 216714 601832 216815
rect 601654 216708 601706 216714
rect 601654 216650 601706 216656
rect 601792 216708 601844 216714
rect 601792 216650 601844 216656
rect 602526 216472 602582 216481
rect 602526 216407 602582 216416
rect 601240 213648 601292 213654
rect 601240 213590 601292 213596
rect 601252 210202 601280 213590
rect 601792 213512 601844 213518
rect 601792 213454 601844 213460
rect 601804 210202 601832 213454
rect 602540 213382 602568 216407
rect 603092 213586 603120 217058
rect 603080 213580 603132 213586
rect 603080 213522 603132 213528
rect 602344 213376 602396 213382
rect 602344 213318 602396 213324
rect 602528 213376 602580 213382
rect 602528 213318 602580 213324
rect 602356 210202 602384 213318
rect 603080 213240 603132 213246
rect 603080 213182 603132 213188
rect 603092 210202 603120 213182
rect 603460 210202 603488 221070
rect 605656 218884 605708 218890
rect 605656 218826 605708 218832
rect 605668 217462 605696 218826
rect 605840 217728 605892 217734
rect 605840 217670 605892 217676
rect 604000 217456 604052 217462
rect 604000 217398 604052 217404
rect 605656 217456 605708 217462
rect 605656 217398 605708 217404
rect 604012 210202 604040 217398
rect 605852 216714 605880 217670
rect 605104 216708 605156 216714
rect 605104 216650 605156 216656
rect 605840 216708 605892 216714
rect 605840 216650 605892 216656
rect 604552 213580 604604 213586
rect 604552 213522 604604 213528
rect 604564 210202 604592 213522
rect 605116 210202 605144 216650
rect 606036 210202 606064 221410
rect 607772 221264 607824 221270
rect 607772 221206 607824 221212
rect 606206 218920 606262 218929
rect 606206 218855 606262 218864
rect 606220 217734 606248 218855
rect 606758 218648 606814 218657
rect 606758 218583 606814 218592
rect 606772 218113 606800 218583
rect 607496 218408 607548 218414
rect 607496 218350 607548 218356
rect 606758 218104 606814 218113
rect 606758 218039 606814 218048
rect 606208 217728 606260 217734
rect 606208 217670 606260 217676
rect 607312 217592 607364 217598
rect 607312 217534 607364 217540
rect 606208 217252 606260 217258
rect 606208 217194 606260 217200
rect 599320 210174 599380 210202
rect 600424 210174 600484 210202
rect 600608 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602356 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605116 210174 605452 210202
rect 606004 210174 606064 210202
rect 606220 210202 606248 217194
rect 606760 216708 606812 216714
rect 606760 216650 606812 216656
rect 606772 210202 606800 216650
rect 607324 210202 607352 217534
rect 607508 216714 607536 218350
rect 607496 216708 607548 216714
rect 607496 216650 607548 216656
rect 607784 210202 607812 221206
rect 608796 214470 608824 221546
rect 608784 214464 608836 214470
rect 608784 214406 608836 214412
rect 608980 210202 609008 221682
rect 609152 217864 609204 217870
rect 609152 217806 609204 217812
rect 606220 210174 606556 210202
rect 606772 210174 607108 210202
rect 607324 210174 607660 210202
rect 607784 210174 608212 210202
rect 608764 210174 609008 210202
rect 609164 210202 609192 217806
rect 609520 214464 609572 214470
rect 609520 214406 609572 214412
rect 609532 210202 609560 214406
rect 609992 210202 610020 221818
rect 618258 221776 618314 221785
rect 618258 221711 618314 221720
rect 616878 221504 616934 221513
rect 616878 221439 616934 221448
rect 611450 220960 611506 220969
rect 611450 220895 611506 220904
rect 611636 220924 611688 220930
rect 610624 217116 610676 217122
rect 610624 217058 610676 217064
rect 610636 210202 610664 217058
rect 611464 214470 611492 220895
rect 611636 220866 611688 220872
rect 611452 214464 611504 214470
rect 611452 214406 611504 214412
rect 611648 210202 611676 220866
rect 613292 220516 613344 220522
rect 613292 220458 613344 220464
rect 612924 220244 612976 220250
rect 612924 220186 612976 220192
rect 612738 218920 612794 218929
rect 612738 218855 612794 218864
rect 612280 215280 612332 215286
rect 612280 215222 612332 215228
rect 611820 214464 611872 214470
rect 611820 214406 611872 214412
rect 609164 210174 609316 210202
rect 609532 210174 609868 210202
rect 609992 210174 610420 210202
rect 610636 210174 610972 210202
rect 611524 210174 611676 210202
rect 611832 210202 611860 214406
rect 612292 210202 612320 215222
rect 612752 213926 612780 218855
rect 612740 213920 612792 213926
rect 612740 213862 612792 213868
rect 612936 211682 612964 220186
rect 613304 219502 613332 220458
rect 613108 219496 613160 219502
rect 613108 219438 613160 219444
rect 613292 219496 613344 219502
rect 613292 219438 613344 219444
rect 612924 211676 612976 211682
rect 612924 211618 612976 211624
rect 613120 210202 613148 219438
rect 616144 218204 616196 218210
rect 616144 218146 616196 218152
rect 615684 217728 615736 217734
rect 615684 217670 615736 217676
rect 614488 216844 614540 216850
rect 614488 216786 614540 216792
rect 614120 216708 614172 216714
rect 614120 216650 614172 216656
rect 613384 211676 613436 211682
rect 613384 211618 613436 211624
rect 613396 210202 613424 211618
rect 614132 210202 614160 216650
rect 614500 210202 614528 216786
rect 615040 213920 615092 213926
rect 615040 213862 615092 213868
rect 615052 210202 615080 213862
rect 615696 210202 615724 217670
rect 616156 210202 616184 218146
rect 616892 214742 616920 221439
rect 617524 220788 617576 220794
rect 617524 220730 617576 220736
rect 617338 219192 617394 219201
rect 617338 219127 617394 219136
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616880 214736 616932 214742
rect 616880 214678 616932 214684
rect 616708 214470 616736 214678
rect 616696 214464 616748 214470
rect 616696 214406 616748 214412
rect 611832 210174 612076 210202
rect 612292 210174 612628 210202
rect 613120 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 599216 210112 599268 210118
rect 599216 210054 599268 210060
rect 599584 210112 599636 210118
rect 617352 210066 617380 219127
rect 617536 210202 617564 220730
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 221711
rect 618812 220652 618864 220658
rect 618812 220594 618864 220600
rect 618824 210202 618852 220594
rect 620468 220380 620520 220386
rect 620468 220322 620520 220328
rect 619640 216096 619692 216102
rect 619640 216038 619692 216044
rect 619652 210202 619680 216038
rect 620008 215144 620060 215150
rect 620008 215086 620060 215092
rect 620020 210202 620048 215086
rect 620480 210202 620508 220322
rect 621572 219904 621624 219910
rect 621572 219846 621624 219852
rect 621112 216368 621164 216374
rect 621112 216310 621164 216316
rect 621124 210202 621152 216310
rect 621584 210202 621612 219846
rect 623056 215966 623084 244258
rect 631324 241528 631376 241534
rect 631324 241470 631376 241476
rect 631336 229094 631364 241470
rect 632716 229094 632744 246298
rect 648632 242214 648660 277366
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 633624 235272 633676 235278
rect 633624 235214 633676 235220
rect 631336 229066 631456 229094
rect 632716 229066 632928 229094
rect 627092 220108 627144 220114
rect 627092 220050 627144 220056
rect 623780 219768 623832 219774
rect 623780 219710 623832 219716
rect 623320 216504 623372 216510
rect 623320 216446 623372 216452
rect 623044 215960 623096 215966
rect 623044 215902 623096 215908
rect 622400 215008 622452 215014
rect 622400 214950 622452 214956
rect 622412 210202 622440 214950
rect 622768 213376 622820 213382
rect 622768 213318 622820 213324
rect 622780 210202 622808 213318
rect 623332 210202 623360 216446
rect 623792 210202 623820 219710
rect 625436 219632 625488 219638
rect 625436 219574 625488 219580
rect 623962 218376 624018 218385
rect 623962 218311 624018 218320
rect 623976 213246 624004 218311
rect 625252 216980 625304 216986
rect 625252 216922 625304 216928
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 623964 213240 624016 213246
rect 623964 213182 624016 213188
rect 624436 210202 624464 214406
rect 625264 210202 625292 216922
rect 625448 210202 625476 219574
rect 626630 216200 626686 216209
rect 626630 216135 626686 216144
rect 626080 214872 626132 214878
rect 626080 214814 626132 214820
rect 626092 210202 626120 214814
rect 626644 210202 626672 216135
rect 627104 210202 627132 220050
rect 630770 219736 630826 219745
rect 630770 219671 630826 219680
rect 628104 219496 628156 219502
rect 628104 219438 628156 219444
rect 627734 218648 627790 218657
rect 627734 218583 627790 218592
rect 627748 214198 627776 218583
rect 627920 217456 627972 217462
rect 627920 217398 627972 217404
rect 627736 214192 627788 214198
rect 627736 214134 627788 214140
rect 627932 210202 627960 217398
rect 628116 214690 628144 219438
rect 629392 218068 629444 218074
rect 629392 218010 629444 218016
rect 628116 214662 628788 214690
rect 628288 214600 628340 214606
rect 628288 214542 628340 214548
rect 628300 210202 628328 214542
rect 628760 210202 628788 214662
rect 629404 210202 629432 218010
rect 629944 213240 629996 213246
rect 629944 213182 629996 213188
rect 629956 210202 629984 213182
rect 630784 210202 630812 219671
rect 631230 219464 631286 219473
rect 631230 219399 631286 219408
rect 631048 214192 631100 214198
rect 631048 214134 631100 214140
rect 631060 210202 631088 214134
rect 631244 210338 631272 219399
rect 631428 214606 631456 229066
rect 631416 214600 631468 214606
rect 631416 214542 631468 214548
rect 632704 214600 632756 214606
rect 632704 214542 632756 214548
rect 631244 210310 631548 210338
rect 631520 210202 631548 210310
rect 632716 210202 632744 214542
rect 632900 212906 632928 229066
rect 632888 212900 632940 212906
rect 632888 212842 632940 212848
rect 633636 210202 633664 235214
rect 652036 232558 652064 378111
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652024 232552 652076 232558
rect 652024 232494 652076 232500
rect 640246 231432 640302 231441
rect 640246 231367 640302 231376
rect 639602 230208 639658 230217
rect 639602 230143 639658 230152
rect 637486 229800 637542 229809
rect 637486 229735 637542 229744
rect 637500 219434 637528 229735
rect 637670 220144 637726 220153
rect 637670 220079 637726 220088
rect 637684 219434 637712 220079
rect 637316 219406 637528 219434
rect 637592 219406 637712 219434
rect 633808 215960 633860 215966
rect 633808 215902 633860 215908
rect 617536 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618824 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620480 210174 620908 210202
rect 621124 210174 621460 210202
rect 621584 210174 622012 210202
rect 622412 210174 622564 210202
rect 622780 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624436 210174 624772 210202
rect 625264 210174 625324 210202
rect 625448 210174 625876 210202
rect 626092 210174 626428 210202
rect 626644 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628760 210174 629188 210202
rect 629404 210174 629740 210202
rect 629956 210174 630292 210202
rect 630784 210174 630844 210202
rect 631060 210174 631396 210202
rect 631520 210174 631948 210202
rect 632716 210174 633052 210202
rect 633604 210174 633664 210202
rect 633820 210202 633848 215902
rect 635556 213376 635608 213382
rect 635556 213318 635608 213324
rect 634360 212900 634412 212906
rect 634360 212842 634412 212848
rect 634372 210202 634400 212842
rect 635568 210202 635596 213318
rect 636660 212832 636712 212838
rect 636660 212774 636712 212780
rect 636672 210202 636700 212774
rect 637316 210202 637344 219406
rect 637592 213926 637620 219406
rect 637580 213920 637632 213926
rect 637580 213862 637632 213868
rect 638224 213920 638276 213926
rect 638224 213862 638276 213868
rect 638040 213784 638092 213790
rect 638040 213726 638092 213732
rect 638052 210202 638080 213726
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637344 210202
rect 638020 210174 638080 210202
rect 638236 210202 638264 213862
rect 639616 212838 639644 230143
rect 639972 213920 640024 213926
rect 639972 213862 640024 213868
rect 639604 212832 639656 212838
rect 639604 212774 639656 212780
rect 639984 210202 640012 213862
rect 640260 210202 640288 231367
rect 650642 225584 650698 225593
rect 650642 225519 650698 225528
rect 643190 220416 643246 220425
rect 643190 220351 643246 220360
rect 640430 218920 640486 218929
rect 640430 218855 640486 218864
rect 640444 213790 640472 218855
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 640432 213784 640484 213790
rect 640432 213726 640484 213732
rect 641628 213648 641680 213654
rect 641628 213590 641680 213596
rect 641640 210202 641668 213590
rect 642180 213512 642232 213518
rect 642180 213454 642232 213460
rect 642192 210202 642220 213454
rect 643020 210202 643048 215863
rect 643204 213926 643232 220351
rect 647332 220108 647384 220114
rect 647332 220050 647384 220056
rect 645490 218648 645546 218657
rect 645490 218583 645546 218592
rect 643192 213920 643244 213926
rect 643192 213862 643244 213868
rect 644940 213784 644992 213790
rect 644940 213726 644992 213732
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 643848 210202 643876 213182
rect 644952 210202 644980 213726
rect 645504 210202 645532 218583
rect 646870 217560 646926 217569
rect 646870 217495 646926 217504
rect 646594 216472 646650 216481
rect 646594 216407 646650 216416
rect 646608 210202 646636 216407
rect 646884 213790 646912 217495
rect 646872 213784 646924 213790
rect 646872 213726 646924 213732
rect 647146 213208 647202 213217
rect 647146 213143 647202 213152
rect 647160 210202 647188 213143
rect 647344 210338 647372 220050
rect 649906 217832 649962 217841
rect 649906 217767 649962 217776
rect 648526 214568 648582 214577
rect 648526 214503 648582 214512
rect 647344 210310 647556 210338
rect 638236 210174 638572 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647528 210202 647556 210310
rect 648540 210202 648568 214503
rect 649920 210202 649948 217767
rect 650656 213654 650684 225519
rect 651286 223136 651342 223145
rect 651286 223071 651342 223080
rect 651102 216200 651158 216209
rect 651102 216135 651158 216144
rect 650644 213648 650696 213654
rect 650644 213590 650696 213596
rect 650460 213036 650512 213042
rect 650460 212978 650512 212984
rect 650472 210202 650500 212978
rect 647528 210174 647956 210202
rect 648508 210174 648568 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 216135
rect 651300 213042 651328 223071
rect 651838 222864 651894 222873
rect 651838 222799 651894 222808
rect 651852 213382 651880 222799
rect 652024 213648 652076 213654
rect 652024 213590 652076 213596
rect 651840 213376 651892 213382
rect 651840 213318 651892 213324
rect 651288 213036 651340 213042
rect 651288 212978 651340 212984
rect 652036 210202 652064 213590
rect 651116 210174 651268 210202
rect 651820 210174 652064 210202
rect 599636 210060 599932 210066
rect 599584 210054 599932 210060
rect 599596 210038 599932 210054
rect 617044 210038 617380 210066
rect 581736 209840 581788 209846
rect 581736 209782 581788 209788
rect 580448 207664 580500 207670
rect 580448 207606 580500 207612
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 581748 206310 581776 209782
rect 652220 209574 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 405657 660344 550598
rect 663076 538801 663104 656882
rect 664456 579737 664484 709310
rect 665836 626113 665864 749362
rect 666282 742520 666338 742529
rect 666282 742455 666338 742464
rect 666296 665553 666324 742455
rect 666480 711657 666508 778359
rect 666466 711648 666522 711657
rect 666466 711583 666522 711592
rect 666466 699816 666522 699825
rect 666466 699751 666522 699760
rect 666282 665544 666338 665553
rect 666282 665479 666338 665488
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 666480 621217 666508 699751
rect 667216 671129 667244 803150
rect 667860 750825 667888 866623
rect 668584 789404 668636 789410
rect 668584 789346 668636 789352
rect 668214 782504 668270 782513
rect 668214 782439 668270 782448
rect 667846 750816 667902 750825
rect 667846 750751 667902 750760
rect 667846 743200 667902 743209
rect 667846 743135 667902 743144
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 667860 665281 667888 743135
rect 668228 710433 668256 782439
rect 668400 775600 668452 775606
rect 668400 775542 668452 775548
rect 668412 734777 668440 775542
rect 668398 734768 668454 734777
rect 668398 734703 668454 734712
rect 668398 733136 668454 733145
rect 668398 733071 668454 733080
rect 668214 710424 668270 710433
rect 668214 710359 668270 710368
rect 668030 686216 668086 686225
rect 668030 686151 668086 686160
rect 667846 665272 667902 665281
rect 667846 665207 667902 665216
rect 667846 661056 667902 661065
rect 667846 660991 667902 661000
rect 667204 629332 667256 629338
rect 667204 629274 667256 629280
rect 666466 621208 666522 621217
rect 666466 621143 666522 621152
rect 666466 608832 666522 608841
rect 666466 608767 666522 608776
rect 664628 603152 664680 603158
rect 664628 603094 664680 603100
rect 664442 579728 664498 579737
rect 664442 579663 664498 579672
rect 663062 538792 663118 538801
rect 663062 538727 663118 538736
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661684 416832 661736 416838
rect 661684 416774 661736 416780
rect 660302 405648 660358 405657
rect 660302 405583 660358 405592
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 661696 268161 661724 416774
rect 661880 406337 661908 522990
rect 664640 491745 664668 603094
rect 666008 576904 666060 576910
rect 666008 576846 666060 576852
rect 665824 494760 665876 494766
rect 665824 494702 665876 494708
rect 664626 491736 664682 491745
rect 664626 491671 664682 491680
rect 663064 470620 663116 470626
rect 663064 470562 663116 470568
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 663076 315489 663104 470562
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663248 364404 663300 364410
rect 663248 364346 663300 364352
rect 663062 315480 663118 315489
rect 663062 315415 663118 315424
rect 661682 268152 661738 268161
rect 661682 268087 661738 268096
rect 663260 234161 663288 364346
rect 664456 271153 664484 404330
rect 665836 358737 665864 494702
rect 666020 494057 666048 576846
rect 666480 531457 666508 608767
rect 667216 534449 667244 629274
rect 667202 534440 667258 534449
rect 667202 534375 667258 534384
rect 666466 531448 666522 531457
rect 666466 531383 666522 531392
rect 666006 494048 666062 494057
rect 666006 493983 666062 493992
rect 667204 456816 667256 456822
rect 667204 456758 667256 456764
rect 665822 358728 665878 358737
rect 665822 358663 665878 358672
rect 666376 338156 666428 338162
rect 666376 338098 666428 338104
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 666190 236192 666246 236201
rect 666190 236127 666246 236136
rect 663246 234152 663302 234161
rect 663246 234087 663302 234096
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 662328 232416 662380 232422
rect 662328 232358 662380 232364
rect 660946 229528 661002 229537
rect 660946 229463 661002 229472
rect 652758 226400 652814 226409
rect 652758 226335 652814 226344
rect 652772 220114 652800 226335
rect 660210 225312 660266 225321
rect 660210 225247 660266 225256
rect 655426 225040 655482 225049
rect 655426 224975 655482 224984
rect 653034 220688 653090 220697
rect 653034 220623 653090 220632
rect 652760 220108 652812 220114
rect 652760 220050 652812 220056
rect 652852 213376 652904 213382
rect 652852 213318 652904 213324
rect 652864 210202 652892 213318
rect 653048 210202 653076 220623
rect 655242 219192 655298 219201
rect 655242 219127 655298 219136
rect 654876 213920 654928 213926
rect 654876 213862 654928 213868
rect 654888 210202 654916 213862
rect 655256 210202 655284 219127
rect 655440 213926 655468 224975
rect 658186 224496 658242 224505
rect 658186 224431 658242 224440
rect 656622 223680 656678 223689
rect 656622 223615 656678 223624
rect 655428 213920 655480 213926
rect 655428 213862 655480 213868
rect 656636 210202 656664 223615
rect 658002 221504 658058 221513
rect 658002 221439 658058 221448
rect 656808 214600 656860 214606
rect 656808 214542 656860 214548
rect 656820 210202 656848 214542
rect 658016 213654 658044 221439
rect 658004 213648 658056 213654
rect 658004 213590 658056 213596
rect 658200 210202 658228 224431
rect 658922 223952 658978 223961
rect 658922 223887 658978 223896
rect 658740 214736 658792 214742
rect 658740 214678 658792 214684
rect 658752 210202 658780 214678
rect 658936 214606 658964 223887
rect 659382 221232 659438 221241
rect 659382 221167 659438 221176
rect 658924 214600 658976 214606
rect 658924 214542 658976 214548
rect 659396 213518 659424 221167
rect 659568 213648 659620 213654
rect 659568 213590 659620 213596
rect 659384 213512 659436 213518
rect 659384 213454 659436 213460
rect 659580 210202 659608 213590
rect 660224 213382 660252 225247
rect 660960 213926 660988 229463
rect 661682 229256 661738 229265
rect 661682 229191 661738 229200
rect 661696 214742 661724 229191
rect 661684 214736 661736 214742
rect 661684 214678 661736 214684
rect 662052 214600 662104 214606
rect 662052 214542 662104 214548
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 660212 213376 660264 213382
rect 660212 213318 660264 213324
rect 660408 210202 660436 213862
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660960 210202 660988 213726
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 214542
rect 662340 210202 662368 232358
rect 665088 232212 665140 232218
rect 665088 232154 665140 232160
rect 663062 231704 663118 231713
rect 663062 231639 663118 231648
rect 663076 215294 663104 231639
rect 663246 230888 663302 230897
rect 663246 230823 663302 230832
rect 662984 215266 663104 215294
rect 662984 213790 663012 215266
rect 663260 214606 663288 230823
rect 664442 230616 664498 230625
rect 664442 230551 664498 230560
rect 663708 227792 663760 227798
rect 663708 227734 663760 227740
rect 663430 220416 663486 220425
rect 663430 220351 663486 220360
rect 663444 219609 663472 220351
rect 663430 219600 663486 219609
rect 663430 219535 663486 219544
rect 663524 214940 663576 214946
rect 663524 214882 663576 214888
rect 663248 214600 663300 214606
rect 663248 214542 663300 214548
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 662972 213784 663024 213790
rect 662972 213726 663024 213732
rect 663168 210202 663196 213862
rect 663536 210202 663564 214882
rect 663720 213926 663748 227734
rect 664456 214946 664484 230551
rect 664902 215112 664958 215121
rect 664902 215047 664958 215056
rect 664444 214940 664496 214946
rect 664444 214882 664496 214888
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664718 213752 664774 213761
rect 664718 213687 664774 213696
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664732 210202 664760 213687
rect 664916 213654 664944 215047
rect 664904 213648 664956 213654
rect 664904 213590 664956 213596
rect 665100 213042 665128 232154
rect 665270 231160 665326 231169
rect 665270 231095 665326 231104
rect 665284 227798 665312 231095
rect 665272 227792 665324 227798
rect 665272 227734 665324 227740
rect 665270 222048 665326 222057
rect 665270 221983 665326 221992
rect 665284 213246 665312 221983
rect 665272 213240 665324 213246
rect 665272 213182 665324 213188
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654580 210174 654916 210202
rect 655132 210174 655284 210202
rect 656236 210174 656664 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664760 210202
rect 632152 209568 632204 209574
rect 652208 209568 652260 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652208 209510 652260 209516
rect 632164 209494 632500 209510
rect 591304 208684 591356 208690
rect 591304 208626 591356 208632
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 207664 589516 207670
rect 589464 207606 589516 207612
rect 589476 206417 589504 207606
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 581736 206304 581788 206310
rect 581736 206246 581788 206252
rect 589648 206304 589700 206310
rect 589648 206246 589700 206252
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 589660 204785 589688 206246
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 589648 186312 589700 186318
rect 579580 186280 579582 186289
rect 589648 186254 589700 186260
rect 579526 186215 579582 186224
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 578804 180169 578832 180746
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 578804 175137 578832 178026
rect 589660 177954 589688 180231
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 583208 175296 583260 175302
rect 583208 175238 583260 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 579526 171048 579582 171057
rect 579526 170983 579528 170992
rect 579580 170983 579582 170992
rect 579528 170954 579580 170960
rect 580920 169726 580948 172518
rect 581644 171148 581696 171154
rect 581644 171090 581696 171096
rect 578332 169720 578384 169726
rect 578332 169662 578384 169668
rect 580908 169720 580960 169726
rect 580908 169662 580960 169668
rect 578344 169289 578372 169662
rect 578330 169280 578386 169289
rect 578330 169215 578386 169224
rect 579620 168428 579672 168434
rect 579620 168370 579672 168376
rect 578976 167204 579028 167210
rect 578976 167146 579028 167152
rect 578988 166977 579016 167146
rect 578974 166968 579030 166977
rect 578974 166903 579030 166912
rect 578884 165572 578936 165578
rect 578884 165514 578936 165520
rect 578896 164529 578924 165514
rect 578882 164520 578938 164529
rect 578882 164455 578938 164464
rect 579434 162480 579490 162489
rect 579632 162466 579660 168370
rect 581656 167210 581684 171090
rect 583220 171018 583248 175238
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 583208 171012 583260 171018
rect 583208 170954 583260 170960
rect 589462 170504 589518 170513
rect 589462 170439 589518 170448
rect 589476 169794 589504 170439
rect 582380 169788 582432 169794
rect 582380 169730 582432 169736
rect 589464 169788 589516 169794
rect 589464 169730 589516 169736
rect 581644 167204 581696 167210
rect 581644 167146 581696 167152
rect 581644 167068 581696 167074
rect 581644 167010 581696 167016
rect 579490 162438 579660 162466
rect 579434 162415 579490 162424
rect 580448 161492 580500 161498
rect 580448 161434 580500 161440
rect 579252 160064 579304 160070
rect 579252 160006 579304 160012
rect 579264 159905 579292 160006
rect 579250 159896 579306 159905
rect 579250 159831 579306 159840
rect 579160 158704 579212 158710
rect 579160 158646 579212 158652
rect 579172 158273 579200 158646
rect 579158 158264 579214 158273
rect 579158 158199 579214 158208
rect 579526 155952 579582 155961
rect 579526 155887 579528 155896
rect 579580 155887 579582 155896
rect 579528 155858 579580 155864
rect 580460 154562 580488 161434
rect 581656 160070 581684 167010
rect 582392 165578 582420 169730
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589462 165608 589518 165617
rect 582380 165572 582432 165578
rect 589462 165543 589518 165552
rect 582380 165514 582432 165520
rect 589476 164286 589504 165543
rect 585968 164280 586020 164286
rect 585968 164222 586020 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 584404 162920 584456 162926
rect 584404 162862 584456 162868
rect 582380 160132 582432 160138
rect 582380 160074 582432 160080
rect 581644 160064 581696 160070
rect 581644 160006 581696 160012
rect 581828 158840 581880 158846
rect 581828 158782 581880 158788
rect 578240 154556 578292 154562
rect 578240 154498 578292 154504
rect 580448 154556 580500 154562
rect 580448 154498 580500 154504
rect 578252 154057 578280 154498
rect 578238 154048 578294 154057
rect 578238 153983 578294 153992
rect 580264 153264 580316 153270
rect 580264 153206 580316 153212
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 578252 151745 578280 152730
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 147416 579580 147422
rect 579528 147358 579580 147364
rect 579540 147257 579568 147358
rect 579526 147248 579582 147257
rect 579526 147183 579582 147192
rect 578884 145580 578936 145586
rect 578884 145522 578936 145528
rect 578516 143336 578568 143342
rect 578516 143278 578568 143284
rect 578528 143041 578556 143278
rect 578514 143032 578570 143041
rect 578514 142967 578570 142976
rect 578700 139392 578752 139398
rect 578700 139334 578752 139340
rect 578712 138825 578740 139334
rect 578698 138816 578754 138825
rect 578698 138751 578754 138760
rect 578896 136649 578924 145522
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 580276 143342 580304 153206
rect 581840 150618 581868 158782
rect 582392 152794 582420 160074
rect 584416 155922 584444 162862
rect 585980 158710 586008 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158846 589504 159015
rect 589464 158840 589516 158846
rect 589464 158782 589516 158788
rect 585968 158704 586020 158710
rect 585968 158646 586020 158652
rect 589462 157448 589518 157457
rect 585784 157412 585836 157418
rect 589462 157383 589464 157392
rect 585784 157354 585836 157360
rect 589516 157383 589518 157392
rect 589464 157354 589516 157360
rect 584404 155916 584456 155922
rect 584404 155858 584456 155864
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 582380 152788 582432 152794
rect 582380 152730 582432 152736
rect 583024 151836 583076 151842
rect 583024 151778 583076 151784
rect 581828 150612 581880 150618
rect 581828 150554 581880 150560
rect 581644 150476 581696 150482
rect 581644 150418 581696 150424
rect 580264 143336 580316 143342
rect 580264 143278 580316 143284
rect 580448 142180 580500 142186
rect 580448 142122 580500 142128
rect 579528 140616 579580 140622
rect 579526 140584 579528 140593
rect 579580 140584 579582 140593
rect 579526 140519 579582 140528
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 578332 135924 578384 135930
rect 578332 135866 578384 135872
rect 578344 134473 578372 135866
rect 578330 134464 578386 134473
rect 578330 134399 578386 134408
rect 578240 134292 578292 134298
rect 578240 134234 578292 134240
rect 578252 132297 578280 134234
rect 579252 133204 579304 133210
rect 579252 133146 579304 133152
rect 578238 132288 578294 132297
rect 578238 132223 578294 132232
rect 578332 128308 578384 128314
rect 578332 128250 578384 128256
rect 578344 127809 578372 128250
rect 578330 127800 578386 127809
rect 578330 127735 578386 127744
rect 579264 125361 579292 133146
rect 579528 129736 579580 129742
rect 579526 129704 579528 129713
rect 579580 129704 579582 129713
rect 579526 129639 579582 129648
rect 580460 128314 580488 142122
rect 581656 139398 581684 150418
rect 583036 140622 583064 151778
rect 584416 144702 584444 154566
rect 585796 147422 585824 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 589462 150920 589518 150929
rect 589462 150855 589518 150864
rect 589476 150482 589504 150855
rect 589464 150476 589516 150482
rect 589464 150418 589516 150424
rect 589186 149288 589242 149297
rect 589186 149223 589242 149232
rect 585784 147416 585836 147422
rect 585784 147358 585836 147364
rect 587348 146328 587400 146334
rect 587348 146270 587400 146276
rect 585784 144968 585836 144974
rect 585784 144910 585836 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 140616 583076 140622
rect 583024 140558 583076 140564
rect 584404 139460 584456 139466
rect 584404 139402 584456 139408
rect 581644 139392 581696 139398
rect 581644 139334 581696 139340
rect 581644 136672 581696 136678
rect 581644 136614 581696 136620
rect 580448 128308 580500 128314
rect 580448 128250 580500 128256
rect 580264 127016 580316 127022
rect 580264 126958 580316 126964
rect 579250 125352 579306 125361
rect 579250 125287 579306 125296
rect 579252 124160 579304 124166
rect 579252 124102 579304 124108
rect 579264 123593 579292 124102
rect 579250 123584 579306 123593
rect 579250 123519 579306 123528
rect 579252 122868 579304 122874
rect 579252 122810 579304 122816
rect 579068 121168 579120 121174
rect 579066 121136 579068 121145
rect 579120 121136 579122 121145
rect 579066 121071 579122 121080
rect 578516 118652 578568 118658
rect 578516 118594 578568 118600
rect 578528 118425 578556 118594
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 579068 115252 579120 115258
rect 579068 115194 579120 115200
rect 578332 108384 578384 108390
rect 578330 108352 578332 108361
rect 578384 108352 578386 108361
rect 578330 108287 578386 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578332 106956 578384 106962
rect 578332 106898 578384 106904
rect 578344 105913 578372 106898
rect 578330 105904 578386 105913
rect 578330 105839 578386 105848
rect 577504 99340 577556 99346
rect 577504 99282 577556 99288
rect 577504 97300 577556 97306
rect 577504 97242 577556 97248
rect 575480 57248 575532 57254
rect 575480 57190 575532 57196
rect 574928 56160 574980 56166
rect 574928 56102 574980 56108
rect 574560 56024 574612 56030
rect 574560 55966 574612 55972
rect 574008 55616 574060 55622
rect 574008 55558 574060 55564
rect 574020 53854 574048 55558
rect 574572 54262 574600 55966
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 55214 574784 55830
rect 574744 55208 574796 55214
rect 574744 55150 574796 55156
rect 574560 54256 574612 54262
rect 574560 54198 574612 54204
rect 574940 53990 574968 56102
rect 575492 54126 575520 57190
rect 577516 54398 577544 97242
rect 578700 95056 578752 95062
rect 578698 95024 578700 95033
rect 578752 95024 578754 95033
rect 578698 94959 578754 94968
rect 578608 86624 578660 86630
rect 578608 86566 578660 86572
rect 578620 86465 578648 86566
rect 578606 86456 578662 86465
rect 578606 86391 578662 86400
rect 578896 84194 578924 107578
rect 579080 90953 579108 115194
rect 579264 101833 579292 122810
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579526 114472 579582 114481
rect 579526 114407 579528 114416
rect 579580 114407 579582 114416
rect 579528 114378 579580 114384
rect 579528 113144 579580 113150
rect 579528 113086 579580 113092
rect 579540 112713 579568 113086
rect 579526 112704 579582 112713
rect 579526 112639 579582 112648
rect 579436 110288 579488 110294
rect 579434 110256 579436 110265
rect 579488 110256 579490 110265
rect 579434 110191 579490 110200
rect 580276 106962 580304 126958
rect 581656 121174 581684 136614
rect 582380 131776 582432 131782
rect 582380 131718 582432 131724
rect 582392 129742 582420 131718
rect 582380 129736 582432 129742
rect 582380 129678 582432 129684
rect 583024 128376 583076 128382
rect 583024 128318 583076 128324
rect 581644 121168 581696 121174
rect 581644 121110 581696 121116
rect 582012 120760 582064 120766
rect 582012 120702 582064 120708
rect 582024 110294 582052 120702
rect 582012 110288 582064 110294
rect 582012 110230 582064 110236
rect 581828 109744 581880 109750
rect 581828 109686 581880 109692
rect 580632 107092 580684 107098
rect 580632 107034 580684 107040
rect 580264 106956 580316 106962
rect 580264 106898 580316 106904
rect 580448 106956 580500 106962
rect 580448 106898 580500 106904
rect 579528 103352 579580 103358
rect 579526 103320 579528 103329
rect 579580 103320 579582 103329
rect 579526 103255 579582 103264
rect 579250 101824 579306 101833
rect 579250 101759 579306 101768
rect 579526 99240 579582 99249
rect 579526 99175 579528 99184
rect 579580 99175 579582 99184
rect 579528 99146 579580 99152
rect 579528 97504 579580 97510
rect 579526 97472 579528 97481
rect 579580 97472 579582 97481
rect 579526 97407 579582 97416
rect 579528 93288 579580 93294
rect 579528 93230 579580 93236
rect 579540 93129 579568 93230
rect 580264 93152 580316 93158
rect 579526 93120 579582 93129
rect 580264 93094 580316 93100
rect 579526 93055 579582 93064
rect 579066 90944 579122 90953
rect 579066 90879 579122 90888
rect 579528 88324 579580 88330
rect 579528 88266 579580 88272
rect 579540 88097 579568 88266
rect 579526 88088 579582 88097
rect 579526 88023 579582 88032
rect 578804 84166 578924 84194
rect 579252 84176 579304 84182
rect 578804 80073 578832 84166
rect 579252 84118 579304 84124
rect 579264 84017 579292 84118
rect 579250 84008 579306 84017
rect 579250 83943 579306 83952
rect 579252 82816 579304 82822
rect 579252 82758 579304 82764
rect 579264 82249 579292 82758
rect 579250 82240 579306 82249
rect 579250 82175 579306 82184
rect 578976 80708 579028 80714
rect 578976 80650 579028 80656
rect 578790 80064 578846 80073
rect 578790 79999 578846 80008
rect 578988 77897 579016 80650
rect 579160 80096 579212 80102
rect 579160 80038 579212 80044
rect 578974 77888 579030 77897
rect 578974 77823 579030 77832
rect 578884 75948 578936 75954
rect 578884 75890 578936 75896
rect 578700 75472 578752 75478
rect 578698 75440 578700 75449
rect 578752 75440 578754 75449
rect 578698 75375 578754 75384
rect 578516 73160 578568 73166
rect 578514 73128 578516 73137
rect 578568 73128 578570 73137
rect 578514 73063 578570 73072
rect 578516 62076 578568 62082
rect 578516 62018 578568 62024
rect 578528 61849 578556 62018
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 577688 58676 577740 58682
rect 577688 58618 577740 58624
rect 577504 54392 577556 54398
rect 577504 54334 577556 54340
rect 577700 54233 577728 58618
rect 578896 55078 578924 75890
rect 579172 71369 579200 80038
rect 580276 73166 580304 93094
rect 580460 86630 580488 106898
rect 580644 95062 580672 107034
rect 581644 104916 581696 104922
rect 581644 104858 581696 104864
rect 580632 95056 580684 95062
rect 580632 94998 580684 95004
rect 580448 86624 580500 86630
rect 580448 86566 580500 86572
rect 581656 75478 581684 104858
rect 581840 84182 581868 109686
rect 583036 103358 583064 128318
rect 584416 124166 584444 139402
rect 585796 134298 585824 144910
rect 587360 135930 587388 146270
rect 589200 145586 589228 149223
rect 589370 147656 589426 147665
rect 589370 147591 589426 147600
rect 589384 146334 589412 147591
rect 589372 146328 589424 146334
rect 589372 146270 589424 146276
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589188 145580 589240 145586
rect 589188 145522 589240 145528
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589922 144392 589978 144401
rect 589922 144327 589978 144336
rect 589462 142760 589518 142769
rect 589462 142695 589518 142704
rect 589476 142186 589504 142695
rect 589464 142180 589516 142186
rect 589464 142122 589516 142128
rect 589094 141128 589150 141137
rect 589094 141063 589150 141072
rect 587348 135924 587400 135930
rect 587348 135866 587400 135872
rect 587164 135312 587216 135318
rect 587164 135254 587216 135260
rect 585784 134292 585836 134298
rect 585784 134234 585836 134240
rect 585968 133952 586020 133958
rect 585968 133894 586020 133900
rect 585784 124228 585836 124234
rect 585784 124170 585836 124176
rect 584404 124160 584456 124166
rect 584404 124102 584456 124108
rect 584404 121508 584456 121514
rect 584404 121450 584456 121456
rect 583208 117360 583260 117366
rect 583208 117302 583260 117308
rect 583024 103352 583076 103358
rect 583024 103294 583076 103300
rect 583220 93294 583248 117302
rect 584416 97510 584444 121450
rect 585140 115388 585192 115394
rect 585140 115330 585192 115336
rect 585152 108390 585180 115330
rect 585140 108384 585192 108390
rect 585140 108326 585192 108332
rect 585796 99210 585824 124170
rect 585980 116958 586008 133894
rect 587176 118658 587204 135254
rect 589108 133210 589136 141063
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589278 136232 589334 136241
rect 589278 136167 589334 136176
rect 589292 135318 589320 136167
rect 589280 135312 589332 135318
rect 589280 135254 589332 135260
rect 589462 134600 589518 134609
rect 589462 134535 589518 134544
rect 589476 133958 589504 134535
rect 589464 133952 589516 133958
rect 589464 133894 589516 133900
rect 589096 133204 589148 133210
rect 589096 133146 589148 133152
rect 588542 132968 588598 132977
rect 588542 132903 588598 132912
rect 587164 118652 587216 118658
rect 587164 118594 587216 118600
rect 585968 116952 586020 116958
rect 585968 116894 586020 116900
rect 587808 116000 587860 116006
rect 587808 115942 587860 115948
rect 587820 115258 587848 115942
rect 587808 115252 587860 115258
rect 587808 115194 587860 115200
rect 587164 114572 587216 114578
rect 587164 114514 587216 114520
rect 585968 100768 586020 100774
rect 585968 100710 586020 100716
rect 585784 99204 585836 99210
rect 585784 99146 585836 99152
rect 584404 97504 584456 97510
rect 584404 97446 584456 97452
rect 583208 93288 583260 93294
rect 583208 93230 583260 93236
rect 581828 84176 581880 84182
rect 581828 84118 581880 84124
rect 585980 80102 586008 100710
rect 587176 88330 587204 114514
rect 588556 113150 588584 132903
rect 589936 131782 589964 144327
rect 589924 131776 589976 131782
rect 589924 131718 589976 131724
rect 590106 131336 590162 131345
rect 590106 131271 590162 131280
rect 589462 129704 589518 129713
rect 589462 129639 589518 129648
rect 589476 128382 589504 129639
rect 589464 128376 589516 128382
rect 589464 128318 589516 128324
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589922 126440 589978 126449
rect 589922 126375 589978 126384
rect 589462 124808 589518 124817
rect 589462 124743 589518 124752
rect 589476 124234 589504 124743
rect 589464 124228 589516 124234
rect 589464 124170 589516 124176
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589462 121544 589518 121553
rect 589462 121479 589464 121488
rect 589516 121479 589518 121488
rect 589464 121450 589516 121456
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589936 115394 589964 126375
rect 590120 120766 590148 131271
rect 590108 120760 590160 120766
rect 590108 120702 590160 120708
rect 590106 119912 590162 119921
rect 590106 119847 590162 119856
rect 589924 115388 589976 115394
rect 589924 115330 589976 115336
rect 589830 115016 589886 115025
rect 589830 114951 589886 114960
rect 589844 114578 589872 114951
rect 589832 114572 589884 114578
rect 589832 114514 589884 114520
rect 588544 113144 588596 113150
rect 588544 113086 588596 113092
rect 589370 111752 589426 111761
rect 589370 111687 589426 111696
rect 588544 110492 588596 110498
rect 588544 110434 588596 110440
rect 587164 88324 587216 88330
rect 587164 88266 587216 88272
rect 588556 82822 588584 110434
rect 589384 109750 589412 111687
rect 589646 110120 589702 110129
rect 589646 110055 589702 110064
rect 589372 109744 589424 109750
rect 589372 109686 589424 109692
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589660 106962 589688 110055
rect 590120 107098 590148 119847
rect 591316 114442 591344 208626
rect 666204 160177 666232 236127
rect 666388 209774 666416 338098
rect 666652 324352 666704 324358
rect 666652 324294 666704 324300
rect 666388 209746 666508 209774
rect 666480 186969 666508 209746
rect 666466 186960 666522 186969
rect 666466 186895 666522 186904
rect 666664 178809 666692 324294
rect 667216 313721 667244 456758
rect 667860 456113 667888 660991
rect 668044 621761 668072 686151
rect 668412 659705 668440 733071
rect 668596 670449 668624 789346
rect 668780 755993 668808 877639
rect 668950 783864 669006 783873
rect 668950 783799 669006 783808
rect 668766 755984 668822 755993
rect 668766 755919 668822 755928
rect 668766 731504 668822 731513
rect 668766 731439 668822 731448
rect 668582 670440 668638 670449
rect 668582 670375 668638 670384
rect 668780 664601 668808 731439
rect 668964 708801 668992 783799
rect 669240 753545 669268 879135
rect 670514 874032 670570 874041
rect 670514 873967 670570 873976
rect 669594 872264 669650 872273
rect 669594 872199 669650 872208
rect 669608 755449 669636 872199
rect 669964 841832 670016 841838
rect 669964 841774 670016 841780
rect 669778 789440 669834 789449
rect 669778 789375 669834 789384
rect 669594 755440 669650 755449
rect 669594 755375 669650 755384
rect 669226 753536 669282 753545
rect 669226 753471 669282 753480
rect 669410 741840 669466 741849
rect 669410 741775 669466 741784
rect 669134 734496 669190 734505
rect 669134 734431 669190 734440
rect 669148 721754 669176 734431
rect 669056 721726 669176 721754
rect 669056 708914 669084 721726
rect 669056 708886 669176 708914
rect 668950 708792 669006 708801
rect 668950 708727 669006 708736
rect 669148 707954 669176 708886
rect 669056 707926 669176 707954
rect 668766 664592 668822 664601
rect 668766 664527 668822 664536
rect 669056 662561 669084 707926
rect 669226 701176 669282 701185
rect 669226 701111 669282 701120
rect 669042 662552 669098 662561
rect 669042 662487 669098 662496
rect 668398 659696 668454 659705
rect 668398 659631 668454 659640
rect 668214 647320 668270 647329
rect 668214 647255 668270 647264
rect 668030 621752 668086 621761
rect 668030 621687 668086 621696
rect 668228 574841 668256 647255
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668398 608016 668454 608025
rect 668398 607951 668454 607960
rect 668214 574832 668270 574841
rect 668214 574767 668270 574776
rect 668214 557560 668270 557569
rect 668214 557495 668270 557504
rect 668228 486033 668256 557495
rect 668412 530641 668440 607951
rect 668596 535945 668624 643078
rect 668950 638752 669006 638761
rect 668950 638687 669006 638696
rect 668766 593600 668822 593609
rect 668766 593535 668822 593544
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668398 530632 668454 530641
rect 668398 530567 668454 530576
rect 668780 528601 668808 593535
rect 668964 574433 668992 638687
rect 669240 622033 669268 701111
rect 669424 663377 669452 741775
rect 669594 738576 669650 738585
rect 669594 738511 669650 738520
rect 669608 666369 669636 738511
rect 669792 709617 669820 789375
rect 669976 715737 670004 841774
rect 670330 780056 670386 780065
rect 670330 779991 670386 780000
rect 670146 778968 670202 778977
rect 670146 778903 670202 778912
rect 670160 777073 670188 778903
rect 670146 777064 670202 777073
rect 670146 776999 670202 777008
rect 670146 775024 670202 775033
rect 670146 774959 670202 774968
rect 669962 715728 670018 715737
rect 669962 715663 670018 715672
rect 669778 709608 669834 709617
rect 669778 709543 669834 709552
rect 670160 705945 670188 774959
rect 670344 707169 670372 779991
rect 670528 754225 670556 873967
rect 670514 754216 670570 754225
rect 670514 754151 670570 754160
rect 670712 734097 670740 929455
rect 671344 895688 671396 895694
rect 671344 895630 671396 895636
rect 671158 867232 671214 867241
rect 671158 867167 671214 867176
rect 670974 778424 671030 778433
rect 670974 778359 671030 778368
rect 670988 776529 671016 778359
rect 670974 776520 671030 776529
rect 670974 776455 671030 776464
rect 670882 757480 670938 757489
rect 670882 757415 670938 757424
rect 670698 734088 670754 734097
rect 670698 734023 670754 734032
rect 670698 728512 670754 728521
rect 670698 728447 670700 728456
rect 670752 728447 670754 728456
rect 670700 728418 670752 728424
rect 670896 721754 670924 757415
rect 671172 753409 671200 867167
rect 671356 763065 671384 895630
rect 671342 763056 671398 763065
rect 671342 762991 671398 763000
rect 671632 760345 671660 937751
rect 671618 760336 671674 760345
rect 671618 760271 671674 760280
rect 671618 759928 671674 759937
rect 671618 759863 671674 759872
rect 671158 753400 671214 753409
rect 671158 753335 671214 753344
rect 671066 751360 671122 751369
rect 671066 751295 671122 751304
rect 671080 728113 671108 751295
rect 671434 750136 671490 750145
rect 671434 750071 671490 750080
rect 671250 737080 671306 737089
rect 671250 737015 671306 737024
rect 671066 728104 671122 728113
rect 671066 728039 671122 728048
rect 670896 721726 671108 721754
rect 670882 713280 670938 713289
rect 670882 713215 670938 713224
rect 670330 707160 670386 707169
rect 670330 707095 670386 707104
rect 670146 705936 670202 705945
rect 670146 705871 670202 705880
rect 669778 696960 669834 696969
rect 669778 696895 669834 696904
rect 669594 666360 669650 666369
rect 669594 666295 669650 666304
rect 669410 663368 669466 663377
rect 669410 663303 669466 663312
rect 669226 622024 669282 622033
rect 669226 621959 669282 621968
rect 669792 620673 669820 696895
rect 670422 690432 670478 690441
rect 670422 690367 670478 690376
rect 670238 685400 670294 685409
rect 670238 685335 670294 685344
rect 669964 683188 670016 683194
rect 669964 683130 670016 683136
rect 669778 620664 669834 620673
rect 669778 620599 669834 620608
rect 669778 616176 669834 616185
rect 669778 616111 669834 616120
rect 669226 608560 669282 608569
rect 669226 608495 669282 608504
rect 668950 574424 669006 574433
rect 668950 574359 669006 574368
rect 669042 564496 669098 564505
rect 669042 564431 669098 564440
rect 668766 528592 668822 528601
rect 668766 528527 668822 528536
rect 668214 486024 668270 486033
rect 668214 485959 668270 485968
rect 669056 485081 669084 564431
rect 669240 529009 669268 608495
rect 669594 554704 669650 554713
rect 669594 554639 669650 554648
rect 669226 529000 669282 529009
rect 669226 528935 669282 528944
rect 669042 485072 669098 485081
rect 669042 485007 669098 485016
rect 669608 482769 669636 554639
rect 669594 482760 669650 482769
rect 669594 482695 669650 482704
rect 667846 456104 667902 456113
rect 667846 456039 667902 456048
rect 669792 455161 669820 616111
rect 669976 580145 670004 683130
rect 670252 615777 670280 685335
rect 670436 620265 670464 690367
rect 670896 668273 670924 713215
rect 671080 712881 671108 721726
rect 671066 712872 671122 712881
rect 671066 712807 671122 712816
rect 671066 712464 671122 712473
rect 671066 712399 671122 712408
rect 670882 668264 670938 668273
rect 670882 668199 670938 668208
rect 670882 667992 670938 668001
rect 670882 667927 670938 667936
rect 670606 659968 670662 659977
rect 670606 659903 670662 659912
rect 670422 620256 670478 620265
rect 670422 620191 670478 620200
rect 670238 615768 670294 615777
rect 670238 615703 670294 615712
rect 670422 614952 670478 614961
rect 670422 614887 670478 614896
rect 670238 600672 670294 600681
rect 670238 600607 670294 600616
rect 669962 580136 670018 580145
rect 669962 580071 670018 580080
rect 670054 554024 670110 554033
rect 670054 553959 670110 553968
rect 670068 551585 670096 553959
rect 670054 551576 670110 551585
rect 670054 551511 670110 551520
rect 669964 536852 670016 536858
rect 669964 536794 670016 536800
rect 669778 455152 669834 455161
rect 669778 455087 669834 455096
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667388 350600 667440 350606
rect 667388 350542 667440 350548
rect 667202 313712 667258 313721
rect 667202 313647 667258 313656
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 666836 229628 666888 229634
rect 666836 229570 666888 229576
rect 666848 222873 666876 229570
rect 667020 225480 667072 225486
rect 667020 225422 667072 225428
rect 667032 225321 667060 225422
rect 667018 225312 667074 225321
rect 667018 225247 667074 225256
rect 667018 224224 667074 224233
rect 667018 224159 667020 224168
rect 667072 224159 667074 224168
rect 667020 224130 667072 224136
rect 666834 222864 666890 222873
rect 666834 222799 666890 222808
rect 666834 217288 666890 217297
rect 666834 217223 666890 217232
rect 666848 198393 666876 217223
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 198384 666890 198393
rect 666834 198319 666890 198328
rect 666650 178800 666706 178809
rect 666650 178735 666706 178744
rect 666190 160168 666246 160177
rect 666190 160103 666246 160112
rect 667032 133113 667060 209034
rect 667216 134609 667244 310490
rect 667400 181393 667428 350542
rect 668596 311953 668624 444382
rect 669976 403753 670004 536794
rect 670252 530097 670280 600607
rect 670238 530088 670294 530097
rect 670238 530023 670294 530032
rect 670148 484424 670200 484430
rect 670148 484366 670200 484372
rect 669962 403744 670018 403753
rect 669962 403679 670018 403688
rect 670160 360913 670188 484366
rect 670436 455433 670464 614887
rect 670620 455841 670648 659903
rect 670896 623529 670924 667927
rect 671080 666641 671108 712399
rect 671066 666632 671122 666641
rect 671066 666567 671122 666576
rect 671264 661337 671292 737015
rect 671448 728385 671476 750071
rect 671434 728376 671490 728385
rect 671434 728311 671490 728320
rect 671632 715329 671660 759863
rect 671816 759529 671844 938023
rect 672446 936456 672502 936465
rect 672446 936391 672502 936400
rect 672460 765914 672488 936391
rect 672630 935776 672686 935785
rect 672630 935711 672686 935720
rect 672644 794894 672672 935711
rect 673104 933201 673132 943906
rect 673090 933192 673146 933201
rect 673090 933127 673146 933136
rect 673288 933042 673316 943906
rect 673196 933014 673316 933042
rect 673196 930753 673224 933014
rect 673380 932929 673408 966583
rect 675128 966090 675156 966583
rect 675680 966521 675708 966723
rect 675666 966512 675722 966521
rect 675666 966447 675722 966456
rect 675128 966062 675418 966090
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675298 964744 675354 964753
rect 675298 964679 675354 964688
rect 675312 963254 675340 964679
rect 675496 963393 675524 963595
rect 675482 963384 675538 963393
rect 675482 963319 675538 963328
rect 675220 963226 675340 963254
rect 674286 962840 674342 962849
rect 674286 962775 674342 962784
rect 674102 957128 674158 957137
rect 674102 957063 674158 957072
rect 673366 932920 673422 932929
rect 673366 932855 673422 932864
rect 673182 930744 673238 930753
rect 673182 930679 673238 930688
rect 674116 930209 674144 957063
rect 674300 932657 674328 962775
rect 675220 962418 675248 963226
rect 675496 962849 675524 963016
rect 675482 962840 675538 962849
rect 675482 962775 675538 962784
rect 675220 962390 675418 962418
rect 675128 961741 675418 961769
rect 675128 960809 675156 961741
rect 675114 960800 675170 960809
rect 675114 960735 675170 960744
rect 674484 959262 675418 959290
rect 674484 933881 674512 959262
rect 674930 959168 674986 959177
rect 674930 959103 674986 959112
rect 674654 958760 674710 958769
rect 674654 958695 674710 958704
rect 674470 933872 674526 933881
rect 674470 933807 674526 933816
rect 674286 932648 674342 932657
rect 674286 932583 674342 932592
rect 674668 930481 674696 958695
rect 674944 953594 674972 959103
rect 675206 958760 675262 958769
rect 675262 958718 675418 958746
rect 675206 958695 675262 958704
rect 675772 957817 675800 958052
rect 675298 957808 675354 957817
rect 675298 957743 675354 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 675312 955482 675340 957743
rect 675496 957137 675524 957440
rect 675482 957128 675538 957137
rect 675482 957063 675538 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675206 954680 675262 954689
rect 675206 954615 675262 954624
rect 674944 953566 675156 953594
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 930472 674710 930481
rect 674654 930407 674710 930416
rect 674102 930200 674158 930209
rect 674102 930135 674158 930144
rect 674852 928792 674880 953391
rect 675128 934153 675156 953566
rect 675220 943934 675248 954615
rect 675312 954366 675418 954394
rect 675312 949498 675340 954366
rect 675496 953465 675524 953768
rect 675482 953456 675538 953465
rect 675482 953391 675538 953400
rect 675588 952241 675616 952544
rect 675574 952232 675630 952241
rect 675574 952167 675630 952176
rect 683302 950736 683358 950745
rect 683302 950671 683358 950680
rect 679622 949512 679678 949521
rect 675312 949482 675892 949498
rect 675312 949476 675904 949482
rect 675312 949470 675852 949476
rect 679622 949447 679678 949456
rect 682384 949476 682436 949482
rect 675852 949418 675904 949424
rect 675220 943906 675340 943934
rect 675312 934697 675340 943906
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676494 937680 676550 937689
rect 676494 937615 676550 937624
rect 676508 936873 676536 937615
rect 676494 936864 676550 936873
rect 676494 936799 676550 936808
rect 679636 935649 679664 949447
rect 682384 949418 682436 949424
rect 679622 935640 679678 935649
rect 679622 935575 679678 935584
rect 682396 935241 682424 949418
rect 683118 947336 683174 947345
rect 683118 947271 683174 947280
rect 683132 939729 683160 947271
rect 683118 939720 683174 939729
rect 683118 939655 683174 939664
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 675298 934688 675354 934697
rect 675298 934623 675354 934632
rect 675114 934144 675170 934153
rect 675114 934079 675170 934088
rect 683316 932385 683344 950671
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683302 932376 683358 932385
rect 683302 932311 683358 932320
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 673366 928296 673422 928305
rect 673366 928231 673422 928240
rect 673090 868456 673146 868465
rect 673090 868391 673146 868400
rect 672644 794866 672764 794894
rect 672736 785234 672764 794866
rect 672736 785206 672856 785234
rect 672630 784272 672686 784281
rect 672630 784207 672686 784216
rect 672644 775574 672672 784207
rect 672828 780450 672856 785206
rect 672368 765886 672488 765914
rect 672552 775546 672672 775574
rect 672736 780422 672856 780450
rect 672172 761932 672224 761938
rect 672172 761874 672224 761880
rect 671802 759520 671858 759529
rect 671802 759455 671858 759464
rect 671802 758296 671858 758305
rect 671802 758231 671858 758240
rect 671618 715320 671674 715329
rect 671618 715255 671674 715264
rect 671618 714912 671674 714921
rect 671618 714847 671674 714856
rect 671434 714096 671490 714105
rect 671434 714031 671490 714040
rect 671448 669905 671476 714031
rect 671632 670177 671660 714847
rect 671816 713697 671844 758231
rect 672184 757897 672212 761874
rect 672368 758713 672396 765886
rect 672354 758704 672410 758713
rect 672354 758639 672410 758648
rect 672170 757888 672226 757897
rect 672170 757823 672226 757832
rect 672262 743472 672318 743481
rect 672262 743407 672318 743416
rect 672078 741160 672134 741169
rect 672078 741095 672134 741104
rect 672092 731414 672120 741095
rect 672092 731386 672212 731414
rect 671986 730552 672042 730561
rect 671986 730487 672042 730496
rect 671802 713688 671858 713697
rect 671802 713623 671858 713632
rect 671802 687440 671858 687449
rect 671802 687375 671858 687384
rect 671618 670168 671674 670177
rect 671618 670103 671674 670112
rect 671434 669896 671490 669905
rect 671434 669831 671490 669840
rect 671618 669488 671674 669497
rect 671618 669423 671674 669432
rect 671434 668672 671490 668681
rect 671434 668607 671490 668616
rect 671250 661328 671306 661337
rect 671250 661263 671306 661272
rect 671448 630674 671476 668607
rect 671264 630646 671476 630674
rect 671066 624744 671122 624753
rect 671066 624679 671122 624688
rect 670882 623520 670938 623529
rect 670882 623455 670938 623464
rect 670882 622840 670938 622849
rect 670882 622775 670938 622784
rect 670896 577697 670924 622775
rect 671080 621014 671108 624679
rect 671264 624345 671292 630646
rect 671632 625161 671660 669423
rect 671816 647234 671844 687375
rect 672000 666097 672028 730487
rect 672184 721754 672212 731386
rect 672092 721726 672212 721754
rect 672092 673454 672120 721726
rect 672092 673426 672212 673454
rect 671986 666088 672042 666097
rect 671986 666023 672042 666032
rect 672184 665938 672212 673426
rect 672092 665910 672212 665938
rect 672092 663921 672120 665910
rect 672276 665825 672304 743407
rect 672552 709209 672580 775546
rect 672736 761938 672764 780422
rect 672906 773800 672962 773809
rect 672906 773735 672962 773744
rect 672724 761932 672776 761938
rect 672724 761874 672776 761880
rect 672722 759112 672778 759121
rect 672722 759047 672778 759056
rect 672736 714513 672764 759047
rect 672722 714504 672778 714513
rect 672722 714439 672778 714448
rect 672920 710025 672948 773735
rect 673104 751777 673132 868391
rect 673090 751768 673146 751777
rect 673090 751703 673146 751712
rect 673090 733680 673146 733689
rect 673090 733615 673146 733624
rect 672906 710016 672962 710025
rect 672906 709951 672962 709960
rect 672538 709200 672594 709209
rect 672538 709135 672594 709144
rect 672446 685944 672502 685953
rect 672446 685879 672502 685888
rect 672262 665816 672318 665825
rect 672262 665751 672318 665760
rect 672078 663912 672134 663921
rect 672078 663847 672134 663856
rect 671986 654256 672042 654265
rect 671986 654191 672042 654200
rect 672000 649994 672028 654191
rect 671724 647206 671844 647234
rect 671908 649966 672028 649994
rect 671908 647234 671936 649966
rect 671908 647206 672120 647234
rect 671724 637574 671752 647206
rect 671894 643512 671950 643521
rect 671894 643447 671950 643456
rect 671724 637546 671844 637574
rect 671618 625152 671674 625161
rect 671618 625087 671674 625096
rect 671816 625002 671844 637546
rect 671448 624974 671844 625002
rect 671250 624336 671306 624345
rect 671250 624271 671306 624280
rect 671080 620986 671292 621014
rect 671264 611354 671292 620986
rect 671448 618225 671476 624974
rect 671618 622432 671674 622441
rect 671618 622367 671674 622376
rect 671434 618216 671490 618225
rect 671434 618151 671490 618160
rect 671632 611354 671660 622367
rect 671264 611326 671476 611354
rect 671632 611326 671752 611354
rect 671066 594824 671122 594833
rect 671066 594759 671122 594768
rect 670882 577688 670938 577697
rect 670882 577623 670938 577632
rect 670882 552120 670938 552129
rect 670882 552055 670938 552064
rect 670896 483993 670924 552055
rect 671080 525745 671108 594759
rect 671448 580553 671476 611326
rect 671434 580544 671490 580553
rect 671434 580479 671490 580488
rect 671342 578912 671398 578921
rect 671342 578847 671398 578856
rect 671356 577810 671384 578847
rect 671526 578096 671582 578105
rect 671526 578031 671582 578040
rect 671172 577782 671384 577810
rect 671172 567194 671200 577782
rect 671342 576872 671398 576881
rect 671342 576807 671398 576816
rect 671172 567166 671292 567194
rect 671264 534857 671292 567166
rect 671356 557534 671384 576807
rect 671540 557534 671568 578031
rect 671724 577289 671752 611326
rect 671710 577280 671766 577289
rect 671710 577215 671766 577224
rect 671908 576854 671936 643447
rect 672092 637574 672120 647206
rect 671816 576826 671936 576854
rect 672000 637546 672120 637574
rect 671816 571169 671844 576826
rect 672000 574161 672028 637546
rect 672262 623928 672318 623937
rect 672262 623863 672318 623872
rect 672276 618390 672304 623863
rect 672460 619857 672488 685879
rect 672630 667040 672686 667049
rect 672630 666975 672686 666984
rect 672644 635497 672672 666975
rect 673104 661609 673132 733615
rect 673380 728618 673408 928231
rect 675022 879200 675078 879209
rect 675022 879135 675078 879144
rect 675036 877305 675064 879135
rect 675482 877704 675538 877713
rect 675482 877639 675538 877648
rect 675496 877540 675524 877639
rect 675022 877296 675078 877305
rect 675022 877231 675078 877240
rect 675390 877296 675446 877305
rect 675390 877231 675446 877240
rect 675404 876860 675432 877231
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675680 874041 675708 874412
rect 675482 874032 675538 874041
rect 675482 873967 675538 873976
rect 675666 874032 675722 874041
rect 675666 873967 675722 873976
rect 675496 873868 675524 873967
rect 674484 873174 675418 873202
rect 674010 868048 674066 868057
rect 674010 867983 674066 867992
rect 673734 779240 673790 779249
rect 673734 779175 673790 779184
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673368 728612 673420 728618
rect 673368 728554 673420 728560
rect 673366 728376 673422 728385
rect 673366 728311 673368 728320
rect 673420 728311 673422 728320
rect 673368 728282 673420 728288
rect 673368 728136 673420 728142
rect 673366 728104 673368 728113
rect 673420 728104 673422 728113
rect 673366 728039 673422 728048
rect 673564 708393 673592 777407
rect 673748 725121 673776 779175
rect 674024 775574 674052 867983
rect 674484 854321 674512 873174
rect 675588 872273 675616 872576
rect 675114 872264 675170 872273
rect 675114 872199 675170 872208
rect 675574 872264 675630 872273
rect 675574 872199 675630 872208
rect 675128 870074 675156 872199
rect 675128 870046 675418 870074
rect 675114 869544 675170 869553
rect 675170 869502 675418 869530
rect 675114 869479 675170 869488
rect 675128 868861 675418 868889
rect 675128 868057 675156 868861
rect 675298 868728 675354 868737
rect 675298 868663 675354 868672
rect 675114 868048 675170 868057
rect 675114 867983 675170 867992
rect 674930 866688 674986 866697
rect 674930 866623 674986 866632
rect 674654 864784 674710 864793
rect 674654 864719 674710 864728
rect 674470 854312 674526 854321
rect 674470 854247 674526 854256
rect 674470 788080 674526 788089
rect 674470 788015 674526 788024
rect 674286 783048 674342 783057
rect 674286 782983 674342 782992
rect 674300 778818 674328 782983
rect 674300 778790 674420 778818
rect 674194 778696 674250 778705
rect 674194 778631 674250 778640
rect 673932 775546 674052 775574
rect 673932 770681 673960 775546
rect 673918 770672 673974 770681
rect 673918 770607 673974 770616
rect 674208 731414 674236 778631
rect 674392 775574 674420 778790
rect 674116 731386 674236 731414
rect 674300 775546 674420 775574
rect 674116 726889 674144 731386
rect 674300 727977 674328 775546
rect 674286 727968 674342 727977
rect 674286 727903 674342 727912
rect 674102 726880 674158 726889
rect 674102 726815 674158 726824
rect 674484 726594 674512 788015
rect 674668 787250 674696 864719
rect 674944 864566 674972 866623
rect 675312 865858 675340 868663
rect 675482 868456 675538 868465
rect 675482 868391 675538 868400
rect 675496 868224 675524 868391
rect 675482 867232 675538 867241
rect 675482 867167 675538 867176
rect 675496 867035 675524 867167
rect 675312 865830 675418 865858
rect 675220 865181 675418 865209
rect 675220 864793 675248 865181
rect 675206 864784 675262 864793
rect 675206 864719 675262 864728
rect 674944 864538 675418 864566
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675220 863314 675340 863342
rect 675404 863328 675432 863382
rect 675220 794894 675248 863314
rect 674852 794866 675248 794894
rect 674852 787273 674880 794866
rect 675206 789440 675262 789449
rect 675206 789375 675262 789384
rect 675220 787693 675248 789375
rect 675404 788089 675432 788324
rect 675390 788080 675446 788089
rect 675390 788015 675446 788024
rect 675220 787665 675418 787693
rect 674576 787222 674696 787250
rect 674838 787264 674894 787273
rect 674576 782898 674604 787222
rect 674838 787199 674894 787208
rect 675404 786729 675432 787032
rect 675390 786720 675446 786729
rect 675390 786655 675446 786664
rect 675404 784938 675432 785196
rect 675128 784910 675432 784938
rect 675128 783442 675156 784910
rect 675496 784281 675524 784652
rect 675482 784272 675538 784281
rect 675482 784207 675538 784216
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 674760 783414 675156 783442
rect 674760 783170 674788 783414
rect 674930 783320 674986 783329
rect 674930 783255 674986 783264
rect 674760 783142 674880 783170
rect 674576 782870 674788 782898
rect 674760 772041 674788 782870
rect 674852 780314 674880 783142
rect 674944 780450 674972 783255
rect 675404 783057 675432 783360
rect 675390 783048 675446 783057
rect 675390 782983 675446 782992
rect 675114 782776 675170 782785
rect 675114 782711 675170 782720
rect 675128 780745 675156 782711
rect 675298 782504 675354 782513
rect 675298 782439 675354 782448
rect 675312 781402 675340 782439
rect 675312 781374 675432 781402
rect 675404 780844 675432 781374
rect 675114 780736 675170 780745
rect 675114 780671 675170 780680
rect 674944 780422 675156 780450
rect 674852 780286 675064 780314
rect 675036 772814 675064 780286
rect 674944 772786 675064 772814
rect 674746 772032 674802 772041
rect 674746 771967 674802 771976
rect 674944 771882 674972 772786
rect 675128 772562 675156 780422
rect 675496 780065 675524 780300
rect 675482 780056 675538 780065
rect 675482 779991 675538 780000
rect 675312 779674 675418 779702
rect 675312 779249 675340 779674
rect 675298 779240 675354 779249
rect 675298 779175 675354 779184
rect 675496 778705 675524 779008
rect 675482 778696 675538 778705
rect 675482 778631 675538 778640
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675390 777064 675446 777073
rect 675390 776999 675446 777008
rect 675404 776628 675432 776999
rect 675482 776520 675538 776529
rect 675482 776455 675538 776464
rect 675496 776016 675524 776455
rect 675496 775033 675524 775336
rect 675482 775024 675538 775033
rect 675482 774959 675538 774968
rect 675496 773809 675524 774180
rect 675482 773800 675538 773809
rect 675482 773735 675538 773744
rect 682382 772712 682438 772721
rect 682382 772647 682438 772656
rect 675128 772534 675248 772562
rect 674852 771854 674972 771882
rect 674852 765105 674880 771854
rect 675220 766601 675248 772534
rect 681002 768768 681058 768777
rect 681002 768703 681058 768712
rect 675206 766592 675262 766601
rect 675206 766527 675262 766536
rect 674838 765096 674894 765105
rect 674838 765031 674894 765040
rect 676034 763056 676090 763065
rect 676034 762991 676090 763000
rect 676048 760753 676076 762991
rect 676954 761832 677010 761841
rect 676586 761788 676642 761797
rect 676954 761767 677010 761776
rect 676586 761723 676642 761732
rect 676034 760744 676090 760753
rect 676034 760679 676090 760688
rect 676600 757178 676628 761723
rect 676036 757172 676088 757178
rect 676036 757114 676088 757120
rect 676588 757172 676640 757178
rect 676588 757114 676640 757120
rect 675850 754760 675906 754769
rect 675850 754695 675906 754704
rect 675864 754322 675892 754695
rect 675852 754316 675904 754322
rect 675852 754258 675904 754264
rect 676048 752593 676076 757114
rect 676968 755041 676996 761767
rect 681016 757081 681044 768703
rect 681002 757072 681058 757081
rect 681002 757007 681058 757016
rect 682396 755857 682424 772647
rect 683210 772032 683266 772041
rect 683210 771967 683266 771976
rect 683224 756673 683252 771967
rect 683394 770672 683450 770681
rect 683394 770607 683450 770616
rect 683210 756664 683266 756673
rect 683210 756599 683266 756608
rect 682382 755848 682438 755857
rect 682382 755783 682438 755792
rect 676954 755032 677010 755041
rect 676954 754967 677010 754976
rect 683120 754316 683172 754322
rect 683120 754258 683172 754264
rect 676034 752584 676090 752593
rect 676034 752519 676090 752528
rect 683132 752185 683160 754258
rect 683408 753001 683436 770607
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683394 752992 683450 753001
rect 683394 752927 683450 752936
rect 683118 752176 683174 752185
rect 683118 752111 683174 752120
rect 674930 743472 674986 743481
rect 674930 743407 674986 743416
rect 674944 742710 674972 743407
rect 675128 743294 675418 743322
rect 675128 743209 675156 743294
rect 675114 743200 675170 743209
rect 675114 743135 675170 743144
rect 674944 742682 675340 742710
rect 675312 742642 675340 742682
rect 675404 742642 675432 742696
rect 675312 742614 675432 742642
rect 675022 742520 675078 742529
rect 675022 742455 675078 742464
rect 674838 741840 674894 741849
rect 674838 741775 674894 741784
rect 674852 741282 674880 741775
rect 675036 741690 675064 742455
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 674944 741662 675064 741690
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 674944 741418 674972 741662
rect 675128 741577 675156 742002
rect 675114 741568 675170 741577
rect 675114 741503 675170 741512
rect 674944 741390 675156 741418
rect 674760 741254 674880 741282
rect 674760 741010 674788 741254
rect 674930 741160 674986 741169
rect 674930 741095 674986 741104
rect 674760 740982 674880 741010
rect 674852 739038 674880 740982
rect 674944 739650 674972 741095
rect 675128 740194 675156 741390
rect 675128 740166 675418 740194
rect 674944 739622 675418 739650
rect 674852 739010 675340 739038
rect 675312 738970 675340 739010
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675298 738576 675354 738585
rect 675298 738511 675354 738520
rect 675114 737080 675170 737089
rect 675114 737015 675170 737024
rect 675128 735333 675156 737015
rect 675312 735842 675340 738511
rect 675496 738177 675524 738344
rect 675482 738168 675538 738177
rect 675482 738103 675538 738112
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675128 735305 675418 735333
rect 674930 734768 674986 734777
rect 674930 734703 674986 734712
rect 674654 733136 674710 733145
rect 674710 733094 674880 733122
rect 674654 733071 674710 733080
rect 674852 731626 674880 733094
rect 674944 732714 674972 734703
rect 675128 734658 675418 734686
rect 675128 734505 675156 734658
rect 675114 734496 675170 734505
rect 675114 734431 675170 734440
rect 675128 734017 675418 734045
rect 675128 733689 675156 734017
rect 675114 733680 675170 733689
rect 675114 733615 675170 733624
rect 675114 732864 675170 732873
rect 675170 732822 675418 732850
rect 675114 732799 675170 732808
rect 674944 732686 675064 732714
rect 675036 731626 675064 732686
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674852 731598 674972 731626
rect 675036 731598 675340 731626
rect 675404 731612 675432 731734
rect 674654 731504 674710 731513
rect 674710 731462 674880 731490
rect 674654 731439 674710 731448
rect 674852 729178 674880 731462
rect 674944 730365 674972 731598
rect 675128 730986 675418 731014
rect 675128 730561 675156 730986
rect 675114 730552 675170 730561
rect 675114 730487 675170 730496
rect 674944 730337 675418 730365
rect 674852 729150 675418 729178
rect 683762 727968 683818 727977
rect 683762 727903 683818 727912
rect 683210 726744 683266 726753
rect 683210 726679 683266 726688
rect 674746 726608 674802 726617
rect 674484 726566 674746 726594
rect 674746 726543 674802 726552
rect 682382 725792 682438 725801
rect 682382 725727 682438 725736
rect 673734 725112 673790 725121
rect 673734 725047 673790 725056
rect 682396 710841 682424 725727
rect 682382 710832 682438 710841
rect 682382 710767 682438 710776
rect 673550 708384 673606 708393
rect 673550 708319 673606 708328
rect 683224 706761 683252 726679
rect 683394 726472 683450 726481
rect 683394 726407 683450 726416
rect 683408 711249 683436 726407
rect 683578 725112 683634 725121
rect 683578 725047 683634 725056
rect 683394 711240 683450 711249
rect 683394 711175 683450 711184
rect 683592 707985 683620 725047
rect 683578 707976 683634 707985
rect 683578 707911 683634 707920
rect 683776 707577 683804 727903
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683762 707568 683818 707577
rect 683762 707503 683818 707512
rect 683210 706752 683266 706761
rect 683210 706687 683266 706696
rect 674378 706344 674434 706353
rect 674378 706279 674434 706288
rect 674010 693152 674066 693161
rect 674010 693087 674066 693096
rect 673458 690160 673514 690169
rect 673458 690095 673514 690104
rect 673274 689072 673330 689081
rect 673274 689007 673330 689016
rect 673090 661600 673146 661609
rect 673090 661535 673146 661544
rect 673090 648680 673146 648689
rect 673090 648615 673146 648624
rect 672814 647864 672870 647873
rect 672814 647799 672870 647808
rect 672630 635488 672686 635497
rect 672630 635423 672686 635432
rect 672828 630674 672856 647799
rect 672828 630646 672948 630674
rect 672920 627914 672948 630646
rect 673104 627914 673132 648615
rect 673288 627914 673316 689007
rect 673472 636857 673500 690095
rect 673826 644600 673882 644609
rect 673826 644535 673882 644544
rect 673642 641744 673698 641753
rect 673642 641679 673698 641688
rect 673458 636848 673514 636857
rect 673458 636783 673514 636792
rect 672920 627886 673040 627914
rect 673104 627886 673224 627914
rect 673288 627886 673408 627914
rect 672630 621888 672686 621897
rect 672630 621823 672686 621832
rect 672644 621217 672672 621823
rect 672630 621208 672686 621217
rect 672630 621143 672686 621152
rect 673012 621042 673040 627886
rect 672632 621036 672684 621042
rect 672632 620978 672684 620984
rect 673000 621036 673052 621042
rect 673000 620978 673052 620984
rect 672446 619848 672502 619857
rect 672446 619783 672502 619792
rect 672264 618384 672316 618390
rect 672264 618326 672316 618332
rect 672644 618254 672672 620978
rect 672908 618384 672960 618390
rect 673196 618338 673224 627886
rect 673380 624034 673408 627886
rect 673368 624028 673420 624034
rect 673368 623970 673420 623976
rect 673368 623892 673420 623898
rect 673368 623834 673420 623840
rect 672908 618326 672960 618332
rect 672920 618254 672948 618326
rect 673104 618310 673224 618338
rect 672644 618226 672856 618254
rect 672920 618226 673040 618254
rect 672630 597408 672686 597417
rect 672630 597343 672686 597352
rect 672446 578640 672502 578649
rect 672446 578575 672502 578584
rect 671986 574152 672042 574161
rect 671986 574087 672042 574096
rect 671802 571160 671858 571169
rect 671802 571095 671858 571104
rect 671710 570344 671766 570353
rect 671710 570279 671766 570288
rect 671356 557506 671476 557534
rect 671540 557506 671660 557534
rect 671250 534848 671306 534857
rect 671250 534783 671306 534792
rect 671448 533497 671476 557506
rect 671434 533488 671490 533497
rect 671434 533423 671490 533432
rect 671632 533338 671660 557506
rect 671540 533310 671660 533338
rect 671540 532681 671568 533310
rect 671526 532672 671582 532681
rect 671526 532607 671582 532616
rect 671526 529408 671582 529417
rect 671526 529343 671582 529352
rect 671540 528601 671568 529343
rect 671526 528592 671582 528601
rect 671526 528527 671582 528536
rect 671066 525736 671122 525745
rect 671066 525671 671122 525680
rect 671724 500993 671752 570279
rect 671986 569528 672042 569537
rect 671986 569463 672042 569472
rect 671710 500984 671766 500993
rect 671710 500919 671766 500928
rect 670882 483984 670938 483993
rect 670882 483919 670938 483928
rect 670606 455832 670662 455841
rect 670606 455767 670662 455776
rect 670422 455424 670478 455433
rect 670422 455359 670478 455368
rect 672000 455274 672028 569463
rect 672262 559464 672318 559473
rect 672262 559399 672318 559408
rect 672276 485774 672304 559399
rect 672460 534585 672488 578575
rect 672446 534576 672502 534585
rect 672446 534511 672502 534520
rect 672644 534018 672672 597343
rect 672828 571985 672856 618226
rect 673012 579193 673040 618226
rect 673104 611354 673132 618310
rect 673380 618254 673408 623834
rect 673288 618226 673408 618254
rect 673288 616593 673316 618226
rect 673274 616584 673330 616593
rect 673274 616519 673330 616528
rect 673104 611326 673224 611354
rect 672998 579184 673054 579193
rect 672998 579119 673054 579128
rect 673196 576854 673224 611326
rect 673366 604344 673422 604353
rect 673366 604279 673422 604288
rect 673380 601694 673408 604279
rect 673104 576826 673224 576854
rect 673288 601666 673408 601694
rect 673104 573209 673132 576826
rect 673090 573200 673146 573209
rect 673090 573135 673146 573144
rect 672814 571976 672870 571985
rect 672814 571911 672870 571920
rect 673090 553480 673146 553489
rect 673090 553415 673146 553424
rect 672814 534304 672870 534313
rect 672814 534239 672870 534248
rect 672828 534074 672856 534239
rect 672828 534046 672948 534074
rect 672368 533990 672672 534018
rect 672368 532114 672396 533990
rect 672724 532160 672776 532166
rect 672368 532086 672580 532114
rect 672724 532102 672776 532108
rect 672552 532046 672580 532086
rect 672552 532018 672672 532046
rect 672446 531856 672502 531865
rect 672446 531791 672502 531800
rect 672460 488481 672488 531791
rect 672644 531434 672672 532018
rect 672552 531406 672672 531434
rect 672552 531314 672580 531406
rect 672552 531286 672672 531314
rect 672644 528193 672672 531286
rect 672736 528306 672764 532102
rect 672736 528278 672856 528306
rect 672630 528184 672686 528193
rect 672630 528119 672686 528128
rect 672828 524414 672856 528278
rect 672736 524386 672856 524414
rect 672736 489297 672764 524386
rect 672920 490929 672948 534046
rect 672906 490920 672962 490929
rect 672906 490855 672962 490864
rect 672906 489696 672962 489705
rect 672906 489631 672962 489640
rect 672722 489288 672778 489297
rect 672722 489223 672778 489232
rect 672446 488472 672502 488481
rect 672446 488407 672502 488416
rect 672446 488064 672502 488073
rect 672446 487999 672502 488008
rect 672184 485746 672304 485774
rect 672184 484809 672212 485746
rect 672170 484800 672226 484809
rect 672170 484735 672226 484744
rect 672000 455258 672120 455274
rect 672000 455252 672132 455258
rect 672000 455246 672080 455252
rect 672080 455194 672132 455200
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 671344 430636 671396 430642
rect 671344 430578 671396 430584
rect 670146 360904 670202 360913
rect 670146 360839 670202 360848
rect 670146 348528 670202 348537
rect 670146 348463 670202 348472
rect 669962 347304 670018 347313
rect 669962 347239 670018 347248
rect 668582 311944 668638 311953
rect 668582 311879 668638 311888
rect 669226 302288 669282 302297
rect 669226 302223 669282 302232
rect 667572 284368 667624 284374
rect 667572 284310 667624 284316
rect 667386 181384 667442 181393
rect 667386 181319 667442 181328
rect 667584 135969 667612 284310
rect 668768 237244 668820 237250
rect 668768 237186 668820 237192
rect 668124 235340 668176 235346
rect 668124 235282 668176 235288
rect 667940 234116 667992 234122
rect 667940 234058 667992 234064
rect 667952 229094 667980 234058
rect 668136 231690 668164 235282
rect 668400 234456 668452 234462
rect 668400 234398 668452 234404
rect 668044 231662 668164 231690
rect 668044 230466 668072 231662
rect 668216 231600 668268 231606
rect 668216 231542 668268 231548
rect 668228 230625 668256 231542
rect 668214 230616 668270 230625
rect 668214 230551 668270 230560
rect 668044 230438 668348 230466
rect 667952 229066 668072 229094
rect 667848 226092 667900 226098
rect 667848 226034 667900 226040
rect 667860 223145 667888 226034
rect 667846 223136 667902 223145
rect 667846 223071 667902 223080
rect 667846 220960 667902 220969
rect 667846 220895 667902 220904
rect 667860 176497 667888 220895
rect 668044 197441 668072 229066
rect 668030 197432 668086 197441
rect 668030 197367 668086 197376
rect 668124 194200 668176 194206
rect 668122 194168 668124 194177
rect 668176 194168 668178 194177
rect 668122 194103 668178 194112
rect 668032 192568 668084 192574
rect 668030 192536 668032 192545
rect 668084 192536 668086 192545
rect 668030 192471 668086 192480
rect 668122 192264 668178 192273
rect 668122 192199 668178 192208
rect 668136 187649 668164 192199
rect 668122 187640 668178 187649
rect 668122 187575 668178 187584
rect 668032 184408 668084 184414
rect 668030 184376 668032 184385
rect 668084 184376 668086 184385
rect 668030 184311 668086 184320
rect 668320 182753 668348 230438
rect 668412 229094 668440 234398
rect 668582 230480 668638 230489
rect 668582 230415 668638 230424
rect 668596 229265 668624 230415
rect 668582 229256 668638 229265
rect 668582 229191 668638 229200
rect 668412 229066 668532 229094
rect 668306 182744 668362 182753
rect 668306 182679 668362 182688
rect 667846 176488 667902 176497
rect 667846 176423 667902 176432
rect 667940 174888 667992 174894
rect 667940 174830 667992 174836
rect 667952 174593 667980 174830
rect 667938 174584 667994 174593
rect 667938 174519 667994 174528
rect 668032 164824 668084 164830
rect 668030 164792 668032 164801
rect 668084 164792 668086 164801
rect 668030 164727 668086 164736
rect 668504 148481 668532 229066
rect 668780 153377 668808 237186
rect 668952 230716 669004 230722
rect 668952 230658 669004 230664
rect 668964 230466 668992 230658
rect 668872 230438 668992 230466
rect 668872 224954 668900 230438
rect 669044 230376 669096 230382
rect 669044 230318 669096 230324
rect 669056 229094 669084 230318
rect 669056 229066 669176 229094
rect 668872 224926 669084 224954
rect 669056 222194 669084 224926
rect 668872 222166 669084 222194
rect 668872 211426 668900 222166
rect 669148 219434 669176 229066
rect 669056 219406 669176 219434
rect 669056 211857 669084 219406
rect 669240 212401 669268 302223
rect 669780 235544 669832 235550
rect 669780 235486 669832 235492
rect 669596 233368 669648 233374
rect 669596 233310 669648 233316
rect 669412 231600 669464 231606
rect 669410 231568 669412 231577
rect 669464 231568 669466 231577
rect 669410 231503 669466 231512
rect 669412 229764 669464 229770
rect 669412 229706 669464 229712
rect 669226 212392 669282 212401
rect 669226 212327 669282 212336
rect 669226 211984 669282 211993
rect 669226 211919 669282 211928
rect 669042 211848 669098 211857
rect 669042 211783 669098 211792
rect 668872 211398 669176 211426
rect 668950 211304 669006 211313
rect 668950 211239 669006 211248
rect 668964 200114 668992 211239
rect 669148 209774 669176 211398
rect 668872 200086 668992 200114
rect 669056 209746 669176 209774
rect 668872 190454 668900 200086
rect 669056 192574 669084 209746
rect 669044 192568 669096 192574
rect 669044 192510 669096 192516
rect 668872 190426 668992 190454
rect 668964 171134 668992 190426
rect 669240 190369 669268 211919
rect 669226 190360 669282 190369
rect 669226 190295 669282 190304
rect 669136 189304 669188 189310
rect 669134 189272 669136 189281
rect 669188 189272 669190 189281
rect 669134 189207 669190 189216
rect 669134 185600 669190 185609
rect 669134 185535 669190 185544
rect 669148 171134 669176 185535
rect 668872 171106 668992 171134
rect 669056 171106 669176 171134
rect 668872 163282 668900 171106
rect 669056 169810 669084 171106
rect 668964 169782 669084 169810
rect 668964 168178 668992 169782
rect 669134 169688 669190 169697
rect 669424 169674 669452 229706
rect 669608 184414 669636 233310
rect 669596 184408 669648 184414
rect 669596 184350 669648 184356
rect 669792 174894 669820 235486
rect 669780 174888 669832 174894
rect 669780 174830 669832 174836
rect 669190 169646 669452 169674
rect 669134 169623 669190 169632
rect 669778 169552 669834 169561
rect 669778 169487 669834 169496
rect 669594 168328 669650 168337
rect 669594 168263 669650 168272
rect 668964 168150 669084 168178
rect 669056 168065 669084 168150
rect 669042 168056 669098 168065
rect 669042 167991 669098 168000
rect 669136 166116 669188 166122
rect 669136 166058 669188 166064
rect 668872 163254 668992 163282
rect 668964 163169 668992 163254
rect 668950 163160 669006 163169
rect 668950 163095 669006 163104
rect 668766 153368 668822 153377
rect 668766 153303 668822 153312
rect 668676 150272 668728 150278
rect 668676 150214 668728 150220
rect 668688 150113 668716 150214
rect 668674 150104 668730 150113
rect 668674 150039 668730 150048
rect 668490 148472 668546 148481
rect 668490 148407 668546 148416
rect 668766 147792 668822 147801
rect 668766 147727 668822 147736
rect 667940 136468 667992 136474
rect 667940 136410 667992 136416
rect 667570 135960 667626 135969
rect 667570 135895 667626 135904
rect 667952 135425 667980 136410
rect 667938 135416 667994 135425
rect 667938 135351 667994 135360
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 667018 133104 667074 133113
rect 667018 133039 667074 133048
rect 668582 128208 668638 128217
rect 668582 128143 668638 128152
rect 668596 120737 668624 128143
rect 668780 125633 668808 147727
rect 669148 138689 669176 166058
rect 669134 138680 669190 138689
rect 669134 138615 669190 138624
rect 669608 128354 669636 168263
rect 669792 152697 669820 169487
rect 669778 152688 669834 152697
rect 669778 152623 669834 152632
rect 669976 136474 670004 347239
rect 670160 166122 670188 348463
rect 671356 269793 671384 430578
rect 672262 400480 672318 400489
rect 672262 400415 672318 400424
rect 672276 355881 672304 400415
rect 672460 400081 672488 487999
rect 672920 470594 672948 489631
rect 673104 482361 673132 553415
rect 673288 528737 673316 601666
rect 673458 598496 673514 598505
rect 673458 598431 673514 598440
rect 673274 528728 673330 528737
rect 673274 528663 673330 528672
rect 673472 526561 673500 598431
rect 673656 593201 673684 641679
rect 673642 593192 673698 593201
rect 673642 593127 673698 593136
rect 673840 591297 673868 644535
rect 674024 617409 674052 693087
rect 674194 692880 674250 692889
rect 674194 692815 674250 692824
rect 674208 683114 674236 692815
rect 674392 683114 674420 706279
rect 675114 701176 675170 701185
rect 675114 701111 675170 701120
rect 674838 699816 674894 699825
rect 674838 699751 674894 699760
rect 674562 697232 674618 697241
rect 674562 697167 674618 697176
rect 674576 689761 674604 697167
rect 674852 697049 674880 699751
rect 675128 698337 675156 701111
rect 675128 698309 675418 698337
rect 675128 697666 675418 697694
rect 675128 697241 675156 697666
rect 675114 697232 675170 697241
rect 675114 697167 675170 697176
rect 674852 697021 675418 697049
rect 674746 696960 674802 696969
rect 674802 696918 674972 696946
rect 674746 696895 674802 696904
rect 674944 695209 674972 696918
rect 674944 695181 675418 695209
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 675128 693994 675418 694022
rect 675128 692889 675156 693994
rect 675496 693161 675524 693328
rect 675482 693152 675538 693161
rect 675482 693087 675538 693096
rect 675114 692880 675170 692889
rect 675114 692815 675170 692824
rect 675128 690866 675418 690894
rect 675128 690441 675156 690866
rect 675114 690432 675170 690441
rect 675114 690367 675170 690376
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 674562 689752 674618 689761
rect 674562 689687 674618 689696
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 674760 689642 675340 689670
rect 675404 689656 675432 689710
rect 674760 689194 674788 689642
rect 674930 689344 674986 689353
rect 674930 689279 674986 689288
rect 674116 683086 674236 683114
rect 674300 683086 674420 683114
rect 674484 689166 674788 689194
rect 674116 650026 674144 683086
rect 674300 656894 674328 683086
rect 674300 656866 674420 656894
rect 674392 655514 674420 656866
rect 674300 655486 674420 655514
rect 674300 650321 674328 655486
rect 674286 650312 674342 650321
rect 674286 650247 674342 650256
rect 674116 649998 674420 650026
rect 674194 649632 674250 649641
rect 674194 649567 674250 649576
rect 674208 645153 674236 649567
rect 674194 645144 674250 645153
rect 674194 645079 674250 645088
rect 674392 640334 674420 649998
rect 674208 640306 674420 640334
rect 674208 635769 674236 640306
rect 674194 635760 674250 635769
rect 674194 635695 674250 635704
rect 674484 623257 674512 689166
rect 674746 688800 674802 688809
rect 674746 688735 674802 688744
rect 674760 687698 674788 688735
rect 674576 687670 674788 687698
rect 674576 683114 674604 687670
rect 674944 686678 674972 689279
rect 675114 689072 675170 689081
rect 675170 689030 675418 689058
rect 675114 689007 675170 689016
rect 675128 687806 675418 687834
rect 675128 687449 675156 687806
rect 675114 687440 675170 687449
rect 675114 687375 675170 687384
rect 674944 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675114 686216 675170 686225
rect 675114 686151 675170 686160
rect 675128 685998 675156 686151
rect 675128 685970 675418 685998
rect 674930 685944 674986 685953
rect 674930 685879 674986 685888
rect 674944 684162 674972 685879
rect 675114 685400 675170 685409
rect 675170 685358 675340 685386
rect 675114 685335 675170 685344
rect 675312 685250 675340 685358
rect 675404 685250 675432 685372
rect 675312 685222 675432 685250
rect 674944 684134 675418 684162
rect 674576 683086 674696 683114
rect 674470 623248 674526 623257
rect 674470 623183 674526 623192
rect 674668 623098 674696 683086
rect 683210 682408 683266 682417
rect 683210 682343 683266 682352
rect 676494 673160 676550 673169
rect 676494 673095 676550 673104
rect 676508 671129 676536 673095
rect 676494 671120 676550 671129
rect 676494 671055 676550 671064
rect 676494 669896 676550 669905
rect 676494 669831 676550 669840
rect 676508 669497 676536 669831
rect 676494 669488 676550 669497
rect 676494 669423 676550 669432
rect 674838 667448 674894 667457
rect 674838 667383 674894 667392
rect 674852 666641 674880 667383
rect 683224 667049 683252 682343
rect 683394 681048 683450 681057
rect 683394 680983 683450 680992
rect 683210 667040 683266 667049
rect 683210 666975 683266 666984
rect 674838 666632 674894 666641
rect 674838 666567 674894 666576
rect 683408 663377 683436 680983
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683394 663368 683450 663377
rect 683394 663303 683450 663312
rect 674838 661872 674894 661881
rect 674838 661807 674894 661816
rect 674852 661337 674880 661807
rect 674838 661328 674894 661337
rect 674838 661263 674894 661272
rect 675298 660240 675354 660249
rect 675298 660175 675354 660184
rect 675312 659705 675340 660175
rect 675298 659696 675354 659705
rect 675298 659631 675354 659640
rect 675206 654256 675262 654265
rect 675206 654191 675262 654200
rect 675220 652746 675248 654191
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675220 652718 675432 652746
rect 675404 652460 675432 652718
rect 675496 651545 675524 651848
rect 675482 651536 675538 651545
rect 675482 651471 675538 651480
rect 675404 649994 675432 650012
rect 674944 649966 675432 649994
rect 674944 629785 674972 649966
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675128 648774 675418 648802
rect 675128 648689 675156 648774
rect 675114 648680 675170 648689
rect 675114 648615 675170 648624
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675114 647320 675170 647329
rect 675114 647255 675170 647264
rect 675128 645674 675156 647255
rect 675128 645646 675418 645674
rect 675128 645102 675418 645130
rect 675128 644609 675156 645102
rect 675758 644736 675814 644745
rect 675758 644671 675814 644680
rect 675114 644600 675170 644609
rect 675114 644535 675170 644544
rect 675772 644475 675800 644671
rect 675114 643920 675170 643929
rect 675114 643855 675170 643864
rect 675128 641458 675156 643855
rect 675404 643521 675432 643824
rect 675390 643512 675446 643521
rect 675390 643447 675446 643456
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675404 640529 675432 640795
rect 675390 640520 675446 640529
rect 675390 640455 675446 640464
rect 675036 640138 675418 640166
rect 675036 631122 675064 640138
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675758 638072 675814 638081
rect 675758 638007 675814 638016
rect 675574 637800 675630 637809
rect 675574 637735 675630 637744
rect 675206 637664 675262 637673
rect 675206 637599 675262 637608
rect 675220 631394 675248 637599
rect 675588 633049 675616 637735
rect 675574 633040 675630 633049
rect 675574 632975 675630 632984
rect 675772 631417 675800 638007
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 675758 631408 675814 631417
rect 675220 631366 675340 631394
rect 675036 631094 675248 631122
rect 674930 629776 674986 629785
rect 674930 629711 674986 629720
rect 674300 623070 674696 623098
rect 674300 619449 674328 623070
rect 674470 622160 674526 622169
rect 674470 622095 674526 622104
rect 674484 620945 674512 622095
rect 674470 620936 674526 620945
rect 674470 620871 674526 620880
rect 674286 619440 674342 619449
rect 674286 619375 674342 619384
rect 674010 617400 674066 617409
rect 674010 617335 674066 617344
rect 674838 608832 674894 608841
rect 674838 608767 674894 608776
rect 674852 607209 674880 608767
rect 675022 608560 675078 608569
rect 675022 608495 675078 608504
rect 675036 607753 675064 608495
rect 675022 607744 675078 607753
rect 675022 607679 675078 607688
rect 674838 607200 674894 607209
rect 674838 607135 674894 607144
rect 674654 604616 674710 604625
rect 674654 604551 674710 604560
rect 674010 603528 674066 603537
rect 674010 603463 674066 603472
rect 673826 591288 673882 591297
rect 673826 591223 673882 591232
rect 673826 580816 673882 580825
rect 673826 580751 673882 580760
rect 673840 579737 673868 580751
rect 673826 579728 673882 579737
rect 673826 579663 673882 579672
rect 673826 558376 673882 558385
rect 673826 558311 673882 558320
rect 673642 548448 673698 548457
rect 673642 548383 673698 548392
rect 673458 526552 673514 526561
rect 673458 526487 673514 526496
rect 673656 485625 673684 548383
rect 673642 485616 673698 485625
rect 673642 485551 673698 485560
rect 673840 484401 673868 558311
rect 674024 547097 674052 603463
rect 674286 600128 674342 600137
rect 674286 600063 674342 600072
rect 674010 547088 674066 547097
rect 674010 547023 674066 547032
rect 674300 545737 674328 600063
rect 674470 599040 674526 599049
rect 674470 598975 674526 598984
rect 674286 545728 674342 545737
rect 674286 545663 674342 545672
rect 674194 533216 674250 533225
rect 674194 533151 674250 533160
rect 674010 532944 674066 532953
rect 674010 532879 674066 532888
rect 674024 532166 674052 532879
rect 674012 532160 674064 532166
rect 674012 532102 674064 532108
rect 674208 490113 674236 533151
rect 674484 527785 674512 598975
rect 674668 530369 674696 604551
rect 674838 602304 674894 602313
rect 674838 602239 674894 602248
rect 674852 598890 674880 602239
rect 675220 600930 675248 631094
rect 675312 602426 675340 631366
rect 675758 631343 675814 631352
rect 675850 627872 675906 627881
rect 675850 627807 675906 627816
rect 675864 626618 675892 627807
rect 675852 626612 675904 626618
rect 675852 626554 675904 626560
rect 676496 626612 676548 626618
rect 676496 626554 676548 626560
rect 676508 625705 676536 626554
rect 676494 625696 676550 625705
rect 676494 625631 676550 625640
rect 683118 623248 683174 623257
rect 683118 623183 683174 623192
rect 683132 617953 683160 623183
rect 683118 617944 683174 617953
rect 683118 617879 683174 617888
rect 683408 617137 683436 636783
rect 683578 635760 683634 635769
rect 683578 635695 683634 635704
rect 683592 618769 683620 635695
rect 683762 635488 683818 635497
rect 683762 635423 683818 635432
rect 683776 622849 683804 635423
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683762 622840 683818 622849
rect 683762 622775 683818 622784
rect 683578 618760 683634 618769
rect 683578 618695 683634 618704
rect 683394 617128 683450 617137
rect 683394 617063 683450 617072
rect 675496 608025 675524 608124
rect 675482 608016 675538 608025
rect 675482 607951 675538 607960
rect 675482 607744 675538 607753
rect 675482 607679 675538 607688
rect 675496 607479 675524 607679
rect 675482 607200 675538 607209
rect 675482 607135 675538 607144
rect 675496 606832 675524 607135
rect 675496 604625 675524 604996
rect 675482 604616 675538 604625
rect 675482 604551 675538 604560
rect 675496 604353 675524 604452
rect 675482 604344 675538 604353
rect 675482 604279 675538 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675496 602993 675524 603160
rect 675482 602984 675538 602993
rect 675482 602919 675538 602928
rect 675312 602398 675432 602426
rect 675404 602313 675432 602398
rect 675390 602304 675446 602313
rect 675390 602239 675446 602248
rect 674760 598862 674880 598890
rect 674944 600902 675248 600930
rect 674760 596442 674788 598862
rect 674944 596737 674972 600902
rect 675312 600766 675432 600794
rect 675114 600672 675170 600681
rect 675312 600658 675340 600766
rect 675170 600630 675340 600658
rect 675404 600644 675432 600766
rect 675114 600607 675170 600616
rect 675312 600222 675432 600250
rect 675114 600128 675170 600137
rect 675312 600114 675340 600222
rect 675170 600086 675340 600114
rect 675404 600100 675432 600222
rect 675114 600063 675170 600072
rect 675114 599584 675170 599593
rect 675114 599519 675170 599528
rect 674930 596728 674986 596737
rect 674930 596663 674986 596672
rect 675128 596442 675156 599519
rect 675312 599474 675418 599502
rect 675312 599049 675340 599474
rect 675298 599040 675354 599049
rect 675298 598975 675354 598984
rect 675496 598505 675524 598808
rect 675482 598496 675538 598505
rect 675482 598431 675538 598440
rect 675404 597417 675432 597652
rect 675390 597408 675446 597417
rect 675390 597343 675446 597352
rect 674760 596414 674972 596442
rect 675128 596414 675418 596442
rect 674944 594425 674972 596414
rect 675128 595802 675340 595830
rect 674930 594416 674986 594425
rect 674930 594351 674986 594360
rect 675128 594266 675156 595802
rect 675312 595762 675340 595802
rect 675404 595762 675432 595816
rect 675312 595734 675432 595762
rect 675312 595122 675418 595150
rect 675312 594833 675340 595122
rect 675298 594824 675354 594833
rect 675298 594759 675354 594768
rect 675128 594238 675248 594266
rect 675022 593872 675078 593881
rect 675022 593807 675078 593816
rect 674838 580544 674894 580553
rect 674838 580479 674894 580488
rect 674852 579873 674880 580479
rect 674838 579864 674894 579873
rect 674838 579799 674894 579808
rect 674838 579456 674894 579465
rect 674838 579391 674894 579400
rect 674852 578921 674880 579391
rect 674838 578912 674894 578921
rect 674838 578847 674894 578856
rect 675036 576854 675064 593807
rect 675220 589274 675248 594238
rect 675404 593609 675432 593980
rect 675390 593600 675446 593609
rect 675390 593535 675446 593544
rect 675850 592920 675906 592929
rect 675850 592855 675906 592864
rect 683486 592920 683542 592929
rect 683486 592855 683542 592864
rect 674944 576826 675064 576854
rect 675128 589246 675248 589274
rect 674944 575385 674972 576826
rect 674930 575376 674986 575385
rect 674930 575311 674986 575320
rect 674838 559736 674894 559745
rect 674838 559671 674894 559680
rect 674852 557682 674880 559671
rect 674760 557654 674880 557682
rect 674760 550634 674788 557654
rect 674930 557560 674986 557569
rect 674930 557495 674986 557504
rect 674944 555801 674972 557495
rect 674930 555792 674986 555801
rect 674930 555727 674986 555736
rect 675128 555642 675156 589246
rect 675482 578368 675538 578377
rect 675482 578303 675538 578312
rect 675298 577688 675354 577697
rect 675298 577623 675354 577632
rect 675312 576881 675340 577623
rect 675496 577017 675524 578303
rect 675482 577008 675538 577017
rect 675482 576943 675538 576952
rect 675298 576872 675354 576881
rect 675298 576807 675354 576816
rect 675864 576609 675892 592855
rect 683302 592648 683358 592657
rect 683302 592583 683358 592592
rect 676034 592376 676090 592385
rect 676034 592311 676090 592320
rect 676048 591394 676076 592311
rect 676036 591388 676088 591394
rect 676036 591330 676088 591336
rect 682384 591388 682436 591394
rect 682384 591330 682436 591336
rect 681002 590608 681058 590617
rect 681002 590543 681058 590552
rect 675850 576600 675906 576609
rect 675850 576535 675906 576544
rect 681016 576065 681044 590543
rect 681002 576056 681058 576065
rect 681002 575991 681058 576000
rect 682396 570761 682424 591330
rect 683118 591288 683174 591297
rect 683118 591223 683174 591232
rect 683132 571985 683160 591223
rect 683316 574025 683344 592583
rect 683302 574016 683358 574025
rect 683302 573951 683358 573960
rect 683500 573209 683528 592855
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683486 573200 683542 573209
rect 683486 573135 683542 573144
rect 683118 571976 683174 571985
rect 683118 571911 683174 571920
rect 682382 570752 682438 570761
rect 682382 570687 682438 570696
rect 675298 564496 675354 564505
rect 675298 564431 675354 564440
rect 675312 562306 675340 564431
rect 675496 562737 675524 562904
rect 675482 562728 675538 562737
rect 675482 562663 675538 562672
rect 675312 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675312 559830 675432 559858
rect 675312 559745 675340 559830
rect 675404 559776 675432 559830
rect 675298 559736 675354 559745
rect 675298 559671 675354 559680
rect 675390 559464 675446 559473
rect 675390 559399 675446 559408
rect 675404 559232 675432 559399
rect 675404 558385 675432 558620
rect 675390 558376 675446 558385
rect 675390 558311 675446 558320
rect 675772 557705 675800 557940
rect 675758 557696 675814 557705
rect 675758 557631 675814 557640
rect 675482 555792 675538 555801
rect 675482 555727 675538 555736
rect 674852 555614 675156 555642
rect 674852 551970 674880 555614
rect 675496 555492 675524 555727
rect 675404 554713 675432 554919
rect 675390 554704 675446 554713
rect 675390 554639 675446 554648
rect 675772 554033 675800 554268
rect 675758 554024 675814 554033
rect 675758 553959 675814 553968
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 674852 551942 675064 551970
rect 674760 550606 674880 550634
rect 674852 550202 674880 550606
rect 675036 550497 675064 551942
rect 675390 551576 675446 551585
rect 675390 551511 675446 551520
rect 675404 551239 675432 551511
rect 675022 550488 675078 550497
rect 675022 550423 675078 550432
rect 675772 550225 675800 550596
rect 675758 550216 675814 550225
rect 674852 550174 675248 550202
rect 675220 545850 675248 550174
rect 675758 550151 675814 550160
rect 675312 549937 675418 549965
rect 675312 545986 675340 549937
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675944 547664 675996 547670
rect 675942 547632 675944 547641
rect 678244 547664 678296 547670
rect 675996 547632 675998 547641
rect 675942 547567 675998 547576
rect 677414 547632 677470 547641
rect 678244 547606 678296 547612
rect 677414 547567 677470 547576
rect 675312 545958 675524 545986
rect 675220 545822 675340 545850
rect 675312 545306 675340 545822
rect 675128 545278 675340 545306
rect 674838 544504 674894 544513
rect 674838 544439 674894 544448
rect 674852 544218 674880 544439
rect 674852 544190 675064 544218
rect 674838 543960 674894 543969
rect 674838 543895 674894 543904
rect 674852 539594 674880 543895
rect 674852 539566 674972 539594
rect 674654 530360 674710 530369
rect 674654 530295 674710 530304
rect 674470 527776 674526 527785
rect 674470 527711 674526 527720
rect 674194 490104 674250 490113
rect 674194 490039 674250 490048
rect 673826 484392 673882 484401
rect 673826 484327 673882 484336
rect 674944 483041 674972 539566
rect 675036 505094 675064 544190
rect 675128 540974 675156 545278
rect 675298 544912 675354 544921
rect 675298 544847 675354 544856
rect 675128 540946 675248 540974
rect 675220 505094 675248 540946
rect 675312 524414 675340 544847
rect 675496 543969 675524 545958
rect 675482 543960 675538 543969
rect 675482 543895 675538 543904
rect 676034 538792 676090 538801
rect 676034 538727 676090 538736
rect 676048 535741 676076 538727
rect 676034 535732 676090 535741
rect 676034 535667 676090 535676
rect 675758 534576 675814 534585
rect 675758 534511 675814 534520
rect 675772 534109 675800 534511
rect 675758 534100 675814 534109
rect 675758 534035 675814 534044
rect 675758 533692 675814 533701
rect 675758 533627 675814 533636
rect 675772 533225 675800 533627
rect 675758 533216 675814 533225
rect 675758 533151 675814 533160
rect 676862 525736 676918 525745
rect 676862 525671 676918 525680
rect 675312 524386 675892 524414
rect 675482 513768 675538 513777
rect 675482 513703 675538 513712
rect 675496 505094 675524 513703
rect 675036 505066 675156 505094
rect 675220 505066 675340 505094
rect 675496 505066 675616 505094
rect 675128 502625 675156 505066
rect 675114 502616 675170 502625
rect 675114 502551 675170 502560
rect 675312 486441 675340 505066
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 675588 485774 675616 505066
rect 675864 503674 675892 524386
rect 676036 518832 676088 518838
rect 676036 518774 676088 518780
rect 676048 513777 676076 518774
rect 676034 513768 676090 513777
rect 676034 513703 676090 513712
rect 675852 503668 675904 503674
rect 675852 503610 675904 503616
rect 675850 502616 675906 502625
rect 675850 502551 675906 502560
rect 675864 499594 675892 502551
rect 676402 500984 676458 500993
rect 676402 500919 676458 500928
rect 675852 499588 675904 499594
rect 675852 499530 675904 499536
rect 676416 495434 676444 500919
rect 676416 495406 676720 495434
rect 675850 494048 675906 494057
rect 675850 493983 675906 493992
rect 675864 492726 675892 493983
rect 675852 492720 675904 492726
rect 675852 492662 675904 492668
rect 676034 490512 676090 490521
rect 676034 490447 676090 490456
rect 675496 485746 675616 485774
rect 674930 483032 674986 483041
rect 674930 482967 674986 482976
rect 673090 482352 673146 482361
rect 673090 482287 673146 482296
rect 673274 474872 673330 474881
rect 673274 474807 673330 474816
rect 673288 470594 673316 474807
rect 672644 470566 672948 470594
rect 673196 470566 673316 470594
rect 672644 401985 672672 470566
rect 673196 456822 673224 470566
rect 673184 456816 673236 456822
rect 673184 456758 673236 456764
rect 674838 456376 674894 456385
rect 674838 456311 674894 456320
rect 673458 456104 673514 456113
rect 673458 456039 673514 456048
rect 673826 456104 673882 456113
rect 673826 456039 673828 456048
rect 673472 455598 673500 456039
rect 673880 456039 673882 456048
rect 673828 456010 673880 456016
rect 673736 455864 673788 455870
rect 673734 455832 673736 455841
rect 673788 455832 673790 455841
rect 673734 455767 673790 455776
rect 673460 455592 673512 455598
rect 673460 455534 673512 455540
rect 673504 455424 673560 455433
rect 673504 455359 673506 455368
rect 673558 455359 673560 455368
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673386 455152 673388 455161
rect 673440 455152 673442 455161
rect 673386 455087 673442 455096
rect 673550 455152 673606 455161
rect 673550 455087 673606 455096
rect 673564 455002 673592 455087
rect 673176 454986 673592 455002
rect 673164 454980 673592 454986
rect 673216 454974 673592 454980
rect 673164 454922 673216 454928
rect 673044 454880 673100 454889
rect 673044 454815 673046 454824
rect 673098 454815 673100 454824
rect 673046 454786 673098 454792
rect 672814 454472 672870 454481
rect 672814 454407 672816 454416
rect 672868 454407 672870 454416
rect 672816 454378 672868 454384
rect 672954 454232 673006 454238
rect 672952 454200 672954 454209
rect 673006 454200 673008 454209
rect 672952 454135 673008 454144
rect 674852 453937 674880 456311
rect 675496 454889 675524 485746
rect 675850 483032 675906 483041
rect 675850 482967 675906 482976
rect 675666 480720 675722 480729
rect 675666 480655 675722 480664
rect 675482 454880 675538 454889
rect 675482 454815 675538 454824
rect 675680 454481 675708 480655
rect 675864 480418 675892 482967
rect 675852 480412 675904 480418
rect 675852 480354 675904 480360
rect 675852 476128 675904 476134
rect 675852 476070 675904 476076
rect 675864 456385 675892 476070
rect 676048 466454 676076 490447
rect 676048 466426 676168 466454
rect 676140 457502 676168 466426
rect 676128 457496 676180 457502
rect 676128 457438 676180 457444
rect 676312 457496 676364 457502
rect 676312 457438 676364 457444
rect 676324 457314 676352 457438
rect 675956 457286 676352 457314
rect 675956 456794 675984 457286
rect 676128 457224 676180 457230
rect 676128 457166 676180 457172
rect 675956 456766 676076 456794
rect 675850 456376 675906 456385
rect 675850 456311 675906 456320
rect 675852 456136 675904 456142
rect 675850 456104 675852 456113
rect 675904 456104 675906 456113
rect 675850 456039 675906 456048
rect 675666 454472 675722 454481
rect 675666 454407 675722 454416
rect 676048 454322 676076 456766
rect 675956 454294 676076 454322
rect 675956 454209 675984 454294
rect 675942 454200 675998 454209
rect 675942 454135 675998 454144
rect 674838 453928 674894 453937
rect 674838 453863 674894 453872
rect 676140 453801 676168 457166
rect 676692 455161 676720 495406
rect 676876 457502 676904 525671
rect 677428 483177 677456 547567
rect 678256 531457 678284 547606
rect 683394 547088 683450 547097
rect 683394 547023 683450 547032
rect 683210 545728 683266 545737
rect 683210 545663 683266 545672
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 683224 526969 683252 545663
rect 683408 528601 683436 547023
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683578 533896 683634 533905
rect 683578 533831 683634 533840
rect 683394 528592 683450 528601
rect 683394 528527 683450 528536
rect 683592 527377 683620 533831
rect 683578 527368 683634 527377
rect 683578 527303 683634 527312
rect 683210 526960 683266 526969
rect 683210 526895 683266 526904
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 677888 518838 677916 524447
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683578 503704 683634 503713
rect 681004 503668 681056 503674
rect 683578 503639 683634 503648
rect 681004 503610 681056 503616
rect 679624 499588 679676 499594
rect 679624 499530 679676 499536
rect 679636 487665 679664 499530
rect 679622 487656 679678 487665
rect 679622 487591 679678 487600
rect 681016 486849 681044 503610
rect 683394 503432 683450 503441
rect 683394 503367 683450 503376
rect 683120 492720 683172 492726
rect 683120 492662 683172 492668
rect 683132 491337 683160 492662
rect 683118 491328 683174 491337
rect 683118 491263 683174 491272
rect 681002 486840 681058 486849
rect 681002 486775 681058 486784
rect 683408 483585 683436 503367
rect 683592 487257 683620 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 487248 683634 487257
rect 683578 487183 683634 487192
rect 683394 483576 683450 483585
rect 683394 483511 683450 483520
rect 677414 483168 677470 483177
rect 677414 483103 677470 483112
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 680372 476134 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 680360 476128 680412 476134
rect 680360 476070 680412 476076
rect 677138 475416 677194 475425
rect 677138 475351 677194 475360
rect 676864 457496 676916 457502
rect 676864 457438 676916 457444
rect 677152 456142 677180 475351
rect 677140 456136 677192 456142
rect 677140 456078 677192 456084
rect 676678 455152 676734 455161
rect 676678 455087 676734 455096
rect 676126 453792 676182 453801
rect 676126 453727 676182 453736
rect 676034 410544 676090 410553
rect 676034 410479 676090 410488
rect 675850 405648 675906 405657
rect 675850 405583 675906 405592
rect 675864 403481 675892 405583
rect 675850 403472 675906 403481
rect 675850 403407 675906 403416
rect 676048 402665 676076 410479
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 683132 403345 683160 406263
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 676034 402656 676090 402665
rect 676034 402591 676090 402600
rect 674838 402248 674894 402257
rect 674838 402183 674894 402192
rect 672630 401976 672686 401985
rect 672630 401911 672686 401920
rect 674852 401713 674880 402183
rect 672998 401704 673054 401713
rect 672998 401639 673054 401648
rect 674838 401704 674894 401713
rect 674838 401639 674894 401648
rect 672446 400072 672502 400081
rect 672446 400007 672502 400016
rect 673012 394694 673040 401639
rect 673182 401296 673238 401305
rect 673182 401231 673238 401240
rect 673012 394666 673132 394694
rect 672722 392592 672778 392601
rect 672722 392527 672778 392536
rect 672262 355872 672318 355881
rect 672262 355807 672318 355816
rect 672538 354648 672594 354657
rect 672538 354583 672594 354592
rect 672170 349752 672226 349761
rect 672170 349687 672226 349696
rect 671986 348936 672042 348945
rect 671986 348871 672042 348880
rect 672000 332353 672028 348871
rect 672184 333985 672212 349687
rect 672354 347712 672410 347721
rect 672354 347647 672410 347656
rect 672170 333976 672226 333985
rect 672170 333911 672226 333920
rect 671986 332344 672042 332353
rect 671986 332279 672042 332288
rect 672368 327593 672396 347647
rect 672354 327584 672410 327593
rect 672354 327519 672410 327528
rect 672552 310049 672580 354583
rect 672538 310040 672594 310049
rect 672538 309975 672594 309984
rect 672446 301472 672502 301481
rect 672446 301407 672502 301416
rect 671342 269784 671398 269793
rect 671342 269719 671398 269728
rect 671986 264072 672042 264081
rect 671986 264007 672042 264016
rect 671710 262168 671766 262177
rect 671710 262103 671766 262112
rect 671526 259720 671582 259729
rect 671526 259655 671582 259664
rect 671342 258904 671398 258913
rect 671342 258839 671398 258848
rect 670606 257680 670662 257689
rect 670606 257615 670662 257624
rect 670620 235929 670648 257615
rect 671356 241505 671384 258839
rect 671540 245857 671568 259655
rect 671526 245848 671582 245857
rect 671526 245783 671582 245792
rect 671724 245585 671752 262103
rect 671710 245576 671766 245585
rect 671710 245511 671766 245520
rect 672000 244274 672028 264007
rect 672262 257272 672318 257281
rect 672262 257207 672318 257216
rect 672276 244274 672304 257207
rect 671908 244246 672028 244274
rect 672092 244246 672304 244274
rect 671342 241496 671398 241505
rect 671342 241431 671398 241440
rect 671908 238241 671936 244246
rect 671894 238232 671950 238241
rect 671894 238167 671950 238176
rect 671896 237856 671948 237862
rect 671896 237798 671948 237804
rect 671528 237040 671580 237046
rect 671528 236982 671580 236988
rect 670606 235920 670662 235929
rect 670606 235855 670662 235864
rect 671344 234592 671396 234598
rect 671344 234534 671396 234540
rect 670792 233912 670844 233918
rect 670792 233854 670844 233860
rect 670608 233504 670660 233510
rect 670608 233446 670660 233452
rect 670620 232914 670648 233446
rect 670804 233186 670832 233854
rect 671356 233374 671384 234534
rect 671344 233368 671396 233374
rect 671344 233310 671396 233316
rect 671344 233232 671396 233238
rect 670804 233158 670924 233186
rect 671344 233174 671396 233180
rect 670620 232886 670740 232914
rect 670514 232656 670570 232665
rect 670514 232591 670570 232600
rect 670330 232112 670386 232121
rect 670330 232047 670386 232056
rect 670148 166116 670200 166122
rect 670148 166058 670200 166064
rect 670146 165608 670202 165617
rect 670146 165543 670202 165552
rect 669964 136468 670016 136474
rect 669964 136410 670016 136416
rect 669424 128326 669636 128354
rect 668766 125624 668822 125633
rect 668766 125559 668822 125568
rect 669424 125474 669452 128326
rect 669240 125446 669452 125474
rect 668582 120728 668638 120737
rect 668582 120663 668638 120672
rect 668674 120184 668730 120193
rect 668674 120119 668730 120128
rect 668032 118380 668084 118386
rect 668032 118322 668084 118328
rect 668044 117473 668072 118322
rect 668030 117464 668086 117473
rect 668030 117399 668086 117408
rect 591304 114436 591356 114442
rect 591304 114378 591356 114384
rect 668688 114209 668716 120119
rect 669240 119105 669268 125446
rect 669962 122768 670018 122777
rect 669962 122703 670018 122712
rect 669226 119096 669282 119105
rect 669226 119031 669282 119040
rect 668674 114200 668730 114209
rect 668124 114164 668176 114170
rect 669976 114170 670004 122703
rect 670160 118386 670188 165543
rect 670344 164830 670372 232047
rect 670528 229770 670556 232591
rect 670516 229764 670568 229770
rect 670516 229706 670568 229712
rect 670516 227656 670568 227662
rect 670516 227598 670568 227604
rect 670528 227225 670556 227598
rect 670514 227216 670570 227225
rect 670514 227151 670570 227160
rect 670516 227044 670568 227050
rect 670516 226986 670568 226992
rect 670528 226817 670556 226986
rect 670514 226808 670570 226817
rect 670514 226743 670570 226752
rect 670514 226128 670570 226137
rect 670514 226063 670570 226072
rect 670528 225282 670556 226063
rect 670516 225276 670568 225282
rect 670516 225218 670568 225224
rect 670712 224954 670740 232886
rect 670712 224926 670832 224954
rect 670516 224664 670568 224670
rect 670436 224612 670516 224618
rect 670436 224606 670568 224612
rect 670436 224590 670556 224606
rect 670436 223802 670464 224590
rect 670608 224460 670660 224466
rect 670608 224402 670660 224408
rect 670620 223961 670648 224402
rect 670606 223952 670662 223961
rect 670606 223887 670662 223896
rect 670436 223774 670556 223802
rect 670528 223689 670556 223774
rect 670514 223680 670570 223689
rect 670514 223615 670570 223624
rect 670606 218920 670662 218929
rect 670606 218855 670662 218864
rect 670620 218385 670648 218855
rect 670606 218376 670662 218385
rect 670606 218311 670662 218320
rect 670606 215792 670662 215801
rect 670606 215727 670662 215736
rect 670620 201385 670648 215727
rect 670606 201376 670662 201385
rect 670606 201311 670662 201320
rect 670804 199073 670832 224926
rect 670896 222194 670924 233158
rect 671160 233096 671212 233102
rect 671160 233038 671212 233044
rect 671172 231854 671200 233038
rect 671080 231826 671200 231854
rect 670896 222166 671016 222194
rect 670790 199064 670846 199073
rect 670790 198999 670846 199008
rect 670988 194290 671016 222166
rect 671080 215294 671108 231826
rect 671356 228426 671384 233174
rect 671172 228398 671384 228426
rect 671172 225298 671200 228398
rect 671344 228268 671396 228274
rect 671344 228210 671396 228216
rect 671356 225865 671384 228210
rect 671342 225856 671398 225865
rect 671342 225791 671398 225800
rect 671344 225684 671396 225690
rect 671344 225626 671396 225632
rect 671356 225457 671384 225626
rect 671342 225448 671398 225457
rect 671342 225383 671398 225392
rect 671172 225270 671476 225298
rect 671252 225072 671304 225078
rect 671250 225040 671252 225049
rect 671304 225040 671306 225049
rect 671250 224975 671306 224984
rect 671250 224768 671306 224777
rect 671250 224703 671252 224712
rect 671304 224703 671306 224712
rect 671252 224674 671304 224680
rect 671250 220688 671306 220697
rect 671250 220623 671306 220632
rect 671264 219881 671292 220623
rect 671250 219872 671306 219881
rect 671250 219807 671306 219816
rect 671250 219600 671306 219609
rect 671250 219535 671306 219544
rect 671264 218929 671292 219535
rect 671250 218920 671306 218929
rect 671250 218855 671306 218864
rect 671448 215294 671476 225270
rect 671080 215266 671200 215294
rect 670804 194262 671016 194290
rect 670804 194206 670832 194262
rect 670792 194200 670844 194206
rect 670792 194142 670844 194148
rect 671172 190454 671200 215266
rect 670804 190426 671200 190454
rect 671356 215266 671476 215294
rect 670804 189310 670832 190426
rect 670792 189304 670844 189310
rect 670792 189246 670844 189252
rect 670606 172000 670662 172009
rect 670606 171935 670662 171944
rect 670332 164824 670384 164830
rect 670332 164766 670384 164772
rect 670620 149025 670648 171935
rect 671356 157334 671384 215266
rect 671540 158273 671568 236982
rect 671712 236088 671764 236094
rect 671712 236030 671764 236036
rect 671724 172961 671752 236030
rect 671908 234462 671936 237798
rect 671896 234456 671948 234462
rect 671896 234398 671948 234404
rect 671896 228064 671948 228070
rect 671896 228006 671948 228012
rect 671908 227089 671936 228006
rect 671894 227080 671950 227089
rect 671894 227015 671950 227024
rect 671896 226840 671948 226846
rect 671896 226782 671948 226788
rect 671908 226681 671936 226782
rect 671894 226672 671950 226681
rect 672092 226658 672120 244246
rect 672264 237652 672316 237658
rect 672264 237594 672316 237600
rect 672276 233209 672304 237594
rect 672460 236314 672488 301407
rect 672368 236286 672488 236314
rect 672368 234614 672396 236286
rect 672540 236224 672592 236230
rect 672540 236166 672592 236172
rect 672368 234586 672488 234614
rect 672262 233200 672318 233209
rect 672262 233135 672318 233144
rect 672264 232348 672316 232354
rect 672264 232290 672316 232296
rect 672276 232014 672304 232290
rect 672264 232008 672316 232014
rect 672264 231950 672316 231956
rect 672262 228848 672318 228857
rect 672262 228783 672318 228792
rect 672276 228478 672304 228783
rect 672264 228472 672316 228478
rect 672264 228414 672316 228420
rect 672264 227384 672316 227390
rect 672264 227326 672316 227332
rect 672276 226817 672304 227326
rect 672460 227202 672488 234586
rect 672368 227174 672488 227202
rect 672552 227202 672580 236166
rect 672736 235770 672764 392527
rect 673104 389858 673132 394666
rect 672828 389830 673132 389858
rect 672828 376754 672856 389830
rect 672998 385248 673054 385257
rect 672998 385183 673054 385192
rect 673012 385034 673040 385183
rect 673012 385006 673132 385034
rect 673104 379409 673132 385006
rect 673196 379514 673224 401231
rect 674654 399800 674710 399809
rect 674654 399735 674710 399744
rect 674286 397352 674342 397361
rect 674286 397287 674342 397296
rect 673366 396672 673422 396681
rect 673366 396607 673422 396616
rect 673380 382265 673408 396607
rect 673918 396128 673974 396137
rect 673918 396063 673974 396072
rect 673734 395720 673790 395729
rect 673734 395655 673790 395664
rect 673550 394360 673606 394369
rect 673550 394295 673606 394304
rect 673564 385257 673592 394295
rect 673550 385248 673606 385257
rect 673550 385183 673606 385192
rect 673366 382256 673422 382265
rect 673366 382191 673422 382200
rect 673196 379486 673408 379514
rect 673090 379400 673146 379409
rect 673090 379335 673146 379344
rect 672828 376726 672948 376754
rect 672920 373994 672948 376726
rect 673380 373994 673408 379486
rect 673748 375465 673776 395655
rect 673932 381449 673960 396063
rect 674102 393680 674158 393689
rect 674102 393615 674158 393624
rect 673918 381440 673974 381449
rect 673918 381375 673974 381384
rect 673734 375456 673790 375465
rect 673734 375391 673790 375400
rect 672920 373966 673040 373994
rect 673012 357513 673040 373966
rect 673196 373966 673408 373994
rect 672998 357504 673054 357513
rect 672998 357439 673054 357448
rect 673196 356697 673224 373966
rect 673366 357096 673422 357105
rect 673366 357031 673422 357040
rect 673182 356688 673238 356697
rect 673182 356623 673238 356632
rect 673090 355464 673146 355473
rect 673090 355399 673146 355408
rect 672906 351384 672962 351393
rect 672906 351319 672962 351328
rect 672920 338065 672948 351319
rect 672906 338056 672962 338065
rect 672906 337991 672962 338000
rect 672906 312080 672962 312089
rect 672906 312015 672962 312024
rect 672920 267345 672948 312015
rect 673104 311894 673132 355399
rect 673380 331214 673408 357031
rect 673918 356280 673974 356289
rect 673918 356215 673974 356224
rect 673550 352608 673606 352617
rect 673550 352543 673606 352552
rect 673564 336705 673592 352543
rect 673734 350568 673790 350577
rect 673734 350503 673790 350512
rect 673550 336696 673606 336705
rect 673550 336631 673606 336640
rect 673288 331186 673408 331214
rect 673288 312497 673316 331186
rect 673748 331129 673776 350503
rect 673734 331120 673790 331129
rect 673734 331055 673790 331064
rect 673274 312488 673330 312497
rect 673274 312423 673330 312432
rect 673104 311866 673316 311894
rect 673090 311264 673146 311273
rect 673090 311199 673146 311208
rect 672906 267336 672962 267345
rect 672906 267271 672962 267280
rect 673104 266529 673132 311199
rect 673288 310865 673316 311866
rect 673932 311681 673960 356215
rect 673918 311672 673974 311681
rect 673918 311607 673974 311616
rect 673274 310856 673330 310865
rect 673274 310791 673330 310800
rect 673826 310448 673882 310457
rect 673826 310383 673882 310392
rect 673840 309134 673868 310383
rect 674116 309134 674144 393615
rect 674300 378049 674328 397287
rect 674470 394088 674526 394097
rect 674470 394023 674526 394032
rect 674286 378040 674342 378049
rect 674286 377975 674342 377984
rect 674484 376689 674512 394023
rect 674470 376680 674526 376689
rect 674470 376615 674526 376624
rect 674668 355065 674696 399735
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675298 379400 675354 379409
rect 675298 379335 675354 379344
rect 675312 377618 675340 379335
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675114 376680 675170 376689
rect 675114 376615 675170 376624
rect 675128 376462 675156 376615
rect 675128 376434 675340 376462
rect 675312 376394 675340 376434
rect 675404 376394 675432 376448
rect 675312 376366 675432 376394
rect 675114 375456 675170 375465
rect 675114 375391 675170 375400
rect 675128 375238 675156 375391
rect 675128 375210 675418 375238
rect 675298 375048 675354 375057
rect 675298 374983 675354 374992
rect 675312 373402 675340 374983
rect 675312 373374 675418 373402
rect 675758 373008 675814 373017
rect 675758 372943 675814 372952
rect 675772 372776 675800 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 355056 674710 355065
rect 674654 354991 674710 355000
rect 676034 353832 676090 353841
rect 676090 353790 676260 353818
rect 676034 353767 676090 353776
rect 674746 353424 674802 353433
rect 674746 353359 674802 353368
rect 674562 352200 674618 352209
rect 674562 352135 674618 352144
rect 674378 349480 674434 349489
rect 674378 349415 674434 349424
rect 674392 332761 674420 349415
rect 674576 340874 674604 352135
rect 674576 340846 674696 340874
rect 674378 332752 674434 332761
rect 674378 332687 674434 332696
rect 674668 326346 674696 340846
rect 674760 340558 674788 353359
rect 675942 349208 675998 349217
rect 676232 349194 676260 353790
rect 675998 349166 676260 349194
rect 675942 349143 675998 349152
rect 674760 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675404 339017 675432 339252
rect 675390 339008 675446 339017
rect 675390 338943 675446 338952
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675128 336829 675418 336857
rect 675114 336696 675170 336705
rect 675114 336631 675170 336640
rect 675758 336696 675814 336705
rect 675758 336631 675814 336640
rect 675128 333078 675156 336631
rect 675772 336192 675800 336631
rect 675404 335186 675432 335580
rect 675312 335158 675432 335186
rect 675312 333985 675340 335158
rect 675298 333976 675354 333985
rect 675298 333911 675354 333920
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675114 332344 675170 332353
rect 675114 332279 675170 332288
rect 675758 332344 675814 332353
rect 675758 332279 675814 332288
rect 675128 331242 675156 332279
rect 675772 331875 675800 332279
rect 675128 331214 675418 331242
rect 675114 331120 675170 331129
rect 675114 331055 675170 331064
rect 675128 330049 675156 331055
rect 675128 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675114 327584 675170 327593
rect 675170 327542 675418 327570
rect 675114 327519 675170 327528
rect 675312 326454 675432 326482
rect 675312 326346 675340 326454
rect 674668 326318 675340 326346
rect 675404 326332 675432 326454
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 309632 674710 309641
rect 674654 309567 674710 309576
rect 673656 309106 673868 309134
rect 673932 309106 674144 309134
rect 673366 304328 673422 304337
rect 673366 304263 673422 304272
rect 673380 287881 673408 304263
rect 673656 299474 673684 309106
rect 673932 301866 673960 309106
rect 674470 305552 674526 305561
rect 674470 305487 674526 305496
rect 674194 303920 674250 303929
rect 674194 303855 674250 303864
rect 673840 301838 673960 301866
rect 673840 301594 673868 301838
rect 673840 301566 674144 301594
rect 673656 299446 673960 299474
rect 673366 287872 673422 287881
rect 673366 287807 673422 287816
rect 673090 266520 673146 266529
rect 673090 266455 673146 266464
rect 673090 266112 673146 266121
rect 673090 266047 673146 266056
rect 672906 263800 672962 263809
rect 672906 263735 672962 263744
rect 672920 236910 672948 263735
rect 673104 240009 673132 266047
rect 673932 265849 673960 299446
rect 673918 265840 673974 265849
rect 673918 265775 673974 265784
rect 673366 260536 673422 260545
rect 673366 260471 673422 260480
rect 673380 245313 673408 260471
rect 673642 259312 673698 259321
rect 673642 259247 673698 259256
rect 673366 245304 673422 245313
rect 673366 245239 673422 245248
rect 673656 242865 673684 259247
rect 673918 258496 673974 258505
rect 673918 258431 673974 258440
rect 673642 242856 673698 242865
rect 673642 242791 673698 242800
rect 673090 240000 673146 240009
rect 673090 239935 673146 239944
rect 673092 237516 673144 237522
rect 673092 237458 673144 237464
rect 672908 236904 672960 236910
rect 672908 236846 672960 236852
rect 672644 235742 672764 235770
rect 672908 235748 672960 235754
rect 672644 228698 672672 235742
rect 672908 235690 672960 235696
rect 672920 234954 672948 235690
rect 672920 234926 672994 234954
rect 672816 234864 672868 234870
rect 672816 234806 672868 234812
rect 672966 234818 672994 234926
rect 672828 234410 672856 234806
rect 672966 234790 673040 234818
rect 672756 234382 672856 234410
rect 672756 234308 672784 234382
rect 672736 234280 672784 234308
rect 672736 228834 672764 234280
rect 673012 234274 673040 234790
rect 672966 234246 673040 234274
rect 672966 234240 672994 234246
rect 672920 234212 672994 234240
rect 672920 231962 672948 234212
rect 673104 233238 673132 237458
rect 673302 237144 673358 237153
rect 673302 237079 673304 237088
rect 673356 237079 673358 237088
rect 673304 237050 673356 237056
rect 673276 236904 673328 236910
rect 673276 236846 673328 236852
rect 673288 233617 673316 236846
rect 673526 236736 673582 236745
rect 673526 236671 673528 236680
rect 673580 236671 673582 236680
rect 673528 236642 673580 236648
rect 673460 236564 673512 236570
rect 673460 236506 673512 236512
rect 673274 233608 673330 233617
rect 673274 233543 673330 233552
rect 673092 233232 673144 233238
rect 673092 233174 673144 233180
rect 672874 231934 672948 231962
rect 672874 231854 672902 231934
rect 672874 231826 672948 231854
rect 672920 228993 672948 231826
rect 673472 231690 673500 236506
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 673764 236178 673792 236234
rect 673564 236150 673792 236178
rect 673564 232234 673592 236150
rect 673736 235952 673788 235958
rect 673736 235894 673788 235900
rect 673748 232665 673776 235894
rect 673734 232656 673790 232665
rect 673734 232591 673790 232600
rect 673564 232206 673684 232234
rect 673656 232121 673684 232206
rect 673642 232112 673698 232121
rect 673642 232047 673698 232056
rect 673472 231662 673684 231690
rect 673460 231532 673512 231538
rect 673460 231474 673512 231480
rect 673276 230852 673328 230858
rect 673276 230794 673328 230800
rect 673288 229537 673316 230794
rect 673472 230722 673500 231474
rect 673460 230716 673512 230722
rect 673460 230658 673512 230664
rect 673656 230382 673684 231662
rect 673644 230376 673696 230382
rect 673644 230318 673696 230324
rect 673458 230208 673514 230217
rect 673458 230143 673514 230152
rect 673734 230208 673790 230217
rect 673734 230143 673790 230152
rect 673274 229528 673330 229537
rect 673472 229514 673500 230143
rect 673598 230104 673650 230110
rect 673426 229498 673500 229514
rect 673274 229463 673330 229472
rect 673414 229492 673500 229498
rect 673466 229486 673500 229492
rect 673564 230052 673598 230058
rect 673564 230046 673650 230052
rect 673564 230030 673638 230046
rect 673414 229434 673466 229440
rect 673386 229256 673442 229265
rect 673380 229200 673386 229242
rect 673380 229191 673442 229200
rect 673380 229094 673408 229191
rect 673380 229090 673428 229094
rect 673380 229084 673440 229090
rect 673380 229066 673388 229084
rect 673388 229026 673440 229032
rect 673564 228993 673592 230030
rect 673748 229974 673776 230143
rect 673736 229968 673788 229974
rect 673736 229910 673788 229916
rect 673734 229800 673790 229809
rect 673734 229735 673790 229744
rect 673748 229294 673776 229735
rect 673736 229288 673788 229294
rect 673736 229230 673788 229236
rect 672906 228984 672962 228993
rect 672906 228919 672962 228928
rect 673550 228984 673606 228993
rect 673550 228919 673606 228928
rect 672736 228806 672856 228834
rect 672828 228698 672856 228806
rect 673506 228744 673558 228750
rect 672644 228670 672764 228698
rect 672828 228670 673132 228698
rect 673506 228686 673558 228692
rect 672736 228614 672764 228670
rect 672724 228608 672776 228614
rect 672908 228608 672960 228614
rect 672724 228550 672776 228556
rect 672906 228576 672908 228585
rect 672960 228576 672962 228585
rect 672906 228511 672962 228520
rect 673104 228426 673132 228670
rect 673386 228576 673442 228585
rect 673386 228511 673388 228520
rect 673440 228511 673442 228520
rect 673388 228482 673440 228488
rect 673518 228426 673546 228686
rect 673104 228398 673408 228426
rect 673518 228398 673868 228426
rect 672954 227792 673006 227798
rect 673006 227752 673132 227780
rect 672954 227734 673006 227740
rect 672724 227384 672776 227390
rect 672724 227326 672776 227332
rect 672736 227202 672764 227326
rect 672552 227174 672644 227202
rect 672736 227174 672856 227202
rect 672368 226930 672396 227174
rect 672616 226930 672644 227174
rect 672368 226902 672488 226930
rect 672262 226808 672318 226817
rect 672262 226743 672318 226752
rect 672092 226630 672304 226658
rect 671894 226607 671950 226616
rect 672032 226536 672088 226545
rect 672276 226522 672304 226630
rect 672032 226471 672088 226480
rect 672156 226500 672208 226506
rect 671894 226400 671950 226409
rect 671894 226335 671896 226344
rect 671948 226335 671950 226344
rect 671896 226306 671948 226312
rect 672046 226302 672074 226471
rect 672276 226494 672396 226522
rect 672156 226442 672208 226448
rect 672034 226296 672086 226302
rect 672034 226238 672086 226244
rect 672168 225978 672196 226442
rect 672000 225950 672196 225978
rect 671820 225752 671872 225758
rect 671818 225720 671820 225729
rect 671872 225720 671874 225729
rect 671818 225655 671874 225664
rect 672000 224954 672028 225950
rect 672170 225720 672226 225729
rect 672170 225655 672226 225664
rect 671908 224926 672028 224954
rect 672184 224954 672212 225655
rect 672184 224926 672304 224954
rect 671908 224505 671936 224926
rect 672078 224768 672134 224777
rect 672078 224703 672134 224712
rect 671894 224496 671950 224505
rect 671894 224431 671950 224440
rect 671894 219464 671950 219473
rect 671894 219399 671950 219408
rect 671908 174865 671936 219399
rect 672092 219201 672120 224703
rect 672078 219192 672134 219201
rect 672078 219127 672134 219136
rect 672276 216322 672304 224926
rect 672184 216294 672304 216322
rect 672184 216209 672212 216294
rect 672170 216200 672226 216209
rect 672170 216135 672226 216144
rect 672368 215294 672396 226494
rect 672276 215266 672396 215294
rect 672078 214160 672134 214169
rect 672078 214095 672134 214104
rect 672092 201113 672120 214095
rect 672276 203017 672304 215266
rect 672460 210497 672488 226902
rect 672552 226902 672644 226930
rect 672552 210610 672580 226902
rect 672828 226794 672856 227174
rect 672736 226766 672856 226794
rect 672736 225706 672764 226766
rect 673104 226658 673132 227752
rect 673104 226630 673224 226658
rect 673196 226545 673224 226630
rect 673182 226536 673238 226545
rect 673182 226471 673238 226480
rect 673380 226386 673408 228398
rect 673288 226358 673408 226386
rect 672860 225720 672916 225729
rect 672736 225678 672860 225706
rect 672860 225655 672916 225664
rect 672906 224904 672962 224913
rect 672906 224839 672962 224848
rect 672722 211984 672778 211993
rect 672722 211919 672778 211928
rect 672736 211177 672764 211919
rect 672722 211168 672778 211177
rect 672722 211103 672778 211112
rect 672552 210582 672672 210610
rect 672446 210488 672502 210497
rect 672446 210423 672502 210432
rect 672644 210338 672672 210582
rect 672552 210310 672672 210338
rect 672262 203008 672318 203017
rect 672262 202943 672318 202952
rect 672078 201104 672134 201113
rect 672078 201039 672134 201048
rect 672552 185609 672580 210310
rect 672722 210216 672778 210225
rect 672722 210151 672778 210160
rect 672538 185600 672594 185609
rect 672538 185535 672594 185544
rect 672262 183560 672318 183569
rect 672262 183495 672318 183504
rect 672078 182064 672134 182073
rect 672078 181999 672134 182008
rect 671894 174856 671950 174865
rect 671894 174791 671950 174800
rect 671710 172952 671766 172961
rect 671710 172887 671766 172896
rect 671894 169960 671950 169969
rect 671894 169895 671950 169904
rect 671710 166968 671766 166977
rect 671710 166903 671766 166912
rect 671526 158264 671582 158273
rect 671526 158199 671582 158208
rect 670804 157306 671384 157334
rect 670804 150278 670832 157306
rect 670792 150272 670844 150278
rect 670792 150214 670844 150220
rect 670606 149016 670662 149025
rect 670606 148951 670662 148960
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670148 118380 670200 118386
rect 670148 118322 670200 118328
rect 668674 114135 668730 114144
rect 669964 114164 670016 114170
rect 668124 114106 668176 114112
rect 669964 114106 670016 114112
rect 590566 113384 590622 113393
rect 590566 113319 590622 113328
rect 590580 110498 590608 113319
rect 668136 112577 668164 114106
rect 671356 113174 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670712 113146 671384 113174
rect 668122 112568 668178 112577
rect 668122 112503 668178 112512
rect 668306 111888 668362 111897
rect 668306 111823 668362 111832
rect 590568 110492 590620 110498
rect 590568 110434 590620 110440
rect 668030 109304 668086 109313
rect 668030 109239 668086 109248
rect 590108 107092 590160 107098
rect 590108 107034 590160 107040
rect 589648 106956 589700 106962
rect 589648 106898 589700 106904
rect 589922 106856 589978 106865
rect 589922 106791 589978 106800
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100774 589504 101895
rect 589464 100768 589516 100774
rect 589464 100710 589516 100716
rect 588544 82816 588596 82822
rect 588544 82758 588596 82764
rect 589936 80714 589964 106791
rect 667204 106208 667256 106214
rect 667204 106150 667256 106156
rect 667216 106049 667244 106150
rect 666650 106040 666706 106049
rect 666650 105975 666706 105984
rect 667202 106040 667258 106049
rect 667202 105975 667258 105984
rect 590106 103592 590162 103601
rect 590106 103527 590162 103536
rect 590120 93158 590148 103527
rect 613272 100150 613608 100178
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596468 100014 597080 100042
rect 597572 100014 597816 100042
rect 597940 100014 598552 100042
rect 599136 100014 599288 100042
rect 599688 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 595272 99346 595300 100014
rect 595260 99340 595312 99346
rect 595260 99282 595312 99288
rect 594064 95940 594116 95946
rect 594064 95882 594116 95888
rect 590108 93152 590160 93158
rect 590108 93094 590160 93100
rect 589924 80708 589976 80714
rect 589924 80650 589976 80656
rect 585968 80096 586020 80102
rect 585968 80038 586020 80044
rect 585782 77888 585838 77897
rect 585782 77823 585838 77832
rect 581644 75472 581696 75478
rect 581644 75414 581696 75420
rect 580264 73160 580316 73166
rect 580264 73102 580316 73108
rect 579158 71360 579214 71369
rect 579158 71295 579214 71304
rect 579526 68096 579582 68105
rect 579526 68031 579582 68040
rect 579540 67658 579568 68031
rect 579528 67652 579580 67658
rect 579528 67594 579580 67600
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 60716 579580 60722
rect 579528 60658 579580 60664
rect 579540 60353 579568 60658
rect 579526 60344 579582 60353
rect 579526 60279 579582 60288
rect 581644 60036 581696 60042
rect 581644 59978 581696 59984
rect 580264 58812 580316 58818
rect 580264 58754 580316 58760
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 579528 56568 579580 56574
rect 579528 56510 579580 56516
rect 579540 56137 579568 56510
rect 579526 56128 579582 56137
rect 579526 56063 579582 56072
rect 578884 55072 578936 55078
rect 578884 55014 578936 55020
rect 580276 54777 580304 58754
rect 581656 55049 581684 59978
rect 581642 55040 581698 55049
rect 581642 54975 581698 54984
rect 585796 54942 585824 77823
rect 588544 74860 588596 74866
rect 588544 74802 588596 74808
rect 588556 56574 588584 74802
rect 588544 56568 588596 56574
rect 588544 56510 588596 56516
rect 585784 54936 585836 54942
rect 585784 54878 585836 54884
rect 580262 54768 580318 54777
rect 580262 54703 580318 54712
rect 594076 54505 594104 95882
rect 595272 93854 595300 99282
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 596192 54806 596220 100014
rect 596468 55622 596496 100014
rect 596456 55616 596508 55622
rect 596456 55558 596508 55564
rect 596180 54800 596232 54806
rect 596180 54742 596232 54748
rect 597572 54670 597600 100014
rect 597940 56166 597968 100014
rect 598940 96960 598992 96966
rect 598940 96902 598992 96908
rect 597928 56160 597980 56166
rect 597928 56102 597980 56108
rect 598952 56030 598980 96902
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 599136 55894 599164 100014
rect 599688 96966 599716 100014
rect 600424 97306 600452 100014
rect 600412 97300 600464 97306
rect 600412 97242 600464 97248
rect 599676 96960 599728 96966
rect 599676 96902 599728 96908
rect 600884 84194 600912 100014
rect 601896 95946 601924 100014
rect 601884 95940 601936 95946
rect 601884 95882 601936 95888
rect 602356 84194 602384 100014
rect 600332 84166 600912 84194
rect 601896 84166 602384 84194
rect 600332 57254 600360 84166
rect 601896 58818 601924 84166
rect 603092 60042 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 607168 100042
rect 607384 100014 607720 100042
rect 608120 100014 608456 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 604426 99742 604500 99770
rect 603080 60036 603132 60042
rect 603080 59978 603132 59984
rect 601884 58812 601936 58818
rect 601884 58754 601936 58760
rect 604472 58682 604500 99742
rect 605484 97986 605512 100014
rect 605472 97980 605524 97986
rect 605472 97922 605524 97928
rect 606220 96830 606248 100014
rect 606484 97980 606536 97986
rect 606484 97922 606536 97928
rect 606208 96824 606260 96830
rect 606208 96766 606260 96772
rect 606496 76566 606524 97922
rect 607140 93854 607168 100014
rect 607692 96082 607720 100014
rect 607680 96076 607732 96082
rect 607680 96018 607732 96024
rect 608428 94518 608456 100014
rect 609164 96218 609192 100014
rect 609152 96212 609204 96218
rect 609152 96154 609204 96160
rect 608416 94512 608468 94518
rect 608416 94454 608468 94460
rect 607140 93826 607260 93854
rect 607232 88330 607260 93826
rect 607220 88324 607272 88330
rect 607220 88266 607272 88272
rect 609900 85542 609928 100014
rect 610636 96354 610664 100014
rect 610624 96348 610676 96354
rect 610624 96290 610676 96296
rect 611280 91050 611308 100014
rect 612108 96966 612136 100014
rect 612660 97306 612688 100014
rect 613384 100020 613436 100026
rect 613384 99962 613436 99968
rect 612648 97300 612700 97306
rect 612648 97242 612700 97248
rect 612096 96960 612148 96966
rect 612096 96902 612148 96908
rect 612648 96960 612700 96966
rect 612648 96902 612700 96908
rect 612004 96824 612056 96830
rect 612004 96766 612056 96772
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 612016 76702 612044 96766
rect 612660 77994 612688 96902
rect 612648 77988 612700 77994
rect 612648 77930 612700 77936
rect 612004 76696 612056 76702
rect 612004 76638 612056 76644
rect 606484 76560 606536 76566
rect 606484 76502 606536 76508
rect 605840 66292 605892 66298
rect 605840 66234 605892 66240
rect 605852 58682 605880 66234
rect 613396 64870 613424 99962
rect 613580 95946 613608 100150
rect 615224 100156 615276 100162
rect 615224 100098 615276 100104
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 613994 99742 614068 99770
rect 613568 95940 613620 95946
rect 613568 95882 613620 95888
rect 614040 80850 614068 99742
rect 615052 97578 615080 100014
rect 615040 97572 615092 97578
rect 615040 97514 615092 97520
rect 615236 84194 615264 100098
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 615788 96830 615816 100014
rect 616144 97572 616196 97578
rect 616144 97514 616196 97520
rect 615776 96824 615828 96830
rect 615776 96766 615828 96772
rect 614868 84166 615264 84194
rect 614028 80844 614080 80850
rect 614028 80786 614080 80792
rect 613384 64864 613436 64870
rect 613384 64806 613436 64812
rect 614868 60722 614896 84166
rect 616156 79354 616184 97514
rect 616524 94654 616552 100014
rect 617260 96966 617288 100014
rect 617248 96960 617300 96966
rect 617248 96902 617300 96908
rect 616512 94648 616564 94654
rect 616512 94590 616564 94596
rect 617996 92478 618024 100014
rect 618732 97850 618760 100014
rect 618720 97844 618772 97850
rect 618720 97786 618772 97792
rect 618168 96960 618220 96966
rect 618168 96902 618220 96908
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96902
rect 618904 96824 618956 96830
rect 618904 96766 618956 96772
rect 617340 91044 617392 91050
rect 617340 90986 617392 90992
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 617352 88194 617380 90986
rect 617340 88188 617392 88194
rect 617340 88130 617392 88136
rect 616144 79348 616196 79354
rect 616144 79290 616196 79296
rect 618916 75206 618944 96766
rect 619560 93838 619588 100014
rect 620204 97986 620232 100014
rect 620192 97980 620244 97986
rect 620192 97922 620244 97928
rect 620284 97300 620336 97306
rect 620284 97242 620336 97248
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 620296 76838 620324 97242
rect 620940 96082 620968 100014
rect 621676 97714 621704 100014
rect 622320 98802 622348 100014
rect 622308 98796 622360 98802
rect 622308 98738 622360 98744
rect 621664 97708 621716 97714
rect 621664 97650 621716 97656
rect 623148 97578 623176 100014
rect 623700 99074 623728 100014
rect 624620 99346 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628236 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635504 100042
rect 625034 99742 625108 99770
rect 624608 99340 624660 99346
rect 624608 99282 624660 99288
rect 623688 99068 623740 99074
rect 623688 99010 623740 99016
rect 625080 98666 625108 99742
rect 625068 98660 625120 98666
rect 625068 98602 625120 98608
rect 625436 97844 625488 97850
rect 625436 97786 625488 97792
rect 623136 97572 623188 97578
rect 623136 97514 623188 97520
rect 623044 96348 623096 96354
rect 623044 96290 623096 96296
rect 621664 96212 621716 96218
rect 621664 96154 621716 96160
rect 620744 96076 620796 96082
rect 620744 96018 620796 96024
rect 620928 96076 620980 96082
rect 620928 96018 620980 96024
rect 620756 89690 620784 96018
rect 620744 89684 620796 89690
rect 620744 89626 620796 89632
rect 621676 84182 621704 96154
rect 623056 86494 623084 96290
rect 624424 94512 624476 94518
rect 624424 94454 624476 94460
rect 623044 86488 623096 86494
rect 623044 86430 623096 86436
rect 621664 84176 621716 84182
rect 621664 84118 621716 84124
rect 624436 82929 624464 94454
rect 625448 93129 625476 97786
rect 626092 96898 626120 100014
rect 626828 99210 626856 100014
rect 626816 99204 626868 99210
rect 626816 99146 626868 99152
rect 626264 97980 626316 97986
rect 626264 97922 626316 97928
rect 626080 96892 626132 96898
rect 626080 96834 626132 96840
rect 625804 94648 625856 94654
rect 625804 94590 625856 94596
rect 625434 93120 625490 93129
rect 625434 93055 625490 93064
rect 625436 92472 625488 92478
rect 625436 92414 625488 92420
rect 625448 91633 625476 92414
rect 625434 91624 625490 91633
rect 625434 91559 625490 91568
rect 625816 89729 625844 94590
rect 626276 94489 626304 97922
rect 627564 97442 627592 100014
rect 627552 97436 627604 97442
rect 627552 97378 627604 97384
rect 628208 96762 628236 100014
rect 628380 97708 628432 97714
rect 628380 97650 628432 97656
rect 628196 96756 628248 96762
rect 628196 96698 628248 96704
rect 626448 96076 626500 96082
rect 626448 96018 626500 96024
rect 626460 95441 626488 96018
rect 628392 95826 628420 97650
rect 629036 97306 629064 100014
rect 629772 98938 629800 100014
rect 629760 98932 629812 98938
rect 629760 98874 629812 98880
rect 630508 98802 630536 100014
rect 629484 98796 629536 98802
rect 629484 98738 629536 98744
rect 630496 98796 630548 98802
rect 630496 98738 630548 98744
rect 629024 97300 629076 97306
rect 629024 97242 629076 97248
rect 629496 95826 629524 98738
rect 630680 97572 630732 97578
rect 630680 97514 630732 97520
rect 630692 95826 630720 97514
rect 631244 96626 631272 100014
rect 631980 97578 632008 100014
rect 632152 99068 632204 99074
rect 632152 99010 632204 99016
rect 631968 97572 632020 97578
rect 631968 97514 632020 97520
rect 631232 96620 631284 96626
rect 631232 96562 631284 96568
rect 632164 95826 632192 99010
rect 632716 97986 632744 100014
rect 632980 99340 633032 99346
rect 632980 99282 633032 99288
rect 632704 97980 632756 97986
rect 632704 97922 632756 97928
rect 628392 95798 628728 95826
rect 629496 95798 629832 95826
rect 630692 95798 631028 95826
rect 632132 95798 632192 95826
rect 632992 95826 633020 99282
rect 633360 97714 633388 100014
rect 633348 97708 633400 97714
rect 633348 97650 633400 97656
rect 634188 97170 634216 100014
rect 634452 98660 634504 98666
rect 634452 98602 634504 98608
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 632992 95798 633328 95826
rect 634464 95690 634492 98602
rect 634740 97034 634768 100014
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635280 96892 635332 96898
rect 635280 96834 635332 96840
rect 635292 95826 635320 96834
rect 635476 95946 635504 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 637560 100014 637896 100042
rect 638296 100014 638632 100042
rect 639032 100014 639368 100042
rect 639768 100014 640104 100042
rect 640504 100014 640840 100042
rect 641240 100014 641576 100042
rect 641976 100014 642588 100042
rect 642712 100014 643048 100042
rect 643448 100014 643784 100042
rect 644184 100014 644336 100042
rect 644920 100014 645256 100042
rect 645656 100014 645808 100042
rect 646392 100014 646728 100042
rect 635752 96937 635780 100014
rect 636384 99204 636436 99210
rect 636384 99146 636436 99152
rect 635738 96928 635794 96937
rect 635738 96863 635794 96872
rect 635464 95940 635516 95946
rect 635464 95882 635516 95888
rect 636396 95826 636424 99146
rect 637040 96937 637068 100014
rect 637868 98666 637896 100014
rect 637856 98660 637908 98666
rect 637856 98602 637908 98608
rect 637580 97436 637632 97442
rect 637580 97378 637632 97384
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 95826 637620 97378
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637592 95798 637928 95826
rect 638604 95810 638632 100014
rect 639052 96756 639104 96762
rect 639052 96698 639104 96704
rect 639064 95826 639092 96698
rect 639340 96354 639368 100014
rect 639880 97436 639932 97442
rect 639880 97378 639932 97384
rect 639328 96348 639380 96354
rect 639328 96290 639380 96296
rect 638592 95804 638644 95810
rect 639032 95798 639092 95826
rect 639892 95826 639920 97378
rect 640076 96490 640104 100014
rect 640064 96484 640116 96490
rect 640064 96426 640116 96432
rect 640812 96218 640840 100014
rect 640984 98932 641036 98938
rect 640984 98874 641036 98880
rect 640800 96212 640852 96218
rect 640800 96154 640852 96160
rect 640996 95826 641024 98874
rect 641548 96082 641576 100014
rect 642180 98796 642232 98802
rect 642180 98738 642232 98744
rect 641536 96076 641588 96082
rect 641536 96018 641588 96024
rect 642192 95826 642220 98738
rect 642560 96098 642588 100014
rect 643020 97170 643048 100014
rect 643756 97850 643784 100014
rect 644020 97980 644072 97986
rect 644020 97922 644072 97928
rect 643744 97844 643796 97850
rect 643744 97786 643796 97792
rect 643468 97708 643520 97714
rect 643468 97650 643520 97656
rect 643008 97164 643060 97170
rect 643008 97106 643060 97112
rect 643192 96620 643244 96626
rect 643192 96562 643244 96568
rect 642560 96070 642680 96098
rect 639892 95798 640228 95826
rect 640996 95798 641332 95826
rect 642192 95798 642528 95826
rect 638592 95746 638644 95752
rect 634432 95662 634492 95690
rect 626446 95432 626502 95441
rect 626446 95367 626502 95376
rect 642652 95266 642680 96070
rect 642824 95804 642876 95810
rect 642824 95746 642876 95752
rect 642836 95538 642864 95746
rect 642824 95532 642876 95538
rect 642824 95474 642876 95480
rect 642640 95260 642692 95266
rect 642640 95202 642692 95208
rect 643204 95169 643232 96562
rect 643190 95160 643246 95169
rect 643190 95095 643246 95104
rect 626262 94480 626318 94489
rect 626262 94415 626318 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626460 93537 626488 93774
rect 626446 93528 626502 93537
rect 626446 93463 626502 93472
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90681 626488 90986
rect 626446 90672 626502 90681
rect 626446 90607 626502 90616
rect 625802 89720 625858 89729
rect 625802 89655 625858 89664
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626460 88913 626488 89626
rect 626446 88904 626502 88913
rect 626446 88839 626502 88848
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 625620 88188 625672 88194
rect 625620 88130 625672 88136
rect 625632 87009 625660 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 643480 87145 643508 97650
rect 643744 97028 643796 97034
rect 643744 96970 643796 96976
rect 643466 87136 643522 87145
rect 643466 87071 643522 87080
rect 625618 87000 625674 87009
rect 625618 86935 625674 86944
rect 626448 86488 626500 86494
rect 626448 86430 626500 86436
rect 626460 86057 626488 86430
rect 626446 86048 626502 86057
rect 626446 85983 626502 85992
rect 626448 85536 626500 85542
rect 626448 85478 626500 85484
rect 626460 85105 626488 85478
rect 626446 85096 626502 85105
rect 626446 85031 626502 85040
rect 625620 84176 625672 84182
rect 625618 84144 625620 84153
rect 625672 84144 625674 84153
rect 625618 84079 625674 84088
rect 624422 82920 624478 82929
rect 624422 82855 624478 82864
rect 643756 82793 643784 96970
rect 644032 89729 644060 97922
rect 644308 97442 644336 100014
rect 644940 97572 644992 97578
rect 644940 97514 644992 97520
rect 644296 97436 644348 97442
rect 644296 97378 644348 97384
rect 644756 97300 644808 97306
rect 644756 97242 644808 97248
rect 644480 95260 644532 95266
rect 644480 95202 644532 95208
rect 644492 93838 644520 95202
rect 644480 93832 644532 93838
rect 644480 93774 644532 93780
rect 644018 89720 644074 89729
rect 644018 89655 644074 89664
rect 644768 84697 644796 97242
rect 644952 92177 644980 97514
rect 645228 97102 645256 100014
rect 645216 97096 645268 97102
rect 645216 97038 645268 97044
rect 644938 92168 644994 92177
rect 644938 92103 644994 92112
rect 645780 88806 645808 100014
rect 646700 96966 646728 100014
rect 647114 99770 647142 100028
rect 647864 100014 648200 100042
rect 648600 100014 648936 100042
rect 649336 100014 649672 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 647114 99742 647188 99770
rect 647160 97578 647188 99742
rect 647148 97572 647200 97578
rect 647148 97514 647200 97520
rect 646688 96960 646740 96966
rect 646688 96902 646740 96908
rect 647884 96960 647936 96966
rect 647884 96902 647936 96908
rect 647700 96484 647752 96490
rect 647700 96426 647752 96432
rect 647712 95946 647740 96426
rect 646044 95940 646096 95946
rect 646044 95882 646096 95888
rect 647700 95940 647752 95946
rect 647700 95882 647752 95888
rect 645768 88800 645820 88806
rect 645768 88742 645820 88748
rect 644754 84688 644810 84697
rect 644754 84623 644810 84632
rect 643742 82784 643798 82793
rect 643742 82719 643798 82728
rect 628654 81696 628710 81705
rect 628654 81631 628710 81640
rect 628668 80986 628696 81631
rect 628656 80980 628708 80986
rect 628656 80922 628708 80928
rect 631520 80974 631856 81002
rect 639064 80974 639308 81002
rect 642456 80980 642508 80986
rect 629206 80880 629262 80889
rect 629206 80815 629262 80824
rect 629220 79490 629248 80815
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 623044 77308 623096 77314
rect 623044 77250 623096 77256
rect 628380 77308 628432 77314
rect 628380 77250 628432 77256
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 618904 75200 618956 75206
rect 618904 75142 618956 75148
rect 614856 60716 614908 60722
rect 614856 60658 614908 60664
rect 604460 58676 604512 58682
rect 604460 58618 604512 58624
rect 605840 58676 605892 58682
rect 605840 58618 605892 58624
rect 600320 57248 600372 57254
rect 600320 57190 600372 57196
rect 599124 55888 599176 55894
rect 599124 55830 599176 55836
rect 597560 54664 597612 54670
rect 597560 54606 597612 54612
rect 623056 54534 623084 77250
rect 628392 75290 628420 77250
rect 631060 75954 631088 78066
rect 631520 77314 631548 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 80472 633954 80481
rect 633898 80407 633954 80416
rect 633912 77450 633940 80407
rect 633900 77444 633952 77450
rect 633900 77386 633952 77392
rect 631508 77308 631560 77314
rect 631508 77250 631560 77256
rect 631048 75948 631100 75954
rect 631048 75890 631100 75896
rect 631060 75290 631088 75890
rect 633912 75290 633940 77386
rect 636120 77294 636148 80650
rect 638868 79484 638920 79490
rect 638868 79426 638920 79432
rect 638880 78334 638908 79426
rect 638868 78328 638920 78334
rect 638868 78270 638920 78276
rect 639064 78130 639092 80974
rect 642456 80922 642508 80928
rect 639052 78124 639104 78130
rect 639052 78066 639104 78072
rect 639602 77888 639658 77897
rect 639602 77823 639658 77832
rect 636120 77266 636332 77294
rect 628176 75276 628420 75290
rect 628162 75262 628420 75276
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 628162 74882 628190 75262
rect 636304 75154 636332 77266
rect 639616 75290 639644 77823
rect 642468 75290 642496 80922
rect 645308 78328 645360 78334
rect 645308 78270 645360 78276
rect 645320 75290 645348 78270
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 628024 74868 628190 74882
rect 628024 74866 628176 74868
rect 628012 74860 628176 74866
rect 628064 74854 628176 74860
rect 628012 74802 628064 74808
rect 624424 67652 624476 67658
rect 624424 67594 624476 67600
rect 624436 55894 624464 67594
rect 646056 64874 646084 95882
rect 646228 95668 646280 95674
rect 646228 95610 646280 95616
rect 646240 68921 646268 95610
rect 647896 87174 647924 96902
rect 648172 96490 648200 100014
rect 648160 96484 648212 96490
rect 648160 96426 648212 96432
rect 648908 95810 648936 100014
rect 649264 97096 649316 97102
rect 649264 97038 649316 97044
rect 648896 95804 648948 95810
rect 648896 95746 648948 95752
rect 648528 95532 648580 95538
rect 648528 95474 648580 95480
rect 648540 92478 648568 95474
rect 648528 92472 648580 92478
rect 648528 92414 648580 92420
rect 647884 87168 647936 87174
rect 647884 87110 647936 87116
rect 649276 87038 649304 97038
rect 649644 96626 649672 100014
rect 650380 97170 650408 100014
rect 651116 97986 651144 100014
rect 651104 97980 651156 97986
rect 651104 97922 651156 97928
rect 651852 97850 651880 100014
rect 650644 97844 650696 97850
rect 650644 97786 650696 97792
rect 651840 97844 651892 97850
rect 651840 97786 651892 97792
rect 650368 97164 650420 97170
rect 650368 97106 650420 97112
rect 649632 96620 649684 96626
rect 649632 96562 649684 96568
rect 649264 87032 649316 87038
rect 649264 86974 649316 86980
rect 650656 86630 650684 97786
rect 652588 96626 652616 100014
rect 650828 96620 650880 96626
rect 650828 96562 650880 96568
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 650840 86902 650868 96562
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 650828 86896 650880 86902
rect 650828 86838 650880 86844
rect 652036 86766 652064 96426
rect 653324 96354 653352 100014
rect 653968 97306 653996 100014
rect 653956 97300 654008 97306
rect 653956 97242 654008 97248
rect 654796 96966 654824 100014
rect 655440 97986 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655060 97980 655112 97986
rect 655060 97922 655112 97928
rect 655428 97980 655480 97986
rect 655428 97922 655480 97928
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 653864 96484 653916 96490
rect 653864 96426 653916 96432
rect 653312 96348 653364 96354
rect 653312 96290 653364 96296
rect 653404 95940 653456 95946
rect 653404 95882 653456 95888
rect 652024 86760 652076 86766
rect 652024 86702 652076 86708
rect 650644 86624 650696 86630
rect 650644 86566 650696 86572
rect 653416 86358 653444 95882
rect 653876 90794 653904 96426
rect 654876 93832 654928 93838
rect 654876 93774 654928 93780
rect 654888 92585 654916 93774
rect 655072 93401 655100 97922
rect 655244 97300 655296 97306
rect 655244 97242 655296 97248
rect 655256 94217 655284 97242
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655242 94208 655298 94217
rect 655242 94143 655298 94152
rect 655058 93392 655114 93401
rect 655058 93327 655114 93336
rect 655440 92698 655468 96902
rect 655072 92670 655468 92698
rect 654874 92576 654930 92585
rect 654874 92511 654930 92520
rect 653876 90766 654180 90794
rect 654152 90681 654180 90766
rect 654138 90672 654194 90681
rect 654138 90607 654194 90616
rect 655072 88330 655100 92670
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655808 89865 655836 100014
rect 656820 97306 656848 100014
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97578 658228 99742
rect 659212 97714 659240 100014
rect 659948 97850 659976 100014
rect 660396 98660 660448 98666
rect 660396 98602 660448 98608
rect 659568 97844 659620 97850
rect 659568 97786 659620 97792
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659200 97708 659252 97714
rect 659200 97650 659252 97656
rect 658004 97572 658056 97578
rect 658004 97514 658056 97520
rect 658188 97572 658240 97578
rect 658188 97514 658240 97520
rect 658016 97034 658044 97514
rect 658832 97436 658884 97442
rect 658832 97378 658884 97384
rect 658280 97164 658332 97170
rect 658280 97106 658332 97112
rect 658004 97028 658056 97034
rect 658004 96970 658056 96976
rect 658292 95132 658320 97106
rect 658844 95132 658872 97378
rect 659580 95132 659608 97786
rect 660120 96824 660172 96830
rect 660120 96766 660172 96772
rect 660132 95132 660160 96766
rect 660408 95146 660436 98602
rect 660684 96762 660712 100014
rect 662512 97980 662564 97986
rect 662512 97922 662564 97928
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660672 96756 660724 96762
rect 660672 96698 660724 96704
rect 660408 95118 660698 95146
rect 661420 95132 661448 97242
rect 661960 97028 662012 97034
rect 661960 96970 662012 96976
rect 661972 95132 662000 96970
rect 662524 95132 662552 97922
rect 665548 97844 665600 97850
rect 665548 97786 665600 97792
rect 663892 97708 663944 97714
rect 663892 97650 663944 97656
rect 663064 97572 663116 97578
rect 663064 97514 663116 97520
rect 663076 95132 663104 97514
rect 663248 96756 663300 96762
rect 663248 96698 663300 96704
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 657452 88800 657504 88806
rect 662328 88800 662380 88806
rect 657504 88748 657754 88754
rect 657452 88742 657754 88748
rect 657464 88726 657754 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 655060 88324 655112 88330
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 655060 88266 655112 88272
rect 658464 88266 658516 88272
rect 657188 87174 657216 88196
rect 657176 87168 657228 87174
rect 657176 87110 657228 87116
rect 658844 86902 658872 88196
rect 659580 86902 659608 88196
rect 658832 86896 658884 86902
rect 658832 86838 658884 86844
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86358 660160 88196
rect 660684 87038 660712 88196
rect 660672 87032 660724 87038
rect 660672 86974 660724 86980
rect 661420 86630 661448 88196
rect 662524 86766 662552 88196
rect 663260 86902 663288 96698
rect 663708 96212 663760 96218
rect 663708 96154 663760 96160
rect 663720 96098 663748 96154
rect 663720 96070 663840 96098
rect 663812 92154 663840 96070
rect 663720 92126 663840 92154
rect 663720 92041 663748 92126
rect 663706 92032 663762 92041
rect 663706 91967 663762 91976
rect 663904 88806 663932 97650
rect 665364 96620 665416 96626
rect 665364 96562 665416 96568
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89049 664208 96290
rect 665180 96076 665232 96082
rect 665180 96018 665232 96024
rect 664628 95940 664680 95946
rect 664628 95882 664680 95888
rect 664444 92540 664496 92546
rect 664444 92482 664496 92488
rect 664166 89040 664222 89049
rect 664166 88975 664222 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663248 86896 663300 86902
rect 663248 86838 663300 86844
rect 662512 86760 662564 86766
rect 662512 86702 662564 86708
rect 661408 86624 661460 86630
rect 661408 86566 661460 86572
rect 653404 86352 653456 86358
rect 653404 86294 653456 86300
rect 660120 86352 660172 86358
rect 660120 86294 660172 86300
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 647056 76696 647108 76702
rect 647056 76638 647108 76644
rect 646872 75200 646924 75206
rect 646872 75142 646924 75148
rect 646884 73001 646912 75142
rect 647068 74497 647096 76638
rect 647054 74488 647110 74497
rect 647054 74423 647110 74432
rect 646870 72992 646926 73001
rect 646870 72927 646926 72936
rect 647344 70009 647372 80786
rect 648988 79348 649040 79354
rect 648988 79290 649040 79296
rect 647516 77988 647568 77994
rect 647516 77930 647568 77936
rect 647330 70000 647386 70009
rect 647330 69935 647386 69944
rect 646226 68912 646282 68921
rect 646226 68847 646282 68856
rect 647528 65521 647556 77930
rect 649000 71505 649028 79290
rect 649172 76832 649224 76838
rect 649172 76774 649224 76780
rect 648986 71496 649042 71505
rect 648986 71431 649042 71440
rect 649184 67017 649212 76774
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 649170 67008 649226 67017
rect 649170 66943 649226 66952
rect 647514 65512 647570 65521
rect 647514 65447 647570 65456
rect 646056 64846 646176 64874
rect 646148 64433 646176 64846
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 624424 55888 624476 55894
rect 624424 55830 624476 55836
rect 623044 54528 623096 54534
rect 594062 54496 594118 54505
rect 623044 54470 623096 54476
rect 594062 54431 594118 54440
rect 577686 54224 577742 54233
rect 577686 54159 577742 54168
rect 575480 54120 575532 54126
rect 575480 54062 575532 54068
rect 574928 53984 574980 53990
rect 574928 53926 574980 53932
rect 574008 53848 574060 53854
rect 574008 53790 574060 53796
rect 460754 53680 460810 53689
rect 459468 53644 459520 53650
rect 459468 53586 459520 53592
rect 460388 53644 460440 53650
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 462594 53680 462650 53689
rect 462274 53644 462326 53650
rect 461674 53615 461730 53624
rect 460388 53586 460440 53592
rect 129004 53372 129056 53378
rect 129004 53314 129056 53320
rect 126888 51740 126940 51746
rect 126888 51682 126940 51688
rect 126900 50794 126928 51682
rect 126888 50788 126940 50794
rect 126888 50730 126940 50736
rect 129016 50674 129044 53314
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 129464 51876 129516 51882
rect 129464 51818 129516 51824
rect 129280 50788 129332 50794
rect 129280 50730 129332 50736
rect 129016 50646 129228 50674
rect 128636 50516 128688 50522
rect 128636 50458 128688 50464
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 128452 49156 128504 49162
rect 128452 49098 128504 49104
rect 47584 49020 47636 49026
rect 47584 48962 47636 48968
rect 128464 44674 128492 49098
rect 128648 48142 128676 50458
rect 129004 50380 129056 50386
rect 129004 50322 129056 50328
rect 128636 48136 128688 48142
rect 128636 48078 128688 48084
rect 128452 44668 128504 44674
rect 128452 44610 128504 44616
rect 129016 44198 129044 50322
rect 129200 47734 129228 50646
rect 129292 48314 129320 50730
rect 129292 48286 129412 48314
rect 129188 47728 129240 47734
rect 129188 47670 129240 47676
rect 129384 44538 129412 48286
rect 129476 47682 129504 51818
rect 129648 49020 129700 49026
rect 129648 48962 129700 48968
rect 129660 48314 129688 48962
rect 129660 48286 129780 48314
rect 129476 47654 129596 47682
rect 129568 45082 129596 47654
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129752 44946 129780 48286
rect 129740 44940 129792 44946
rect 129740 44882 129792 44888
rect 129372 44532 129424 44538
rect 129372 44474 129424 44480
rect 129004 44192 129056 44198
rect 129004 44134 129056 44140
rect 130396 43926 130424 53178
rect 312360 53168 312412 53174
rect 130568 53100 130620 53106
rect 130568 53042 130620 53048
rect 130580 44062 130608 53042
rect 306024 52494 306052 53108
rect 145380 52488 145432 52494
rect 145380 52430 145432 52436
rect 306012 52488 306064 52494
rect 306012 52430 306064 52436
rect 130752 52012 130804 52018
rect 130752 51954 130804 51960
rect 130764 44334 130792 51954
rect 145392 50810 145420 52430
rect 145084 50782 145420 50810
rect 308048 50289 308076 53108
rect 309704 53094 310040 53122
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 309704 49745 309732 53094
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53586
rect 459926 53408 459982 53417
rect 459926 53343 459982 53352
rect 459940 52578 459968 53343
rect 460400 52578 460428 53586
rect 460768 52578 460796 53615
rect 461308 53508 461360 53514
rect 461308 53450 461360 53456
rect 461320 52578 461348 53450
rect 461688 52578 461716 53615
rect 462148 53604 462274 53632
rect 462148 52578 462176 53604
rect 463698 53680 463754 53689
rect 463666 53650 463698 53666
rect 462594 53615 462650 53624
rect 462964 53644 463016 53650
rect 462274 53586 462326 53592
rect 462608 52578 462636 53615
rect 462964 53586 463016 53592
rect 463148 53644 463200 53650
rect 463148 53586 463200 53592
rect 463654 53644 463698 53650
rect 472254 53680 472310 53689
rect 463706 53615 463754 53624
rect 465172 53644 465224 53650
rect 463654 53586 463706 53592
rect 465172 53586 465224 53592
rect 465356 53644 465408 53650
rect 465356 53586 465408 53592
rect 465540 53644 465592 53650
rect 465540 53586 465592 53592
rect 465724 53644 465776 53650
rect 465724 53586 465776 53592
rect 471888 53644 471940 53650
rect 472254 53615 472256 53624
rect 471888 53586 471940 53592
rect 472308 53615 472310 53624
rect 472440 53644 472492 53650
rect 472256 53586 472308 53592
rect 472440 53586 472492 53592
rect 472624 53644 472676 53650
rect 472624 53586 472676 53592
rect 462976 53281 463004 53586
rect 462962 53272 463018 53281
rect 462962 53207 463018 53216
rect 463160 52578 463188 53586
rect 464528 53372 464580 53378
rect 464528 53314 464580 53320
rect 463608 53236 463660 53242
rect 463608 53178 463660 53184
rect 463620 52578 463648 53178
rect 463746 52828 463798 52834
rect 463746 52770 463798 52776
rect 459172 52550 459508 52578
rect 459632 52550 459968 52578
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462176 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463758 52564 463786 52770
rect 464540 52578 464568 53314
rect 464988 53100 465040 53106
rect 464988 53042 465040 53048
rect 465000 52578 465028 53042
rect 465184 52578 465212 53586
rect 465368 53106 465396 53586
rect 465552 53378 465580 53586
rect 465540 53372 465592 53378
rect 465540 53314 465592 53320
rect 465356 53100 465408 53106
rect 465356 53042 465408 53048
rect 465736 52578 465764 53586
rect 471900 53281 471928 53586
rect 471886 53272 471942 53281
rect 472452 53242 472480 53586
rect 471886 53207 471942 53216
rect 472440 53236 472492 53242
rect 472440 53178 472492 53184
rect 472636 52834 472664 53586
rect 472624 52828 472676 52834
rect 472624 52770 472676 52776
rect 464232 52550 464568 52578
rect 464692 52550 465028 52578
rect 465152 52550 465212 52578
rect 465612 52550 465764 52578
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 309690 49736 309746 49745
rect 309690 49671 309746 49680
rect 132132 48136 132184 48142
rect 132132 48078 132184 48084
rect 131856 47728 131908 47734
rect 131856 47670 131908 47676
rect 131868 44606 131896 47670
rect 131856 44600 131908 44606
rect 131856 44542 131908 44548
rect 132144 44506 132172 48078
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132132 44500 132184 44506
rect 132132 44442 132184 44448
rect 132408 44464 132460 44470
rect 132236 44412 132408 44418
rect 132236 44406 132460 44412
rect 132236 44390 132448 44406
rect 130752 44328 130804 44334
rect 130752 44270 130804 44276
rect 132236 44198 132264 44390
rect 132224 44192 132276 44198
rect 132224 44134 132276 44140
rect 130568 44056 130620 44062
rect 130568 43998 130620 44004
rect 130384 43920 130436 43926
rect 130384 43862 130436 43868
rect 43444 42832 43496 42838
rect 43444 42774 43496 42780
rect 142632 40497 142660 46702
rect 458362 46679 458418 46688
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 310426 44160 310482 44169
rect 310426 44095 310482 44104
rect 364890 44160 364946 44169
rect 364890 44095 364946 44104
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 187344 42092 187372 43522
rect 308954 42800 309010 42809
rect 307300 42764 307352 42770
rect 308954 42735 309010 42744
rect 307300 42706 307352 42712
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 42706
rect 308968 42231 308996 42735
rect 308956 42225 309008 42231
rect 308956 42167 309008 42173
rect 310440 42106 310468 44095
rect 361764 42492 361816 42498
rect 361764 42434 361816 42440
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 42434
rect 364904 42092 364932 44095
rect 431236 43654 431264 44775
rect 431224 43648 431276 43654
rect 431224 43590 431276 43596
rect 369400 42764 369452 42770
rect 369400 42706 369452 42712
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 369412 42498 369440 42706
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 369400 42492 369452 42498
rect 369400 42434 369452 42440
rect 416594 42392 416650 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 416594 42327 416650 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 194322 42055 194378 42064
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415766 42120 415822 42129
rect 405200 42078 405582 42106
rect 415426 42078 415766 42106
rect 416608 42092 416636 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 415766 42055 415822 42064
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42090 427124 42570
rect 431236 42090 431264 42706
rect 455880 42628 455932 42634
rect 455880 42570 455932 42576
rect 443550 42256 443606 42265
rect 443550 42191 443606 42200
rect 427084 42084 427136 42090
rect 427084 42026 427136 42032
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 443564 41585 443592 42191
rect 455892 41954 455920 42570
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 455880 41948 455932 41954
rect 455880 41890 455932 41896
rect 443550 41576 443606 41585
rect 443550 41511 443606 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460860 43489 460888 47654
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461964 44441 461992 47654
rect 462378 47410 462406 47668
rect 462332 47382 462406 47410
rect 462516 47654 462852 47682
rect 462976 47654 463312 47682
rect 461950 44432 462006 44441
rect 461950 44367 462006 44376
rect 462332 43217 462360 47382
rect 462516 44441 462544 47654
rect 462502 44432 462558 44441
rect 462502 44367 462558 44376
rect 462976 43897 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463988 47654 464232 47682
rect 464356 47654 464692 47682
rect 463712 44169 463740 47382
rect 463698 44160 463754 44169
rect 463698 44095 463754 44104
rect 462962 43888 463018 43897
rect 462962 43823 463018 43832
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 463698 42936 463754 42945
rect 463698 42871 463754 42880
rect 463712 42378 463740 42871
rect 463988 42634 464016 47654
rect 464356 42770 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 662432 47433 662460 76502
rect 664456 62082 664484 92482
rect 664640 89865 664668 95882
rect 665192 92585 665220 96018
rect 665178 92576 665234 92585
rect 665178 92511 665234 92520
rect 665376 90681 665404 96562
rect 665560 93401 665588 97786
rect 665546 93392 665602 93401
rect 665546 93327 665602 93336
rect 665362 90672 665418 90681
rect 665362 90607 665418 90616
rect 664626 89856 664682 89865
rect 664626 89791 664682 89800
rect 666664 84194 666692 105975
rect 668044 100162 668072 109239
rect 668320 104417 668348 111823
rect 670712 106214 670740 113146
rect 671540 107681 671568 130863
rect 671724 115841 671752 166903
rect 671908 151745 671936 169895
rect 671894 151736 671950 151745
rect 671894 151671 671950 151680
rect 672092 133793 672120 181999
rect 672276 140321 672304 183495
rect 672262 140312 672318 140321
rect 672262 140247 672318 140256
rect 672078 133784 672134 133793
rect 672078 133719 672134 133728
rect 672736 124001 672764 210151
rect 672920 177857 672948 224839
rect 673288 222194 673316 226358
rect 673642 225448 673698 225457
rect 673642 225383 673698 225392
rect 673458 223952 673514 223961
rect 673458 223887 673514 223896
rect 673104 222166 673316 222194
rect 673104 215294 673132 222166
rect 673472 222057 673500 223887
rect 673458 222048 673514 222057
rect 673458 221983 673514 221992
rect 673656 221513 673684 225383
rect 673840 224954 673868 228398
rect 673748 224926 673868 224954
rect 673748 221626 673776 224926
rect 673932 223689 673960 258431
rect 674116 226273 674144 301566
rect 674208 296714 674236 303855
rect 674484 303770 674512 305487
rect 674668 304858 674696 309567
rect 675022 309224 675078 309233
rect 675022 309159 675078 309168
rect 674300 303742 674512 303770
rect 674576 304830 674696 304858
rect 674300 296970 674328 303742
rect 674576 302234 674604 304830
rect 674746 304736 674802 304745
rect 674746 304671 674802 304680
rect 674760 302234 674788 304671
rect 674484 302206 674604 302234
rect 674668 302206 674788 302234
rect 674300 296942 674420 296970
rect 674208 296686 674328 296714
rect 674300 286521 674328 296686
rect 674392 288946 674420 296942
rect 674484 292574 674512 302206
rect 674668 296714 674696 302206
rect 674838 302016 674894 302025
rect 674838 301951 674894 301960
rect 674576 296686 674696 296714
rect 674576 294893 674604 296686
rect 674852 295905 674880 301951
rect 674838 295896 674894 295905
rect 674838 295831 674894 295840
rect 675036 294893 675064 309159
rect 676034 308408 676090 308417
rect 676090 308366 676352 308394
rect 676034 308343 676090 308352
rect 676034 308000 676090 308009
rect 676090 307958 676260 307986
rect 676034 307935 676090 307944
rect 676232 305130 676260 307958
rect 675864 305102 676260 305130
rect 675206 303784 675262 303793
rect 675206 303719 675262 303728
rect 675220 302025 675248 303719
rect 675206 302016 675262 302025
rect 675206 301951 675262 301960
rect 675864 301594 675892 305102
rect 676324 304910 676352 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 676494 305960 676550 305969
rect 676494 305895 676550 305904
rect 676036 304904 676088 304910
rect 676036 304846 676088 304852
rect 676312 304904 676364 304910
rect 676312 304846 676364 304852
rect 676048 303793 676076 304846
rect 676034 303784 676090 303793
rect 676034 303719 676090 303728
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 674576 294865 674696 294893
rect 674668 292574 674696 294865
rect 674944 294865 675064 294893
rect 675128 301566 675892 301594
rect 674944 294545 674972 294865
rect 674930 294536 674986 294545
rect 674930 294471 674986 294480
rect 675128 294386 675156 301566
rect 676048 301481 676076 303447
rect 676508 301617 676536 305895
rect 676678 305144 676734 305153
rect 676678 305079 676734 305088
rect 676494 301608 676550 301617
rect 676494 301543 676550 301552
rect 676692 301481 676720 305079
rect 676034 301472 676090 301481
rect 676034 301407 676090 301416
rect 676678 301472 676734 301481
rect 676678 301407 676734 301416
rect 675852 298104 675904 298110
rect 678256 298081 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 675852 298046 675904 298052
rect 678242 298072 678298 298081
rect 675864 296714 675892 298046
rect 678980 298046 679032 298052
rect 678242 298007 678298 298016
rect 681016 297090 681044 307527
rect 676036 297084 676088 297090
rect 676036 297026 676088 297032
rect 681004 297084 681056 297090
rect 681004 297026 681056 297032
rect 675588 296686 675892 296714
rect 675390 296576 675446 296585
rect 675390 296511 675446 296520
rect 675404 296426 675432 296511
rect 675036 294358 675156 294386
rect 675220 296398 675432 296426
rect 675036 292777 675064 294358
rect 675022 292768 675078 292777
rect 675022 292703 675078 292712
rect 674484 292546 674604 292574
rect 674668 292546 674788 292574
rect 674576 289814 674604 292546
rect 674760 291009 674788 292546
rect 674746 291000 674802 291009
rect 674746 290935 674802 290944
rect 674576 289786 674880 289814
rect 674392 288918 674512 288946
rect 674286 286512 674342 286521
rect 674286 286447 674342 286456
rect 674484 285569 674512 288918
rect 674470 285560 674526 285569
rect 674470 285495 674526 285504
rect 674852 280154 674880 289786
rect 675220 288062 675248 296398
rect 675588 296290 675616 296686
rect 676048 296585 676076 297026
rect 676034 296576 676090 296585
rect 676034 296511 676090 296520
rect 675312 296262 675616 296290
rect 675312 291870 675340 296262
rect 675482 295896 675538 295905
rect 675482 295831 675538 295840
rect 675496 295528 675524 295831
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675482 294536 675538 294545
rect 675482 294471 675538 294480
rect 675496 294236 675524 294471
rect 675482 292768 675538 292777
rect 675482 292703 675538 292712
rect 675496 292400 675524 292703
rect 675312 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675390 291000 675446 291009
rect 675390 290935 675446 290944
rect 675404 290564 675432 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 675220 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675482 285560 675538 285569
rect 675482 285495 675538 285504
rect 675496 285056 675524 285495
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 674484 280126 674880 280154
rect 674484 265033 674512 280126
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 676034 269784 676090 269793
rect 676034 269719 676090 269728
rect 676048 268297 676076 269719
rect 676034 268288 676090 268297
rect 676034 268223 676090 268232
rect 683132 268161 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 675022 267064 675078 267073
rect 675022 266999 675078 267008
rect 674470 265024 674526 265033
rect 674470 264959 674526 264968
rect 674838 264480 674894 264489
rect 674838 264415 674894 264424
rect 674852 263809 674880 264415
rect 674838 263800 674894 263809
rect 674838 263735 674894 263744
rect 674562 263120 674618 263129
rect 674562 263055 674618 263064
rect 674378 260944 674434 260953
rect 674378 260879 674434 260888
rect 674392 253934 674420 260879
rect 674576 260834 674604 263055
rect 675036 260834 675064 266999
rect 675390 265432 675446 265441
rect 675390 265367 675446 265376
rect 675404 263129 675432 265367
rect 676494 264072 676550 264081
rect 676494 264007 676550 264016
rect 676508 263673 676536 264007
rect 676494 263664 676550 263673
rect 676494 263599 676550 263608
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 675390 263120 675446 263129
rect 675390 263055 675446 263064
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 674576 260806 674696 260834
rect 674668 258754 674696 260806
rect 674300 253906 674420 253934
rect 674484 258726 674696 258754
rect 674760 260806 675064 260834
rect 674300 246945 674328 253906
rect 674286 246936 674342 246945
rect 674286 246871 674342 246880
rect 674312 235000 674364 235006
rect 674300 234948 674312 234954
rect 674300 234942 674364 234948
rect 674300 234926 674352 234942
rect 674300 233832 674328 234926
rect 674484 234841 674512 258726
rect 674760 253934 674788 260806
rect 676232 259570 676260 262783
rect 676140 259542 676260 259570
rect 676140 255377 676168 259542
rect 675390 255368 675446 255377
rect 675390 255303 675446 255312
rect 676126 255368 676182 255377
rect 676126 255303 676182 255312
rect 674668 253906 674788 253934
rect 674470 234832 674526 234841
rect 674470 234767 674526 234776
rect 674668 234614 674696 253906
rect 675114 251832 675170 251841
rect 675114 251767 675170 251776
rect 674930 249928 674986 249937
rect 674930 249863 674986 249872
rect 674944 243085 674972 249863
rect 675128 247058 675156 251767
rect 675404 251682 675432 255303
rect 676036 252408 676088 252414
rect 676036 252350 676088 252356
rect 675852 252272 675904 252278
rect 675220 251654 675432 251682
rect 675496 252220 675852 252226
rect 675496 252214 675904 252220
rect 675496 252198 675892 252214
rect 675220 247398 675248 251654
rect 675496 251410 675524 252198
rect 676048 251841 676076 252350
rect 678256 252278 678284 263191
rect 678426 261216 678482 261225
rect 678426 261151 678482 261160
rect 678440 252414 678468 261151
rect 678428 252408 678480 252414
rect 678428 252350 678480 252356
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 676034 251832 676090 251841
rect 676034 251767 676090 251776
rect 675312 251382 675524 251410
rect 675312 250526 675340 251382
rect 675312 250498 675418 250526
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249656 675446 249665
rect 675390 249591 675446 249600
rect 675404 249220 675432 249591
rect 675220 247370 675418 247398
rect 675128 247030 675340 247058
rect 675114 246936 675170 246945
rect 675114 246871 675170 246880
rect 675128 246213 675156 246871
rect 675312 246854 675340 247030
rect 675312 246826 675418 246854
rect 675128 246185 675418 246213
rect 675298 245848 675354 245857
rect 675298 245783 675354 245792
rect 675312 245562 675340 245783
rect 675312 245534 675418 245562
rect 674944 243057 675418 243085
rect 675298 242856 675354 242865
rect 675298 242791 675354 242800
rect 675312 242533 675340 242791
rect 675312 242505 675418 242533
rect 675666 242312 675722 242321
rect 675666 242247 675722 242256
rect 675680 241876 675708 242247
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675114 238232 675170 238241
rect 675170 238190 675418 238218
rect 675114 238167 675170 238176
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 674944 237510 675340 237538
rect 675404 237524 675432 237646
rect 674944 235929 674972 237510
rect 675114 237280 675170 237289
rect 675114 237215 675170 237224
rect 675128 236382 675156 237215
rect 675128 236354 675418 236382
rect 674930 235920 674986 235929
rect 674930 235855 674986 235864
rect 676034 235240 676090 235249
rect 676034 235175 676090 235184
rect 675850 234832 675906 234841
rect 675850 234767 675906 234776
rect 674208 233804 674328 233832
rect 674576 234586 674696 234614
rect 675864 234598 675892 234767
rect 675852 234592 675904 234598
rect 674208 230194 674236 233804
rect 674576 230874 674604 234586
rect 675852 234534 675904 234540
rect 674748 234524 674800 234530
rect 674748 234466 674800 234472
rect 674760 234410 674788 234466
rect 674668 234382 674788 234410
rect 674668 231554 674696 234382
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674898 234002 674926 234262
rect 674760 233974 674926 234002
rect 674760 233322 674788 233974
rect 675236 233912 675288 233918
rect 675288 233860 675892 233866
rect 675236 233854 675892 233860
rect 675248 233850 675892 233854
rect 675248 233844 675904 233850
rect 675248 233838 675852 233844
rect 675852 233786 675904 233792
rect 675850 233608 675906 233617
rect 675850 233543 675852 233552
rect 675904 233543 675906 233552
rect 675852 233514 675904 233520
rect 674760 233294 674880 233322
rect 676048 233306 676076 235175
rect 678244 234592 678296 234598
rect 678244 234534 678296 234540
rect 677784 233844 677836 233850
rect 677784 233786 677836 233792
rect 674852 233102 674880 233294
rect 676036 233300 676088 233306
rect 676036 233242 676088 233248
rect 674840 233096 674892 233102
rect 674840 233038 674892 233044
rect 675484 232552 675536 232558
rect 675536 232500 675892 232506
rect 675484 232494 675892 232500
rect 675496 232478 675892 232494
rect 675864 232422 675892 232478
rect 675852 232416 675904 232422
rect 675852 232358 675904 232364
rect 675178 231840 675234 231849
rect 675178 231775 675180 231784
rect 675232 231775 675234 231784
rect 675180 231746 675232 231752
rect 675070 231600 675122 231606
rect 675068 231568 675070 231577
rect 675122 231568 675124 231577
rect 674668 231538 674788 231554
rect 674668 231532 674800 231538
rect 674668 231526 674748 231532
rect 675068 231503 675124 231512
rect 674748 231474 674800 231480
rect 674956 231328 675008 231334
rect 675008 231276 675892 231282
rect 674956 231270 675892 231276
rect 674968 231266 675892 231270
rect 674840 231260 674892 231266
rect 674968 231260 675904 231266
rect 674968 231254 675852 231260
rect 674840 231202 674892 231208
rect 675852 231202 675904 231208
rect 677600 231260 677652 231266
rect 677600 231202 677652 231208
rect 674730 231160 674786 231169
rect 674730 231095 674786 231104
rect 674744 230994 674772 231095
rect 674732 230988 674784 230994
rect 674732 230930 674784 230936
rect 674852 230897 674880 231202
rect 674838 230888 674894 230897
rect 674576 230846 674696 230874
rect 674668 230704 674696 230846
rect 674838 230823 674894 230832
rect 674668 230676 674788 230704
rect 674396 230648 674448 230654
rect 674300 230596 674396 230602
rect 674300 230590 674448 230596
rect 674516 230616 674572 230625
rect 674300 230574 674436 230590
rect 674300 230330 674328 230574
rect 674516 230551 674518 230560
rect 674570 230551 674572 230560
rect 674518 230522 674570 230528
rect 674394 230480 674450 230489
rect 674394 230415 674396 230424
rect 674448 230415 674450 230424
rect 674396 230386 674448 230392
rect 674300 230302 674604 230330
rect 674208 230166 674420 230194
rect 674102 226264 674158 226273
rect 674102 226199 674158 226208
rect 674102 225992 674158 226001
rect 674102 225927 674158 225936
rect 674116 225298 674144 225927
rect 674024 225270 674144 225298
rect 674024 224954 674052 225270
rect 674194 225176 674250 225185
rect 674194 225111 674250 225120
rect 674024 224926 674144 224954
rect 673918 223680 673974 223689
rect 673918 223615 673974 223624
rect 673748 221598 673868 221626
rect 673642 221504 673698 221513
rect 673642 221439 673698 221448
rect 673840 220561 673868 221598
rect 673826 220552 673882 220561
rect 673826 220487 673882 220496
rect 673550 220280 673606 220289
rect 673550 220215 673606 220224
rect 673104 215266 673316 215294
rect 673090 213752 673146 213761
rect 673090 213687 673146 213696
rect 673104 196489 673132 213687
rect 673090 196480 673146 196489
rect 673090 196415 673146 196424
rect 673288 192273 673316 215266
rect 673274 192264 673330 192273
rect 673274 192199 673330 192208
rect 672906 177848 672962 177857
rect 672906 177783 672962 177792
rect 673366 176896 673422 176905
rect 673366 176831 673422 176840
rect 673182 176080 673238 176089
rect 673182 176015 673238 176024
rect 672998 169144 673054 169153
rect 672998 169079 673054 169088
rect 673012 153105 673040 169079
rect 672998 153096 673054 153105
rect 672998 153031 673054 153040
rect 673196 131345 673224 176015
rect 673380 132161 673408 176831
rect 673564 175681 673592 220215
rect 673918 219872 673974 219881
rect 674116 219858 674144 224926
rect 673974 219830 674144 219858
rect 673918 219807 673974 219816
rect 674208 215294 674236 225111
rect 674392 215294 674420 230166
rect 674576 229945 674604 230302
rect 674562 229936 674618 229945
rect 674562 229871 674618 229880
rect 674760 222329 674788 230676
rect 676862 230616 676918 230625
rect 676862 230551 676918 230560
rect 676586 230208 676642 230217
rect 676586 230143 676642 230152
rect 675114 229936 675170 229945
rect 675170 229906 675892 229922
rect 675170 229900 675904 229906
rect 675170 229894 675852 229900
rect 675114 229871 675170 229880
rect 675852 229842 675904 229848
rect 675114 229256 675170 229265
rect 675170 229214 675892 229242
rect 675114 229191 675170 229200
rect 675864 229090 675892 229214
rect 675852 229084 675904 229090
rect 675852 229026 675904 229032
rect 676220 229084 676272 229090
rect 676220 229026 676272 229032
rect 674930 227080 674986 227089
rect 674930 227015 674986 227024
rect 674746 222320 674802 222329
rect 674746 222255 674802 222264
rect 674654 221912 674710 221921
rect 674654 221847 674710 221856
rect 674668 216322 674696 221847
rect 674944 221241 674972 227015
rect 675666 225720 675722 225729
rect 675666 225655 675722 225664
rect 675206 224496 675262 224505
rect 675206 224431 675262 224440
rect 674930 221232 674986 221241
rect 674930 221167 674986 221176
rect 675022 219056 675078 219065
rect 675022 218991 675078 219000
rect 674838 217832 674894 217841
rect 674838 217767 674894 217776
rect 674668 216294 674788 216322
rect 674562 216200 674618 216209
rect 674562 216135 674618 216144
rect 674576 215294 674604 216135
rect 674760 215294 674788 216294
rect 674116 215266 674236 215294
rect 674300 215266 674420 215294
rect 674484 215266 674604 215294
rect 674668 215266 674788 215294
rect 674116 212945 674144 215266
rect 674102 212936 674158 212945
rect 674102 212871 674158 212880
rect 674102 212120 674158 212129
rect 674102 212055 674158 212064
rect 673918 209672 673974 209681
rect 673918 209607 673974 209616
rect 673734 206952 673790 206961
rect 673734 206887 673790 206896
rect 673748 201657 673776 206887
rect 673932 203289 673960 209607
rect 673918 203280 673974 203289
rect 673918 203215 673974 203224
rect 673734 201648 673790 201657
rect 673734 201583 673790 201592
rect 673550 175672 673606 175681
rect 673550 175607 673606 175616
rect 673918 168736 673974 168745
rect 673918 168671 673974 168680
rect 673932 151065 673960 168671
rect 673918 151056 673974 151065
rect 673918 150991 673974 151000
rect 673366 132152 673422 132161
rect 673366 132087 673422 132096
rect 673182 131336 673238 131345
rect 673182 131271 673238 131280
rect 674116 128217 674144 212055
rect 674300 179489 674328 215266
rect 674484 201929 674512 215266
rect 674470 201920 674526 201929
rect 674470 201855 674526 201864
rect 674286 179480 674342 179489
rect 674286 179415 674342 179424
rect 674668 177313 674696 215266
rect 674852 202209 674880 217767
rect 675036 204049 675064 218991
rect 675220 214577 675248 224431
rect 675390 224224 675446 224233
rect 675390 224159 675446 224168
rect 675404 216889 675432 224159
rect 675680 217569 675708 225655
rect 675850 218376 675906 218385
rect 676232 218362 676260 229026
rect 676600 224954 676628 230143
rect 675906 218334 676260 218362
rect 676324 224926 676628 224954
rect 675850 218311 675906 218320
rect 676324 218226 676352 224926
rect 676232 218198 676352 218226
rect 675666 217560 675722 217569
rect 675666 217495 675722 217504
rect 675390 216880 675446 216889
rect 675390 216815 675446 216824
rect 675390 216608 675446 216617
rect 675390 216543 675446 216552
rect 675206 214568 675262 214577
rect 675206 214503 675262 214512
rect 675404 210474 675432 216543
rect 676232 215294 676260 218198
rect 676404 218136 676456 218142
rect 676404 218078 676456 218084
rect 675864 215266 676260 215294
rect 675666 214568 675722 214577
rect 675666 214503 675722 214512
rect 675680 211449 675708 214503
rect 675666 211440 675722 211449
rect 675666 211375 675722 211384
rect 675128 210446 675432 210474
rect 675128 204694 675156 210446
rect 675864 207233 675892 215266
rect 676220 215144 676272 215150
rect 676034 215112 676090 215121
rect 676090 215092 676220 215098
rect 676090 215086 676272 215092
rect 676090 215070 676260 215086
rect 676034 215047 676090 215056
rect 676034 213480 676090 213489
rect 676416 213466 676444 218078
rect 676680 217864 676732 217870
rect 676680 217806 676732 217812
rect 676090 213438 676444 213466
rect 676034 213415 676090 213424
rect 676220 213240 676272 213246
rect 676034 213208 676090 213217
rect 676090 213188 676220 213194
rect 676090 213182 676272 213188
rect 676090 213166 676260 213182
rect 676034 213143 676090 213152
rect 676692 209681 676720 217806
rect 676876 213246 676904 230551
rect 677232 229900 677284 229906
rect 677232 229842 677284 229848
rect 677046 228576 677102 228585
rect 677046 228511 677102 228520
rect 677060 217870 677088 228511
rect 677048 217864 677100 217870
rect 677048 217806 677100 217812
rect 677244 215150 677272 229842
rect 677612 218142 677640 231202
rect 677600 218136 677652 218142
rect 677600 218078 677652 218084
rect 677232 215144 677284 215150
rect 677232 215086 677284 215092
rect 676864 213240 676916 213246
rect 676864 213182 676916 213188
rect 676678 209672 676734 209681
rect 676678 209607 676734 209616
rect 675850 207224 675906 207233
rect 675850 207159 675906 207168
rect 677796 206961 677824 233786
rect 678256 220697 678284 234534
rect 683210 234152 683266 234161
rect 683210 234087 683266 234096
rect 678428 233300 678480 233306
rect 678428 233242 678480 233248
rect 678440 221513 678468 233242
rect 679256 232416 679308 232422
rect 679256 232358 679308 232364
rect 679268 223825 679296 232358
rect 679254 223816 679310 223825
rect 679254 223751 679310 223760
rect 683224 222737 683252 234087
rect 683670 233880 683726 233889
rect 683670 233815 683726 233824
rect 683488 233572 683540 233578
rect 683488 233514 683540 233520
rect 683210 222728 683266 222737
rect 683210 222663 683266 222672
rect 678426 221504 678482 221513
rect 678426 221439 678482 221448
rect 678242 220688 678298 220697
rect 678242 220623 678298 220632
rect 683500 219881 683528 233514
rect 683684 223145 683712 233815
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683670 223136 683726 223145
rect 683670 223071 683726 223080
rect 683486 219872 683542 219881
rect 683486 219807 683542 219816
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 677782 206952 677838 206961
rect 677782 206887 677838 206896
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675128 204666 675418 204694
rect 675036 204021 675418 204049
rect 674852 202181 675418 202209
rect 675390 201920 675446 201929
rect 675390 201855 675446 201864
rect 675404 201620 675432 201855
rect 675390 201376 675446 201385
rect 675390 201311 675446 201320
rect 674838 201104 674894 201113
rect 674838 201039 674894 201048
rect 674852 197577 674880 201039
rect 675404 201008 675432 201311
rect 675758 200832 675814 200841
rect 675758 200767 675814 200776
rect 675772 200328 675800 200767
rect 675390 198384 675446 198393
rect 675390 198319 675446 198328
rect 675404 197880 675432 198319
rect 674838 197568 674894 197577
rect 674838 197503 674894 197512
rect 675482 197568 675538 197577
rect 675482 197503 675538 197512
rect 675496 197336 675524 197503
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675390 196480 675446 196489
rect 675390 196415 675446 196424
rect 675404 196044 675432 196415
rect 675666 195256 675722 195265
rect 675666 195191 675722 195200
rect 675680 194820 675708 195191
rect 675666 193216 675722 193225
rect 675666 193151 675722 193160
rect 675680 192984 675708 193151
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190369 675340 191950
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675298 190360 675354 190369
rect 675298 190295 675354 190304
rect 683118 186960 683174 186969
rect 683118 186895 683174 186904
rect 676494 181384 676550 181393
rect 676494 181319 676550 181328
rect 676034 178120 676090 178129
rect 676508 178106 676536 181319
rect 683132 178809 683160 186895
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 178800 683174 178809
rect 683118 178735 683174 178744
rect 676090 178078 676536 178106
rect 676034 178055 676090 178064
rect 674654 177304 674710 177313
rect 674654 177239 674710 177248
rect 674654 175264 674710 175273
rect 674654 175199 674710 175208
rect 674378 174448 674434 174457
rect 674378 174383 674434 174392
rect 674392 129713 674420 174383
rect 674668 130529 674696 175199
rect 681002 173224 681058 173233
rect 681002 173159 681058 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674852 157593 674880 172751
rect 678242 171592 678298 171601
rect 678242 171527 678298 171536
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 676048 165617 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162858 678284 171527
rect 679622 171184 679678 171193
rect 679622 171119 679678 171128
rect 675852 162852 675904 162858
rect 675852 162794 675904 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675864 161945 675892 162794
rect 679636 162654 679664 171119
rect 676036 162648 676088 162654
rect 676036 162590 676088 162596
rect 679624 162648 679676 162654
rect 679624 162590 679676 162596
rect 675206 161936 675262 161945
rect 675206 161871 675262 161880
rect 675850 161936 675906 161945
rect 675850 161871 675906 161880
rect 675220 159678 675248 161871
rect 675852 161764 675904 161770
rect 675852 161706 675904 161712
rect 675864 161242 675892 161706
rect 676048 161401 676076 162590
rect 681016 161770 681044 173159
rect 681004 161764 681056 161770
rect 681004 161706 681056 161712
rect 676034 161392 676090 161401
rect 676034 161327 676090 161336
rect 675312 161214 675892 161242
rect 675312 160290 675340 161214
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 675758 159488 675814 159497
rect 675758 159423 675814 159432
rect 675772 159052 675800 159423
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675574 157040 675630 157049
rect 675574 156975 675630 156984
rect 675588 156643 675616 156975
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675404 154986 675432 155380
rect 675312 154958 675432 154986
rect 675114 153096 675170 153105
rect 675114 153031 675170 153040
rect 675128 152334 675156 153031
rect 675312 152697 675340 154958
rect 675758 153096 675814 153105
rect 675758 153031 675814 153040
rect 675772 152864 675800 153031
rect 675298 152688 675354 152697
rect 675298 152623 675354 152632
rect 675128 152306 675418 152334
rect 675114 151736 675170 151745
rect 675170 151680 675418 151689
rect 675114 151671 675418 151680
rect 675128 151661 675418 151671
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675758 150376 675814 150385
rect 675758 150311 675814 150320
rect 675772 149835 675800 150311
rect 675298 149016 675354 149025
rect 675298 148951 675354 148960
rect 675312 146690 675340 148951
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 683132 132705 683160 135895
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674654 130520 674710 130529
rect 674654 130455 674710 130464
rect 675942 130112 675998 130121
rect 675942 130047 675998 130056
rect 674378 129704 674434 129713
rect 674378 129639 674434 129648
rect 674470 129296 674526 129305
rect 674470 129231 674526 129240
rect 674286 128344 674342 128353
rect 674286 128279 674342 128288
rect 674102 128208 674158 128217
rect 674102 128143 674158 128152
rect 672998 126032 673054 126041
rect 672998 125967 673054 125976
rect 672722 123992 672778 124001
rect 672722 123927 672778 123936
rect 672538 123720 672594 123729
rect 672538 123655 672594 123664
rect 672354 123176 672410 123185
rect 672354 123111 672410 123120
rect 672368 120193 672396 123111
rect 672354 120184 672410 120193
rect 672354 120119 672410 120128
rect 671710 115832 671766 115841
rect 671710 115767 671766 115776
rect 671526 107672 671582 107681
rect 671526 107607 671582 107616
rect 672552 106321 672580 123655
rect 672722 121408 672778 121417
rect 672722 121343 672778 121352
rect 672736 110945 672764 121343
rect 673012 111489 673040 125967
rect 674102 125216 674158 125225
rect 674102 125151 674158 125160
rect 673182 124400 673238 124409
rect 673182 124335 673238 124344
rect 672998 111480 673054 111489
rect 672998 111415 673054 111424
rect 672722 110936 672778 110945
rect 672722 110871 672778 110880
rect 673196 110401 673224 124335
rect 673366 123584 673422 123593
rect 673366 123519 673422 123528
rect 673182 110392 673238 110401
rect 673182 110327 673238 110336
rect 672538 106312 672594 106321
rect 672538 106247 672594 106256
rect 670700 106208 670752 106214
rect 670700 106150 670752 106156
rect 673380 105641 673408 123519
rect 673366 105632 673422 105641
rect 673366 105567 673422 105576
rect 674116 104689 674144 125151
rect 674102 104680 674158 104689
rect 674102 104615 674158 104624
rect 668306 104408 668362 104417
rect 668306 104343 668362 104352
rect 668032 100156 668084 100162
rect 668032 100098 668084 100104
rect 668320 92546 668348 104343
rect 674300 102241 674328 128279
rect 674484 111897 674512 129231
rect 675956 128353 675984 130047
rect 675942 128344 675998 128353
rect 675942 128279 675998 128288
rect 682382 127800 682438 127809
rect 682382 127735 682438 127744
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 125624 674710 125633
rect 674654 125559 674710 125568
rect 674470 111888 674526 111897
rect 674470 111823 674526 111832
rect 674668 110786 674696 125559
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 682396 117298 682424 127735
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 682384 117292 682436 117298
rect 682384 117234 682436 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 675114 111480 675170 111489
rect 675170 111438 675418 111466
rect 675114 111415 675170 111424
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 674668 110758 675340 110786
rect 675404 110772 675432 110894
rect 675114 110392 675170 110401
rect 675114 110327 675170 110336
rect 675128 110174 675156 110327
rect 675128 110146 675418 110174
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675772 106185 675800 106488
rect 675758 106176 675814 106185
rect 675758 106111 675814 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 675128 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 105641 675156 105794
rect 675114 105632 675170 105641
rect 675114 105567 675170 105576
rect 675114 104680 675170 104689
rect 675170 104638 675340 104666
rect 675114 104615 675170 104624
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 668490 102232 668546 102241
rect 668490 102167 668546 102176
rect 674286 102232 674342 102241
rect 674286 102167 674342 102176
rect 668504 100026 668532 102167
rect 675680 102136 675708 102575
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668492 100020 668544 100026
rect 668492 99962 668544 99968
rect 668308 92540 668360 92546
rect 668308 92482 668360 92488
rect 666572 84166 666692 84194
rect 664444 62076 664496 62082
rect 664444 62018 664496 62024
rect 663800 58676 663852 58682
rect 663800 58618 663852 58624
rect 663812 47841 663840 58618
rect 666572 57934 666600 84166
rect 666560 57928 666612 57934
rect 666560 57870 666612 57876
rect 663984 55888 664036 55894
rect 663984 55830 664036 55836
rect 663996 48521 664024 55830
rect 663982 48512 664038 48521
rect 663982 48447 664038 48456
rect 663798 47832 663854 47841
rect 663798 47767 663854 47776
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464344 42764 464396 42770
rect 464344 42706 464396 42712
rect 463976 42628 464028 42634
rect 463976 42570 464028 42576
rect 465828 42500 465856 43143
rect 463712 42350 464036 42378
rect 461122 42256 461178 42265
rect 461122 42191 461178 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42364 518848 42735
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40488 141754 40497
rect 141698 40423 141754 40432
rect 142618 40488 142674 40497
rect 142618 40423 142674 40432
rect 141712 39984 141740 40423
<< via2 >>
rect 431682 1007140 431738 1007176
rect 431682 1007120 431684 1007140
rect 431684 1007120 431736 1007140
rect 431736 1007120 431738 1007140
rect 428002 1007004 428058 1007040
rect 428002 1006984 428004 1007004
rect 428004 1006984 428056 1007004
rect 428056 1006984 428058 1007004
rect 359738 1006884 359740 1006904
rect 359740 1006884 359792 1006904
rect 359792 1006884 359794 1006904
rect 359738 1006848 359794 1006884
rect 359370 1006748 359372 1006768
rect 359372 1006748 359424 1006768
rect 359424 1006748 359426 1006768
rect 101126 1006460 101182 1006496
rect 101126 1006440 101128 1006460
rect 101128 1006440 101180 1006460
rect 101180 1006440 101182 1006460
rect 80426 995696 80482 995752
rect 85946 995696 86002 995752
rect 86590 995696 86646 995752
rect 87878 995696 87934 995752
rect 77022 995016 77078 995072
rect 81990 994744 82046 994800
rect 88982 995424 89038 995480
rect 90270 995424 90326 995480
rect 92938 996920 92994 996976
rect 92570 995424 92626 995480
rect 85302 994472 85358 994528
rect 93490 997192 93546 997248
rect 93582 996920 93638 996976
rect 94502 996920 94558 996976
rect 93306 995968 93362 996024
rect 101954 1006324 102010 1006360
rect 101954 1006304 101956 1006324
rect 101956 1006304 102008 1006324
rect 102008 1006304 102010 1006324
rect 108486 1006324 108542 1006360
rect 108486 1006304 108488 1006324
rect 108488 1006304 108540 1006324
rect 108540 1006304 108542 1006324
rect 99470 1006188 99526 1006224
rect 99470 1006168 99472 1006188
rect 99472 1006168 99524 1006188
rect 99524 1006168 99526 1006188
rect 104806 1006188 104862 1006224
rect 104806 1006168 104808 1006188
rect 104808 1006168 104860 1006188
rect 104860 1006168 104862 1006188
rect 106830 1006188 106886 1006224
rect 106830 1006168 106832 1006188
rect 106832 1006168 106884 1006188
rect 106884 1006168 106886 1006188
rect 98274 1006052 98330 1006088
rect 98274 1006032 98276 1006052
rect 98276 1006032 98328 1006052
rect 98328 1006032 98330 1006052
rect 94686 995968 94742 996024
rect 93582 994472 93638 994528
rect 84474 994200 84530 994256
rect 42154 967544 42210 967600
rect 42614 967544 42670 967600
rect 41786 967136 41842 967192
rect 42154 967136 42210 967192
rect 42430 964688 42486 964744
rect 42430 963872 42486 963928
rect 42430 963328 42486 963384
rect 42430 963056 42486 963112
rect 41786 962104 41842 962160
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42430 958704 42486 958760
rect 41786 957752 41842 957808
rect 41786 955440 41842 955496
rect 41786 954624 41842 954680
rect 41786 954352 41842 954408
rect 35162 952856 35218 952912
rect 31758 946600 31814 946656
rect 28722 942656 28778 942712
rect 33782 938168 33838 938224
rect 37922 952448 37978 952504
rect 35806 943064 35862 943120
rect 35806 941840 35862 941896
rect 35806 940208 35862 940264
rect 36542 938984 36598 939040
rect 39302 952176 39358 952232
rect 37922 938576 37978 938632
rect 35162 937760 35218 937816
rect 40038 951632 40094 951688
rect 39762 943744 39818 943800
rect 39302 937352 39358 937408
rect 39762 935720 39818 935776
rect 40038 934496 40094 934552
rect 42062 940616 42118 940672
rect 42062 939800 42118 939856
rect 41786 935584 41842 935640
rect 43442 967136 43498 967192
rect 43442 964688 43498 964744
rect 43258 963872 43314 963928
rect 43074 963328 43130 963384
rect 42798 936944 42854 937000
rect 43074 934904 43130 934960
rect 44270 963056 44326 963112
rect 43442 935312 43498 935368
rect 44454 958704 44510 958760
rect 46202 946600 46258 946656
rect 45558 943472 45614 943528
rect 44822 941432 44878 941488
rect 44638 941024 44694 941080
rect 44454 936264 44510 936320
rect 44270 934088 44326 934144
rect 43258 933680 43314 933736
rect 43626 933272 43682 933328
rect 42338 932864 42394 932920
rect 41602 911920 41658 911976
rect 41418 911648 41474 911704
rect 42936 892472 42992 892528
rect 43074 892254 43130 892256
rect 43074 892202 43076 892254
rect 43076 892202 43128 892254
rect 43128 892202 43130 892254
rect 43074 892200 43130 892202
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 35806 817264 35862 817320
rect 35806 816448 35862 816504
rect 42062 884584 42118 884640
rect 35806 814816 35862 814872
rect 41326 812776 41382 812832
rect 40958 812368 41014 812424
rect 35162 811552 35218 811608
rect 35898 811144 35954 811200
rect 40774 808288 40830 808344
rect 40590 805296 40646 805352
rect 40774 805024 40830 805080
rect 41142 811960 41198 812016
rect 41970 809104 42026 809160
rect 41786 808696 41842 808752
rect 42154 806656 42210 806712
rect 41970 805432 42026 805488
rect 41142 804752 41198 804808
rect 40958 804480 41014 804536
rect 41694 802460 41750 802496
rect 41694 802440 41696 802460
rect 41696 802440 41748 802460
rect 41748 802440 41750 802460
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 43074 810736 43130 810792
rect 42798 809920 42854 809976
rect 42522 802440 42578 802496
rect 42522 799176 42578 799232
rect 42430 796728 42486 796784
rect 42154 796184 42210 796240
rect 42430 794280 42486 794336
rect 41786 794144 41842 794200
rect 42246 792512 42302 792568
rect 42890 790744 42946 790800
rect 42522 788704 42578 788760
rect 41786 788568 41842 788624
rect 42706 788568 42762 788624
rect 42430 788296 42486 788352
rect 42246 788160 42302 788216
rect 43442 809512 43498 809568
rect 43258 807472 43314 807528
rect 43074 788296 43130 788352
rect 35806 773472 35862 773528
rect 35346 769392 35402 769448
rect 35530 769004 35586 769040
rect 35530 768984 35532 769004
rect 35532 768984 35584 769004
rect 35584 768984 35586 769004
rect 35806 768984 35862 769040
rect 31022 768168 31078 768224
rect 35530 767760 35586 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 37094 763292 37150 763328
rect 37094 763272 37096 763292
rect 37096 763272 37148 763292
rect 37148 763272 37150 763292
rect 41326 765720 41382 765776
rect 40038 764496 40094 764552
rect 36542 757696 36598 757752
rect 39302 757968 39358 758024
rect 42890 766264 42946 766320
rect 42706 765720 42762 765776
rect 41694 758784 41750 758840
rect 42246 758784 42302 758840
rect 41694 758276 41696 758296
rect 41696 758276 41748 758296
rect 41748 758276 41750 758296
rect 41694 758240 41750 758276
rect 42430 758240 42486 758296
rect 42246 757968 42302 758024
rect 39118 757288 39174 757344
rect 41786 757016 41842 757072
rect 41878 756608 41934 756664
rect 42430 754432 42486 754488
rect 41970 754024 42026 754080
rect 42246 753888 42302 753944
rect 42246 752120 42302 752176
rect 42062 751712 42118 751768
rect 41786 751032 41842 751088
rect 42246 749400 42302 749456
rect 42430 749264 42486 749320
rect 43074 763000 43130 763056
rect 42890 753888 42946 753944
rect 42890 753480 42946 753536
rect 42890 751712 42946 751768
rect 42430 745048 42486 745104
rect 42246 744776 42302 744832
rect 41786 743688 41842 743744
rect 42706 743008 42762 743064
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 33782 725192 33838 725248
rect 33046 723968 33102 724024
rect 31666 723152 31722 723208
rect 36542 724784 36598 724840
rect 40682 724376 40738 724432
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41878 722336 41934 722392
rect 41694 719616 41750 719672
rect 42154 720296 42210 720352
rect 41878 718528 41934 718584
rect 41142 715808 41198 715864
rect 41694 715828 41750 715864
rect 41694 715808 41696 715828
rect 41696 715808 41748 715828
rect 41748 715808 41750 715828
rect 40682 714720 40738 714776
rect 41970 714584 42026 714640
rect 42522 719616 42578 719672
rect 42706 715808 42762 715864
rect 42246 711048 42302 711104
rect 41970 709824 42026 709880
rect 42246 709144 42302 709200
rect 41786 708464 41842 708520
rect 41786 706696 41842 706752
rect 42154 706696 42210 706752
rect 42246 705472 42302 705528
rect 41786 704248 41842 704304
rect 42062 703024 42118 703080
rect 42890 715536 42946 715592
rect 42706 706696 42762 706752
rect 42706 703024 42762 703080
rect 42338 701800 42394 701856
rect 41786 700440 41842 700496
rect 42614 701528 42670 701584
rect 41694 697856 41750 697912
rect 35622 691328 35678 691384
rect 41326 687656 41382 687712
rect 35622 687248 35678 687304
rect 41326 683188 41382 683224
rect 41326 683168 41328 683188
rect 41328 683168 41380 683188
rect 41380 683168 41382 683188
rect 41326 682352 41382 682408
rect 40038 681944 40094 682000
rect 36726 681536 36782 681592
rect 36542 681128 36598 681184
rect 35162 680720 35218 680776
rect 41694 681844 41696 681864
rect 41696 681844 41748 681864
rect 41748 681844 41750 681864
rect 41694 681808 41750 681844
rect 42614 681808 42670 681864
rect 42798 679904 42854 679960
rect 41694 677320 41750 677376
rect 39946 677048 40002 677104
rect 40130 671200 40186 671256
rect 36542 670928 36598 670984
rect 42706 677320 42762 677376
rect 42246 667800 42302 667856
rect 42430 667528 42486 667584
rect 42246 667120 42302 667176
rect 42246 666032 42302 666088
rect 41786 665352 41842 665408
rect 41970 663992 42026 664048
rect 42154 663448 42210 663504
rect 42246 662904 42302 662960
rect 42890 667120 42946 667176
rect 42246 662632 42302 662688
rect 42890 663448 42946 663504
rect 42614 658552 42670 658608
rect 42430 658280 42486 658336
rect 41786 657192 41842 657248
rect 35806 646720 35862 646776
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35622 639784 35678 639840
rect 35806 639376 35862 639432
rect 35806 638560 35862 638616
rect 40038 638560 40094 638616
rect 32402 638152 32458 638208
rect 35806 636520 35862 636576
rect 41786 638152 41842 638208
rect 41786 637540 41842 637596
rect 42246 633800 42302 633856
rect 42246 624960 42302 625016
rect 42798 635704 42854 635760
rect 42062 624416 42118 624472
rect 41786 622104 41842 622160
rect 42154 621560 42210 621616
rect 42062 620744 42118 620800
rect 41970 620200 42026 620256
rect 42430 619248 42486 619304
rect 42614 618976 42670 619032
rect 42246 615984 42302 616040
rect 41786 615712 41842 615768
rect 42890 615576 42946 615632
rect 41786 612720 41842 612776
rect 43442 796184 43498 796240
rect 43442 633392 43498 633448
rect 43074 612312 43130 612368
rect 43810 932048 43866 932104
rect 44086 892764 44142 892800
rect 44086 892744 44088 892764
rect 44088 892744 44140 892764
rect 44140 892744 44142 892764
rect 44086 891948 44142 891984
rect 44086 891928 44088 891948
rect 44088 891928 44140 891948
rect 44140 891928 44142 891948
rect 44454 816040 44510 816096
rect 44270 810328 44326 810384
rect 43994 806248 44050 806304
rect 44270 790744 44326 790800
rect 48962 940072 49018 940128
rect 51722 942248 51778 942304
rect 50342 939800 50398 939856
rect 47582 891928 47638 891984
rect 44638 815632 44694 815688
rect 45006 815224 45062 815280
rect 44638 814408 44694 814464
rect 44454 773200 44510 773256
rect 44454 772792 44510 772848
rect 44270 771976 44326 772032
rect 44822 813592 44878 813648
rect 44638 771568 44694 771624
rect 45190 807880 45246 807936
rect 45190 796728 45246 796784
rect 45006 772384 45062 772440
rect 44822 771160 44878 771216
rect 44638 770752 44694 770808
rect 44638 770344 44694 770400
rect 44454 730088 44510 730144
rect 44270 729272 44326 729328
rect 44454 728864 44510 728920
rect 44270 728048 44326 728104
rect 45098 766672 45154 766728
rect 45282 764768 45338 764824
rect 46018 764224 46074 764280
rect 45282 753480 45338 753536
rect 45098 749264 45154 749320
rect 45006 729680 45062 729736
rect 44822 728456 44878 728512
rect 44638 727640 44694 727696
rect 44638 727368 44694 727424
rect 44454 686024 44510 686080
rect 44270 685208 44326 685264
rect 44362 684800 44418 684856
rect 44178 679496 44234 679552
rect 44178 666576 44234 666632
rect 44822 722744 44878 722800
rect 44822 709416 44878 709472
rect 45190 723560 45246 723616
rect 45190 705472 45246 705528
rect 45006 686840 45062 686896
rect 44822 686432 44878 686488
rect 44638 684392 44694 684448
rect 44546 680312 44602 680368
rect 44546 662904 44602 662960
rect 45006 685616 45062 685672
rect 44822 643592 44878 643648
rect 44638 643320 44694 643376
rect 44362 642232 44418 642288
rect 44178 635296 44234 635352
rect 44362 634480 44418 634536
rect 44178 620744 44234 620800
rect 44178 614080 44234 614136
rect 43718 612332 43774 612368
rect 43718 612312 43720 612332
rect 43720 612312 43772 612332
rect 43772 612312 43774 612332
rect 44270 610972 44326 611008
rect 44270 610952 44272 610972
rect 44272 610952 44324 610972
rect 44324 610952 44326 610972
rect 45374 683984 45430 684040
rect 45006 643048 45062 643104
rect 44822 642504 44878 642560
rect 44638 600480 44694 600536
rect 44638 600072 44694 600128
rect 42982 596944 43038 597000
rect 42430 596808 42486 596864
rect 41234 595992 41290 596048
rect 33782 595584 33838 595640
rect 32402 594768 32458 594824
rect 36542 595176 36598 595232
rect 32402 585656 32458 585712
rect 37922 594360 37978 594416
rect 40682 593544 40738 593600
rect 39946 590688 40002 590744
rect 40498 589636 40500 589656
rect 40500 589636 40552 589656
rect 40552 589636 40554 589656
rect 40498 589600 40554 589636
rect 39946 585928 40002 585984
rect 39670 585248 39726 585304
rect 40222 584976 40278 585032
rect 42062 593136 42118 593192
rect 41878 592728 41934 592784
rect 42062 589328 42118 589384
rect 41510 585928 41566 585984
rect 42246 584976 42302 585032
rect 40682 584568 40738 584624
rect 41418 584568 41474 584624
rect 41786 582528 41842 582584
rect 42798 593952 42854 594008
rect 42706 585928 42762 585984
rect 42246 581440 42302 581496
rect 42430 580624 42486 580680
rect 41786 580216 41842 580272
rect 42062 580080 42118 580136
rect 42062 578856 42118 578912
rect 42246 578312 42302 578368
rect 42246 577768 42302 577824
rect 42246 576816 42302 576872
rect 41970 576544 42026 576600
rect 42154 574096 42210 574152
rect 44454 591912 44510 591968
rect 43442 590280 43498 590336
rect 42890 574096 42946 574152
rect 41970 573144 42026 573200
rect 42430 571648 42486 571704
rect 42246 571376 42302 571432
rect 42062 570968 42118 571024
rect 42246 569064 42302 569120
rect 35806 558048 35862 558104
rect 42062 558456 42118 558512
rect 42062 557504 42118 557560
rect 35806 554804 35862 554840
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35622 553968 35678 554024
rect 35806 553580 35862 553616
rect 35806 553560 35808 553580
rect 35808 553560 35860 553580
rect 35860 553560 35862 553580
rect 40866 553152 40922 553208
rect 33782 551928 33838 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41234 551112 41290 551168
rect 41234 549480 41290 549536
rect 41326 548256 41382 548312
rect 41326 546352 41382 546408
rect 41786 553152 41842 553208
rect 43166 552336 43222 552392
rect 42062 550296 42118 550352
rect 41878 549888 41934 549944
rect 41694 549364 41750 549400
rect 41694 549344 41696 549364
rect 41696 549344 41748 549364
rect 41748 549344 41750 549364
rect 41694 547712 41750 547768
rect 42062 545672 42118 545728
rect 41878 545400 41934 545456
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42614 540232 42670 540288
rect 42246 538192 42302 538248
rect 42062 537920 42118 537976
rect 42614 537920 42670 537976
rect 42154 535200 42210 535256
rect 41786 534928 41842 534984
rect 42154 534384 42210 534440
rect 42154 533840 42210 533896
rect 42246 533160 42302 533216
rect 42982 549344 43038 549400
rect 43166 533840 43222 533896
rect 42982 533160 43038 533216
rect 42522 532752 42578 532808
rect 42154 530032 42210 530088
rect 41878 529352 41934 529408
rect 42522 530576 42578 530632
rect 42706 530032 42762 530088
rect 42614 529624 42670 529680
rect 42890 529080 42946 529136
rect 40958 425992 41014 426048
rect 40774 425584 40830 425640
rect 36542 424360 36598 424416
rect 40498 421912 40554 421968
rect 41326 423952 41382 424008
rect 41786 423000 41842 423056
rect 41786 422184 41842 422240
rect 41786 421504 41842 421560
rect 40774 418784 40830 418840
rect 40498 418648 40554 418704
rect 41786 418240 41842 418296
rect 42154 422728 42210 422784
rect 42522 419872 42578 419928
rect 42154 418512 42210 418568
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42430 407088 42486 407144
rect 42430 406816 42486 406872
rect 41786 406272 41842 406328
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 42430 399744 42486 399800
rect 43074 422184 43130 422240
rect 43258 421096 43314 421152
rect 43258 407768 43314 407824
rect 43074 402872 43130 402928
rect 41786 398792 41842 398848
rect 41142 387116 41198 387152
rect 41142 387096 41144 387116
rect 41144 387096 41196 387116
rect 41196 387096 41198 387116
rect 41878 386960 41934 387016
rect 41326 386688 41382 386744
rect 41510 386688 41566 386744
rect 41142 383016 41198 383072
rect 41326 382608 41382 382664
rect 40038 382200 40094 382256
rect 41694 382236 41696 382256
rect 41696 382236 41748 382256
rect 41748 382236 41750 382256
rect 41694 382200 41750 382236
rect 35806 379344 35862 379400
rect 40774 381384 40830 381440
rect 41326 380976 41382 381032
rect 40774 378528 40830 378584
rect 42798 382200 42854 382256
rect 41694 379344 41750 379400
rect 41326 377712 41382 377768
rect 42338 377712 42394 377768
rect 35806 376488 35862 376544
rect 40038 376488 40094 376544
rect 28906 376080 28962 376136
rect 39486 375672 39542 375728
rect 41694 371884 41750 371920
rect 41694 371864 41696 371884
rect 41696 371864 41748 371884
rect 41748 371864 41750 371884
rect 41786 368600 41842 368656
rect 42430 366968 42486 367024
rect 42430 365744 42486 365800
rect 41786 364248 41842 364304
rect 41786 363568 41842 363624
rect 41786 362888 41842 362944
rect 42430 361528 42486 361584
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 41786 358672 41842 358728
rect 42430 357312 42486 357368
rect 44454 578856 44510 578912
rect 45650 677864 45706 677920
rect 45374 641416 45430 641472
rect 45190 641144 45246 641200
rect 45006 640872 45062 640928
rect 44822 599664 44878 599720
rect 44822 599256 44878 599312
rect 44638 557232 44694 557288
rect 45834 637744 45890 637800
rect 45834 615576 45890 615632
rect 46202 756336 46258 756392
rect 46938 721112 46994 721168
rect 45650 610952 45706 611008
rect 46386 636928 46442 636984
rect 46386 619248 46442 619304
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47858 719888 47914 719944
rect 47582 712136 47638 712192
rect 47674 676640 47730 676696
rect 47214 638152 47270 638208
rect 47398 636384 47454 636440
rect 47398 621560 47454 621616
rect 47214 618976 47270 619032
rect 46202 600888 46258 600944
rect 45190 598848 45246 598904
rect 45190 598440 45246 598496
rect 45006 598032 45062 598088
rect 97262 994744 97318 994800
rect 100298 1002652 100354 1002688
rect 100298 1002632 100300 1002652
rect 100300 1002632 100352 1002652
rect 100352 1002632 100354 1002652
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 99102 1002108 99158 1002144
rect 99102 1002088 99104 1002108
rect 99104 1002088 99156 1002108
rect 99156 1002088 99158 1002108
rect 98826 995696 98882 995752
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 101126 1001972 101182 1002008
rect 101126 1001952 101128 1001972
rect 101128 1001952 101180 1001972
rect 101180 1001952 101182 1001972
rect 102322 1002788 102378 1002824
rect 102322 1002768 102324 1002788
rect 102324 1002768 102376 1002788
rect 102376 1002768 102378 1002788
rect 101954 1002244 102010 1002280
rect 101954 1002224 101956 1002244
rect 101956 1002224 102008 1002244
rect 102008 1002224 102010 1002244
rect 101402 995016 101458 995072
rect 100022 994472 100078 994528
rect 103978 1006052 104034 1006088
rect 103978 1006032 103980 1006052
rect 103980 1006032 104032 1006052
rect 104032 1006032 104034 1006052
rect 106002 1006052 106058 1006088
rect 106002 1006032 106004 1006052
rect 106004 1006032 106056 1006052
rect 106056 1006032 106058 1006052
rect 108854 1005252 108856 1005272
rect 108856 1005252 108908 1005272
rect 108908 1005252 108910 1005272
rect 108854 1005216 108910 1005252
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 103150 1002516 103206 1002552
rect 103150 1002496 103152 1002516
rect 103152 1002496 103204 1002516
rect 103204 1002496 103206 1002516
rect 105634 1002244 105690 1002280
rect 105634 1002224 105636 1002244
rect 105636 1002224 105688 1002244
rect 105688 1002224 105690 1002244
rect 103150 1002108 103206 1002144
rect 103150 1002088 103152 1002108
rect 103152 1002088 103204 1002108
rect 103204 1002088 103206 1002108
rect 103978 1002108 104034 1002144
rect 103978 1002088 103980 1002108
rect 103980 1002088 104032 1002108
rect 104032 1002088 104034 1002108
rect 104806 1001952 104862 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 107658 1002380 107714 1002416
rect 107658 1002360 107660 1002380
rect 107660 1002360 107712 1002380
rect 107712 1002360 107714 1002380
rect 108026 1002244 108082 1002280
rect 108026 1002224 108028 1002244
rect 108028 1002224 108080 1002244
rect 108080 1002224 108082 1002244
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 117134 997192 117190 997248
rect 116214 996920 116270 996976
rect 143998 1000592 144054 1000648
rect 143722 997192 143778 997248
rect 126242 996104 126298 996160
rect 138018 995696 138074 995752
rect 141790 995696 141846 995752
rect 144182 996920 144238 996976
rect 124862 995016 124918 995072
rect 133418 994744 133474 994800
rect 133142 994472 133198 994528
rect 137374 995424 137430 995480
rect 140502 995288 140558 995344
rect 138754 994744 138810 994800
rect 138938 994744 138994 994800
rect 135902 994200 135958 994256
rect 143998 995696 144054 995752
rect 140594 994472 140650 994528
rect 140778 994472 140834 994528
rect 138754 993928 138810 993984
rect 144182 994744 144238 994800
rect 144734 995968 144790 996024
rect 144918 995288 144974 995344
rect 144550 994472 144606 994528
rect 359370 1006712 359426 1006748
rect 152094 1006596 152150 1006632
rect 152094 1006576 152096 1006596
rect 152096 1006576 152148 1006596
rect 152148 1006576 152150 1006596
rect 157430 1006596 157486 1006632
rect 360566 1006612 360568 1006632
rect 360568 1006612 360620 1006632
rect 360620 1006612 360622 1006632
rect 157430 1006576 157432 1006596
rect 157432 1006576 157484 1006596
rect 157484 1006576 157486 1006596
rect 360566 1006576 360622 1006612
rect 151266 1006476 151268 1006496
rect 151268 1006476 151320 1006496
rect 151320 1006476 151322 1006496
rect 151266 1006440 151322 1006476
rect 151726 1006440 151782 1006496
rect 158626 1006460 158682 1006496
rect 158626 1006440 158628 1006460
rect 158628 1006440 158680 1006460
rect 158680 1006440 158682 1006460
rect 147126 1006032 147182 1006088
rect 145746 996512 145802 996568
rect 145562 993928 145618 993984
rect 140594 993656 140650 993712
rect 147126 1000592 147182 1000648
rect 158258 1006324 158314 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 159454 1006324 159510 1006360
rect 159454 1006304 159456 1006324
rect 159456 1006304 159508 1006324
rect 159508 1006304 159510 1006324
rect 150898 1006204 150900 1006224
rect 150900 1006204 150952 1006224
rect 150952 1006204 150954 1006224
rect 150898 1006168 150954 1006204
rect 153750 1006188 153806 1006224
rect 153750 1006168 153752 1006188
rect 153752 1006168 153804 1006188
rect 153804 1006168 153806 1006188
rect 148874 1006068 148876 1006088
rect 148876 1006068 148928 1006088
rect 148928 1006068 148930 1006088
rect 148874 1006032 148930 1006068
rect 150070 1006068 150072 1006088
rect 150072 1006068 150124 1006088
rect 150124 1006068 150126 1006088
rect 150070 1006032 150126 1006068
rect 152922 1005100 152978 1005136
rect 152922 1005080 152924 1005100
rect 152924 1005080 152976 1005100
rect 152976 1005080 152978 1005100
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 153750 1004964 153806 1005000
rect 153750 1004944 153752 1004964
rect 153752 1004944 153804 1004964
rect 153804 1004944 153806 1004964
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 152922 1004828 152978 1004864
rect 152922 1004808 152924 1004828
rect 152924 1004808 152976 1004828
rect 152976 1004808 152978 1004828
rect 160282 1006188 160338 1006224
rect 255318 1006460 255374 1006496
rect 255318 1006440 255320 1006460
rect 255320 1006440 255372 1006460
rect 255372 1006440 255374 1006460
rect 361394 1006460 361450 1006496
rect 361394 1006440 361396 1006460
rect 361396 1006440 361448 1006460
rect 361448 1006440 361450 1006460
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 158258 1006052 158314 1006088
rect 158258 1006032 158260 1006052
rect 158260 1006032 158312 1006052
rect 158312 1006032 158314 1006052
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 154118 1004692 154174 1004728
rect 154118 1004672 154120 1004692
rect 154120 1004672 154172 1004692
rect 154172 1004672 154174 1004692
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 154578 1002108 154634 1002144
rect 154578 1002088 154580 1002108
rect 154580 1002088 154632 1002108
rect 154632 1002088 154634 1002108
rect 154302 995696 154358 995752
rect 154302 995016 154358 995072
rect 154946 1001952 155002 1002008
rect 155774 1001972 155830 1002008
rect 155774 1001952 155776 1001972
rect 155776 1001952 155828 1001972
rect 155828 1001952 155830 1001972
rect 156602 1001952 156658 1002008
rect 157798 1001972 157854 1002008
rect 157798 1001952 157800 1001972
rect 157800 1001952 157852 1001972
rect 157852 1001952 157854 1001972
rect 152462 994200 152518 994256
rect 149702 993656 149758 993712
rect 168930 995288 168986 995344
rect 171690 995329 171746 995344
rect 171690 995288 171692 995329
rect 171692 995288 171744 995329
rect 171744 995288 171746 995329
rect 169390 995016 169446 995072
rect 170678 995016 170734 995072
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 208398 1006052 208454 1006088
rect 208398 1006032 208400 1006052
rect 208400 1006032 208452 1006052
rect 208452 1006032 208454 1006052
rect 195058 998280 195114 998336
rect 178866 996376 178922 996432
rect 175922 995696 175978 995752
rect 188066 995696 188122 995752
rect 189446 995696 189502 995752
rect 191746 995696 191802 995752
rect 192482 995696 192538 995752
rect 194322 995696 194378 995752
rect 195058 995696 195114 995752
rect 173162 995016 173218 995072
rect 183834 995424 183890 995480
rect 183650 995288 183706 995344
rect 181442 994744 181498 994800
rect 187606 994472 187662 994528
rect 190366 994200 190422 994256
rect 188802 993928 188858 993984
rect 197818 996920 197874 996976
rect 212078 1005252 212080 1005272
rect 212080 1005252 212132 1005272
rect 212132 1005252 212134 1005272
rect 200210 998316 200212 998336
rect 200212 998316 200264 998336
rect 200264 998316 200266 998336
rect 200210 998280 200266 998316
rect 202694 998588 202696 998608
rect 202696 998588 202748 998608
rect 202748 998588 202750 998608
rect 202694 998552 202750 998588
rect 200670 997892 200726 997928
rect 200670 997872 200672 997892
rect 200672 997872 200724 997892
rect 200724 997872 200726 997892
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 199382 995968 199438 996024
rect 201866 998164 201922 998200
rect 201866 998144 201868 998164
rect 201868 998144 201920 998164
rect 201920 998144 201922 998164
rect 201682 995580 201738 995616
rect 201682 995560 201684 995580
rect 201684 995560 201736 995580
rect 201736 995560 201738 995580
rect 202694 998028 202750 998064
rect 202694 998008 202696 998028
rect 202696 998008 202748 998028
rect 202748 998008 202750 998028
rect 202326 995832 202382 995888
rect 204350 998996 204352 999016
rect 204352 998996 204404 999016
rect 204404 998996 204406 999016
rect 204350 998960 204406 998996
rect 203890 998724 203892 998744
rect 203892 998724 203944 998744
rect 203944 998724 203946 998744
rect 203890 998688 203946 998724
rect 203890 998452 203892 998472
rect 203892 998452 203944 998472
rect 203944 998452 203946 998472
rect 203890 998416 203946 998452
rect 204718 997772 204720 997792
rect 204720 997772 204772 997792
rect 204772 997772 204774 997792
rect 204718 997736 204774 997772
rect 203522 994472 203578 994528
rect 200946 994200 201002 994256
rect 200762 993928 200818 993984
rect 212078 1005216 212134 1005252
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 211250 1004828 211306 1004864
rect 211250 1004808 211252 1004828
rect 211252 1004808 211304 1004828
rect 211304 1004808 211306 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002244 206430 1002280
rect 206374 1002224 206376 1002244
rect 206376 1002224 206428 1002244
rect 206428 1002224 206430 1002244
rect 206742 1002244 206798 1002280
rect 206742 1002224 206744 1002244
rect 206744 1002224 206796 1002244
rect 206796 1002224 206798 1002244
rect 210882 1002244 210938 1002280
rect 210882 1002224 210884 1002244
rect 210884 1002224 210936 1002244
rect 210936 1002224 210938 1002244
rect 207202 1002108 207258 1002144
rect 207202 1002088 207204 1002108
rect 207204 1002088 207256 1002108
rect 207256 1002088 207258 1002108
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 205546 998164 205602 998200
rect 205546 998144 205548 998164
rect 205548 998144 205600 998164
rect 205600 998144 205602 998164
rect 206742 1001952 206798 1002008
rect 207570 1001952 207626 1002008
rect 210882 1001972 210938 1002008
rect 210882 1001952 210884 1001972
rect 210884 1001952 210936 1001972
rect 210936 1001952 210938 1001972
rect 212538 1002108 212594 1002144
rect 212538 1002088 212540 1002108
rect 212540 1002088 212592 1002108
rect 212592 1002088 212594 1002108
rect 207018 994744 207074 994800
rect 246578 996376 246634 996432
rect 240874 995696 240930 995752
rect 236550 995560 236606 995616
rect 231582 994744 231638 994800
rect 238574 995288 238630 995344
rect 234526 993928 234582 993984
rect 242070 995424 242126 995480
rect 239908 995152 239964 995208
rect 243266 994472 243322 994528
rect 243542 994472 243598 994528
rect 247038 995696 247094 995752
rect 243542 993928 243598 993984
rect 248142 995968 248198 996024
rect 248326 995016 248382 995072
rect 254122 1006324 254178 1006360
rect 254122 1006304 254124 1006324
rect 254124 1006304 254176 1006324
rect 254176 1006304 254178 1006324
rect 306930 1006324 306986 1006360
rect 306930 1006304 306932 1006324
rect 306932 1006304 306984 1006324
rect 306984 1006304 306986 1006324
rect 314658 1006324 314714 1006360
rect 314658 1006304 314660 1006324
rect 314660 1006304 314712 1006324
rect 314712 1006304 314714 1006324
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 252466 1006052 252522 1006088
rect 252466 1006032 252468 1006052
rect 252468 1006032 252520 1006052
rect 252520 1006032 252522 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 263046 1004964 263102 1005000
rect 263046 1004944 263048 1004964
rect 263048 1004944 263100 1004964
rect 263100 1004944 263102 1004964
rect 256146 1002652 256202 1002688
rect 256146 1002632 256148 1002652
rect 256148 1002632 256200 1002652
rect 256200 1002632 256202 1002652
rect 249246 995968 249302 996024
rect 252466 997892 252522 997928
rect 252466 997872 252468 997892
rect 252468 997872 252520 997892
rect 252520 997872 252522 997892
rect 252006 995288 252062 995344
rect 253294 998028 253350 998064
rect 253294 998008 253296 998028
rect 253296 998008 253348 998028
rect 253348 998008 253350 998028
rect 255318 1002516 255374 1002552
rect 255318 1002496 255320 1002516
rect 255320 1002496 255372 1002516
rect 255372 1002496 255374 1002516
rect 261022 1002516 261078 1002552
rect 261022 1002496 261024 1002516
rect 261024 1002496 261076 1002516
rect 261076 1002496 261078 1002516
rect 256146 1002380 256202 1002416
rect 256146 1002360 256148 1002380
rect 256148 1002360 256200 1002380
rect 256200 1002360 256202 1002380
rect 254490 1002244 254546 1002280
rect 254490 1002224 254492 1002244
rect 254492 1002224 254544 1002244
rect 254544 1002224 254546 1002244
rect 263506 1002108 263562 1002144
rect 263506 1002088 263508 1002108
rect 263508 1002088 263560 1002108
rect 263560 1002088 263562 1002108
rect 261022 1001972 261078 1002008
rect 261022 1001952 261024 1001972
rect 261024 1001952 261076 1001972
rect 261076 1001952 261078 1001972
rect 263874 1001972 263930 1002008
rect 263874 1001952 263876 1001972
rect 263876 1001952 263928 1001972
rect 263928 1001952 263930 1001972
rect 256974 998572 257030 998608
rect 256974 998552 256976 998572
rect 256976 998552 257028 998572
rect 257028 998552 257030 998572
rect 258998 998436 259054 998472
rect 258998 998416 259000 998436
rect 259000 998416 259052 998436
rect 259052 998416 259054 998436
rect 253662 998300 253718 998336
rect 253662 998280 253664 998300
rect 253664 998280 253716 998300
rect 253716 998280 253718 998300
rect 258170 998164 258226 998200
rect 258170 998144 258172 998164
rect 258172 998144 258224 998164
rect 258224 998144 258226 998164
rect 256514 998028 256570 998064
rect 256514 998008 256516 998028
rect 256516 998008 256568 998028
rect 256568 998008 256570 998028
rect 251822 995016 251878 995072
rect 257342 997892 257398 997928
rect 257342 997872 257344 997892
rect 257344 997872 257396 997892
rect 257396 997872 257398 997892
rect 255778 995560 255834 995616
rect 256054 995288 256110 995344
rect 255778 994744 255834 994800
rect 260194 998044 260196 998064
rect 260196 998044 260248 998064
rect 260248 998044 260250 998064
rect 260194 998008 260250 998044
rect 259826 997908 259828 997928
rect 259828 997908 259880 997928
rect 259880 997908 259882 997928
rect 259826 997872 259882 997908
rect 260194 997772 260196 997792
rect 260196 997772 260248 997792
rect 260248 997772 260250 997792
rect 260194 997736 260250 997772
rect 261850 997736 261906 997792
rect 259458 994472 259514 994528
rect 251454 994200 251510 994256
rect 249062 993928 249118 993984
rect 239586 993656 239642 993712
rect 287978 995696 288034 995752
rect 290554 995696 290610 995752
rect 291106 995696 291162 995752
rect 293590 995696 293646 995752
rect 298282 997192 298338 997248
rect 280802 995016 280858 995072
rect 285954 994744 286010 994800
rect 291382 995288 291438 995344
rect 291750 995288 291806 995344
rect 287150 994472 287206 994528
rect 300306 996648 300362 996704
rect 299570 995696 299626 995752
rect 304906 1006188 304962 1006224
rect 304906 1006168 304908 1006188
rect 304908 1006168 304960 1006188
rect 304960 1006168 304962 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006032 303306 1006088
rect 304078 1006032 304134 1006088
rect 311806 1006052 311862 1006088
rect 311806 1006032 311808 1006052
rect 311808 1006032 311860 1006052
rect 311860 1006032 311862 1006052
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 305274 1002108 305330 1002144
rect 305274 1002088 305276 1002108
rect 305276 1002088 305328 1002108
rect 305328 1002088 305330 1002108
rect 310150 1002108 310206 1002144
rect 310150 1002088 310152 1002108
rect 310152 1002088 310204 1002108
rect 310204 1002088 310206 1002108
rect 310978 1001972 311034 1002008
rect 310978 1001952 310980 1001972
rect 310980 1001952 311032 1001972
rect 311032 1001952 311034 1001972
rect 308954 1000492 308956 1000512
rect 308956 1000492 309008 1000512
rect 309008 1000492 309010 1000512
rect 308954 1000456 309010 1000492
rect 307298 998452 307300 998472
rect 307300 998452 307352 998472
rect 307352 998452 307354 998472
rect 301686 997192 301742 997248
rect 303066 996920 303122 996976
rect 304078 996104 304134 996160
rect 302882 995560 302938 995616
rect 301502 995288 301558 995344
rect 301686 995288 301742 995344
rect 307298 998416 307354 998452
rect 306102 998316 306104 998336
rect 306104 998316 306156 998336
rect 306156 998316 306158 998336
rect 306102 998280 306158 998316
rect 306930 998180 306932 998200
rect 306932 998180 306984 998200
rect 306984 998180 306986 998200
rect 306930 998144 306986 998180
rect 307758 998044 307760 998064
rect 307760 998044 307812 998064
rect 307812 998044 307814 998064
rect 304446 995288 304502 995344
rect 307758 998008 307814 998044
rect 310610 998044 310612 998064
rect 310612 998044 310664 998064
rect 310664 998044 310666 998064
rect 306102 997772 306104 997792
rect 306104 997772 306156 997792
rect 306156 997772 306158 997792
rect 306102 997736 306158 997772
rect 308126 997772 308128 997792
rect 308128 997772 308180 997792
rect 308180 997772 308182 997792
rect 308126 997736 308182 997772
rect 307206 995288 307262 995344
rect 310610 998008 310666 998044
rect 308954 997908 308956 997928
rect 308956 997908 309008 997928
rect 309008 997908 309010 997928
rect 308954 997872 309010 997908
rect 309782 997736 309838 997792
rect 310610 997736 310666 997792
rect 309138 994744 309194 994800
rect 304262 994472 304318 994528
rect 316406 994200 316462 994256
rect 295522 993928 295578 993984
rect 310518 993928 310574 993984
rect 355690 1006188 355746 1006224
rect 355690 1006168 355692 1006188
rect 355692 1006168 355744 1006188
rect 355744 1006168 355746 1006188
rect 365074 1006188 365130 1006224
rect 365074 1006168 365076 1006188
rect 365076 1006168 365128 1006188
rect 365128 1006168 365130 1006188
rect 354862 1006032 354918 1006088
rect 363418 1006052 363474 1006088
rect 363418 1006032 363420 1006052
rect 363420 1006032 363472 1006052
rect 363472 1006032 363474 1006052
rect 360566 1005388 360568 1005408
rect 360568 1005388 360620 1005408
rect 360620 1005388 360622 1005408
rect 360566 1005352 360622 1005388
rect 357714 1005252 357716 1005272
rect 357716 1005252 357768 1005272
rect 357768 1005252 357770 1005272
rect 357714 1005216 357770 1005252
rect 356518 1005100 356574 1005136
rect 356518 1005080 356520 1005100
rect 356520 1005080 356572 1005100
rect 356572 1005080 356574 1005100
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 355690 1004964 355746 1005000
rect 355690 1004944 355692 1004964
rect 355692 1004944 355744 1004964
rect 355744 1004944 355746 1004964
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 358542 1002244 358598 1002280
rect 358542 1002224 358544 1002244
rect 358544 1002224 358596 1002244
rect 358596 1002224 358598 1002244
rect 356518 1002108 356574 1002144
rect 356518 1002088 356520 1002108
rect 356520 1002088 356572 1002108
rect 356572 1002088 356574 1002108
rect 356886 1001952 356942 1002008
rect 357714 1001952 357770 1002008
rect 358542 1001952 358598 1002008
rect 360198 1001972 360254 1002008
rect 360198 1001952 360200 1001972
rect 360200 1001952 360252 1001972
rect 360252 1001952 360254 1001972
rect 365074 1005100 365130 1005136
rect 365074 1005080 365076 1005100
rect 365076 1005080 365128 1005100
rect 365128 1005080 365130 1005100
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 428370 1006868 428426 1006904
rect 428370 1006848 428372 1006868
rect 428372 1006848 428424 1006868
rect 428424 1006848 428426 1006868
rect 429198 1006732 429254 1006768
rect 429198 1006712 429200 1006732
rect 429200 1006712 429252 1006732
rect 429252 1006712 429254 1006732
rect 372710 996956 372712 996976
rect 372712 996956 372764 996976
rect 372764 996956 372766 996976
rect 372710 996920 372766 996956
rect 372526 996648 372582 996704
rect 372342 996376 372398 996432
rect 382094 997192 382150 997248
rect 382094 996376 382150 996432
rect 382278 996240 382334 996296
rect 380898 995152 380954 995208
rect 374826 994744 374882 994800
rect 383290 995968 383346 996024
rect 382922 995424 382978 995480
rect 383106 994472 383162 994528
rect 399942 996920 399998 996976
rect 399850 996240 399906 996296
rect 385038 995696 385094 995752
rect 388626 995696 388682 995752
rect 387890 995424 387946 995480
rect 388166 995424 388222 995480
rect 388442 995016 388498 995072
rect 392122 994744 392178 994800
rect 399850 995424 399906 995480
rect 431682 1006324 431738 1006360
rect 431682 1006304 431684 1006324
rect 431684 1006304 431736 1006324
rect 431736 1006304 431738 1006324
rect 429198 1006188 429254 1006224
rect 505006 1007020 505008 1007040
rect 505008 1007020 505060 1007040
rect 505060 1007020 505062 1007040
rect 505006 1006984 505062 1007020
rect 505374 1006884 505376 1006904
rect 505376 1006884 505428 1006904
rect 505428 1006884 505430 1006904
rect 505374 1006848 505430 1006884
rect 429198 1006168 429200 1006188
rect 429200 1006168 429252 1006188
rect 429252 1006168 429254 1006188
rect 422666 1006032 422722 1006088
rect 425518 1006052 425574 1006088
rect 425518 1006032 425520 1006052
rect 425520 1006032 425572 1006052
rect 425572 1006032 425574 1006052
rect 430026 1006052 430082 1006088
rect 430026 1006032 430028 1006052
rect 430028 1006032 430080 1006052
rect 430080 1006032 430082 1006052
rect 427542 1005660 427544 1005680
rect 427544 1005660 427596 1005680
rect 427596 1005660 427598 1005680
rect 427542 1005624 427598 1005660
rect 428370 1005524 428372 1005544
rect 428372 1005524 428424 1005544
rect 428424 1005524 428426 1005544
rect 428370 1005488 428426 1005524
rect 423494 1005388 423496 1005408
rect 423496 1005388 423548 1005408
rect 423548 1005388 423550 1005408
rect 423494 1005352 423550 1005388
rect 424322 1005252 424324 1005272
rect 424324 1005252 424376 1005272
rect 424376 1005252 424378 1005272
rect 424322 1005216 424378 1005252
rect 423494 1004964 423550 1005000
rect 423494 1004944 423496 1004964
rect 423496 1004944 423548 1004964
rect 423548 1004944 423550 1004964
rect 416134 995696 416190 995752
rect 415398 995444 415454 995480
rect 415398 995424 415400 995444
rect 415400 995424 415452 995444
rect 415452 995424 415454 995444
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 424322 1004572 424324 1004592
rect 424324 1004572 424376 1004592
rect 424376 1004572 424378 1004592
rect 424322 1004536 424378 1004572
rect 425518 1004164 425520 1004184
rect 425520 1004164 425572 1004184
rect 425572 1004164 425574 1004184
rect 425518 1004128 425574 1004164
rect 425150 1004028 425152 1004048
rect 425152 1004028 425204 1004048
rect 425204 1004028 425206 1004048
rect 425150 1003992 425206 1004028
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 426346 1002496 426402 1002552
rect 426346 1002244 426402 1002280
rect 426346 1002224 426348 1002244
rect 426348 1002224 426400 1002244
rect 426400 1002224 426402 1002244
rect 427174 1001972 427230 1002008
rect 427174 1001952 427176 1001972
rect 427176 1001952 427228 1001972
rect 427228 1001952 427230 1001972
rect 430854 1004828 430910 1004864
rect 430854 1004808 430856 1004828
rect 430856 1004808 430908 1004828
rect 430908 1004808 430910 1004828
rect 432050 1004828 432106 1004864
rect 432050 1004808 432052 1004828
rect 432052 1004808 432104 1004828
rect 432104 1004808 432106 1004828
rect 430026 1004692 430082 1004728
rect 430026 1004672 430028 1004692
rect 430028 1004672 430080 1004692
rect 430080 1004672 430082 1004692
rect 432878 1004692 432934 1004728
rect 432878 1004672 432880 1004692
rect 432880 1004672 432932 1004692
rect 432932 1004672 432934 1004692
rect 433338 1001972 433394 1002008
rect 433338 1001952 433340 1001972
rect 433340 1001952 433392 1001972
rect 433392 1001952 433394 1001972
rect 400862 994472 400918 994528
rect 440882 998280 440938 998336
rect 439870 996920 439926 996976
rect 439686 996376 439742 996432
rect 505374 1006612 505376 1006632
rect 505376 1006612 505428 1006632
rect 505428 1006612 505430 1006632
rect 505374 1006576 505430 1006612
rect 446402 995560 446458 995616
rect 454866 995832 454922 995888
rect 464342 994744 464398 994800
rect 465722 994472 465778 994528
rect 449162 994200 449218 994256
rect 507858 1006340 507860 1006360
rect 507860 1006340 507912 1006360
rect 507912 1006340 507914 1006360
rect 507858 1006304 507914 1006340
rect 506202 1006204 506204 1006224
rect 506204 1006204 506256 1006224
rect 506256 1006204 506258 1006224
rect 506202 1006168 506258 1006204
rect 471242 996648 471298 996704
rect 469862 996104 469918 996160
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 500498 1006052 500554 1006088
rect 500498 1006032 500500 1006052
rect 500500 1006032 500552 1006052
rect 500552 1006032 500554 1006052
rect 471426 995288 471482 995344
rect 488906 996920 488962 996976
rect 483754 995696 483810 995752
rect 485594 995696 485650 995752
rect 474738 995560 474794 995616
rect 480718 995560 480774 995616
rect 481270 995560 481326 995616
rect 476486 995288 476542 995344
rect 472254 995016 472310 995072
rect 476946 995016 477002 995072
rect 480718 995016 480774 995072
rect 481638 994744 481694 994800
rect 478602 994472 478658 994528
rect 509054 1005916 509110 1005952
rect 509054 1005896 509056 1005916
rect 509056 1005896 509108 1005916
rect 509108 1005896 509110 1005916
rect 498842 1005252 498844 1005272
rect 498844 1005252 498896 1005272
rect 498896 1005252 498898 1005272
rect 498842 1005216 498898 1005252
rect 499670 1004964 499726 1005000
rect 499670 1004944 499672 1004964
rect 499672 1004944 499724 1004964
rect 499724 1004944 499726 1004964
rect 508226 1004964 508282 1005000
rect 508226 1004944 508228 1004964
rect 508228 1004944 508280 1004964
rect 508280 1004944 508282 1004964
rect 509882 1004944 509938 1005000
rect 501326 1004828 501382 1004864
rect 501326 1004808 501328 1004828
rect 501328 1004808 501380 1004828
rect 501380 1004808 501382 1004828
rect 507030 1004828 507086 1004864
rect 507030 1004808 507032 1004828
rect 507032 1004808 507084 1004828
rect 507084 1004808 507086 1004828
rect 503350 1004692 503406 1004728
rect 503350 1004672 503352 1004692
rect 503352 1004672 503404 1004692
rect 503404 1004672 503406 1004692
rect 508226 1004692 508282 1004728
rect 508226 1004672 508228 1004692
rect 508228 1004672 508280 1004692
rect 508280 1004672 508282 1004692
rect 500498 1004572 500500 1004592
rect 500500 1004572 500552 1004592
rect 500552 1004572 500554 1004592
rect 500498 1004536 500554 1004572
rect 502522 1004028 502524 1004048
rect 502524 1004028 502576 1004048
rect 502576 1004028 502578 1004048
rect 502522 1003992 502578 1004028
rect 501694 1002244 501750 1002280
rect 501694 1002224 501696 1002244
rect 501696 1002224 501748 1002244
rect 501748 1002224 501750 1002244
rect 501694 1001972 501750 1002008
rect 501694 1001952 501696 1001972
rect 501696 1001952 501748 1001972
rect 501748 1001952 501750 1001972
rect 502522 1001952 502578 1002008
rect 503350 1001972 503406 1002008
rect 503350 1001952 503352 1001972
rect 503352 1001952 503404 1001972
rect 503404 1001952 503406 1001972
rect 504178 1001972 504234 1002008
rect 504178 1001952 504180 1001972
rect 504180 1001952 504232 1001972
rect 504232 1001952 504234 1001972
rect 504546 1002108 504602 1002144
rect 504546 1002088 504548 1002108
rect 504548 1002088 504600 1002108
rect 504600 1002088 504602 1002108
rect 504546 998008 504602 998064
rect 506202 995852 506258 995888
rect 506202 995832 506204 995852
rect 506204 995832 506256 995852
rect 506256 995832 506258 995852
rect 510342 1001972 510398 1002008
rect 510342 1001952 510344 1001972
rect 510344 1001952 510396 1001972
rect 510396 1001952 510398 1001972
rect 509054 995016 509110 995072
rect 511078 995016 511134 995072
rect 477958 994200 478014 994256
rect 517058 996920 517114 996976
rect 516874 996648 516930 996704
rect 516690 996376 516746 996432
rect 517518 995016 517574 995072
rect 552294 1007004 552350 1007040
rect 552294 1006984 552296 1007004
rect 552296 1006984 552348 1007004
rect 552348 1006984 552350 1007004
rect 518162 994744 518218 994800
rect 517702 994472 517758 994528
rect 519542 996104 519598 996160
rect 557170 1006748 557172 1006768
rect 557172 1006748 557224 1006768
rect 557224 1006748 557226 1006768
rect 557170 1006712 557226 1006748
rect 553122 1006612 553124 1006632
rect 553124 1006612 553176 1006632
rect 553176 1006612 553178 1006632
rect 553122 1006576 553178 1006612
rect 551098 1006476 551100 1006496
rect 551100 1006476 551152 1006496
rect 551152 1006476 551154 1006496
rect 551098 1006440 551154 1006476
rect 556802 1006476 556804 1006496
rect 556804 1006476 556856 1006496
rect 556856 1006476 556858 1006496
rect 553950 1006204 553952 1006224
rect 553952 1006204 554004 1006224
rect 554004 1006204 554006 1006224
rect 553950 1006168 554006 1006204
rect 554318 1006052 554374 1006088
rect 554318 1006032 554320 1006052
rect 554320 1006032 554372 1006052
rect 554372 1006032 554374 1006052
rect 551466 1005100 551522 1005136
rect 551466 1005080 551468 1005100
rect 551468 1005080 551520 1005100
rect 551520 1005080 551522 1005100
rect 555146 1002396 555148 1002416
rect 555148 1002396 555200 1002416
rect 555200 1002396 555202 1002416
rect 555146 1002360 555202 1002396
rect 554318 1002244 554374 1002280
rect 554318 1002224 554320 1002244
rect 554320 1002224 554372 1002244
rect 554372 1002224 554374 1002244
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 522486 995696 522542 995752
rect 551466 997772 551468 997792
rect 551468 997772 551520 997792
rect 551520 997772 551522 997792
rect 524050 997192 524106 997248
rect 551466 997736 551522 997772
rect 553122 998572 553178 998608
rect 553122 998552 553124 998572
rect 553124 998552 553176 998572
rect 553176 998552 553178 998572
rect 552294 998436 552350 998472
rect 552294 998416 552296 998436
rect 552296 998416 552348 998436
rect 552348 998416 552350 998436
rect 540886 996920 540942 996976
rect 524050 996648 524106 996704
rect 549442 996396 549498 996432
rect 549442 996376 549444 996396
rect 549444 996376 549496 996396
rect 549496 996376 549498 996396
rect 526074 995696 526130 995752
rect 528558 995696 528614 995752
rect 529110 995696 529166 995752
rect 533526 995696 533582 995752
rect 536562 995696 536618 995752
rect 523866 995424 523922 995480
rect 524786 995424 524842 995480
rect 530030 995016 530086 995072
rect 520922 994200 520978 994256
rect 532698 995424 532754 995480
rect 532514 994472 532570 994528
rect 532146 994200 532202 994256
rect 537390 994744 537446 994800
rect 538126 995152 538182 995208
rect 538310 995152 538366 995208
rect 555146 1001952 555202 1002008
rect 555974 1005388 555976 1005408
rect 555976 1005388 556028 1005408
rect 556028 1005388 556030 1005408
rect 555974 1005352 556030 1005388
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 556802 1006440 556858 1006476
rect 558826 1006340 558828 1006360
rect 558828 1006340 558880 1006360
rect 558880 1006340 558882 1006360
rect 558826 1006304 558882 1006340
rect 560850 1004964 560906 1005000
rect 560850 1004944 560852 1004964
rect 560852 1004944 560904 1004964
rect 560904 1004944 560906 1004964
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002516 558054 1002552
rect 557998 1002496 558000 1002516
rect 558000 1002496 558052 1002516
rect 558052 1002496 558054 1002516
rect 557998 1002244 558054 1002280
rect 557998 1002224 558000 1002244
rect 558000 1002224 558052 1002244
rect 558052 1002224 558054 1002244
rect 560850 1004692 560906 1004728
rect 560850 1004672 560852 1004692
rect 560852 1004672 560904 1004692
rect 560904 1004672 560906 1004692
rect 558826 1002380 558882 1002416
rect 558826 1002360 558828 1002380
rect 558828 1002360 558880 1002380
rect 558880 1002360 558882 1002380
rect 560482 1002244 560538 1002280
rect 560482 1002224 560484 1002244
rect 560484 1002224 560536 1002244
rect 560536 1002224 560538 1002244
rect 559654 1002108 559710 1002144
rect 559654 1002088 559656 1002108
rect 559656 1002088 559708 1002108
rect 559708 1002088 559710 1002108
rect 560022 1001972 560078 1002008
rect 560022 1001952 560024 1001972
rect 560024 1001952 560076 1001972
rect 560076 1001952 560078 1001972
rect 561678 1002108 561734 1002144
rect 561678 1002088 561680 1002108
rect 561680 1002088 561732 1002108
rect 561732 1002088 561734 1002108
rect 568210 994200 568266 994256
rect 570234 994744 570290 994800
rect 572902 994472 572958 994528
rect 590566 996920 590622 996976
rect 590566 996684 590568 996704
rect 590568 996684 590620 996704
rect 590620 996684 590622 996704
rect 590566 996648 590622 996684
rect 590566 996376 590622 996432
rect 625618 995968 625674 996024
rect 617154 995288 617210 995344
rect 590566 995016 590622 995072
rect 625802 995696 625858 995752
rect 627182 995696 627238 995752
rect 629758 995696 629814 995752
rect 630862 995696 630918 995752
rect 634542 995696 634598 995752
rect 637670 995696 637726 995752
rect 642086 995696 642142 995752
rect 629574 995560 629630 995616
rect 635830 995288 635886 995344
rect 635186 994744 635242 994800
rect 631506 994472 631562 994528
rect 627918 994200 627974 994256
rect 660578 995035 660634 995072
rect 660578 995016 660580 995035
rect 660580 995016 660632 995035
rect 660632 995016 660634 995035
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 937216 660358 937272
rect 663062 941704 663118 941760
rect 665822 939800 665878 939856
rect 673366 966592 673422 966648
rect 675114 966592 675170 966648
rect 673182 960744 673238 960800
rect 672998 952176 673054 952232
rect 672722 947280 672778 947336
rect 669962 938440 670018 938496
rect 671802 938032 671858 938088
rect 671618 937760 671674 937816
rect 668582 937488 668638 937544
rect 658922 935992 658978 936048
rect 670698 929464 670754 929520
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 55862 892744 55918 892800
rect 54482 892472 54538 892528
rect 53286 892200 53342 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62762 858608 62818 858664
rect 62118 845552 62174 845608
rect 53102 799312 53158 799368
rect 50342 730496 50398 730552
rect 48962 669296 49018 669352
rect 47766 614080 47822 614136
rect 62118 832496 62174 832552
rect 54482 774288 54538 774344
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793620 62174 793656
rect 62118 793600 62120 793620
rect 62120 793600 62172 793620
rect 62172 793600 62174 793620
rect 652390 856296 652446 856352
rect 651838 842968 651894 843024
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 651470 789928 651526 789984
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 55862 772792 55918 772848
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 652390 776600 652446 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62762 743008 62818 743064
rect 62118 741240 62174 741296
rect 53102 730088 53158 730144
rect 51722 691328 51778 691384
rect 51722 646584 51778 646640
rect 652022 736752 652078 736808
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 651470 723424 651526 723480
rect 651470 710232 651526 710288
rect 62762 697856 62818 697912
rect 651470 696940 651472 696960
rect 651472 696940 651524 696960
rect 651524 696940 651526 696960
rect 651470 696904 651526 696940
rect 62118 689152 62174 689208
rect 651654 683576 651710 683632
rect 62118 676096 62174 676152
rect 651470 670384 651526 670440
rect 62118 663040 62174 663096
rect 651470 657056 651526 657112
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 50342 626592 50398 626648
rect 651470 630536 651526 630592
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652022 627816 652078 627872
rect 664442 868672 664498 868728
rect 663062 760416 663118 760472
rect 661682 673104 661738 673160
rect 661682 643728 661738 643784
rect 660302 625232 660358 625288
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 51722 601704 51778 601760
rect 50342 601296 50398 601352
rect 47582 582392 47638 582448
rect 44822 556416 44878 556472
rect 44822 556008 44878 556064
rect 48962 557776 49018 557832
rect 51722 557504 51778 557560
rect 45558 556824 45614 556880
rect 45006 555600 45062 555656
rect 44362 555192 44418 555248
rect 44178 548664 44234 548720
rect 43626 547712 43682 547768
rect 43810 547032 43866 547088
rect 42982 379344 43038 379400
rect 43350 371864 43406 371920
rect 42982 365744 43038 365800
rect 42430 356088 42486 356144
rect 43350 355816 43406 355872
rect 41878 355680 41934 355736
rect 44178 535200 44234 535256
rect 44730 554376 44786 554432
rect 44546 550704 44602 550760
rect 44546 532752 44602 532808
rect 44362 428032 44418 428088
rect 44454 427624 44510 427680
rect 44270 426808 44326 426864
rect 43994 419464 44050 419520
rect 45098 551520 45154 551576
rect 45282 549072 45338 549128
rect 45282 534384 45338 534440
rect 45098 529624 45154 529680
rect 45558 429664 45614 429720
rect 45190 429256 45246 429312
rect 44914 428848 44970 428904
rect 45006 428440 45062 428496
rect 44730 427216 44786 427272
rect 44638 422456 44694 422512
rect 44822 420688 44878 420744
rect 44638 407088 44694 407144
rect 44638 385192 44694 385248
rect 44454 384784 44510 384840
rect 44270 383968 44326 384024
rect 44454 379888 44510 379944
rect 44270 377440 44326 377496
rect 45374 418240 45430 418296
rect 45374 406816 45430 406872
rect 45190 386688 45246 386744
rect 45190 386008 45246 386064
rect 45006 385600 45062 385656
rect 44454 359896 44510 359952
rect 44270 356632 44326 356688
rect 45190 384376 45246 384432
rect 45374 383560 45430 383616
rect 43902 354184 43958 354240
rect 44730 353776 44786 353832
rect 28538 351192 28594 351248
rect 38290 346296 38346 346352
rect 28906 344256 28962 344312
rect 28538 343848 28594 343904
rect 45006 343304 45062 343360
rect 45558 380296 45614 380352
rect 47582 430072 47638 430128
rect 46938 426400 46994 426456
rect 47122 423544 47178 423600
rect 47122 400152 47178 400208
rect 46938 399744 46994 399800
rect 46938 380704 46994 380760
rect 46202 366968 46258 367024
rect 45558 357312 45614 357368
rect 45650 356632 45706 356688
rect 45926 355816 45982 355872
rect 45282 341672 45338 341728
rect 45282 341264 45338 341320
rect 45466 340856 45522 340912
rect 35806 339768 35862 339824
rect 34426 338544 34482 338600
rect 34426 336096 34482 336152
rect 43074 334600 43130 334656
rect 43626 334600 43682 334656
rect 44270 334600 44326 334656
rect 42798 334328 42854 334384
rect 37922 328344 37978 328400
rect 41786 326712 41842 326768
rect 41786 325352 41842 325408
rect 41786 324808 41842 324864
rect 42062 322768 42118 322824
rect 42430 321408 42486 321464
rect 43442 323040 43498 323096
rect 42430 320048 42486 320104
rect 42430 319368 42486 319424
rect 42246 317464 42302 317520
rect 41786 316648 41842 316704
rect 42154 315968 42210 316024
rect 41786 315560 41842 315616
rect 42154 313656 42210 313712
rect 42430 312704 42486 312760
rect 42154 312296 42210 312352
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 42890 299648 42946 299704
rect 41786 296792 41842 296848
rect 41326 295976 41382 296032
rect 32402 294752 32458 294808
rect 41786 292440 41842 292496
rect 41786 290400 41842 290456
rect 41326 290264 41382 290320
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42430 278704 42486 278760
rect 42338 278432 42394 278488
rect 41786 277888 41842 277944
rect 42154 277888 42210 277944
rect 42062 277072 42118 277128
rect 42062 276528 42118 276584
rect 41786 274216 41842 274272
rect 42062 273400 42118 273456
rect 42062 272992 42118 273048
rect 41786 270408 41842 270464
rect 42430 270408 42486 270464
rect 41786 269048 41842 269104
rect 40682 267008 40738 267064
rect 35806 259936 35862 259992
rect 35806 258304 35862 258360
rect 35806 257080 35862 257136
rect 43258 298832 43314 298888
rect 43074 295160 43130 295216
rect 43074 276528 43130 276584
rect 42890 256808 42946 256864
rect 42798 256400 42854 256456
rect 35438 253408 35494 253464
rect 35622 253000 35678 253056
rect 35806 252592 35862 252648
rect 35806 252184 35862 252240
rect 40682 242800 40738 242856
rect 41786 240080 41842 240136
rect 42154 238448 42210 238504
rect 41786 235864 41842 235920
rect 42246 235864 42302 235920
rect 42246 234504 42302 234560
rect 42246 234096 42302 234152
rect 42154 233280 42210 233336
rect 42246 231648 42302 231704
rect 42154 230152 42210 230208
rect 42246 229880 42302 229936
rect 42614 237360 42670 237416
rect 41970 227296 42026 227352
rect 42154 226616 42210 226672
rect 42430 225664 42486 225720
rect 40682 222808 40738 222864
rect 35530 217912 35586 217968
rect 35530 214240 35586 214296
rect 35806 214240 35862 214296
rect 43626 322768 43682 322824
rect 44270 320048 44326 320104
rect 44178 311480 44234 311536
rect 44362 311208 44418 311264
rect 44362 300056 44418 300112
rect 44178 299240 44234 299296
rect 45834 340040 45890 340096
rect 45650 339224 45706 339280
rect 46018 338408 46074 338464
rect 46018 319368 46074 319424
rect 45834 313656 45890 313712
rect 45650 312296 45706 312352
rect 47122 379072 47178 379128
rect 47122 361528 47178 361584
rect 46938 356088 46994 356144
rect 47582 333104 47638 333160
rect 46386 303048 46442 303104
rect 45466 298424 45522 298480
rect 44178 298016 44234 298072
rect 43626 293936 43682 293992
rect 43994 293120 44050 293176
rect 43810 291896 43866 291952
rect 43994 279792 44050 279848
rect 43810 277072 43866 277128
rect 43626 272992 43682 273048
rect 43442 257624 43498 257680
rect 43258 255992 43314 256048
rect 43626 255584 43682 255640
rect 42982 254768 43038 254824
rect 42798 213696 42854 213752
rect 43442 251096 43498 251152
rect 43258 242800 43314 242856
rect 44362 294344 44418 294400
rect 44638 293528 44694 293584
rect 44638 273400 44694 273456
rect 44362 270408 44418 270464
rect 44178 255176 44234 255232
rect 44178 253952 44234 254008
rect 43718 249056 43774 249112
rect 43718 231648 43774 231704
rect 43442 226616 43498 226672
rect 43258 225664 43314 225720
rect 43442 213288 43498 213344
rect 42982 212064 43038 212120
rect 35806 211384 35862 211440
rect 42798 209616 42854 209672
rect 35806 208936 35862 208992
rect 41694 208936 41750 208992
rect 40038 207712 40094 207768
rect 35622 204040 35678 204096
rect 35806 203632 35862 203688
rect 35622 202136 35678 202192
rect 37922 197784 37978 197840
rect 41786 197104 41842 197160
rect 41878 195744 41934 195800
rect 42614 195472 42670 195528
rect 41970 195200 42026 195256
rect 42430 193160 42486 193216
rect 42614 192888 42670 192944
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41786 187176 41842 187232
rect 42338 186224 42394 186280
rect 41786 185816 41842 185872
rect 42430 184864 42486 184920
rect 42430 183096 42486 183152
rect 43258 207984 43314 208040
rect 42982 206352 43038 206408
rect 42982 191120 43038 191176
rect 43626 212880 43682 212936
rect 44638 251912 44694 251968
rect 44546 248648 44602 248704
rect 44362 248240 44418 248296
rect 44362 235864 44418 235920
rect 44454 234096 44510 234152
rect 44638 233280 44694 233336
rect 45006 297200 45062 297256
rect 45190 291624 45246 291680
rect 46202 290672 46258 290728
rect 45190 277888 45246 277944
rect 45006 254360 45062 254416
rect 45558 250688 45614 250744
rect 45834 250280 45890 250336
rect 46018 249464 46074 249520
rect 46018 234504 46074 234560
rect 45834 230152 45890 230208
rect 45558 229880 45614 229936
rect 44822 214920 44878 214976
rect 44178 211248 44234 211304
rect 45006 210840 45062 210896
rect 44178 210432 44234 210488
rect 43626 206760 43682 206816
rect 43442 206216 43498 206272
rect 43442 202136 43498 202192
rect 43258 183096 43314 183152
rect 43810 205536 43866 205592
rect 43626 193160 43682 193216
rect 43994 205128 44050 205184
rect 43994 191664 44050 191720
rect 43810 190440 43866 190496
rect 44362 208528 44418 208584
rect 44546 205944 44602 206000
rect 44362 189896 44418 189952
rect 44822 204720 44878 204776
rect 44546 187584 44602 187640
rect 44178 184864 44234 184920
rect 46938 247016 46994 247072
rect 46938 238448 46994 238504
rect 50342 430888 50398 430944
rect 48962 386960 49018 387016
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 49146 346296 49202 346352
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 212472 48006 212528
rect 48594 194384 48650 194440
rect 47950 192344 48006 192400
rect 49146 289856 49202 289912
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 660302 599528 660358 599584
rect 62118 597896 62174 597952
rect 652390 590708 652446 590744
rect 652390 590688 652392 590708
rect 652392 590688 652444 590708
rect 652444 590688 652446 590708
rect 62118 584840 62174 584896
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 652574 497664 652630 497720
rect 62118 493584 62174 493640
rect 669226 879144 669282 879200
rect 668766 877648 668822 877704
rect 667846 866632 667902 866688
rect 666466 778368 666522 778424
rect 665822 761504 665878 761560
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661866 581032 661922 581088
rect 659106 553968 659162 554024
rect 658922 491952 658978 492008
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 55862 408448 55918 408504
rect 651470 404640 651526 404696
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51722 301280 51778 301336
rect 51722 289856 51778 289912
rect 50342 259936 50398 259992
rect 50526 247696 50582 247752
rect 50342 246472 50398 246528
rect 49514 208936 49570 208992
rect 49330 206216 49386 206272
rect 49514 196424 49570 196480
rect 49330 190440 49386 190496
rect 50710 203224 50766 203280
rect 652574 391448 652630 391504
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 652022 378120 652078 378176
rect 62118 376216 62174 376272
rect 651654 364792 651710 364848
rect 62118 363296 62174 363352
rect 651470 351600 651526 351656
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 55862 278704 55918 278760
rect 651470 338272 651526 338328
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 651470 285232 651526 285288
rect 62946 285096 63002 285152
rect 62762 267008 62818 267064
rect 53102 217912 53158 217968
rect 136546 269728 136602 269784
rect 139950 269764 139952 269784
rect 139952 269764 140004 269784
rect 140004 269764 140006 269784
rect 139950 269728 140006 269764
rect 468758 269184 468814 269240
rect 475382 269456 475438 269512
rect 475750 269728 475806 269784
rect 476302 269456 476358 269512
rect 476026 269184 476082 269240
rect 480258 270680 480314 270736
rect 478878 269728 478934 269784
rect 479062 269356 479064 269376
rect 479064 269356 479116 269376
rect 479116 269356 479118 269376
rect 479062 269320 479118 269356
rect 480350 269356 480352 269376
rect 480352 269356 480404 269376
rect 480404 269356 480406 269376
rect 480350 269320 480406 269356
rect 482282 270036 482284 270056
rect 482284 270036 482336 270056
rect 482336 270036 482338 270056
rect 482282 270000 482338 270036
rect 483110 270680 483166 270736
rect 484582 270000 484638 270056
rect 484306 269456 484362 269512
rect 484858 266756 484914 266792
rect 484858 266736 484860 266756
rect 484860 266736 484912 266756
rect 484912 266736 484914 266756
rect 487434 266736 487490 266792
rect 490010 269492 490012 269512
rect 490012 269492 490064 269512
rect 490064 269492 490066 269512
rect 490010 269456 490066 269492
rect 494242 270272 494298 270328
rect 504914 270544 504970 270600
rect 504730 269728 504786 269784
rect 504914 267416 504970 267472
rect 507858 270544 507914 270600
rect 508042 267436 508098 267472
rect 508042 267416 508044 267436
rect 508044 267416 508096 267436
rect 508096 267416 508098 267436
rect 509238 267028 509294 267064
rect 509238 267008 509240 267028
rect 509240 267008 509292 267028
rect 509292 267008 509294 267028
rect 513194 273944 513250 274000
rect 514114 273964 514170 274000
rect 514114 273944 514116 273964
rect 514116 273944 514168 273964
rect 514168 273944 514170 273964
rect 514298 271260 514300 271280
rect 514300 271260 514352 271280
rect 514352 271260 514354 271280
rect 514298 271224 514354 271260
rect 513838 268388 513894 268424
rect 513838 268368 513840 268388
rect 513840 268368 513892 268388
rect 513892 268368 513894 268388
rect 514942 268368 514998 268424
rect 514666 267280 514722 267336
rect 519726 271632 519782 271688
rect 518346 271224 518402 271280
rect 521106 273944 521162 274000
rect 517518 267044 517520 267064
rect 517520 267044 517572 267064
rect 517572 267044 517574 267064
rect 517518 267008 517574 267044
rect 517334 266736 517390 266792
rect 518898 267552 518954 267608
rect 518990 267280 519046 267336
rect 519174 267008 519230 267064
rect 518714 266736 518770 266792
rect 521474 272448 521530 272504
rect 525522 275732 525578 275768
rect 525522 275712 525524 275732
rect 525524 275712 525576 275732
rect 525576 275712 525578 275732
rect 524050 273964 524106 274000
rect 524050 273944 524052 273964
rect 524052 273944 524104 273964
rect 524104 273944 524106 273964
rect 523498 271360 523554 271416
rect 524142 271088 524198 271144
rect 523498 268252 523554 268288
rect 523498 268232 523500 268252
rect 523500 268232 523552 268252
rect 523552 268232 523554 268252
rect 521658 267552 521714 267608
rect 522670 267280 522726 267336
rect 525890 271632 525946 271688
rect 525706 271360 525762 271416
rect 527178 268524 527234 268560
rect 527178 268504 527180 268524
rect 527180 268504 527232 268524
rect 527232 268504 527234 268524
rect 527730 275732 527786 275768
rect 527730 275712 527732 275732
rect 527732 275712 527784 275732
rect 527784 275712 527786 275732
rect 528512 274372 528568 274408
rect 528512 274352 528514 274372
rect 528514 274352 528566 274372
rect 528566 274352 528568 274372
rect 528098 274080 528154 274136
rect 527914 272856 527970 272912
rect 527546 268232 527602 268288
rect 527454 266736 527510 266792
rect 528650 274100 528706 274136
rect 528650 274080 528652 274100
rect 528652 274080 528704 274100
rect 528704 274080 528706 274100
rect 528650 272892 528652 272912
rect 528652 272892 528704 272912
rect 528704 272892 528706 272912
rect 528650 272856 528706 272892
rect 528374 272448 528430 272504
rect 528558 272484 528560 272504
rect 528560 272484 528612 272504
rect 528612 272484 528614 272504
rect 528558 272448 528614 272484
rect 530766 274896 530822 274952
rect 529846 271360 529902 271416
rect 528926 268524 528982 268560
rect 528926 268504 528928 268524
rect 528928 268504 528980 268524
rect 528980 268504 528982 268524
rect 528558 268252 528614 268288
rect 528558 268232 528566 268252
rect 528566 268232 528614 268252
rect 528558 267552 528614 267608
rect 528650 267300 528706 267336
rect 528650 267280 528652 267300
rect 528652 267280 528704 267300
rect 528704 267280 528706 267300
rect 528466 267028 528522 267064
rect 528466 267008 528468 267028
rect 528468 267008 528520 267028
rect 528520 267008 528522 267028
rect 528742 267028 528798 267064
rect 528742 267008 528744 267028
rect 528744 267008 528796 267028
rect 528796 267008 528798 267028
rect 528742 266620 528798 266656
rect 528742 266600 528744 266620
rect 528744 266600 528796 266620
rect 528796 266600 528798 266620
rect 531318 269728 531374 269784
rect 531686 272448 531742 272504
rect 534170 274916 534226 274952
rect 534170 274896 534172 274916
rect 534172 274896 534224 274916
rect 534224 274896 534226 274916
rect 533710 272176 533766 272232
rect 532790 270000 532846 270056
rect 533066 270000 533122 270056
rect 531870 267572 531926 267608
rect 531870 267552 531872 267572
rect 531872 267552 531924 267572
rect 531924 267552 531926 267572
rect 535274 275324 535330 275360
rect 535274 275304 535276 275324
rect 535276 275304 535328 275324
rect 535328 275304 535330 275324
rect 534722 269728 534778 269784
rect 538218 275032 538274 275088
rect 536102 270544 536158 270600
rect 535642 268232 535698 268288
rect 536378 267008 536434 267064
rect 538218 274624 538274 274680
rect 537942 274352 537998 274408
rect 538126 274080 538182 274136
rect 538310 274080 538366 274136
rect 538218 272720 538274 272776
rect 538310 272176 538366 272232
rect 538034 271360 538090 271416
rect 537850 270544 537906 270600
rect 538034 270580 538036 270600
rect 538036 270580 538088 270600
rect 538088 270580 538090 270600
rect 538034 270544 538090 270580
rect 538862 275324 538918 275360
rect 538862 275304 538864 275324
rect 538864 275304 538916 275324
rect 538916 275304 538918 275324
rect 538862 273808 538918 273864
rect 538034 269728 538090 269784
rect 537850 269456 537906 269512
rect 537574 267552 537630 267608
rect 537390 266600 537446 266656
rect 538402 269456 538458 269512
rect 538218 269048 538274 269104
rect 538310 267572 538366 267608
rect 538310 267552 538312 267572
rect 538312 267552 538364 267572
rect 538364 267552 538366 267572
rect 538218 267280 538274 267336
rect 540702 272448 540758 272504
rect 539598 270544 539654 270600
rect 539230 267960 539286 268016
rect 538862 267008 538918 267064
rect 539690 267552 539746 267608
rect 540242 266736 540298 266792
rect 544198 275032 544254 275088
rect 544382 274896 544438 274952
rect 543186 274624 543242 274680
rect 541438 269320 541494 269376
rect 540886 266736 540942 266792
rect 542174 267008 542230 267064
rect 543554 269356 543556 269376
rect 543556 269356 543608 269376
rect 543608 269356 543610 269376
rect 543554 269320 543610 269356
rect 546038 274916 546094 274952
rect 546038 274896 546040 274916
rect 546040 274896 546092 274916
rect 546092 274896 546094 274916
rect 545118 272720 545174 272776
rect 544382 269048 544438 269104
rect 543692 268388 543748 268424
rect 543692 268368 543694 268388
rect 543694 268368 543746 268388
rect 543746 268368 543748 268388
rect 543830 267960 543886 268016
rect 544014 267824 544070 267880
rect 543830 267280 543886 267336
rect 549442 268368 549498 268424
rect 552662 267824 552718 267880
rect 574926 270272 574982 270328
rect 580262 267280 580318 267336
rect 617982 271088 618038 271144
rect 626446 272448 626502 272504
rect 607862 267008 607918 267064
rect 635646 273808 635702 273864
rect 630678 270000 630734 270056
rect 637578 269728 637634 269784
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553490 255604 553546 255640
rect 553490 255584 553492 255604
rect 553492 255584 553544 255604
rect 553544 255584 553546 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 553858 249056 553914 249112
rect 554410 246880 554466 246936
rect 554502 244704 554558 244760
rect 553950 242528 554006 242584
rect 553858 240352 553914 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 62946 222808 63002 222864
rect 73066 226888 73122 226944
rect 68926 224168 68982 224224
rect 70030 220088 70086 220144
rect 72882 220360 72938 220416
rect 79966 228248 80022 228304
rect 103610 229744 103666 229800
rect 101862 221448 101918 221504
rect 123482 222808 123538 222864
rect 134614 227976 134670 228032
rect 139306 226480 139362 226536
rect 136362 225256 136418 225312
rect 138570 221720 138626 221776
rect 141146 227976 141202 228032
rect 142158 227160 142214 227216
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 142250 225292 142252 225312
rect 142252 225292 142304 225312
rect 142304 225292 142306 225312
rect 142250 225256 142306 225292
rect 143078 227160 143134 227216
rect 142986 225528 143042 225584
rect 141422 223932 141424 223952
rect 141424 223932 141476 223952
rect 141476 223932 141478 223952
rect 141422 223896 141478 223932
rect 141054 220768 141110 220824
rect 140226 218612 140282 218648
rect 140226 218592 140228 218612
rect 140228 218592 140280 218612
rect 140280 218592 140282 218612
rect 142434 221176 142490 221232
rect 145654 229744 145710 229800
rect 146298 229220 146354 229256
rect 146298 229200 146300 229220
rect 146300 229200 146352 229220
rect 146352 229200 146354 229220
rect 145930 227976 145986 228032
rect 145378 223932 145380 223952
rect 145380 223932 145432 223952
rect 145432 223932 145434 223952
rect 145378 223896 145434 223932
rect 144182 221196 144238 221232
rect 144182 221176 144184 221196
rect 144184 221176 144236 221196
rect 144236 221176 144238 221196
rect 143630 218592 143686 218648
rect 146206 223896 146262 223952
rect 147954 229200 148010 229256
rect 147402 225564 147404 225584
rect 147404 225564 147456 225584
rect 147456 225564 147458 225584
rect 147402 225528 147458 225564
rect 147678 223932 147680 223952
rect 147680 223932 147732 223952
rect 147732 223932 147734 223952
rect 147678 223896 147734 223932
rect 147310 222128 147366 222184
rect 146574 221720 146630 221776
rect 147494 221856 147550 221912
rect 146390 220768 146446 220824
rect 147218 220768 147274 220824
rect 148414 220768 148470 220824
rect 151358 229880 151414 229936
rect 150346 227976 150402 228032
rect 150346 226616 150402 226672
rect 149058 221856 149114 221912
rect 149334 218748 149390 218784
rect 149334 218728 149336 218748
rect 149336 218728 149388 218748
rect 149388 218728 149390 218748
rect 150622 220768 150678 220824
rect 152370 229880 152426 229936
rect 151818 227296 151874 227352
rect 151726 223760 151782 223816
rect 150806 220088 150862 220144
rect 152278 226616 152334 226672
rect 152922 226072 152978 226128
rect 152738 224304 152794 224360
rect 152094 222128 152150 222184
rect 154670 227296 154726 227352
rect 155866 227976 155922 228032
rect 155314 226888 155370 226944
rect 153750 220496 153806 220552
rect 154578 223984 154634 223986
rect 154578 223932 154580 223984
rect 154580 223932 154632 223984
rect 154632 223932 154634 223984
rect 154578 223930 154634 223932
rect 153934 218728 153990 218784
rect 155314 222400 155370 222456
rect 157430 228520 157486 228576
rect 157982 228928 158038 228984
rect 157798 227976 157854 228032
rect 157614 226108 157616 226128
rect 157616 226108 157668 226128
rect 157668 226108 157670 226128
rect 157614 226072 157670 226108
rect 156142 220768 156198 220824
rect 156878 223760 156934 223816
rect 157338 224440 157394 224496
rect 157430 224032 157486 224088
rect 157246 223388 157248 223408
rect 157248 223388 157300 223408
rect 157300 223388 157302 223408
rect 157246 223352 157302 223388
rect 157430 223388 157432 223408
rect 157432 223388 157484 223408
rect 157484 223388 157486 223408
rect 157430 223352 157486 223388
rect 157246 222436 157248 222456
rect 157248 222436 157300 222456
rect 157300 222436 157302 222456
rect 157246 222400 157302 222436
rect 157614 220380 157670 220416
rect 157614 220360 157616 220380
rect 157616 220360 157668 220380
rect 157668 220360 157670 220380
rect 158810 228520 158866 228576
rect 159638 227452 159694 227488
rect 159638 227432 159640 227452
rect 159640 227432 159692 227452
rect 159692 227432 159694 227452
rect 160466 228248 160522 228304
rect 158626 223352 158682 223408
rect 161570 225528 161626 225584
rect 161570 220360 161626 220416
rect 161570 218340 161626 218376
rect 161570 218320 161572 218340
rect 161572 218320 161624 218340
rect 161624 218320 161626 218340
rect 162306 218320 162362 218376
rect 163870 228928 163926 228984
rect 162950 224440 163006 224496
rect 163962 223896 164018 223952
rect 165158 220224 165214 220280
rect 166630 228384 166686 228440
rect 166446 227432 166502 227488
rect 166814 225836 166816 225856
rect 166816 225836 166868 225856
rect 166868 225836 166870 225856
rect 166814 225800 166870 225836
rect 166722 225528 166778 225584
rect 166538 225020 166540 225040
rect 166540 225020 166592 225040
rect 166592 225020 166594 225040
rect 166538 224984 166594 225020
rect 166446 223352 166502 223408
rect 166262 223116 166264 223136
rect 166264 223116 166316 223136
rect 166316 223116 166318 223136
rect 166262 223080 166318 223116
rect 165618 222808 165674 222864
rect 166078 222572 166080 222592
rect 166080 222572 166132 222592
rect 166132 222572 166134 222592
rect 166078 222536 166134 222572
rect 166998 222572 167000 222592
rect 167000 222572 167052 222592
rect 167052 222572 167054 222592
rect 166998 222536 167054 222572
rect 166814 222264 166870 222320
rect 168102 222264 168158 222320
rect 167642 220224 167698 220280
rect 169850 225800 169906 225856
rect 171138 228928 171194 228984
rect 170862 225936 170918 225992
rect 171230 225972 171232 225992
rect 171232 225972 171284 225992
rect 171284 225972 171286 225992
rect 171230 225936 171286 225972
rect 171046 225700 171048 225720
rect 171048 225700 171100 225720
rect 171100 225700 171102 225720
rect 171046 225664 171102 225700
rect 171046 225020 171048 225040
rect 171048 225020 171100 225040
rect 171100 225020 171102 225040
rect 171046 224984 171102 225020
rect 170954 224204 170956 224224
rect 170956 224204 171008 224224
rect 171008 224204 171010 224224
rect 170954 224168 171010 224204
rect 172242 228928 172298 228984
rect 172426 228928 172482 228984
rect 171598 228384 171654 228440
rect 171414 224168 171470 224224
rect 170954 223896 171010 223952
rect 170402 223080 170458 223136
rect 171138 222164 171140 222184
rect 171140 222164 171192 222184
rect 171192 222164 171194 222184
rect 171138 222128 171194 222164
rect 170862 221856 170918 221912
rect 171414 221876 171470 221912
rect 171414 221856 171416 221876
rect 171416 221856 171468 221876
rect 171468 221856 171470 221876
rect 174082 228948 174138 228984
rect 174082 228928 174084 228948
rect 174084 228928 174136 228948
rect 174136 228928 174138 228948
rect 174266 228792 174322 228848
rect 174818 222572 174820 222592
rect 174820 222572 174872 222592
rect 174872 222572 174874 222592
rect 174818 222536 174874 222572
rect 175646 228792 175702 228848
rect 176658 226072 176714 226128
rect 176934 225664 176990 225720
rect 176474 225256 176530 225312
rect 176750 225256 176806 225312
rect 175462 222536 175518 222592
rect 177578 222148 177634 222184
rect 177578 222128 177580 222148
rect 177580 222128 177632 222148
rect 177632 222128 177634 222148
rect 178038 221448 178094 221504
rect 178314 221332 178370 221368
rect 178314 221312 178316 221332
rect 178316 221312 178368 221332
rect 178368 221312 178370 221332
rect 180614 228928 180670 228984
rect 181902 228948 181958 228984
rect 181902 228928 181904 228948
rect 181904 228928 181956 228948
rect 181956 228928 181958 228948
rect 180798 226072 180854 226128
rect 181074 226072 181130 226128
rect 184846 225664 184902 225720
rect 185582 225120 185638 225176
rect 186134 226072 186190 226128
rect 186410 225972 186412 225992
rect 186412 225972 186464 225992
rect 186464 225972 186466 225992
rect 186410 225936 186466 225972
rect 186410 225664 186466 225720
rect 186134 225392 186190 225448
rect 187054 225392 187110 225448
rect 185122 221312 185178 221368
rect 188066 225936 188122 225992
rect 190550 229084 190606 229120
rect 190550 229064 190552 229084
rect 190552 229064 190604 229084
rect 190604 229064 190606 229084
rect 190550 225428 190552 225448
rect 190552 225428 190604 225448
rect 190604 225428 190606 225448
rect 190550 225392 190606 225428
rect 192298 229064 192354 229120
rect 194874 225392 194930 225448
rect 195518 225120 195574 225176
rect 194874 220788 194930 220824
rect 194874 220768 194876 220788
rect 194876 220768 194928 220788
rect 194928 220768 194930 220788
rect 196070 220788 196126 220824
rect 196070 220768 196072 220788
rect 196072 220768 196124 220788
rect 196124 220768 196126 220788
rect 202602 225120 202658 225176
rect 203522 222400 203578 222456
rect 205086 225156 205088 225176
rect 205088 225156 205140 225176
rect 205140 225156 205142 225176
rect 205086 225120 205142 225156
rect 205086 222400 205142 222456
rect 484858 219544 484914 219600
rect 487066 220904 487122 220960
rect 487434 219272 487490 219328
rect 488906 217232 488962 217288
rect 489918 218592 489974 218648
rect 491206 218592 491262 218648
rect 490654 218048 490710 218104
rect 494886 219680 494942 219736
rect 494702 217640 494758 217696
rect 495162 217640 495218 217696
rect 497462 218592 497518 218648
rect 500406 218320 500462 218376
rect 498842 217232 498898 217288
rect 501326 217504 501382 217560
rect 501326 216960 501382 217016
rect 503166 219136 503222 219192
rect 502982 217776 503038 217832
rect 501694 217504 501750 217560
rect 503626 217776 503682 217832
rect 505926 221176 505982 221232
rect 505190 218864 505246 218920
rect 505098 217504 505154 217560
rect 507214 219156 507270 219192
rect 507214 219136 507216 219156
rect 507216 219136 507268 219156
rect 507268 219136 507270 219156
rect 507398 219136 507454 219192
rect 509238 219136 509294 219192
rect 509514 219156 509570 219192
rect 509514 219136 509516 219156
rect 509516 219136 509568 219156
rect 509568 219136 509570 219156
rect 509238 218864 509294 218920
rect 508042 217796 508098 217832
rect 508042 217776 508044 217796
rect 508044 217776 508096 217796
rect 508096 217776 508098 217796
rect 508226 217776 508282 217832
rect 509330 217776 509386 217832
rect 509514 217796 509570 217832
rect 509514 217776 509516 217796
rect 509516 217776 509568 217796
rect 509568 217776 509570 217796
rect 517794 221448 517850 221504
rect 517978 221448 518034 221504
rect 518990 219136 519046 219192
rect 519174 219172 519176 219192
rect 519176 219172 519228 219192
rect 519228 219172 519230 219192
rect 519174 219136 519230 219172
rect 518852 218864 518908 218920
rect 518714 218728 518770 218784
rect 518852 218628 518854 218648
rect 518854 218628 518906 218648
rect 518906 218628 518908 218648
rect 518852 218592 518908 218628
rect 518990 217232 519046 217288
rect 519174 217232 519230 217288
rect 519726 221720 519782 221776
rect 528558 218592 528614 218648
rect 528742 218592 528798 218648
rect 528650 217776 528706 217832
rect 528282 217232 528338 217288
rect 528466 217232 528522 217288
rect 529110 217796 529166 217832
rect 529110 217776 529112 217796
rect 529112 217776 529164 217796
rect 529164 217776 529166 217796
rect 532698 220380 532754 220416
rect 532698 220360 532700 220380
rect 532700 220360 532752 220380
rect 532752 220360 532754 220380
rect 534170 220380 534226 220416
rect 534170 220360 534172 220380
rect 534172 220360 534224 220380
rect 534224 220360 534226 220380
rect 534078 218592 534134 218648
rect 534262 218592 534318 218648
rect 534078 217232 534134 217288
rect 534262 217232 534318 217288
rect 495162 216688 495218 216744
rect 543922 220224 543978 220280
rect 544934 219952 544990 220008
rect 543462 217232 543518 217288
rect 543646 217232 543702 217288
rect 547142 220224 547198 220280
rect 548338 220632 548394 220688
rect 552386 220632 552442 220688
rect 552846 220224 552902 220280
rect 553674 220360 553730 220416
rect 554042 220632 554098 220688
rect 553352 219952 553408 220008
rect 554042 218320 554098 218376
rect 554226 218320 554282 218376
rect 554594 220224 554650 220280
rect 562874 222264 562930 222320
rect 562322 221992 562378 222048
rect 562690 222012 562746 222048
rect 562690 221992 562692 222012
rect 562692 221992 562744 222012
rect 562744 221992 562746 222012
rect 563334 222264 563390 222320
rect 563518 222012 563574 222048
rect 563518 221992 563520 222012
rect 563520 221992 563572 222012
rect 563572 221992 563574 222012
rect 564898 222264 564954 222320
rect 565082 221992 565138 222048
rect 563426 220632 563482 220688
rect 563242 220496 563298 220552
rect 563794 220360 563850 220416
rect 563610 220088 563666 220144
rect 540150 216416 540206 216472
rect 557078 216436 557134 216472
rect 557078 216416 557080 216436
rect 557080 216416 557132 216436
rect 557132 216416 557134 216436
rect 557722 216416 557778 216472
rect 558550 216436 558606 216472
rect 564070 219850 564126 219906
rect 564622 220088 564678 220144
rect 567198 222264 567254 222320
rect 570510 222536 570566 222592
rect 571062 221992 571118 222048
rect 570878 219850 570934 219906
rect 558550 216416 558552 216436
rect 558552 216416 558604 216436
rect 558604 216416 558606 216436
rect 572442 222264 572498 222320
rect 572626 220496 572682 220552
rect 572810 220224 572866 220280
rect 573454 220224 573510 220280
rect 573914 220224 573970 220280
rect 573270 219952 573326 220008
rect 572350 218320 572406 218376
rect 572534 218048 572590 218104
rect 571890 217776 571946 217832
rect 572166 217776 572222 217832
rect 572902 217776 572958 217832
rect 574834 222536 574890 222592
rect 575202 220632 575258 220688
rect 576030 221992 576086 222048
rect 591946 222012 592002 222048
rect 591946 221992 591948 222012
rect 591948 221992 592000 222012
rect 592000 221992 592002 222012
rect 578238 220360 578294 220416
rect 592038 220360 592094 220416
rect 582746 220244 582802 220280
rect 582746 220224 582748 220244
rect 582748 220224 582800 220244
rect 582800 220224 582802 220244
rect 591854 220224 591910 220280
rect 582010 219952 582066 220008
rect 582562 219952 582618 220008
rect 592038 219972 592094 220008
rect 592038 219952 592040 219972
rect 592040 219952 592092 219972
rect 592092 219952 592094 219972
rect 582102 218048 582158 218104
rect 582562 218048 582618 218104
rect 582562 217776 582618 217832
rect 582746 217776 582802 217832
rect 591946 217504 592002 217560
rect 590106 216688 590162 216744
rect 578882 213968 578938 214024
rect 578514 211676 578570 211712
rect 578514 211656 578516 211676
rect 578516 211656 578568 211676
rect 578568 211656 578570 211676
rect 579250 209788 579252 209808
rect 579252 209788 579304 209808
rect 579304 209788 579306 209808
rect 579250 209752 579306 209788
rect 599306 222012 599362 222048
rect 599306 221992 599308 222012
rect 599308 221992 599360 222012
rect 599360 221992 599362 222012
rect 597926 221176 597982 221232
rect 596362 217504 596418 217560
rect 594798 213152 594854 213208
rect 596822 217232 596878 217288
rect 597466 216960 597522 217016
rect 599306 220360 599362 220416
rect 601422 218356 601424 218376
rect 601424 218356 601476 218376
rect 601476 218356 601478 218376
rect 601422 218320 601478 218356
rect 601606 218320 601662 218376
rect 601422 218048 601478 218104
rect 600962 216960 601018 217016
rect 601652 217540 601654 217560
rect 601654 217540 601706 217560
rect 601706 217540 601708 217560
rect 601652 217504 601708 217540
rect 603262 217504 603318 217560
rect 601514 217096 601570 217152
rect 601790 217116 601846 217152
rect 601790 217096 601792 217116
rect 601792 217096 601844 217116
rect 601844 217096 601846 217116
rect 601330 216824 601386 216880
rect 601790 216824 601846 216880
rect 602526 216416 602582 216472
rect 606206 218864 606262 218920
rect 606758 218592 606814 218648
rect 606758 218048 606814 218104
rect 618258 221720 618314 221776
rect 616878 221448 616934 221504
rect 611450 220904 611506 220960
rect 612738 218864 612794 218920
rect 617338 219136 617394 219192
rect 623962 218320 624018 218376
rect 626630 216144 626686 216200
rect 630770 219680 630826 219736
rect 627734 218592 627790 218648
rect 631230 219408 631286 219464
rect 652206 298424 652262 298480
rect 640246 231376 640302 231432
rect 639602 230152 639658 230208
rect 637486 229744 637542 229800
rect 637670 220088 637726 220144
rect 650642 225528 650698 225584
rect 643190 220360 643246 220416
rect 640430 218864 640486 218920
rect 643006 215872 643062 215928
rect 645490 218592 645546 218648
rect 646870 217504 646926 217560
rect 646594 216416 646650 216472
rect 647146 213152 647202 213208
rect 649906 217776 649962 217832
rect 648526 214512 648582 214568
rect 651286 223080 651342 223136
rect 651102 216144 651158 216200
rect 651838 222808 651894 222864
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 666282 742464 666338 742520
rect 666466 711592 666522 711648
rect 666466 699760 666522 699816
rect 666282 665488 666338 665544
rect 665822 626048 665878 626104
rect 668214 782448 668270 782504
rect 667846 750760 667902 750816
rect 667846 743144 667902 743200
rect 667202 671064 667258 671120
rect 668398 734712 668454 734768
rect 668398 733080 668454 733136
rect 668214 710368 668270 710424
rect 668030 686160 668086 686216
rect 667846 665216 667902 665272
rect 667846 661000 667902 661056
rect 666466 621152 666522 621208
rect 666466 608776 666522 608832
rect 664442 579672 664498 579728
rect 663062 538736 663118 538792
rect 660302 405592 660358 405648
rect 659106 360032 659162 360088
rect 664626 491680 664682 491736
rect 661866 406272 661922 406328
rect 663062 315424 663118 315480
rect 661682 268096 661738 268152
rect 667202 534384 667258 534440
rect 666466 531392 666522 531448
rect 666006 493992 666062 494048
rect 665822 358672 665878 358728
rect 664442 271088 664498 271144
rect 666190 236136 666246 236192
rect 663246 234096 663302 234152
rect 658922 233824 658978 233880
rect 660946 229472 661002 229528
rect 652758 226344 652814 226400
rect 660210 225256 660266 225312
rect 655426 224984 655482 225040
rect 653034 220632 653090 220688
rect 655242 219136 655298 219192
rect 658186 224440 658242 224496
rect 656622 223624 656678 223680
rect 658002 221448 658058 221504
rect 658922 223896 658978 223952
rect 659382 221176 659438 221232
rect 661682 229200 661738 229256
rect 661498 213424 661554 213480
rect 663062 231648 663118 231704
rect 663246 230832 663302 230888
rect 664442 230560 664498 230616
rect 663430 220360 663486 220416
rect 663430 219544 663486 219600
rect 664902 215056 664958 215112
rect 664718 213696 664774 213752
rect 665270 231104 665326 231160
rect 665270 221992 665326 222048
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 579526 198872 579582 198928
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 579526 192208 579582 192264
rect 589462 191664 589518 191720
rect 579526 190712 579582 190768
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 579526 187992 579582 188048
rect 589462 186768 589518 186824
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 589462 185136 589518 185192
rect 579526 184320 579582 184376
rect 589462 183504 589518 183560
rect 579526 181872 579582 181928
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 578790 180104 578846 180160
rect 589462 178608 589518 178664
rect 579526 177656 579582 177712
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 579526 171012 579582 171048
rect 579526 170992 579528 171012
rect 579528 170992 579580 171012
rect 579580 170992 579582 171012
rect 578330 169224 578386 169280
rect 578974 166912 579030 166968
rect 578882 164464 578938 164520
rect 579434 162424 579490 162480
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589462 170448 589518 170504
rect 579250 159840 579306 159896
rect 579158 158208 579214 158264
rect 579526 155916 579582 155952
rect 579526 155896 579528 155916
rect 579528 155896 579580 155916
rect 579580 155896 579582 155916
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 578238 153992 578294 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147192 579582 147248
rect 578514 142976 578570 143032
rect 578698 138760 578754 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589462 157412 589518 157448
rect 589462 157392 589464 157412
rect 589464 157392 589516 157412
rect 589516 157392 589518 157412
rect 579526 140564 579528 140584
rect 579528 140564 579580 140584
rect 579580 140564 579582 140584
rect 579526 140528 579582 140564
rect 578882 136584 578938 136640
rect 578330 134408 578386 134464
rect 578238 132232 578294 132288
rect 578330 127744 578386 127800
rect 579526 129684 579528 129704
rect 579528 129684 579580 129704
rect 579580 129684 579582 129704
rect 579526 129648 579582 129684
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 589462 150864 589518 150920
rect 589186 149232 589242 149288
rect 579250 125296 579306 125352
rect 579250 123528 579306 123584
rect 579066 121116 579068 121136
rect 579068 121116 579120 121136
rect 579120 121116 579122 121136
rect 579066 121080 579122 121116
rect 578514 118360 578570 118416
rect 578330 108332 578332 108352
rect 578332 108332 578384 108352
rect 578384 108332 578386 108352
rect 578330 108296 578386 108332
rect 578330 105848 578386 105904
rect 578698 95004 578700 95024
rect 578700 95004 578752 95024
rect 578752 95004 578754 95024
rect 578698 94968 578754 95004
rect 578606 86400 578662 86456
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579526 114436 579582 114472
rect 579526 114416 579528 114436
rect 579528 114416 579580 114436
rect 579580 114416 579582 114436
rect 579526 112648 579582 112704
rect 579434 110236 579436 110256
rect 579436 110236 579488 110256
rect 579488 110236 579490 110256
rect 579434 110200 579490 110236
rect 579526 103300 579528 103320
rect 579528 103300 579580 103320
rect 579580 103300 579582 103320
rect 579526 103264 579582 103300
rect 579250 101768 579306 101824
rect 579526 99204 579582 99240
rect 579526 99184 579528 99204
rect 579528 99184 579580 99204
rect 579580 99184 579582 99204
rect 579526 97452 579528 97472
rect 579528 97452 579580 97472
rect 579580 97452 579582 97472
rect 579526 97416 579582 97452
rect 579526 93064 579582 93120
rect 579066 90888 579122 90944
rect 579526 88032 579582 88088
rect 579250 83952 579306 84008
rect 579250 82184 579306 82240
rect 578790 80008 578846 80064
rect 578974 77832 579030 77888
rect 578698 75420 578700 75440
rect 578700 75420 578752 75440
rect 578752 75420 578754 75440
rect 578698 75384 578754 75420
rect 578514 73108 578516 73128
rect 578516 73108 578568 73128
rect 578568 73108 578570 73128
rect 578514 73072 578570 73108
rect 578514 61784 578570 61840
rect 589370 147600 589426 147656
rect 589462 145968 589518 146024
rect 589922 144336 589978 144392
rect 589462 142704 589518 142760
rect 589094 141072 589150 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589278 136176 589334 136232
rect 589462 134544 589518 134600
rect 588542 132912 588598 132968
rect 590106 131280 590162 131336
rect 589462 129648 589518 129704
rect 589462 128016 589518 128072
rect 589922 126384 589978 126440
rect 589462 124752 589518 124808
rect 589462 123120 589518 123176
rect 589462 121508 589518 121544
rect 589462 121488 589464 121508
rect 589464 121488 589516 121508
rect 589516 121488 589518 121508
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 590106 119856 590162 119912
rect 589830 114960 589886 115016
rect 589370 111696 589426 111752
rect 589646 110064 589702 110120
rect 589462 108432 589518 108488
rect 666466 186904 666522 186960
rect 668950 783808 669006 783864
rect 668766 755928 668822 755984
rect 668766 731448 668822 731504
rect 668582 670384 668638 670440
rect 670514 873976 670570 874032
rect 669594 872208 669650 872264
rect 669778 789384 669834 789440
rect 669594 755384 669650 755440
rect 669226 753480 669282 753536
rect 669410 741784 669466 741840
rect 669134 734440 669190 734496
rect 668950 708736 669006 708792
rect 668766 664536 668822 664592
rect 669226 701120 669282 701176
rect 669042 662496 669098 662552
rect 668398 659640 668454 659696
rect 668214 647264 668270 647320
rect 668030 621696 668086 621752
rect 668398 607960 668454 608016
rect 668214 574776 668270 574832
rect 668214 557504 668270 557560
rect 668950 638696 669006 638752
rect 668766 593544 668822 593600
rect 668582 535880 668638 535936
rect 668398 530576 668454 530632
rect 669594 738520 669650 738576
rect 670330 780000 670386 780056
rect 670146 778912 670202 778968
rect 670146 777008 670202 777064
rect 670146 774968 670202 775024
rect 669962 715672 670018 715728
rect 669778 709552 669834 709608
rect 670514 754160 670570 754216
rect 671158 867176 671214 867232
rect 670974 778368 671030 778424
rect 670974 776464 671030 776520
rect 670882 757424 670938 757480
rect 670698 734032 670754 734088
rect 670698 728476 670754 728512
rect 670698 728456 670700 728476
rect 670700 728456 670752 728476
rect 670752 728456 670754 728476
rect 671342 763000 671398 763056
rect 671618 760280 671674 760336
rect 671618 759872 671674 759928
rect 671158 753344 671214 753400
rect 671066 751304 671122 751360
rect 671434 750080 671490 750136
rect 671250 737024 671306 737080
rect 671066 728048 671122 728104
rect 670882 713224 670938 713280
rect 670330 707104 670386 707160
rect 670146 705880 670202 705936
rect 669778 696904 669834 696960
rect 669594 666304 669650 666360
rect 669410 663312 669466 663368
rect 669226 621968 669282 622024
rect 670422 690376 670478 690432
rect 670238 685344 670294 685400
rect 669778 620608 669834 620664
rect 669778 616120 669834 616176
rect 669226 608504 669282 608560
rect 668950 574368 669006 574424
rect 669042 564440 669098 564496
rect 668766 528536 668822 528592
rect 668214 485968 668270 486024
rect 669594 554648 669650 554704
rect 669226 528944 669282 529000
rect 669042 485016 669098 485072
rect 669594 482704 669650 482760
rect 667846 456048 667902 456104
rect 671066 712816 671122 712872
rect 671066 712408 671122 712464
rect 670882 668208 670938 668264
rect 670882 667936 670938 667992
rect 670606 659912 670662 659968
rect 670422 620200 670478 620256
rect 670238 615712 670294 615768
rect 670422 614896 670478 614952
rect 670238 600616 670294 600672
rect 669962 580080 670018 580136
rect 670054 553968 670110 554024
rect 670054 551520 670110 551576
rect 669778 455096 669834 455152
rect 667202 313656 667258 313712
rect 667018 225256 667074 225312
rect 667018 224188 667074 224224
rect 667018 224168 667020 224188
rect 667020 224168 667072 224188
rect 667072 224168 667074 224188
rect 666834 222808 666890 222864
rect 666834 217232 666890 217288
rect 666834 198328 666890 198384
rect 666650 178744 666706 178800
rect 666190 160112 666246 160168
rect 670238 530032 670294 530088
rect 669962 403688 670018 403744
rect 671066 666576 671122 666632
rect 671434 728320 671490 728376
rect 672446 936400 672502 936456
rect 672630 935720 672686 935776
rect 673090 933136 673146 933192
rect 675666 966456 675722 966512
rect 675758 965096 675814 965152
rect 675298 964688 675354 964744
rect 675482 963328 675538 963384
rect 674286 962784 674342 962840
rect 674102 957072 674158 957128
rect 673366 932864 673422 932920
rect 673182 930688 673238 930744
rect 675482 962784 675538 962840
rect 675114 960744 675170 960800
rect 674930 959112 674986 959168
rect 674654 958704 674710 958760
rect 674470 933816 674526 933872
rect 674286 932592 674342 932648
rect 675206 958704 675262 958760
rect 675298 957752 675354 957808
rect 675758 957752 675814 957808
rect 675482 957072 675538 957128
rect 675758 956392 675814 956448
rect 675206 954624 675262 954680
rect 674838 953400 674894 953456
rect 674654 930416 674710 930472
rect 674102 930144 674158 930200
rect 675482 953400 675538 953456
rect 675574 952176 675630 952232
rect 683302 950680 683358 950736
rect 679622 949456 679678 949512
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 676494 937624 676550 937680
rect 676494 936808 676550 936864
rect 679622 935584 679678 935640
rect 683118 947280 683174 947336
rect 683118 939664 683174 939720
rect 682382 935176 682438 935232
rect 675298 934632 675354 934688
rect 675114 934088 675170 934144
rect 683302 932320 683358 932376
rect 683118 929056 683174 929112
rect 673366 928240 673422 928296
rect 673090 868400 673146 868456
rect 672630 784216 672686 784272
rect 671802 759464 671858 759520
rect 671802 758240 671858 758296
rect 671618 715264 671674 715320
rect 671618 714856 671674 714912
rect 671434 714040 671490 714096
rect 672354 758648 672410 758704
rect 672170 757832 672226 757888
rect 672262 743416 672318 743472
rect 672078 741104 672134 741160
rect 671986 730496 672042 730552
rect 671802 713632 671858 713688
rect 671802 687384 671858 687440
rect 671618 670112 671674 670168
rect 671434 669840 671490 669896
rect 671618 669432 671674 669488
rect 671434 668616 671490 668672
rect 671250 661272 671306 661328
rect 671066 624688 671122 624744
rect 670882 623464 670938 623520
rect 670882 622784 670938 622840
rect 671986 666032 672042 666088
rect 672906 773744 672962 773800
rect 672722 759056 672778 759112
rect 672722 714448 672778 714504
rect 673090 751712 673146 751768
rect 673090 733624 673146 733680
rect 672906 709960 672962 710016
rect 672538 709144 672594 709200
rect 672446 685888 672502 685944
rect 672262 665760 672318 665816
rect 672078 663856 672134 663912
rect 671986 654200 672042 654256
rect 671894 643456 671950 643512
rect 671618 625096 671674 625152
rect 671250 624280 671306 624336
rect 671618 622376 671674 622432
rect 671434 618160 671490 618216
rect 671066 594768 671122 594824
rect 670882 577632 670938 577688
rect 670882 552064 670938 552120
rect 671434 580488 671490 580544
rect 671342 578856 671398 578912
rect 671526 578040 671582 578096
rect 671342 576816 671398 576872
rect 671710 577224 671766 577280
rect 672262 623872 672318 623928
rect 672630 666984 672686 667040
rect 675022 879144 675078 879200
rect 675482 877648 675538 877704
rect 675022 877240 675078 877296
rect 675390 877240 675446 877296
rect 675758 875880 675814 875936
rect 675482 873976 675538 874032
rect 675666 873976 675722 874032
rect 674010 867992 674066 868048
rect 673734 779184 673790 779240
rect 673550 777416 673606 777472
rect 673366 728340 673422 728376
rect 673366 728320 673368 728340
rect 673368 728320 673420 728340
rect 673420 728320 673422 728340
rect 673366 728084 673368 728104
rect 673368 728084 673420 728104
rect 673420 728084 673422 728104
rect 673366 728048 673422 728084
rect 675114 872208 675170 872264
rect 675574 872208 675630 872264
rect 675114 869488 675170 869544
rect 675298 868672 675354 868728
rect 675114 867992 675170 868048
rect 674930 866632 674986 866688
rect 674654 864728 674710 864784
rect 674470 854256 674526 854312
rect 674470 788024 674526 788080
rect 674286 782992 674342 783048
rect 674194 778640 674250 778696
rect 673918 770616 673974 770672
rect 674286 727912 674342 727968
rect 674102 726824 674158 726880
rect 675482 868400 675538 868456
rect 675482 867176 675538 867232
rect 675206 864728 675262 864784
rect 675206 789384 675262 789440
rect 675390 788024 675446 788080
rect 674838 787208 674894 787264
rect 675390 786664 675446 786720
rect 675482 784216 675538 784272
rect 675482 783808 675538 783864
rect 674930 783264 674986 783320
rect 675390 782992 675446 783048
rect 675114 782720 675170 782776
rect 675298 782448 675354 782504
rect 675114 780680 675170 780736
rect 674746 771976 674802 772032
rect 675482 780000 675538 780056
rect 675298 779184 675354 779240
rect 675482 778640 675538 778696
rect 675482 777416 675538 777472
rect 675390 777008 675446 777064
rect 675482 776464 675538 776520
rect 675482 774968 675538 775024
rect 675482 773744 675538 773800
rect 682382 772656 682438 772712
rect 681002 768712 681058 768768
rect 675206 766536 675262 766592
rect 674838 765040 674894 765096
rect 676034 763000 676090 763056
rect 676586 761732 676642 761788
rect 676954 761776 677010 761832
rect 676034 760688 676090 760744
rect 675850 754704 675906 754760
rect 681002 757016 681058 757072
rect 683210 771976 683266 772032
rect 683394 770616 683450 770672
rect 683210 756608 683266 756664
rect 682382 755792 682438 755848
rect 676954 754976 677010 755032
rect 676034 752528 676090 752584
rect 683394 752936 683450 752992
rect 683118 752120 683174 752176
rect 674930 743416 674986 743472
rect 675114 743144 675170 743200
rect 675022 742464 675078 742520
rect 674838 741784 674894 741840
rect 675114 741512 675170 741568
rect 674930 741104 674986 741160
rect 675298 738520 675354 738576
rect 675114 737024 675170 737080
rect 675482 738112 675538 738168
rect 674930 734712 674986 734768
rect 674654 733080 674710 733136
rect 675114 734440 675170 734496
rect 675114 733624 675170 733680
rect 675114 732808 675170 732864
rect 674654 731448 674710 731504
rect 675114 730496 675170 730552
rect 683762 727912 683818 727968
rect 683210 726688 683266 726744
rect 674746 726552 674802 726608
rect 682382 725736 682438 725792
rect 673734 725056 673790 725112
rect 682382 710776 682438 710832
rect 673550 708328 673606 708384
rect 683394 726416 683450 726472
rect 683578 725056 683634 725112
rect 683394 711184 683450 711240
rect 683578 707920 683634 707976
rect 683762 707512 683818 707568
rect 683210 706696 683266 706752
rect 674378 706288 674434 706344
rect 674010 693096 674066 693152
rect 673458 690104 673514 690160
rect 673274 689016 673330 689072
rect 673090 661544 673146 661600
rect 673090 648624 673146 648680
rect 672814 647808 672870 647864
rect 672630 635432 672686 635488
rect 673826 644544 673882 644600
rect 673642 641688 673698 641744
rect 673458 636792 673514 636848
rect 672630 621832 672686 621888
rect 672630 621152 672686 621208
rect 672446 619792 672502 619848
rect 672630 597352 672686 597408
rect 672446 578584 672502 578640
rect 671986 574096 672042 574152
rect 671802 571104 671858 571160
rect 671710 570288 671766 570344
rect 671250 534792 671306 534848
rect 671434 533432 671490 533488
rect 671526 532616 671582 532672
rect 671526 529352 671582 529408
rect 671526 528536 671582 528592
rect 671066 525680 671122 525736
rect 671986 569472 672042 569528
rect 671710 500928 671766 500984
rect 670882 483928 670938 483984
rect 670606 455776 670662 455832
rect 670422 455368 670478 455424
rect 672262 559408 672318 559464
rect 672446 534520 672502 534576
rect 673274 616528 673330 616584
rect 672998 579128 673054 579184
rect 673366 604288 673422 604344
rect 673090 573144 673146 573200
rect 672814 571920 672870 571976
rect 673090 553424 673146 553480
rect 672814 534248 672870 534304
rect 672446 531800 672502 531856
rect 672630 528128 672686 528184
rect 672906 490864 672962 490920
rect 672906 489640 672962 489696
rect 672722 489232 672778 489288
rect 672446 488416 672502 488472
rect 672446 488008 672502 488064
rect 672170 484744 672226 484800
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 670146 360848 670202 360904
rect 670146 348472 670202 348528
rect 669962 347248 670018 347304
rect 668582 311888 668638 311944
rect 669226 302232 669282 302288
rect 667386 181328 667442 181384
rect 668214 230560 668270 230616
rect 667846 223080 667902 223136
rect 667846 220904 667902 220960
rect 668030 197376 668086 197432
rect 668122 194148 668124 194168
rect 668124 194148 668176 194168
rect 668176 194148 668178 194168
rect 668122 194112 668178 194148
rect 668030 192516 668032 192536
rect 668032 192516 668084 192536
rect 668084 192516 668086 192536
rect 668030 192480 668086 192516
rect 668122 192208 668178 192264
rect 668122 187584 668178 187640
rect 668030 184356 668032 184376
rect 668032 184356 668084 184376
rect 668084 184356 668086 184376
rect 668030 184320 668086 184356
rect 668582 230424 668638 230480
rect 668582 229200 668638 229256
rect 668306 182688 668362 182744
rect 667846 176432 667902 176488
rect 667938 174528 667994 174584
rect 668030 164772 668032 164792
rect 668032 164772 668084 164792
rect 668084 164772 668086 164792
rect 668030 164736 668086 164772
rect 669410 231548 669412 231568
rect 669412 231548 669464 231568
rect 669464 231548 669466 231568
rect 669410 231512 669466 231548
rect 669226 212336 669282 212392
rect 669226 211928 669282 211984
rect 669042 211792 669098 211848
rect 668950 211248 669006 211304
rect 669226 190304 669282 190360
rect 669134 189252 669136 189272
rect 669136 189252 669188 189272
rect 669188 189252 669190 189272
rect 669134 189216 669190 189252
rect 669134 185544 669190 185600
rect 669134 169632 669190 169688
rect 669778 169496 669834 169552
rect 669594 168272 669650 168328
rect 669042 168000 669098 168056
rect 668950 163104 669006 163160
rect 668766 153312 668822 153368
rect 668674 150048 668730 150104
rect 668490 148416 668546 148472
rect 668766 147736 668822 147792
rect 667570 135904 667626 135960
rect 667938 135360 667994 135416
rect 667202 134544 667258 134600
rect 667018 133048 667074 133104
rect 668582 128152 668638 128208
rect 669134 138624 669190 138680
rect 669778 152632 669834 152688
rect 672262 400424 672318 400480
rect 673458 598440 673514 598496
rect 673274 528672 673330 528728
rect 673642 593136 673698 593192
rect 674194 692824 674250 692880
rect 675114 701120 675170 701176
rect 674838 699760 674894 699816
rect 674562 697176 674618 697232
rect 675114 697176 675170 697232
rect 674746 696904 674802 696960
rect 675666 694320 675722 694376
rect 675482 693096 675538 693152
rect 675114 692824 675170 692880
rect 675114 690376 675170 690432
rect 675390 690104 675446 690160
rect 674562 689696 674618 689752
rect 674930 689288 674986 689344
rect 674286 650256 674342 650312
rect 674194 649576 674250 649632
rect 674194 645088 674250 645144
rect 674194 635704 674250 635760
rect 674746 688744 674802 688800
rect 675114 689016 675170 689072
rect 675114 687384 675170 687440
rect 675114 686160 675170 686216
rect 674930 685888 674986 685944
rect 675114 685344 675170 685400
rect 674470 623192 674526 623248
rect 683210 682352 683266 682408
rect 676494 673104 676550 673160
rect 676494 671064 676550 671120
rect 676494 669840 676550 669896
rect 676494 669432 676550 669488
rect 674838 667392 674894 667448
rect 683394 680992 683450 681048
rect 683210 666984 683266 667040
rect 674838 666576 674894 666632
rect 683394 663312 683450 663368
rect 674838 661816 674894 661872
rect 674838 661272 674894 661328
rect 675298 660184 675354 660240
rect 675298 659640 675354 659696
rect 675206 654200 675262 654256
rect 675390 652840 675446 652896
rect 675482 651480 675538 651536
rect 675390 648896 675446 648952
rect 675114 648624 675170 648680
rect 675390 647808 675446 647864
rect 675114 647264 675170 647320
rect 675758 644680 675814 644736
rect 675114 644544 675170 644600
rect 675114 643864 675170 643920
rect 675390 643456 675446 643512
rect 675298 641688 675354 641744
rect 675390 640464 675446 640520
rect 675482 638696 675538 638752
rect 675758 638016 675814 638072
rect 675574 637744 675630 637800
rect 675206 637608 675262 637664
rect 675574 632984 675630 633040
rect 683394 636792 683450 636848
rect 674930 629720 674986 629776
rect 674470 622104 674526 622160
rect 674470 620880 674526 620936
rect 674286 619384 674342 619440
rect 674010 617344 674066 617400
rect 674838 608776 674894 608832
rect 675022 608504 675078 608560
rect 675022 607688 675078 607744
rect 674838 607144 674894 607200
rect 674654 604560 674710 604616
rect 674010 603472 674066 603528
rect 673826 591232 673882 591288
rect 673826 580760 673882 580816
rect 673826 579672 673882 579728
rect 673826 558320 673882 558376
rect 673642 548392 673698 548448
rect 673458 526496 673514 526552
rect 673642 485560 673698 485616
rect 674286 600072 674342 600128
rect 674010 547032 674066 547088
rect 674470 598984 674526 599040
rect 674286 545672 674342 545728
rect 674194 533160 674250 533216
rect 674010 532888 674066 532944
rect 674838 602248 674894 602304
rect 675758 631352 675814 631408
rect 675850 627816 675906 627872
rect 676494 625640 676550 625696
rect 683118 623192 683174 623248
rect 683118 617888 683174 617944
rect 683578 635704 683634 635760
rect 683762 635432 683818 635488
rect 683762 622784 683818 622840
rect 683578 618704 683634 618760
rect 683394 617072 683450 617128
rect 675482 607960 675538 608016
rect 675482 607688 675538 607744
rect 675482 607144 675538 607200
rect 675482 604560 675538 604616
rect 675482 604288 675538 604344
rect 675482 603472 675538 603528
rect 675482 602928 675538 602984
rect 675390 602248 675446 602304
rect 675114 600616 675170 600672
rect 675114 600072 675170 600128
rect 675114 599528 675170 599584
rect 674930 596672 674986 596728
rect 675298 598984 675354 599040
rect 675482 598440 675538 598496
rect 675390 597352 675446 597408
rect 674930 594360 674986 594416
rect 675298 594768 675354 594824
rect 675022 593816 675078 593872
rect 674838 580488 674894 580544
rect 674838 579808 674894 579864
rect 674838 579400 674894 579456
rect 674838 578856 674894 578912
rect 675390 593544 675446 593600
rect 675850 592864 675906 592920
rect 683486 592864 683542 592920
rect 674930 575320 674986 575376
rect 674838 559680 674894 559736
rect 674930 557504 674986 557560
rect 674930 555736 674986 555792
rect 675482 578312 675538 578368
rect 675298 577632 675354 577688
rect 675482 576952 675538 577008
rect 675298 576816 675354 576872
rect 683302 592592 683358 592648
rect 676034 592320 676090 592376
rect 681002 590552 681058 590608
rect 675850 576544 675906 576600
rect 681002 576000 681058 576056
rect 683118 591232 683174 591288
rect 683302 573960 683358 574016
rect 683486 573144 683542 573200
rect 683118 571920 683174 571976
rect 682382 570696 682438 570752
rect 675298 564440 675354 564496
rect 675482 562672 675538 562728
rect 675482 561176 675538 561232
rect 675298 559680 675354 559736
rect 675390 559408 675446 559464
rect 675390 558320 675446 558376
rect 675758 557640 675814 557696
rect 675482 555736 675538 555792
rect 675390 554648 675446 554704
rect 675758 553968 675814 554024
rect 675390 553424 675446 553480
rect 675390 552064 675446 552120
rect 675390 551520 675446 551576
rect 675022 550432 675078 550488
rect 675758 550160 675814 550216
rect 675482 548392 675538 548448
rect 675942 547612 675944 547632
rect 675944 547612 675996 547632
rect 675996 547612 675998 547632
rect 675942 547576 675998 547612
rect 677414 547576 677470 547632
rect 674838 544448 674894 544504
rect 674838 543904 674894 543960
rect 674654 530304 674710 530360
rect 674470 527720 674526 527776
rect 674194 490048 674250 490104
rect 673826 484336 673882 484392
rect 675298 544856 675354 544912
rect 675482 543904 675538 543960
rect 676034 538736 676090 538792
rect 676034 535676 676090 535732
rect 675758 534520 675814 534576
rect 675758 534044 675814 534100
rect 675758 533636 675814 533692
rect 675758 533160 675814 533216
rect 676862 525680 676918 525736
rect 675482 513712 675538 513768
rect 675114 502560 675170 502616
rect 675298 486376 675354 486432
rect 676034 513712 676090 513768
rect 675850 502560 675906 502616
rect 676402 500928 676458 500984
rect 675850 493992 675906 494048
rect 676034 490456 676090 490512
rect 674930 482976 674986 483032
rect 673090 482296 673146 482352
rect 673274 474816 673330 474872
rect 674838 456320 674894 456376
rect 673458 456048 673514 456104
rect 673826 456068 673882 456104
rect 673826 456048 673828 456068
rect 673828 456048 673880 456068
rect 673880 456048 673882 456068
rect 673734 455812 673736 455832
rect 673736 455812 673788 455832
rect 673788 455812 673790 455832
rect 673734 455776 673790 455812
rect 673504 455388 673560 455424
rect 673504 455368 673506 455388
rect 673506 455368 673558 455388
rect 673558 455368 673560 455388
rect 673386 455132 673388 455152
rect 673388 455132 673440 455152
rect 673440 455132 673442 455152
rect 673386 455096 673442 455132
rect 673550 455096 673606 455152
rect 673044 454844 673100 454880
rect 673044 454824 673046 454844
rect 673046 454824 673098 454844
rect 673098 454824 673100 454844
rect 672814 454436 672870 454472
rect 672814 454416 672816 454436
rect 672816 454416 672868 454436
rect 672868 454416 672870 454436
rect 672952 454180 672954 454200
rect 672954 454180 673006 454200
rect 673006 454180 673008 454200
rect 672952 454144 673008 454180
rect 675850 482976 675906 483032
rect 675666 480664 675722 480720
rect 675482 454824 675538 454880
rect 675850 456320 675906 456376
rect 675850 456084 675852 456104
rect 675852 456084 675904 456104
rect 675904 456084 675906 456104
rect 675850 456048 675906 456084
rect 675666 454416 675722 454472
rect 675942 454144 675998 454200
rect 674838 453872 674894 453928
rect 683394 547032 683450 547088
rect 683210 545672 683266 545728
rect 678242 531392 678298 531448
rect 683578 533840 683634 533896
rect 683394 528536 683450 528592
rect 683578 527312 683634 527368
rect 683210 526904 683266 526960
rect 677874 524456 677930 524512
rect 683578 503648 683634 503704
rect 679622 487600 679678 487656
rect 683394 503376 683450 503432
rect 683118 491272 683174 491328
rect 681002 486784 681058 486840
rect 683578 487192 683634 487248
rect 683394 483520 683450 483576
rect 677414 483112 677470 483168
rect 680358 481888 680414 481944
rect 683118 481072 683174 481128
rect 677138 475360 677194 475416
rect 676678 455096 676734 455152
rect 676126 453736 676182 453792
rect 676034 410488 676090 410544
rect 675850 405592 675906 405648
rect 675850 403416 675906 403472
rect 683118 406272 683174 406328
rect 683118 403280 683174 403336
rect 676034 402600 676090 402656
rect 674838 402192 674894 402248
rect 672630 401920 672686 401976
rect 672998 401648 673054 401704
rect 674838 401648 674894 401704
rect 672446 400016 672502 400072
rect 673182 401240 673238 401296
rect 672722 392536 672778 392592
rect 672262 355816 672318 355872
rect 672538 354592 672594 354648
rect 672170 349696 672226 349752
rect 671986 348880 672042 348936
rect 672354 347656 672410 347712
rect 672170 333920 672226 333976
rect 671986 332288 672042 332344
rect 672354 327528 672410 327584
rect 672538 309984 672594 310040
rect 672446 301416 672502 301472
rect 671342 269728 671398 269784
rect 671986 264016 672042 264072
rect 671710 262112 671766 262168
rect 671526 259664 671582 259720
rect 671342 258848 671398 258904
rect 670606 257624 670662 257680
rect 671526 245792 671582 245848
rect 671710 245520 671766 245576
rect 672262 257216 672318 257272
rect 671342 241440 671398 241496
rect 671894 238176 671950 238232
rect 670606 235864 670662 235920
rect 670514 232600 670570 232656
rect 670330 232056 670386 232112
rect 670146 165552 670202 165608
rect 668766 125568 668822 125624
rect 668582 120672 668638 120728
rect 668674 120128 668730 120184
rect 668030 117408 668086 117464
rect 669962 122712 670018 122768
rect 669226 119040 669282 119096
rect 668674 114144 668730 114200
rect 670514 227160 670570 227216
rect 670514 226752 670570 226808
rect 670514 226072 670570 226128
rect 670606 223896 670662 223952
rect 670514 223624 670570 223680
rect 670606 218864 670662 218920
rect 670606 218320 670662 218376
rect 670606 215736 670662 215792
rect 670606 201320 670662 201376
rect 670790 199008 670846 199064
rect 671342 225800 671398 225856
rect 671342 225392 671398 225448
rect 671250 225020 671252 225040
rect 671252 225020 671304 225040
rect 671304 225020 671306 225040
rect 671250 224984 671306 225020
rect 671250 224732 671306 224768
rect 671250 224712 671252 224732
rect 671252 224712 671304 224732
rect 671304 224712 671306 224732
rect 671250 220632 671306 220688
rect 671250 219816 671306 219872
rect 671250 219544 671306 219600
rect 671250 218864 671306 218920
rect 670606 171944 670662 172000
rect 671894 227024 671950 227080
rect 671894 226616 671950 226672
rect 672262 233144 672318 233200
rect 672262 228792 672318 228848
rect 672998 385192 673054 385248
rect 674654 399744 674710 399800
rect 674286 397296 674342 397352
rect 673366 396616 673422 396672
rect 673918 396072 673974 396128
rect 673734 395664 673790 395720
rect 673550 394304 673606 394360
rect 673550 385192 673606 385248
rect 673366 382200 673422 382256
rect 673090 379344 673146 379400
rect 674102 393624 674158 393680
rect 673918 381384 673974 381440
rect 673734 375400 673790 375456
rect 672998 357448 673054 357504
rect 673366 357040 673422 357096
rect 673182 356632 673238 356688
rect 673090 355408 673146 355464
rect 672906 351328 672962 351384
rect 672906 338000 672962 338056
rect 672906 312024 672962 312080
rect 673918 356224 673974 356280
rect 673550 352552 673606 352608
rect 673734 350512 673790 350568
rect 673550 336640 673606 336696
rect 673734 331064 673790 331120
rect 673274 312432 673330 312488
rect 673090 311208 673146 311264
rect 672906 267280 672962 267336
rect 673918 311616 673974 311672
rect 673274 310800 673330 310856
rect 673826 310392 673882 310448
rect 674470 394032 674526 394088
rect 674286 377984 674342 378040
rect 674470 376624 674526 376680
rect 676034 399336 676090 399392
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675298 379344 675354 379400
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675114 376624 675170 376680
rect 675114 375400 675170 375456
rect 675298 374992 675354 375048
rect 675758 372952 675814 373008
rect 675114 372544 675170 372600
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 355000 674710 355056
rect 676034 353776 676090 353832
rect 674746 353368 674802 353424
rect 674562 352144 674618 352200
rect 674378 349424 674434 349480
rect 674378 332696 674434 332752
rect 675942 349152 675998 349208
rect 675758 340176 675814 340232
rect 675390 338952 675446 339008
rect 675114 338000 675170 338056
rect 675574 337728 675630 337784
rect 675114 336640 675170 336696
rect 675758 336640 675814 336696
rect 675298 333920 675354 333976
rect 675114 332696 675170 332752
rect 675114 332288 675170 332344
rect 675758 332288 675814 332344
rect 675114 331064 675170 331120
rect 675758 328344 675814 328400
rect 675114 327528 675170 327584
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 309576 674710 309632
rect 673366 304272 673422 304328
rect 674470 305496 674526 305552
rect 674194 303864 674250 303920
rect 673366 287816 673422 287872
rect 673090 266464 673146 266520
rect 673090 266056 673146 266112
rect 672906 263744 672962 263800
rect 673918 265784 673974 265840
rect 673366 260480 673422 260536
rect 673642 259256 673698 259312
rect 673366 245248 673422 245304
rect 673918 258440 673974 258496
rect 673642 242800 673698 242856
rect 673090 239944 673146 240000
rect 673302 237108 673358 237144
rect 673302 237088 673304 237108
rect 673304 237088 673356 237108
rect 673356 237088 673358 237108
rect 673526 236700 673582 236736
rect 673526 236680 673528 236700
rect 673528 236680 673580 236700
rect 673580 236680 673582 236700
rect 673274 233552 673330 233608
rect 673734 232600 673790 232656
rect 673642 232056 673698 232112
rect 673458 230152 673514 230208
rect 673734 230152 673790 230208
rect 673274 229472 673330 229528
rect 673386 229200 673442 229256
rect 673734 229744 673790 229800
rect 672906 228928 672962 228984
rect 673550 228928 673606 228984
rect 672906 228556 672908 228576
rect 672908 228556 672960 228576
rect 672960 228556 672962 228576
rect 672906 228520 672962 228556
rect 673386 228540 673442 228576
rect 673386 228520 673388 228540
rect 673388 228520 673440 228540
rect 673440 228520 673442 228540
rect 672262 226752 672318 226808
rect 672032 226480 672088 226536
rect 671894 226364 671950 226400
rect 671894 226344 671896 226364
rect 671896 226344 671948 226364
rect 671948 226344 671950 226364
rect 671818 225700 671820 225720
rect 671820 225700 671872 225720
rect 671872 225700 671874 225720
rect 671818 225664 671874 225700
rect 672170 225664 672226 225720
rect 672078 224712 672134 224768
rect 671894 224440 671950 224496
rect 671894 219408 671950 219464
rect 672078 219136 672134 219192
rect 672170 216144 672226 216200
rect 672078 214104 672134 214160
rect 673182 226480 673238 226536
rect 672860 225664 672916 225720
rect 672906 224848 672962 224904
rect 672722 211928 672778 211984
rect 672722 211112 672778 211168
rect 672446 210432 672502 210488
rect 672262 202952 672318 203008
rect 672078 201048 672134 201104
rect 672722 210160 672778 210216
rect 672538 185544 672594 185600
rect 672262 183504 672318 183560
rect 672078 182008 672134 182064
rect 671894 174800 671950 174856
rect 671710 172896 671766 172952
rect 671894 169904 671950 169960
rect 671710 166912 671766 166968
rect 671526 158208 671582 158264
rect 670606 148960 670662 149016
rect 671342 131688 671398 131744
rect 590566 113328 590622 113384
rect 671526 130872 671582 130928
rect 668122 112512 668178 112568
rect 668306 111832 668362 111888
rect 668030 109248 668086 109304
rect 589922 106800 589978 106856
rect 589462 105168 589518 105224
rect 589462 101904 589518 101960
rect 666650 105984 666706 106040
rect 667202 105984 667258 106040
rect 590106 103536 590162 103592
rect 585782 77832 585838 77888
rect 579158 71304 579214 71360
rect 579526 68040 579582 68096
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579526 64504 579582 64560
rect 579526 60288 579582 60344
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 579526 56072 579582 56128
rect 581642 54984 581698 55040
rect 580262 54712 580318 54768
rect 625434 93064 625490 93120
rect 625434 91568 625490 91624
rect 635738 96872 635794 96928
rect 637026 96872 637082 96928
rect 626446 95376 626502 95432
rect 643190 95104 643246 95160
rect 626262 94424 626318 94480
rect 626446 93472 626502 93528
rect 626446 90616 626502 90672
rect 625802 89664 625858 89720
rect 626446 88848 626502 88904
rect 626446 87896 626502 87952
rect 643466 87080 643522 87136
rect 625618 86944 625674 87000
rect 626446 85992 626502 86048
rect 626446 85040 626502 85096
rect 625618 84124 625620 84144
rect 625620 84124 625672 84144
rect 625672 84124 625674 84144
rect 625618 84088 625674 84124
rect 624422 82864 624478 82920
rect 644018 89664 644074 89720
rect 644938 92112 644994 92168
rect 644754 84632 644810 84688
rect 643742 82728 643798 82784
rect 628654 81640 628710 81696
rect 629206 80824 629262 80880
rect 633898 80416 633954 80472
rect 639602 77832 639658 77888
rect 655242 94152 655298 94208
rect 655058 93336 655114 93392
rect 654874 92520 654930 92576
rect 654138 90616 654194 90672
rect 655426 91432 655482 91488
rect 655794 89800 655850 89856
rect 663706 91976 663762 92032
rect 664166 88984 664222 89040
rect 647054 74432 647110 74488
rect 646870 72936 646926 72992
rect 647330 69944 647386 70000
rect 646226 68856 646282 68912
rect 648986 71440 649042 71496
rect 649170 66952 649226 67008
rect 647514 65456 647570 65512
rect 646134 64368 646190 64424
rect 594062 54440 594118 54496
rect 577686 54168 577742 54224
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 308034 50224 308090 50280
rect 459926 53352 459982 53408
rect 462594 53624 462650 53680
rect 463698 53644 463754 53680
rect 463698 53624 463706 53644
rect 463706 53624 463754 53644
rect 472254 53644 472310 53680
rect 472254 53624 472256 53644
rect 472256 53624 472308 53644
rect 472308 53624 472310 53644
rect 462962 53216 463018 53272
rect 471886 53216 471942 53272
rect 309690 49680 309746 49736
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 458362 46688 458418 46744
rect 431222 44784 431278 44840
rect 310426 44104 310482 44160
rect 364890 44104 364946 44160
rect 308954 42744 309010 42800
rect 194322 42064 194378 42120
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 419906 41792 419962 41848
rect 443550 42200 443606 42256
rect 443550 41520 443606 41576
rect 460110 44784 460166 44840
rect 460846 43424 460902 43480
rect 461950 44376 462006 44432
rect 462502 44376 462558 44432
rect 463698 44104 463754 44160
rect 462962 43832 463018 43888
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463698 42880 463754 42936
rect 549994 48864 550050 48920
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 665178 92520 665234 92576
rect 665546 93336 665602 93392
rect 665362 90616 665418 90672
rect 664626 89800 664682 89856
rect 671894 151680 671950 151736
rect 672262 140256 672318 140312
rect 672078 133728 672134 133784
rect 673642 225392 673698 225448
rect 673458 223896 673514 223952
rect 673458 221992 673514 222048
rect 675022 309168 675078 309224
rect 674746 304680 674802 304736
rect 674838 301960 674894 302016
rect 674838 295840 674894 295896
rect 676034 308352 676090 308408
rect 676034 307944 676090 308000
rect 675206 303728 675262 303784
rect 675206 301960 675262 302016
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 676494 305904 676550 305960
rect 676034 303728 676090 303784
rect 676034 303456 676090 303512
rect 674930 294480 674986 294536
rect 676678 305088 676734 305144
rect 676494 301552 676550 301608
rect 676034 301416 676090 301472
rect 676678 301416 676734 301472
rect 678978 306312 679034 306368
rect 678242 298016 678298 298072
rect 675390 296520 675446 296576
rect 675022 292712 675078 292768
rect 674746 290944 674802 291000
rect 674286 286456 674342 286512
rect 674470 285504 674526 285560
rect 676034 296520 676090 296576
rect 675482 295840 675538 295896
rect 675758 295160 675814 295216
rect 675482 294480 675538 294536
rect 675482 292712 675538 292768
rect 675758 291488 675814 291544
rect 675390 290944 675446 291000
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 675482 285504 675538 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 683118 271088 683174 271144
rect 676034 269728 676090 269784
rect 676034 268232 676090 268288
rect 683118 268096 683174 268152
rect 675022 267008 675078 267064
rect 674470 264968 674526 265024
rect 674838 264424 674894 264480
rect 674838 263744 674894 263800
rect 674562 263064 674618 263120
rect 674378 260888 674434 260944
rect 675390 265376 675446 265432
rect 676494 264016 676550 264072
rect 676494 263608 676550 263664
rect 678242 263200 678298 263256
rect 675390 263064 675446 263120
rect 676218 262792 676274 262848
rect 674286 246880 674342 246936
rect 675390 255312 675446 255368
rect 676126 255312 676182 255368
rect 674470 234776 674526 234832
rect 675114 251776 675170 251832
rect 674930 249872 674986 249928
rect 678426 261160 678482 261216
rect 676034 251776 676090 251832
rect 675758 250280 675814 250336
rect 675390 249600 675446 249656
rect 675114 246880 675170 246936
rect 675298 245792 675354 245848
rect 675298 242800 675354 242856
rect 675666 242256 675722 242312
rect 675114 241440 675170 241496
rect 675390 240216 675446 240272
rect 675114 238176 675170 238232
rect 675114 237224 675170 237280
rect 674930 235864 674986 235920
rect 676034 235184 676090 235240
rect 675850 234776 675906 234832
rect 675850 233572 675906 233608
rect 675850 233552 675852 233572
rect 675852 233552 675904 233572
rect 675904 233552 675906 233572
rect 675178 231804 675234 231840
rect 675178 231784 675180 231804
rect 675180 231784 675232 231804
rect 675232 231784 675234 231804
rect 675068 231548 675070 231568
rect 675070 231548 675122 231568
rect 675122 231548 675124 231568
rect 675068 231512 675124 231548
rect 674730 231104 674786 231160
rect 674838 230832 674894 230888
rect 674516 230580 674572 230616
rect 674516 230560 674518 230580
rect 674518 230560 674570 230580
rect 674570 230560 674572 230580
rect 674394 230444 674450 230480
rect 674394 230424 674396 230444
rect 674396 230424 674448 230444
rect 674448 230424 674450 230444
rect 674102 226208 674158 226264
rect 674102 225936 674158 225992
rect 674194 225120 674250 225176
rect 673918 223624 673974 223680
rect 673642 221448 673698 221504
rect 673826 220496 673882 220552
rect 673550 220224 673606 220280
rect 673090 213696 673146 213752
rect 673090 196424 673146 196480
rect 673274 192208 673330 192264
rect 672906 177792 672962 177848
rect 673366 176840 673422 176896
rect 673182 176024 673238 176080
rect 672998 169088 673054 169144
rect 672998 153040 673054 153096
rect 673918 219816 673974 219872
rect 674562 229880 674618 229936
rect 676862 230560 676918 230616
rect 676586 230152 676642 230208
rect 675114 229880 675170 229936
rect 675114 229200 675170 229256
rect 674930 227024 674986 227080
rect 674746 222264 674802 222320
rect 674654 221856 674710 221912
rect 675666 225664 675722 225720
rect 675206 224440 675262 224496
rect 674930 221176 674986 221232
rect 675022 219000 675078 219056
rect 674838 217776 674894 217832
rect 674562 216144 674618 216200
rect 674102 212880 674158 212936
rect 674102 212064 674158 212120
rect 673918 209616 673974 209672
rect 673734 206896 673790 206952
rect 673918 203224 673974 203280
rect 673734 201592 673790 201648
rect 673550 175616 673606 175672
rect 673918 168680 673974 168736
rect 673918 151000 673974 151056
rect 673366 132096 673422 132152
rect 673182 131280 673238 131336
rect 674470 201864 674526 201920
rect 674286 179424 674342 179480
rect 675390 224168 675446 224224
rect 675850 218320 675906 218376
rect 675666 217504 675722 217560
rect 675390 216824 675446 216880
rect 675390 216552 675446 216608
rect 675206 214512 675262 214568
rect 675666 214512 675722 214568
rect 675666 211384 675722 211440
rect 676034 215056 676090 215112
rect 676034 213424 676090 213480
rect 676034 213152 676090 213208
rect 677046 228520 677102 228576
rect 676678 209616 676734 209672
rect 675850 207168 675906 207224
rect 683210 234096 683266 234152
rect 679254 223760 679310 223816
rect 683670 233824 683726 233880
rect 683210 222672 683266 222728
rect 678426 221448 678482 221504
rect 678242 220632 678298 220688
rect 683670 223080 683726 223136
rect 683486 219816 683542 219872
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 677782 206896 677838 206952
rect 675758 205536 675814 205592
rect 675390 201864 675446 201920
rect 675390 201320 675446 201376
rect 674838 201048 674894 201104
rect 675758 200776 675814 200832
rect 675390 198328 675446 198384
rect 674838 197512 674894 197568
rect 675482 197512 675538 197568
rect 675758 197104 675814 197160
rect 675390 196424 675446 196480
rect 675666 195200 675722 195256
rect 675666 193160 675722 193216
rect 675758 191528 675814 191584
rect 675298 190304 675354 190360
rect 683118 186904 683174 186960
rect 676494 181328 676550 181384
rect 676034 178064 676090 178120
rect 683118 178744 683174 178800
rect 674654 177248 674710 177304
rect 674654 175208 674710 175264
rect 674378 174392 674434 174448
rect 681002 173168 681058 173224
rect 674838 172760 674894 172816
rect 678242 171536 678298 171592
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 676586 166368 676642 166424
rect 676034 165552 676090 165608
rect 679622 171128 679678 171184
rect 675206 161880 675262 161936
rect 675850 161880 675906 161936
rect 676034 161336 676090 161392
rect 675758 159432 675814 159488
rect 674838 157528 674894 157584
rect 675482 157528 675538 157584
rect 675574 156984 675630 157040
rect 675758 156304 675814 156360
rect 675114 153040 675170 153096
rect 675758 153040 675814 153096
rect 675298 152632 675354 152688
rect 675114 151680 675170 151736
rect 675114 151000 675170 151056
rect 675758 150320 675814 150376
rect 675298 148960 675354 149016
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 683118 135904 683174 135960
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 683118 132640 683174 132696
rect 674654 130464 674710 130520
rect 675942 130056 675998 130112
rect 674378 129648 674434 129704
rect 674470 129240 674526 129296
rect 674286 128288 674342 128344
rect 674102 128152 674158 128208
rect 672998 125976 673054 126032
rect 672722 123936 672778 123992
rect 672538 123664 672594 123720
rect 672354 123120 672410 123176
rect 672354 120128 672410 120184
rect 671710 115776 671766 115832
rect 671526 107616 671582 107672
rect 672722 121352 672778 121408
rect 674102 125160 674158 125216
rect 673182 124344 673238 124400
rect 672998 111424 673054 111480
rect 672722 110880 672778 110936
rect 673366 123528 673422 123584
rect 673182 110336 673238 110392
rect 672538 106256 672594 106312
rect 673366 105576 673422 105632
rect 674102 104624 674158 104680
rect 668306 104352 668362 104408
rect 675942 128288 675998 128344
rect 682382 127744 682438 127800
rect 674838 127608 674894 127664
rect 674654 125568 674710 125624
rect 674470 111832 674526 111888
rect 675022 126384 675078 126440
rect 675298 113056 675354 113112
rect 675114 111424 675170 111480
rect 675114 110336 675170 110392
rect 675666 108024 675722 108080
rect 675114 106256 675170 106312
rect 675758 106120 675814 106176
rect 675114 105576 675170 105632
rect 675114 104624 675170 104680
rect 675758 103128 675814 103184
rect 675666 102584 675722 102640
rect 668490 102176 668546 102232
rect 674286 102176 674342 102232
rect 675758 101360 675814 101416
rect 663982 48456 664038 48512
rect 663798 47776 663854 47832
rect 662418 47368 662474 47424
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40432 141754 40488
rect 142618 40432 142674 40488
<< metal3 >>
rect 431677 1007178 431743 1007181
rect 431480 1007176 431743 1007178
rect 431480 1007120 431682 1007176
rect 431738 1007120 431743 1007176
rect 431480 1007118 431743 1007120
rect 431677 1007115 431743 1007118
rect 427997 1007042 428063 1007045
rect 505001 1007042 505067 1007045
rect 427800 1007040 428063 1007042
rect 427800 1006984 428002 1007040
rect 428058 1006984 428063 1007040
rect 427800 1006982 428063 1006984
rect 504804 1007040 505067 1007042
rect 504804 1006984 505006 1007040
rect 505062 1006984 505067 1007040
rect 504804 1006982 505067 1006984
rect 427997 1006979 428063 1006982
rect 505001 1006979 505067 1006982
rect 552289 1007042 552355 1007045
rect 552289 1007040 552552 1007042
rect 552289 1006984 552294 1007040
rect 552350 1006984 552552 1007040
rect 552289 1006982 552552 1006984
rect 552289 1006979 552355 1006982
rect 359733 1006906 359799 1006909
rect 428365 1006906 428431 1006909
rect 505369 1006906 505435 1006909
rect 359628 1006904 359799 1006906
rect 359628 1006848 359738 1006904
rect 359794 1006848 359799 1006904
rect 359628 1006846 359799 1006848
rect 428260 1006904 428431 1006906
rect 428260 1006848 428370 1006904
rect 428426 1006848 428431 1006904
rect 428260 1006846 428431 1006848
rect 505172 1006904 505435 1006906
rect 505172 1006848 505374 1006904
rect 505430 1006848 505435 1006904
rect 505172 1006846 505435 1006848
rect 359733 1006843 359799 1006846
rect 428365 1006843 428431 1006846
rect 505369 1006843 505435 1006846
rect 359365 1006770 359431 1006773
rect 429193 1006770 429259 1006773
rect 557165 1006770 557231 1006773
rect 359168 1006768 359431 1006770
rect 359168 1006712 359370 1006768
rect 359426 1006712 359431 1006768
rect 359168 1006710 359431 1006712
rect 428996 1006768 429259 1006770
rect 428996 1006712 429198 1006768
rect 429254 1006712 429259 1006768
rect 428996 1006710 429259 1006712
rect 557060 1006768 557231 1006770
rect 557060 1006712 557170 1006768
rect 557226 1006712 557231 1006768
rect 557060 1006710 557231 1006712
rect 359365 1006707 359431 1006710
rect 429193 1006707 429259 1006710
rect 557165 1006707 557231 1006710
rect 152089 1006634 152155 1006637
rect 157425 1006634 157491 1006637
rect 152089 1006632 152352 1006634
rect 152089 1006576 152094 1006632
rect 152150 1006576 152352 1006632
rect 152089 1006574 152352 1006576
rect 157228 1006632 157491 1006634
rect 157228 1006576 157430 1006632
rect 157486 1006576 157491 1006632
rect 157228 1006574 157491 1006576
rect 152089 1006571 152155 1006574
rect 157425 1006571 157491 1006574
rect 360561 1006634 360627 1006637
rect 505369 1006634 505435 1006637
rect 553117 1006634 553183 1006637
rect 360561 1006632 360824 1006634
rect 360561 1006576 360566 1006632
rect 360622 1006576 360824 1006632
rect 360561 1006574 360824 1006576
rect 505369 1006632 505632 1006634
rect 505369 1006576 505374 1006632
rect 505430 1006576 505632 1006632
rect 505369 1006574 505632 1006576
rect 553117 1006632 553380 1006634
rect 553117 1006576 553122 1006632
rect 553178 1006576 553380 1006632
rect 553117 1006574 553380 1006576
rect 360561 1006571 360627 1006574
rect 505369 1006571 505435 1006574
rect 553117 1006571 553183 1006574
rect 101121 1006498 101187 1006501
rect 100924 1006496 101187 1006498
rect 100924 1006440 101126 1006496
rect 101182 1006440 101187 1006496
rect 100924 1006438 101187 1006440
rect 101121 1006435 101187 1006438
rect 151261 1006498 151327 1006501
rect 151721 1006498 151787 1006501
rect 158621 1006498 158687 1006501
rect 255313 1006498 255379 1006501
rect 361389 1006498 361455 1006501
rect 551093 1006498 551159 1006501
rect 556797 1006498 556863 1006501
rect 151261 1006496 151524 1006498
rect 151261 1006440 151266 1006496
rect 151322 1006440 151524 1006496
rect 151261 1006438 151524 1006440
rect 151721 1006496 151892 1006498
rect 151721 1006440 151726 1006496
rect 151782 1006440 151892 1006496
rect 151721 1006438 151892 1006440
rect 158621 1006496 158884 1006498
rect 158621 1006440 158626 1006496
rect 158682 1006440 158884 1006496
rect 158621 1006438 158884 1006440
rect 255313 1006496 255576 1006498
rect 255313 1006440 255318 1006496
rect 255374 1006440 255576 1006496
rect 255313 1006438 255576 1006440
rect 361192 1006496 361455 1006498
rect 361192 1006440 361394 1006496
rect 361450 1006440 361455 1006496
rect 361192 1006438 361455 1006440
rect 550436 1006496 551159 1006498
rect 550436 1006440 551098 1006496
rect 551154 1006440 551159 1006496
rect 550436 1006438 551159 1006440
rect 556600 1006496 556863 1006498
rect 556600 1006440 556802 1006496
rect 556858 1006440 556863 1006496
rect 556600 1006438 556863 1006440
rect 151261 1006435 151327 1006438
rect 151721 1006435 151787 1006438
rect 158621 1006435 158687 1006438
rect 255313 1006435 255379 1006438
rect 361389 1006435 361455 1006438
rect 551093 1006435 551159 1006438
rect 556797 1006435 556863 1006438
rect 101949 1006362 102015 1006365
rect 108481 1006362 108547 1006365
rect 101949 1006360 102212 1006362
rect 101949 1006304 101954 1006360
rect 102010 1006304 102212 1006360
rect 101949 1006302 102212 1006304
rect 108284 1006360 108547 1006362
rect 108284 1006304 108486 1006360
rect 108542 1006304 108547 1006360
rect 108284 1006302 108547 1006304
rect 101949 1006299 102015 1006302
rect 108481 1006299 108547 1006302
rect 158253 1006362 158319 1006365
rect 159449 1006362 159515 1006365
rect 254117 1006362 254183 1006365
rect 306925 1006362 306991 1006365
rect 314653 1006362 314719 1006365
rect 158253 1006360 158516 1006362
rect 158253 1006304 158258 1006360
rect 158314 1006304 158516 1006360
rect 158253 1006302 158516 1006304
rect 159449 1006360 159712 1006362
rect 159449 1006304 159454 1006360
rect 159510 1006304 159712 1006360
rect 159449 1006302 159712 1006304
rect 254117 1006360 254380 1006362
rect 254117 1006304 254122 1006360
rect 254178 1006304 254380 1006360
rect 254117 1006302 254380 1006304
rect 306728 1006360 306991 1006362
rect 306728 1006304 306930 1006360
rect 306986 1006304 306991 1006360
rect 306728 1006302 306991 1006304
rect 314548 1006360 314719 1006362
rect 314548 1006304 314658 1006360
rect 314714 1006304 314719 1006360
rect 314548 1006302 314719 1006304
rect 158253 1006299 158319 1006302
rect 159449 1006299 159515 1006302
rect 254117 1006299 254183 1006302
rect 306925 1006299 306991 1006302
rect 314653 1006299 314719 1006302
rect 431677 1006362 431743 1006365
rect 507853 1006362 507919 1006365
rect 558821 1006362 558887 1006365
rect 431677 1006360 431940 1006362
rect 431677 1006304 431682 1006360
rect 431738 1006304 431940 1006360
rect 431677 1006302 431940 1006304
rect 507656 1006360 507919 1006362
rect 507656 1006304 507858 1006360
rect 507914 1006304 507919 1006360
rect 507656 1006302 507919 1006304
rect 558624 1006360 558887 1006362
rect 558624 1006304 558826 1006360
rect 558882 1006304 558887 1006360
rect 558624 1006302 558887 1006304
rect 431677 1006299 431743 1006302
rect 507853 1006299 507919 1006302
rect 558821 1006299 558887 1006302
rect 99465 1006226 99531 1006229
rect 104801 1006226 104867 1006229
rect 106825 1006226 106891 1006229
rect 99465 1006224 99728 1006226
rect 99465 1006168 99470 1006224
rect 99526 1006168 99728 1006224
rect 99465 1006166 99728 1006168
rect 104604 1006224 104867 1006226
rect 104604 1006168 104806 1006224
rect 104862 1006168 104867 1006224
rect 104604 1006166 104867 1006168
rect 106628 1006224 106891 1006226
rect 106628 1006168 106830 1006224
rect 106886 1006168 106891 1006224
rect 106628 1006166 106891 1006168
rect 99465 1006163 99531 1006166
rect 104801 1006163 104867 1006166
rect 106825 1006163 106891 1006166
rect 150893 1006226 150959 1006229
rect 153745 1006226 153811 1006229
rect 160277 1006226 160343 1006229
rect 210417 1006226 210483 1006229
rect 262673 1006226 262739 1006229
rect 150893 1006224 151156 1006226
rect 150893 1006168 150898 1006224
rect 150954 1006168 151156 1006224
rect 150893 1006166 151156 1006168
rect 153548 1006224 153811 1006226
rect 153548 1006168 153750 1006224
rect 153806 1006168 153811 1006224
rect 153548 1006166 153811 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 210220 1006224 210483 1006226
rect 210220 1006168 210422 1006224
rect 210478 1006168 210483 1006224
rect 210220 1006166 210483 1006168
rect 262476 1006224 262739 1006226
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 150893 1006163 150959 1006166
rect 153745 1006163 153811 1006166
rect 160277 1006163 160343 1006166
rect 210417 1006163 210483 1006166
rect 262673 1006163 262739 1006166
rect 304901 1006226 304967 1006229
rect 355685 1006226 355751 1006229
rect 365069 1006226 365135 1006229
rect 304901 1006224 305164 1006226
rect 304901 1006168 304906 1006224
rect 304962 1006168 305164 1006224
rect 304901 1006166 305164 1006168
rect 355685 1006224 355948 1006226
rect 355685 1006168 355690 1006224
rect 355746 1006168 355948 1006224
rect 355685 1006166 355948 1006168
rect 364872 1006224 365135 1006226
rect 364872 1006168 365074 1006224
rect 365130 1006168 365135 1006224
rect 364872 1006166 365135 1006168
rect 304901 1006163 304967 1006166
rect 355685 1006163 355751 1006166
rect 365069 1006163 365135 1006166
rect 429193 1006226 429259 1006229
rect 506197 1006226 506263 1006229
rect 553945 1006226 554011 1006229
rect 429193 1006224 429456 1006226
rect 429193 1006168 429198 1006224
rect 429254 1006168 429456 1006224
rect 429193 1006166 429456 1006168
rect 506000 1006224 506263 1006226
rect 506000 1006168 506202 1006224
rect 506258 1006168 506263 1006224
rect 506000 1006166 506263 1006168
rect 553748 1006224 554011 1006226
rect 553748 1006168 553950 1006224
rect 554006 1006168 554011 1006224
rect 553748 1006166 554011 1006168
rect 429193 1006163 429259 1006166
rect 506197 1006163 506263 1006166
rect 553945 1006163 554011 1006166
rect 98269 1006090 98335 1006093
rect 103973 1006090 104039 1006093
rect 105997 1006090 106063 1006093
rect 98269 1006088 98900 1006090
rect 98269 1006032 98274 1006088
rect 98330 1006032 98900 1006088
rect 98269 1006030 98900 1006032
rect 103973 1006088 104236 1006090
rect 103973 1006032 103978 1006088
rect 104034 1006032 104236 1006088
rect 103973 1006030 104236 1006032
rect 105892 1006088 106063 1006090
rect 105892 1006032 106002 1006088
rect 106058 1006032 106063 1006088
rect 105892 1006030 106063 1006032
rect 98269 1006027 98335 1006030
rect 103973 1006027 104039 1006030
rect 105997 1006027 106063 1006030
rect 147121 1006090 147187 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 158253 1006090 158319 1006093
rect 147121 1006088 148935 1006090
rect 147121 1006032 147126 1006088
rect 147182 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 147121 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 158056 1006088 158319 1006090
rect 158056 1006032 158258 1006088
rect 158314 1006032 158319 1006088
rect 158056 1006030 158319 1006032
rect 147121 1006027 147187 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 158253 1006027 158319 1006030
rect 201033 1006090 201099 1006093
rect 208393 1006090 208459 1006093
rect 252461 1006090 252527 1006093
rect 261845 1006090 261911 1006093
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 208393 1006088 208656 1006090
rect 208393 1006032 208398 1006088
rect 208454 1006032 208656 1006088
rect 208393 1006030 208656 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 201033 1006027 201099 1006030
rect 208393 1006027 208459 1006030
rect 252461 1006027 252527 1006030
rect 261845 1006027 261911 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 354857 1006090 354923 1006093
rect 363413 1006090 363479 1006093
rect 422661 1006090 422727 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314653 1006088 314916 1006090
rect 314653 1006032 314658 1006088
rect 314714 1006032 314916 1006088
rect 314653 1006030 314916 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 363308 1006088 363479 1006090
rect 363308 1006032 363418 1006088
rect 363474 1006032 363479 1006088
rect 363308 1006030 363479 1006032
rect 422096 1006088 422727 1006090
rect 422096 1006032 422666 1006088
rect 422722 1006032 422727 1006088
rect 422096 1006030 422727 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 354857 1006027 354923 1006030
rect 363413 1006027 363479 1006030
rect 422661 1006027 422727 1006030
rect 425513 1006090 425579 1006093
rect 430021 1006090 430087 1006093
rect 425513 1006088 425776 1006090
rect 425513 1006032 425518 1006088
rect 425574 1006032 425776 1006088
rect 425513 1006030 425776 1006032
rect 429824 1006088 430087 1006090
rect 429824 1006032 430026 1006088
rect 430082 1006032 430087 1006088
rect 429824 1006030 430087 1006032
rect 425513 1006027 425579 1006030
rect 430021 1006027 430087 1006030
rect 498837 1006090 498903 1006093
rect 500493 1006090 500559 1006093
rect 554313 1006090 554379 1006093
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 500493 1006088 500756 1006090
rect 500493 1006032 500498 1006088
rect 500554 1006032 500756 1006088
rect 500493 1006030 500756 1006032
rect 554116 1006088 554379 1006090
rect 554116 1006032 554318 1006088
rect 554374 1006032 554379 1006088
rect 554116 1006030 554379 1006032
rect 498837 1006027 498903 1006030
rect 500493 1006027 500559 1006030
rect 554313 1006027 554379 1006030
rect 509049 1005954 509115 1005957
rect 509049 1005952 509312 1005954
rect 509049 1005896 509054 1005952
rect 509110 1005896 509312 1005952
rect 509049 1005894 509312 1005896
rect 509049 1005891 509115 1005894
rect 427537 1005682 427603 1005685
rect 427340 1005680 427603 1005682
rect 427340 1005624 427542 1005680
rect 427598 1005624 427603 1005680
rect 427340 1005622 427603 1005624
rect 427537 1005619 427603 1005622
rect 428365 1005546 428431 1005549
rect 428365 1005544 428628 1005546
rect 428365 1005488 428370 1005544
rect 428426 1005488 428628 1005544
rect 428365 1005486 428628 1005488
rect 428365 1005483 428431 1005486
rect 360561 1005410 360627 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 360561 1005347 360627 1005350
rect 423489 1005410 423555 1005413
rect 555969 1005410 556035 1005413
rect 423489 1005408 423752 1005410
rect 423489 1005352 423494 1005408
rect 423550 1005352 423752 1005408
rect 423489 1005350 423752 1005352
rect 555969 1005408 556232 1005410
rect 555969 1005352 555974 1005408
rect 556030 1005352 556232 1005408
rect 555969 1005350 556232 1005352
rect 423489 1005347 423555 1005350
rect 555969 1005347 556035 1005350
rect 108849 1005274 108915 1005277
rect 212073 1005274 212139 1005277
rect 108849 1005272 109112 1005274
rect 108849 1005216 108854 1005272
rect 108910 1005216 109112 1005272
rect 108849 1005214 109112 1005216
rect 211876 1005272 212139 1005274
rect 211876 1005216 212078 1005272
rect 212134 1005216 212139 1005272
rect 211876 1005214 212139 1005216
rect 108849 1005211 108915 1005214
rect 212073 1005211 212139 1005214
rect 357709 1005274 357775 1005277
rect 424317 1005274 424383 1005277
rect 498837 1005274 498903 1005277
rect 357709 1005272 357972 1005274
rect 357709 1005216 357714 1005272
rect 357770 1005216 357972 1005272
rect 357709 1005214 357972 1005216
rect 424120 1005272 424383 1005274
rect 424120 1005216 424322 1005272
rect 424378 1005216 424383 1005272
rect 424120 1005214 424383 1005216
rect 498732 1005272 498903 1005274
rect 498732 1005216 498842 1005272
rect 498898 1005216 498903 1005272
rect 498732 1005214 498903 1005216
rect 357709 1005211 357775 1005214
rect 424317 1005211 424383 1005214
rect 498837 1005211 498903 1005214
rect 152917 1005138 152983 1005141
rect 356513 1005138 356579 1005141
rect 152917 1005136 153180 1005138
rect 152917 1005080 152922 1005136
rect 152978 1005080 153180 1005136
rect 152917 1005078 153180 1005080
rect 356316 1005136 356579 1005138
rect 356316 1005080 356518 1005136
rect 356574 1005080 356579 1005136
rect 356316 1005078 356579 1005080
rect 152917 1005075 152983 1005078
rect 356513 1005075 356579 1005078
rect 365069 1005138 365135 1005141
rect 551461 1005138 551527 1005141
rect 365069 1005136 365332 1005138
rect 365069 1005080 365074 1005136
rect 365130 1005080 365332 1005136
rect 365069 1005078 365332 1005080
rect 551356 1005136 551527 1005138
rect 551356 1005080 551466 1005136
rect 551522 1005080 551527 1005136
rect 551356 1005078 551527 1005080
rect 365069 1005075 365135 1005078
rect 551461 1005075 551527 1005078
rect 153745 1005002 153811 1005005
rect 209221 1005002 209287 1005005
rect 263041 1005002 263107 1005005
rect 355685 1005002 355751 1005005
rect 153745 1005000 153916 1005002
rect 153745 1004944 153750 1005000
rect 153806 1004944 153916 1005000
rect 153745 1004942 153916 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 262844 1005000 263107 1005002
rect 262844 1004944 263046 1005000
rect 263102 1004944 263107 1005000
rect 262844 1004942 263107 1004944
rect 355488 1005000 355751 1005002
rect 355488 1004944 355690 1005000
rect 355746 1004944 355751 1005000
rect 355488 1004942 355751 1004944
rect 153745 1004939 153811 1004942
rect 209221 1004939 209287 1004942
rect 263041 1004939 263107 1004942
rect 355685 1004939 355751 1004942
rect 361389 1005002 361455 1005005
rect 423489 1005002 423555 1005005
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 423292 1005000 423555 1005002
rect 423292 1004944 423494 1005000
rect 423550 1004944 423555 1005000
rect 423292 1004942 423555 1004944
rect 361389 1004939 361455 1004942
rect 423489 1004939 423555 1004942
rect 499665 1005002 499731 1005005
rect 508221 1005002 508287 1005005
rect 509877 1005002 509943 1005005
rect 499665 1005000 499928 1005002
rect 499665 1004944 499670 1005000
rect 499726 1004944 499928 1005000
rect 499665 1004942 499928 1004944
rect 508221 1005000 508484 1005002
rect 508221 1004944 508226 1005000
rect 508282 1004944 508484 1005000
rect 508221 1004942 508484 1004944
rect 509680 1005000 509943 1005002
rect 509680 1004944 509882 1005000
rect 509938 1004944 509943 1005000
rect 509680 1004942 509943 1004944
rect 499665 1004939 499731 1004942
rect 508221 1004939 508287 1004942
rect 509877 1004939 509943 1004942
rect 560845 1005002 560911 1005005
rect 560845 1005000 561108 1005002
rect 560845 1004944 560850 1005000
rect 560906 1004944 561108 1005000
rect 560845 1004942 561108 1004944
rect 560845 1004939 560911 1004942
rect 152917 1004866 152983 1004869
rect 160645 1004866 160711 1004869
rect 152720 1004864 152983 1004866
rect 152720 1004808 152922 1004864
rect 152978 1004808 152983 1004864
rect 152720 1004806 152983 1004808
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 152917 1004803 152983 1004806
rect 160645 1004803 160711 1004806
rect 211245 1004866 211311 1004869
rect 313825 1004866 313891 1004869
rect 362585 1004866 362651 1004869
rect 211245 1004864 211508 1004866
rect 211245 1004808 211250 1004864
rect 211306 1004808 211508 1004864
rect 211245 1004806 211508 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 211245 1004803 211311 1004806
rect 313825 1004803 313891 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 430849 1004866 430915 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 430652 1004864 430915 1004866
rect 430652 1004808 430854 1004864
rect 430910 1004808 430915 1004864
rect 430652 1004806 430915 1004808
rect 422661 1004803 422727 1004806
rect 430849 1004803 430915 1004806
rect 432045 1004866 432111 1004869
rect 501321 1004866 501387 1004869
rect 507025 1004866 507091 1004869
rect 555969 1004866 556035 1004869
rect 432045 1004864 432308 1004866
rect 432045 1004808 432050 1004864
rect 432106 1004808 432308 1004864
rect 432045 1004806 432308 1004808
rect 501124 1004864 501387 1004866
rect 501124 1004808 501326 1004864
rect 501382 1004808 501387 1004864
rect 501124 1004806 501387 1004808
rect 506828 1004864 507091 1004866
rect 506828 1004808 507030 1004864
rect 507086 1004808 507091 1004864
rect 506828 1004806 507091 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 432045 1004803 432111 1004806
rect 501321 1004803 501387 1004806
rect 507025 1004803 507091 1004806
rect 555969 1004803 556035 1004806
rect 108481 1004730 108547 1004733
rect 154113 1004730 154179 1004733
rect 161105 1004730 161171 1004733
rect 209221 1004730 209287 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 154113 1004728 154376 1004730
rect 154113 1004672 154118 1004728
rect 154174 1004672 154376 1004728
rect 154113 1004670 154376 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 108481 1004667 108547 1004670
rect 154113 1004667 154179 1004670
rect 161105 1004667 161171 1004670
rect 209221 1004667 209287 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 430021 1004730 430087 1004733
rect 432873 1004730 432939 1004733
rect 503345 1004730 503411 1004733
rect 508221 1004730 508287 1004733
rect 557625 1004730 557691 1004733
rect 560845 1004730 560911 1004733
rect 430021 1004728 430284 1004730
rect 430021 1004672 430026 1004728
rect 430082 1004672 430284 1004728
rect 430021 1004670 430284 1004672
rect 432676 1004728 432939 1004730
rect 432676 1004672 432878 1004728
rect 432934 1004672 432939 1004728
rect 432676 1004670 432939 1004672
rect 503148 1004728 503411 1004730
rect 503148 1004672 503350 1004728
rect 503406 1004672 503411 1004728
rect 503148 1004670 503411 1004672
rect 508116 1004728 508287 1004730
rect 508116 1004672 508226 1004728
rect 508282 1004672 508287 1004728
rect 508116 1004670 508287 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 560740 1004728 560911 1004730
rect 560740 1004672 560850 1004728
rect 560906 1004672 560911 1004728
rect 560740 1004670 560911 1004672
rect 430021 1004667 430087 1004670
rect 432873 1004667 432939 1004670
rect 503345 1004667 503411 1004670
rect 508221 1004667 508287 1004670
rect 557625 1004667 557691 1004670
rect 560845 1004667 560911 1004670
rect 424317 1004594 424383 1004597
rect 500493 1004594 500559 1004597
rect 424317 1004592 424580 1004594
rect 424317 1004536 424322 1004592
rect 424378 1004536 424580 1004592
rect 424317 1004534 424580 1004536
rect 500296 1004592 500559 1004594
rect 500296 1004536 500498 1004592
rect 500554 1004536 500559 1004592
rect 500296 1004534 500559 1004536
rect 424317 1004531 424383 1004534
rect 500493 1004531 500559 1004534
rect 425513 1004186 425579 1004189
rect 425316 1004184 425579 1004186
rect 425316 1004128 425518 1004184
rect 425574 1004128 425579 1004184
rect 425316 1004126 425579 1004128
rect 425513 1004123 425579 1004126
rect 425145 1004050 425211 1004053
rect 502517 1004050 502583 1004053
rect 424948 1004048 425211 1004050
rect 424948 1003992 425150 1004048
rect 425206 1003992 425211 1004048
rect 424948 1003990 425211 1003992
rect 502412 1004048 502583 1004050
rect 502412 1003992 502522 1004048
rect 502578 1003992 502583 1004048
rect 502412 1003990 502583 1003992
rect 425145 1003987 425211 1003990
rect 502517 1003987 502583 1003990
rect 102317 1002826 102383 1002829
rect 102317 1002824 102580 1002826
rect 102317 1002768 102322 1002824
rect 102378 1002768 102580 1002824
rect 102317 1002766 102580 1002768
rect 102317 1002763 102383 1002766
rect 100293 1002690 100359 1002693
rect 100096 1002688 100359 1002690
rect 100096 1002632 100298 1002688
rect 100354 1002632 100359 1002688
rect 100096 1002630 100359 1002632
rect 100293 1002627 100359 1002630
rect 256141 1002690 256207 1002693
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 256141 1002627 256207 1002630
rect 103145 1002554 103211 1002557
rect 255313 1002554 255379 1002557
rect 261017 1002554 261083 1002557
rect 103145 1002552 103408 1002554
rect 103145 1002496 103150 1002552
rect 103206 1002496 103408 1002552
rect 103145 1002494 103408 1002496
rect 255116 1002552 255379 1002554
rect 255116 1002496 255318 1002552
rect 255374 1002496 255379 1002552
rect 255116 1002494 255379 1002496
rect 260820 1002552 261083 1002554
rect 260820 1002496 261022 1002552
rect 261078 1002496 261083 1002552
rect 260820 1002494 261083 1002496
rect 103145 1002491 103211 1002494
rect 255313 1002491 255379 1002494
rect 261017 1002491 261083 1002494
rect 426341 1002554 426407 1002557
rect 557993 1002554 558059 1002557
rect 426341 1002552 426604 1002554
rect 426341 1002496 426346 1002552
rect 426402 1002496 426604 1002552
rect 426341 1002494 426604 1002496
rect 557993 1002552 558256 1002554
rect 557993 1002496 557998 1002552
rect 558054 1002496 558256 1002552
rect 557993 1002494 558256 1002496
rect 426341 1002491 426407 1002494
rect 557993 1002491 558059 1002494
rect 100293 1002418 100359 1002421
rect 107653 1002418 107719 1002421
rect 256141 1002418 256207 1002421
rect 555141 1002418 555207 1002421
rect 100293 1002416 100556 1002418
rect 100293 1002360 100298 1002416
rect 100354 1002360 100556 1002416
rect 100293 1002358 100556 1002360
rect 107456 1002416 107719 1002418
rect 107456 1002360 107658 1002416
rect 107714 1002360 107719 1002416
rect 107456 1002358 107719 1002360
rect 255944 1002416 256207 1002418
rect 255944 1002360 256146 1002416
rect 256202 1002360 256207 1002416
rect 255944 1002358 256207 1002360
rect 555036 1002416 555207 1002418
rect 555036 1002360 555146 1002416
rect 555202 1002360 555207 1002416
rect 555036 1002358 555207 1002360
rect 100293 1002355 100359 1002358
rect 107653 1002355 107719 1002358
rect 256141 1002355 256207 1002358
rect 555141 1002355 555207 1002358
rect 558821 1002418 558887 1002421
rect 558821 1002416 559084 1002418
rect 558821 1002360 558826 1002416
rect 558882 1002360 559084 1002416
rect 558821 1002358 559084 1002360
rect 558821 1002355 558887 1002358
rect 101949 1002282 102015 1002285
rect 105629 1002282 105695 1002285
rect 108021 1002282 108087 1002285
rect 101752 1002280 102015 1002282
rect 101752 1002224 101954 1002280
rect 102010 1002224 102015 1002280
rect 101752 1002222 102015 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 107916 1002280 108087 1002282
rect 107916 1002224 108026 1002280
rect 108082 1002224 108087 1002280
rect 107916 1002222 108087 1002224
rect 101949 1002219 102015 1002222
rect 105629 1002219 105695 1002222
rect 108021 1002219 108087 1002222
rect 155769 1002282 155835 1002285
rect 206369 1002282 206435 1002285
rect 206737 1002282 206803 1002285
rect 155769 1002280 156032 1002282
rect 155769 1002224 155774 1002280
rect 155830 1002224 156032 1002280
rect 155769 1002222 156032 1002224
rect 206172 1002280 206435 1002282
rect 206172 1002224 206374 1002280
rect 206430 1002224 206435 1002280
rect 206172 1002222 206435 1002224
rect 206540 1002280 206803 1002282
rect 206540 1002224 206742 1002280
rect 206798 1002224 206803 1002280
rect 206540 1002222 206803 1002224
rect 155769 1002219 155835 1002222
rect 206369 1002219 206435 1002222
rect 206737 1002219 206803 1002222
rect 210877 1002282 210943 1002285
rect 254485 1002282 254551 1002285
rect 358537 1002282 358603 1002285
rect 426341 1002282 426407 1002285
rect 501689 1002282 501755 1002285
rect 210877 1002280 211140 1002282
rect 210877 1002224 210882 1002280
rect 210938 1002224 211140 1002280
rect 210877 1002222 211140 1002224
rect 254485 1002280 254748 1002282
rect 254485 1002224 254490 1002280
rect 254546 1002224 254748 1002280
rect 254485 1002222 254748 1002224
rect 358537 1002280 358800 1002282
rect 358537 1002224 358542 1002280
rect 358598 1002224 358800 1002280
rect 358537 1002222 358800 1002224
rect 426144 1002280 426407 1002282
rect 426144 1002224 426346 1002280
rect 426402 1002224 426407 1002280
rect 426144 1002222 426407 1002224
rect 501492 1002280 501755 1002282
rect 501492 1002224 501694 1002280
rect 501750 1002224 501755 1002280
rect 501492 1002222 501755 1002224
rect 210877 1002219 210943 1002222
rect 254485 1002219 254551 1002222
rect 358537 1002219 358603 1002222
rect 426341 1002219 426407 1002222
rect 501689 1002219 501755 1002222
rect 554313 1002282 554379 1002285
rect 557993 1002282 558059 1002285
rect 560477 1002282 560543 1002285
rect 554313 1002280 554576 1002282
rect 554313 1002224 554318 1002280
rect 554374 1002224 554576 1002280
rect 554313 1002222 554576 1002224
rect 557796 1002280 558059 1002282
rect 557796 1002224 557998 1002280
rect 558054 1002224 558059 1002280
rect 557796 1002222 558059 1002224
rect 560280 1002280 560543 1002282
rect 560280 1002224 560482 1002280
rect 560538 1002224 560543 1002280
rect 560280 1002222 560543 1002224
rect 554313 1002219 554379 1002222
rect 557993 1002219 558059 1002222
rect 560477 1002219 560543 1002222
rect 99097 1002146 99163 1002149
rect 103145 1002146 103211 1002149
rect 103973 1002146 104039 1002149
rect 99097 1002144 99268 1002146
rect 99097 1002088 99102 1002144
rect 99158 1002088 99268 1002144
rect 99097 1002086 99268 1002088
rect 102948 1002144 103211 1002146
rect 102948 1002088 103150 1002144
rect 103206 1002088 103211 1002144
rect 102948 1002086 103211 1002088
rect 103776 1002144 104039 1002146
rect 103776 1002088 103978 1002144
rect 104034 1002088 104039 1002144
rect 103776 1002086 104039 1002088
rect 99097 1002083 99163 1002086
rect 103145 1002083 103211 1002086
rect 103973 1002083 104039 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 154573 1002146 154639 1002149
rect 207197 1002146 207263 1002149
rect 212533 1002146 212599 1002149
rect 263501 1002146 263567 1002149
rect 154573 1002144 154836 1002146
rect 154573 1002088 154578 1002144
rect 154634 1002088 154836 1002144
rect 154573 1002086 154836 1002088
rect 207197 1002144 207460 1002146
rect 207197 1002088 207202 1002144
rect 207258 1002088 207460 1002144
rect 207197 1002086 207460 1002088
rect 212336 1002144 212599 1002146
rect 212336 1002088 212538 1002144
rect 212594 1002088 212599 1002144
rect 212336 1002086 212599 1002088
rect 263304 1002144 263567 1002146
rect 263304 1002088 263506 1002144
rect 263562 1002088 263567 1002144
rect 263304 1002086 263567 1002088
rect 154573 1002083 154639 1002086
rect 207197 1002083 207263 1002086
rect 212533 1002083 212599 1002086
rect 263501 1002083 263567 1002086
rect 305269 1002146 305335 1002149
rect 310145 1002146 310211 1002149
rect 305269 1002144 305532 1002146
rect 305269 1002088 305274 1002144
rect 305330 1002088 305532 1002144
rect 305269 1002086 305532 1002088
rect 309948 1002144 310211 1002146
rect 309948 1002088 310150 1002144
rect 310206 1002088 310211 1002144
rect 309948 1002086 310211 1002088
rect 305269 1002083 305335 1002086
rect 310145 1002083 310211 1002086
rect 356513 1002146 356579 1002149
rect 504541 1002146 504607 1002149
rect 559649 1002146 559715 1002149
rect 561673 1002146 561739 1002149
rect 356513 1002144 356684 1002146
rect 356513 1002088 356518 1002144
rect 356574 1002088 356684 1002144
rect 356513 1002086 356684 1002088
rect 504436 1002144 504607 1002146
rect 504436 1002088 504546 1002144
rect 504602 1002088 504607 1002144
rect 504436 1002086 504607 1002088
rect 559452 1002144 559715 1002146
rect 559452 1002088 559654 1002144
rect 559710 1002088 559715 1002144
rect 559452 1002086 559715 1002088
rect 561476 1002144 561739 1002146
rect 561476 1002088 561678 1002144
rect 561734 1002088 561739 1002144
rect 561476 1002086 561739 1002088
rect 356513 1002083 356579 1002086
rect 504541 1002083 504607 1002086
rect 559649 1002083 559715 1002086
rect 561673 1002083 561739 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101121 1002010 101187 1002013
rect 104801 1002010 104867 1002013
rect 105997 1002010 106063 1002013
rect 149237 1002010 149303 1002013
rect 154941 1002010 155007 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 157793 1002010 157859 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 104801 1002008 104972 1002010
rect 104801 1001952 104806 1002008
rect 104862 1001952 104972 1002008
rect 104801 1001950 104972 1001952
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 155572 1002008 155835 1002010
rect 155572 1001952 155774 1002008
rect 155830 1001952 155835 1002008
rect 155572 1001950 155835 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 157596 1002008 157859 1002010
rect 157596 1001952 157798 1002008
rect 157854 1001952 157859 1002008
rect 157596 1001950 157859 1001952
rect 101121 1001947 101187 1001950
rect 104801 1001947 104867 1001950
rect 105997 1001947 106063 1001950
rect 149237 1001947 149303 1001950
rect 154941 1001947 155007 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 157793 1001947 157859 1001950
rect 205541 1002010 205607 1002013
rect 206737 1002010 206803 1002013
rect 207565 1002010 207631 1002013
rect 210877 1002010 210943 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 206737 1002008 207000 1002010
rect 206737 1001952 206742 1002008
rect 206798 1001952 207000 1002008
rect 206737 1001950 207000 1001952
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 210680 1002008 210943 1002010
rect 210680 1001952 210882 1002008
rect 210938 1001952 210943 1002008
rect 210680 1001950 210943 1001952
rect 205541 1001947 205607 1001950
rect 206737 1001947 206803 1001950
rect 207565 1001947 207631 1001950
rect 210877 1001947 210943 1001950
rect 261017 1002010 261083 1002013
rect 263869 1002010 263935 1002013
rect 261017 1002008 261280 1002010
rect 261017 1001952 261022 1002008
rect 261078 1001952 261280 1002008
rect 261017 1001950 261280 1001952
rect 263764 1002008 263935 1002010
rect 263764 1001952 263874 1002008
rect 263930 1001952 263935 1002008
rect 263764 1001950 263935 1001952
rect 261017 1001947 261083 1001950
rect 263869 1001947 263935 1001950
rect 310973 1002010 311039 1002013
rect 354029 1002010 354095 1002013
rect 356881 1002010 356947 1002013
rect 357709 1002010 357775 1002013
rect 358537 1002010 358603 1002013
rect 360193 1002010 360259 1002013
rect 365897 1002010 365963 1002013
rect 310973 1002008 311236 1002010
rect 310973 1001952 310978 1002008
rect 311034 1001952 311236 1002008
rect 310973 1001950 311236 1001952
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 356881 1002008 357144 1002010
rect 356881 1001952 356886 1002008
rect 356942 1001952 357144 1002008
rect 356881 1001950 357144 1001952
rect 357604 1002008 357775 1002010
rect 357604 1001952 357714 1002008
rect 357770 1001952 357775 1002008
rect 357604 1001950 357775 1001952
rect 358340 1002008 358603 1002010
rect 358340 1001952 358542 1002008
rect 358598 1001952 358603 1002008
rect 358340 1001950 358603 1001952
rect 359996 1002008 360259 1002010
rect 359996 1001952 360198 1002008
rect 360254 1001952 360259 1002008
rect 359996 1001950 360259 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 310973 1001947 311039 1001950
rect 354029 1001947 354095 1001950
rect 356881 1001947 356947 1001950
rect 357709 1001947 357775 1001950
rect 358537 1001947 358603 1001950
rect 360193 1001947 360259 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 427169 1002010 427235 1002013
rect 433333 1002010 433399 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 426972 1002008 427235 1002010
rect 426972 1001952 427174 1002008
rect 427230 1001952 427235 1002008
rect 426972 1001950 427235 1001952
rect 433136 1002008 433399 1002010
rect 433136 1001952 433338 1002008
rect 433394 1001952 433399 1002008
rect 433136 1001950 433399 1001952
rect 421465 1001947 421531 1001950
rect 427169 1001947 427235 1001950
rect 433333 1001947 433399 1001950
rect 501689 1002010 501755 1002013
rect 502517 1002010 502583 1002013
rect 503345 1002010 503411 1002013
rect 504173 1002010 504239 1002013
rect 510337 1002010 510403 1002013
rect 501689 1002008 501952 1002010
rect 501689 1001952 501694 1002008
rect 501750 1001952 501952 1002008
rect 501689 1001950 501952 1001952
rect 502517 1002008 502780 1002010
rect 502517 1001952 502522 1002008
rect 502578 1001952 502780 1002008
rect 502517 1001950 502780 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 503976 1002008 504239 1002010
rect 503976 1001952 504178 1002008
rect 504234 1001952 504239 1002008
rect 503976 1001950 504239 1001952
rect 510140 1002008 510403 1002010
rect 510140 1001952 510342 1002008
rect 510398 1001952 510403 1002008
rect 510140 1001950 510403 1001952
rect 501689 1001947 501755 1001950
rect 502517 1001947 502583 1001950
rect 503345 1001947 503411 1001950
rect 504173 1001947 504239 1001950
rect 510337 1001947 510403 1001950
rect 555141 1002010 555207 1002013
rect 560017 1002010 560083 1002013
rect 555141 1002008 555404 1002010
rect 555141 1001952 555146 1002008
rect 555202 1001952 555404 1002008
rect 555141 1001950 555404 1001952
rect 559820 1002008 560083 1002010
rect 559820 1001952 560022 1002008
rect 560078 1001952 560083 1002008
rect 559820 1001950 560083 1001952
rect 555141 1001947 555207 1001950
rect 560017 1001947 560083 1001950
rect 550265 1001194 550331 1001197
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 550265 1001131 550331 1001134
rect 143993 1000650 144059 1000653
rect 147121 1000650 147187 1000653
rect 143993 1000648 147187 1000650
rect 143993 1000592 143998 1000648
rect 144054 1000592 147126 1000648
rect 147182 1000592 147187 1000648
rect 143993 1000590 147187 1000592
rect 143993 1000587 144059 1000590
rect 147121 1000587 147187 1000590
rect 308949 1000514 309015 1000517
rect 308752 1000512 309015 1000514
rect 308752 1000456 308954 1000512
rect 309010 1000456 309015 1000512
rect 308752 1000454 309015 1000456
rect 308949 1000451 309015 1000454
rect 204345 999018 204411 999021
rect 204345 999016 204516 999018
rect 204345 998960 204350 999016
rect 204406 998960 204516 999016
rect 204345 998958 204516 998960
rect 204345 998955 204411 998958
rect 203885 998746 203951 998749
rect 203780 998744 203951 998746
rect 203780 998688 203890 998744
rect 203946 998688 203951 998744
rect 203780 998686 203951 998688
rect 203885 998683 203951 998686
rect 202689 998610 202755 998613
rect 256969 998610 257035 998613
rect 553117 998610 553183 998613
rect 202689 998608 202952 998610
rect 202689 998552 202694 998608
rect 202750 998552 202952 998608
rect 202689 998550 202952 998552
rect 256969 998608 257140 998610
rect 256969 998552 256974 998608
rect 257030 998552 257140 998608
rect 256969 998550 257140 998552
rect 552920 998608 553183 998610
rect 552920 998552 553122 998608
rect 553178 998552 553183 998608
rect 552920 998550 553183 998552
rect 202689 998547 202755 998550
rect 256969 998547 257035 998550
rect 553117 998547 553183 998550
rect 203885 998474 203951 998477
rect 258993 998474 259059 998477
rect 203885 998472 204148 998474
rect 203885 998416 203890 998472
rect 203946 998416 204148 998472
rect 203885 998414 204148 998416
rect 258796 998472 259059 998474
rect 258796 998416 258998 998472
rect 259054 998416 259059 998472
rect 258796 998414 259059 998416
rect 203885 998411 203951 998414
rect 258993 998411 259059 998414
rect 307293 998474 307359 998477
rect 552289 998474 552355 998477
rect 307293 998472 307556 998474
rect 307293 998416 307298 998472
rect 307354 998416 307556 998472
rect 307293 998414 307556 998416
rect 552092 998472 552355 998474
rect 552092 998416 552294 998472
rect 552350 998416 552355 998472
rect 552092 998414 552355 998416
rect 307293 998411 307359 998414
rect 552289 998411 552355 998414
rect 195053 998338 195119 998341
rect 200205 998338 200271 998341
rect 195053 998336 200271 998338
rect 195053 998280 195058 998336
rect 195114 998280 200210 998336
rect 200266 998280 200271 998336
rect 195053 998278 200271 998280
rect 195053 998275 195119 998278
rect 200205 998275 200271 998278
rect 253657 998338 253723 998341
rect 306097 998338 306163 998341
rect 440877 998338 440943 998341
rect 253657 998336 253920 998338
rect 253657 998280 253662 998336
rect 253718 998280 253920 998336
rect 253657 998278 253920 998280
rect 306097 998336 306360 998338
rect 306097 998280 306102 998336
rect 306158 998280 306360 998336
rect 306097 998278 306360 998280
rect 440877 998336 451290 998338
rect 440877 998280 440882 998336
rect 440938 998280 451290 998336
rect 440877 998278 451290 998280
rect 253657 998275 253723 998278
rect 306097 998275 306163 998278
rect 440877 998275 440943 998278
rect 201861 998202 201927 998205
rect 205541 998202 205607 998205
rect 258165 998202 258231 998205
rect 201861 998200 202124 998202
rect 201861 998144 201866 998200
rect 201922 998144 202124 998200
rect 201861 998142 202124 998144
rect 205344 998200 205607 998202
rect 205344 998144 205546 998200
rect 205602 998144 205607 998200
rect 205344 998142 205607 998144
rect 257968 998200 258231 998202
rect 257968 998144 258170 998200
rect 258226 998144 258231 998200
rect 257968 998142 258231 998144
rect 201861 998139 201927 998142
rect 205541 998139 205607 998142
rect 258165 998139 258231 998142
rect 306925 998202 306991 998205
rect 451230 998202 451290 998278
rect 306925 998200 307188 998202
rect 306925 998144 306930 998200
rect 306986 998144 307188 998200
rect 306925 998142 307188 998144
rect 451230 998142 470610 998202
rect 306925 998139 306991 998142
rect 202689 998066 202755 998069
rect 202492 998064 202755 998066
rect 202492 998008 202694 998064
rect 202750 998008 202755 998064
rect 202492 998006 202755 998008
rect 202689 998003 202755 998006
rect 253289 998066 253355 998069
rect 256509 998066 256575 998069
rect 260189 998066 260255 998069
rect 253289 998064 253460 998066
rect 253289 998008 253294 998064
rect 253350 998008 253460 998064
rect 253289 998006 253460 998008
rect 256509 998064 256772 998066
rect 256509 998008 256514 998064
rect 256570 998008 256772 998064
rect 256509 998006 256772 998008
rect 260084 998064 260255 998066
rect 260084 998008 260194 998064
rect 260250 998008 260255 998064
rect 260084 998006 260255 998008
rect 253289 998003 253355 998006
rect 256509 998003 256575 998006
rect 260189 998003 260255 998006
rect 307753 998066 307819 998069
rect 310605 998066 310671 998069
rect 307753 998064 307924 998066
rect 307753 998008 307758 998064
rect 307814 998008 307924 998064
rect 307753 998006 307924 998008
rect 310605 998064 310868 998066
rect 310605 998008 310610 998064
rect 310666 998008 310868 998064
rect 310605 998006 310868 998008
rect 307753 998003 307819 998006
rect 310605 998003 310671 998006
rect 200665 997930 200731 997933
rect 252461 997930 252527 997933
rect 200665 997928 200836 997930
rect 200665 997872 200670 997928
rect 200726 997872 200836 997928
rect 200665 997870 200836 997872
rect 252264 997928 252527 997930
rect 252264 997872 252466 997928
rect 252522 997872 252527 997928
rect 252264 997870 252527 997872
rect 200665 997867 200731 997870
rect 252461 997867 252527 997870
rect 257337 997930 257403 997933
rect 259821 997930 259887 997933
rect 257337 997928 257600 997930
rect 257337 997872 257342 997928
rect 257398 997872 257600 997928
rect 257337 997870 257600 997872
rect 259624 997928 259887 997930
rect 259624 997872 259826 997928
rect 259882 997872 259887 997928
rect 259624 997870 259887 997872
rect 257337 997867 257403 997870
rect 259821 997867 259887 997870
rect 308949 997930 309015 997933
rect 308949 997928 309212 997930
rect 308949 997872 308954 997928
rect 309010 997872 309212 997928
rect 308949 997870 309212 997872
rect 308949 997867 309015 997870
rect 417057 997799 417363 997893
rect 418245 997803 418551 997897
rect 204713 997794 204779 997797
rect 260189 997794 260255 997797
rect 261845 997794 261911 997797
rect 306097 997794 306163 997797
rect 204713 997792 204976 997794
rect 204713 997736 204718 997792
rect 204774 997736 204976 997792
rect 204713 997734 204976 997736
rect 260189 997792 260452 997794
rect 260189 997736 260194 997792
rect 260250 997736 260452 997792
rect 260189 997734 260452 997736
rect 261845 997792 262108 997794
rect 261845 997736 261850 997792
rect 261906 997736 262108 997792
rect 261845 997734 262108 997736
rect 305900 997792 306163 997794
rect 305900 997736 306102 997792
rect 306158 997736 306163 997792
rect 305900 997734 306163 997736
rect 204713 997731 204779 997734
rect 260189 997731 260255 997734
rect 261845 997731 261911 997734
rect 306097 997731 306163 997734
rect 308121 997794 308187 997797
rect 309777 997794 309843 997797
rect 310605 997794 310671 997797
rect 308121 997792 308384 997794
rect 308121 997736 308126 997792
rect 308182 997736 308384 997792
rect 308121 997734 308384 997736
rect 309580 997792 309843 997794
rect 309580 997736 309782 997792
rect 309838 997736 309843 997792
rect 309580 997734 309843 997736
rect 310408 997792 310671 997794
rect 310408 997736 310610 997792
rect 310666 997736 310671 997792
rect 310408 997734 310671 997736
rect 308121 997731 308187 997734
rect 309777 997731 309843 997734
rect 310605 997731 310671 997734
rect 93485 997250 93551 997253
rect 89670 997248 93551 997250
rect 89670 997192 93490 997248
rect 93546 997192 93551 997248
rect 89670 997190 93551 997192
rect 89670 996978 89730 997190
rect 93485 997187 93551 997190
rect 117129 997250 117195 997253
rect 143717 997250 143783 997253
rect 117129 997248 143783 997250
rect 117129 997192 117134 997248
rect 117190 997192 143722 997248
rect 143778 997192 143783 997248
rect 117129 997190 143783 997192
rect 117129 997187 117195 997190
rect 143717 997187 143783 997190
rect 192518 997188 192524 997252
rect 192588 997250 192594 997252
rect 200205 997250 200271 997253
rect 192588 997248 200271 997250
rect 192588 997192 200210 997248
rect 200266 997192 200271 997248
rect 192588 997190 200271 997192
rect 192588 997188 192594 997190
rect 200205 997187 200271 997190
rect 298277 997250 298343 997253
rect 301681 997250 301747 997253
rect 298277 997248 301747 997250
rect 298277 997192 298282 997248
rect 298338 997192 301686 997248
rect 301742 997192 301747 997248
rect 298277 997190 301747 997192
rect 298277 997187 298343 997190
rect 301681 997187 301747 997190
rect 382089 997250 382155 997253
rect 388110 997250 388116 997252
rect 382089 997248 388116 997250
rect 382089 997192 382094 997248
rect 382150 997192 388116 997248
rect 382089 997190 388116 997192
rect 382089 997187 382155 997190
rect 388110 997188 388116 997190
rect 388180 997188 388186 997252
rect 470550 997250 470610 998142
rect 504541 998066 504607 998069
rect 504541 998064 504650 998066
rect 504541 998008 504546 998064
rect 504602 998008 504650 998064
rect 504541 998003 504650 998008
rect 504590 997796 504650 998003
rect 504582 997732 504588 997796
rect 504652 997732 504658 997796
rect 551461 997794 551527 997797
rect 551461 997792 551724 997794
rect 551461 997736 551466 997792
rect 551522 997736 551724 997792
rect 551461 997734 551724 997736
rect 551461 997731 551527 997734
rect 476430 997250 476436 997252
rect 470550 997190 476436 997250
rect 476430 997188 476436 997190
rect 476500 997188 476506 997252
rect 524045 997250 524111 997253
rect 529054 997250 529060 997252
rect 524045 997248 529060 997250
rect 524045 997192 524050 997248
rect 524106 997192 529060 997248
rect 524045 997190 529060 997192
rect 524045 997187 524111 997190
rect 529054 997188 529060 997190
rect 529124 997188 529130 997252
rect 80470 996918 89730 996978
rect 80470 995757 80530 996918
rect 89846 996916 89852 996980
rect 89916 996978 89922 996980
rect 92933 996978 92999 996981
rect 89916 996976 92999 996978
rect 89916 996920 92938 996976
rect 92994 996920 92999 996976
rect 89916 996918 92999 996920
rect 89916 996916 89922 996918
rect 92933 996915 92999 996918
rect 93577 996978 93643 996981
rect 94497 996978 94563 996981
rect 93577 996976 94563 996978
rect 93577 996920 93582 996976
rect 93638 996920 94502 996976
rect 94558 996920 94563 996976
rect 93577 996918 94563 996920
rect 93577 996915 93643 996918
rect 94497 996915 94563 996918
rect 116209 996978 116275 996981
rect 144177 996978 144243 996981
rect 197813 996978 197879 996981
rect 303061 996978 303127 996981
rect 116209 996976 144243 996978
rect 116209 996920 116214 996976
rect 116270 996920 144182 996976
rect 144238 996920 144243 996976
rect 116209 996918 144243 996920
rect 116209 996915 116275 996918
rect 144177 996915 144243 996918
rect 190410 996976 197879 996978
rect 190410 996920 197818 996976
rect 197874 996920 197879 996976
rect 190410 996918 197879 996920
rect 89670 996646 92674 996706
rect 89670 996298 89730 996646
rect 86358 996238 89730 996298
rect 92614 996298 92674 996646
rect 140262 996508 140268 996572
rect 140332 996570 140338 996572
rect 145741 996570 145807 996573
rect 190410 996570 190470 996918
rect 197813 996915 197879 996918
rect 288022 996976 303127 996978
rect 288022 996920 303066 996976
rect 303122 996920 303127 996976
rect 288022 996918 303127 996920
rect 140332 996568 145807 996570
rect 140332 996512 145746 996568
rect 145802 996512 145807 996568
rect 140332 996510 145807 996512
rect 140332 996508 140338 996510
rect 145741 996507 145807 996510
rect 188110 996510 190470 996570
rect 178861 996434 178927 996437
rect 183686 996434 183692 996436
rect 178861 996432 183692 996434
rect 178861 996376 178866 996432
rect 178922 996376 183692 996432
rect 178861 996374 183692 996376
rect 178861 996371 178927 996374
rect 183686 996372 183692 996374
rect 183756 996372 183762 996436
rect 92614 996238 93870 996298
rect 80421 995752 80530 995757
rect 80421 995696 80426 995752
rect 80482 995696 80530 995752
rect 80421 995694 80530 995696
rect 85941 995754 86007 995757
rect 86358 995754 86418 996238
rect 93301 996026 93367 996029
rect 87646 996024 93367 996026
rect 87646 995968 93306 996024
rect 93362 995968 93367 996024
rect 87646 995966 93367 995968
rect 93810 996026 93870 996238
rect 137970 996238 147690 996298
rect 126237 996162 126303 996165
rect 137970 996162 138030 996238
rect 126237 996160 138030 996162
rect 126237 996104 126242 996160
rect 126298 996104 138030 996160
rect 126237 996102 138030 996104
rect 126237 996099 126303 996102
rect 94681 996026 94747 996029
rect 144729 996026 144795 996029
rect 93810 996024 94747 996026
rect 93810 995968 94686 996024
rect 94742 995968 94747 996024
rect 93810 995966 94747 995968
rect 85941 995752 86418 995754
rect 85941 995696 85946 995752
rect 86002 995696 86418 995752
rect 85941 995694 86418 995696
rect 86585 995754 86651 995757
rect 87646 995754 87706 995966
rect 93301 995963 93367 995966
rect 94681 995963 94747 995966
rect 138246 996024 144795 996026
rect 138246 995968 144734 996024
rect 144790 995968 144795 996024
rect 138246 995966 144795 995968
rect 86585 995752 87706 995754
rect 86585 995696 86590 995752
rect 86646 995696 87706 995752
rect 86585 995694 87706 995696
rect 87873 995754 87939 995757
rect 98821 995754 98887 995757
rect 87873 995752 98887 995754
rect 87873 995696 87878 995752
rect 87934 995696 98826 995752
rect 98882 995696 98887 995752
rect 87873 995694 98887 995696
rect 80421 995691 80487 995694
rect 85941 995691 86007 995694
rect 86585 995691 86651 995694
rect 87873 995691 87939 995694
rect 98821 995691 98887 995694
rect 138013 995754 138079 995757
rect 138246 995754 138306 995966
rect 144729 995963 144795 995966
rect 138013 995752 138306 995754
rect 138013 995696 138018 995752
rect 138074 995696 138306 995752
rect 138013 995694 138306 995696
rect 141785 995754 141851 995757
rect 143993 995754 144059 995757
rect 141785 995752 144059 995754
rect 141785 995696 141790 995752
rect 141846 995696 143998 995752
rect 144054 995696 144059 995752
rect 141785 995694 144059 995696
rect 138013 995691 138079 995694
rect 141785 995691 141851 995694
rect 143993 995691 144059 995694
rect 88977 995482 89043 995485
rect 89846 995482 89852 995484
rect 88977 995480 89852 995482
rect 88977 995424 88982 995480
rect 89038 995424 89852 995480
rect 88977 995422 89852 995424
rect 88977 995419 89043 995422
rect 89846 995420 89852 995422
rect 89916 995420 89922 995484
rect 90265 995482 90331 995485
rect 92565 995482 92631 995485
rect 90265 995480 92631 995482
rect 90265 995424 90270 995480
rect 90326 995424 92570 995480
rect 92626 995424 92631 995480
rect 90265 995422 92631 995424
rect 90265 995419 90331 995422
rect 92565 995419 92631 995422
rect 137369 995482 137435 995485
rect 140262 995482 140268 995484
rect 137369 995480 140268 995482
rect 137369 995424 137374 995480
rect 137430 995424 140268 995480
rect 137369 995422 140268 995424
rect 137369 995419 137435 995422
rect 140262 995420 140268 995422
rect 140332 995420 140338 995484
rect 147630 995482 147690 996238
rect 154297 995754 154363 995757
rect 156830 995754 156890 996132
rect 154297 995752 156890 995754
rect 154297 995696 154302 995752
rect 154358 995696 156890 995752
rect 154297 995694 156890 995696
rect 154297 995691 154363 995694
rect 159222 995482 159282 996132
rect 187918 995890 187924 995892
rect 184062 995830 187924 995890
rect 175917 995754 175983 995757
rect 184062 995754 184122 995830
rect 187918 995828 187924 995830
rect 187988 995828 187994 995892
rect 188110 995757 188170 996510
rect 238518 996372 238524 996436
rect 238588 996434 238594 996436
rect 246573 996434 246639 996437
rect 238588 996432 246639 996434
rect 238588 996376 246578 996432
rect 246634 996376 246639 996432
rect 238588 996374 246639 996376
rect 238588 996372 238594 996374
rect 246573 996371 246639 996374
rect 175917 995752 184122 995754
rect 175917 995696 175922 995752
rect 175978 995696 184122 995752
rect 175917 995694 184122 995696
rect 188061 995752 188170 995757
rect 188061 995696 188066 995752
rect 188122 995696 188170 995752
rect 188061 995694 188170 995696
rect 188294 996238 200130 996298
rect 175917 995691 175983 995694
rect 188061 995691 188127 995694
rect 147630 995422 159282 995482
rect 183829 995482 183895 995485
rect 188294 995482 188354 996238
rect 199377 996026 199443 996029
rect 190410 996024 199443 996026
rect 190410 995968 199382 996024
rect 199438 995968 199443 996024
rect 190410 995966 199443 995968
rect 189441 995754 189507 995757
rect 190410 995754 190470 995966
rect 199377 995963 199443 995966
rect 200070 995890 200130 996238
rect 202321 995890 202387 995893
rect 200070 995888 202387 995890
rect 200070 995832 202326 995888
rect 202382 995832 202387 995888
rect 200070 995830 202387 995832
rect 202321 995827 202387 995830
rect 191741 995756 191807 995757
rect 192477 995756 192543 995757
rect 191741 995754 191788 995756
rect 189441 995752 190470 995754
rect 189441 995696 189446 995752
rect 189502 995696 190470 995752
rect 189441 995694 190470 995696
rect 191696 995752 191788 995754
rect 191696 995696 191746 995752
rect 191696 995694 191788 995696
rect 189441 995691 189507 995694
rect 191741 995692 191788 995694
rect 191852 995692 191858 995756
rect 192477 995754 192524 995756
rect 192432 995752 192524 995754
rect 192432 995696 192482 995752
rect 192432 995694 192524 995696
rect 192477 995692 192524 995694
rect 192588 995692 192594 995756
rect 194317 995754 194383 995757
rect 195053 995754 195119 995757
rect 194317 995752 195119 995754
rect 194317 995696 194322 995752
rect 194378 995696 195058 995752
rect 195114 995696 195119 995752
rect 194317 995694 195119 995696
rect 191741 995691 191807 995692
rect 192477 995691 192543 995692
rect 194317 995691 194383 995694
rect 195053 995691 195119 995694
rect 201677 995618 201743 995621
rect 203290 995618 203350 996132
rect 201677 995616 203350 995618
rect 201677 995560 201682 995616
rect 201738 995560 203350 995616
rect 201677 995558 203350 995560
rect 201677 995555 201743 995558
rect 183829 995480 188354 995482
rect 183829 995424 183834 995480
rect 183890 995424 188354 995480
rect 183829 995422 188354 995424
rect 183829 995419 183895 995422
rect 140497 995346 140563 995349
rect 144913 995346 144979 995349
rect 140497 995344 144979 995346
rect 140497 995288 140502 995344
rect 140558 995288 144918 995344
rect 144974 995288 144979 995344
rect 140497 995286 144979 995288
rect 140497 995283 140563 995286
rect 144913 995283 144979 995286
rect 168925 995346 168991 995349
rect 171685 995346 171751 995349
rect 183645 995348 183711 995349
rect 183645 995346 183692 995348
rect 168925 995344 171751 995346
rect 168925 995288 168930 995344
rect 168986 995288 171690 995344
rect 171746 995288 171751 995344
rect 168925 995286 171751 995288
rect 183600 995344 183692 995346
rect 183600 995288 183650 995344
rect 183600 995286 183692 995288
rect 168925 995283 168991 995286
rect 171685 995283 171751 995286
rect 183645 995284 183692 995286
rect 183756 995284 183762 995348
rect 188470 995284 188476 995348
rect 188540 995346 188546 995348
rect 208166 995346 208226 996132
rect 188540 995286 208226 995346
rect 188540 995284 188546 995286
rect 183645 995283 183711 995284
rect 77017 995074 77083 995077
rect 101397 995074 101463 995077
rect 77017 995072 101463 995074
rect 77017 995016 77022 995072
rect 77078 995016 101402 995072
rect 101458 995016 101463 995072
rect 77017 995014 101463 995016
rect 77017 995011 77083 995014
rect 101397 995011 101463 995014
rect 124857 995074 124923 995077
rect 154297 995074 154363 995077
rect 124857 995072 154363 995074
rect 124857 995016 124862 995072
rect 124918 995016 154302 995072
rect 154358 995016 154363 995072
rect 124857 995014 154363 995016
rect 124857 995011 124923 995014
rect 154297 995011 154363 995014
rect 169385 995074 169451 995077
rect 170673 995074 170739 995077
rect 169385 995072 170739 995074
rect 169385 995016 169390 995072
rect 169446 995016 170678 995072
rect 170734 995016 170739 995072
rect 169385 995014 170739 995016
rect 169385 995011 169451 995014
rect 170673 995011 170739 995014
rect 173157 995074 173223 995077
rect 209822 995074 209882 996132
rect 248137 996026 248203 996029
rect 249241 996026 249307 996029
rect 238710 996024 248203 996026
rect 238710 995968 248142 996024
rect 248198 995968 248203 996024
rect 238710 995966 248203 995968
rect 236545 995618 236611 995621
rect 238710 995618 238770 995966
rect 248137 995963 248203 995966
rect 248370 996024 249307 996026
rect 248370 995968 249246 996024
rect 249302 995968 249307 996024
rect 248370 995966 249307 995968
rect 240869 995754 240935 995757
rect 247033 995754 247099 995757
rect 240869 995752 247099 995754
rect 240869 995696 240874 995752
rect 240930 995696 247038 995752
rect 247094 995696 247099 995752
rect 240869 995694 247099 995696
rect 240869 995691 240935 995694
rect 247033 995691 247099 995694
rect 248370 995618 248430 995966
rect 249241 995963 249307 995966
rect 236545 995616 238770 995618
rect 236545 995560 236550 995616
rect 236606 995560 238770 995616
rect 236545 995558 238770 995560
rect 247174 995558 248430 995618
rect 255773 995618 255839 995621
rect 258398 995618 258458 996132
rect 255773 995616 258458 995618
rect 255773 995560 255778 995616
rect 255834 995560 258458 995616
rect 255773 995558 258458 995560
rect 236545 995555 236611 995558
rect 242065 995482 242131 995485
rect 247174 995482 247234 995558
rect 255773 995555 255839 995558
rect 242065 995480 247234 995482
rect 242065 995424 242070 995480
rect 242126 995424 247234 995480
rect 242065 995422 247234 995424
rect 242065 995419 242131 995422
rect 238569 995348 238635 995349
rect 238518 995284 238524 995348
rect 238588 995346 238635 995348
rect 252001 995346 252067 995349
rect 238588 995344 238680 995346
rect 238630 995288 238680 995344
rect 238588 995286 238680 995288
rect 248094 995344 252067 995346
rect 248094 995288 252006 995344
rect 252062 995288 252067 995344
rect 248094 995286 252067 995288
rect 238588 995284 238635 995286
rect 238569 995283 238635 995284
rect 239903 995210 239969 995213
rect 248094 995210 248154 995286
rect 252001 995283 252067 995286
rect 256049 995346 256115 995349
rect 259134 995346 259194 996132
rect 288022 995757 288082 996918
rect 303061 996915 303127 996918
rect 372705 996978 372771 996981
rect 399937 996978 400003 996981
rect 372705 996976 400003 996978
rect 372705 996920 372710 996976
rect 372766 996920 399942 996976
rect 399998 996920 400003 996976
rect 372705 996918 400003 996920
rect 372705 996915 372771 996918
rect 399937 996915 400003 996918
rect 439865 996978 439931 996981
rect 488901 996978 488967 996981
rect 439865 996976 488967 996978
rect 439865 996920 439870 996976
rect 439926 996920 488906 996976
rect 488962 996920 488967 996976
rect 439865 996918 488967 996920
rect 439865 996915 439931 996918
rect 488901 996915 488967 996918
rect 517053 996978 517119 996981
rect 540881 996978 540947 996981
rect 517053 996976 540947 996978
rect 517053 996920 517058 996976
rect 517114 996920 540886 996976
rect 540942 996920 540947 996976
rect 517053 996918 540947 996920
rect 517053 996915 517119 996918
rect 540881 996915 540947 996918
rect 590561 996978 590627 996981
rect 630806 996978 630812 996980
rect 590561 996976 630812 996978
rect 590561 996920 590566 996976
rect 590622 996920 630812 996976
rect 590561 996918 630812 996920
rect 590561 996915 590627 996918
rect 630806 996916 630812 996918
rect 630876 996916 630882 996980
rect 291326 996644 291332 996708
rect 291396 996706 291402 996708
rect 300301 996706 300367 996709
rect 291396 996704 300367 996706
rect 291396 996648 300306 996704
rect 300362 996648 300367 996704
rect 291396 996646 300367 996648
rect 291396 996644 291402 996646
rect 300301 996643 300367 996646
rect 372521 996706 372587 996709
rect 384982 996706 384988 996708
rect 372521 996704 384988 996706
rect 372521 996648 372526 996704
rect 372582 996648 384988 996704
rect 372521 996646 384988 996648
rect 372521 996643 372587 996646
rect 384982 996644 384988 996646
rect 385052 996644 385058 996708
rect 471237 996706 471303 996709
rect 476798 996706 476804 996708
rect 471237 996704 476804 996706
rect 471237 996648 471242 996704
rect 471298 996648 476804 996704
rect 471237 996646 476804 996648
rect 471237 996643 471303 996646
rect 476798 996644 476804 996646
rect 476868 996644 476874 996708
rect 516869 996706 516935 996709
rect 524045 996706 524111 996709
rect 516869 996704 524111 996706
rect 516869 996648 516874 996704
rect 516930 996648 524050 996704
rect 524106 996648 524111 996704
rect 516869 996646 524111 996648
rect 516869 996643 516935 996646
rect 524045 996643 524111 996646
rect 590561 996706 590627 996709
rect 629702 996706 629708 996708
rect 590561 996704 629708 996706
rect 590561 996648 590566 996704
rect 590622 996648 629708 996704
rect 590561 996646 629708 996648
rect 590561 996643 590627 996646
rect 629702 996644 629708 996646
rect 629772 996644 629778 996708
rect 372337 996434 372403 996437
rect 382089 996434 382155 996437
rect 372337 996432 382155 996434
rect 372337 996376 372342 996432
rect 372398 996376 382094 996432
rect 382150 996376 382155 996432
rect 372337 996374 382155 996376
rect 372337 996371 372403 996374
rect 382089 996371 382155 996374
rect 439681 996434 439747 996437
rect 481214 996434 481220 996436
rect 439681 996432 481220 996434
rect 439681 996376 439686 996432
rect 439742 996376 481220 996432
rect 439681 996374 481220 996376
rect 439681 996371 439747 996374
rect 481214 996372 481220 996374
rect 481284 996372 481290 996436
rect 516685 996434 516751 996437
rect 549437 996434 549503 996437
rect 516685 996432 528018 996434
rect 516685 996376 516690 996432
rect 516746 996376 528018 996432
rect 516685 996374 528018 996376
rect 516685 996371 516751 996374
rect 382273 996298 382339 996301
rect 399845 996298 399911 996301
rect 290782 996238 301514 996298
rect 287973 995752 288082 995757
rect 287973 995696 287978 995752
rect 288034 995696 288082 995752
rect 287973 995694 288082 995696
rect 290549 995754 290615 995757
rect 290782 995754 290842 996238
rect 293358 995966 299858 996026
rect 290549 995752 290842 995754
rect 290549 995696 290554 995752
rect 290610 995696 290842 995752
rect 290549 995694 290842 995696
rect 291101 995754 291167 995757
rect 293358 995754 293418 995966
rect 291101 995752 293418 995754
rect 291101 995696 291106 995752
rect 291162 995696 293418 995752
rect 291101 995694 293418 995696
rect 293585 995754 293651 995757
rect 299565 995754 299631 995757
rect 293585 995752 299631 995754
rect 293585 995696 293590 995752
rect 293646 995696 299570 995752
rect 299626 995696 299631 995752
rect 293585 995694 299631 995696
rect 287973 995691 288039 995694
rect 290549 995691 290615 995694
rect 291101 995691 291167 995694
rect 293585 995691 293651 995694
rect 299565 995691 299631 995694
rect 299798 995618 299858 995966
rect 301454 995890 301514 996238
rect 382273 996296 399911 996298
rect 382273 996240 382278 996296
rect 382334 996240 399850 996296
rect 399906 996240 399911 996296
rect 382273 996238 399911 996240
rect 382273 996235 382339 996238
rect 399845 996235 399911 996238
rect 304073 996162 304139 996165
rect 303876 996160 304139 996162
rect 303876 996104 304078 996160
rect 304134 996104 304139 996160
rect 469857 996162 469923 996165
rect 519537 996162 519603 996165
rect 469857 996160 489930 996162
rect 303876 996102 304139 996104
rect 304073 996099 304139 996102
rect 301454 995830 306390 995890
rect 302877 995618 302943 995621
rect 299798 995616 302943 995618
rect 299798 995560 302882 995616
rect 302938 995560 302943 995616
rect 299798 995558 302943 995560
rect 302877 995555 302943 995558
rect 291377 995348 291443 995349
rect 256049 995344 259194 995346
rect 256049 995288 256054 995344
rect 256110 995288 259194 995344
rect 256049 995286 259194 995288
rect 256049 995283 256115 995286
rect 291326 995284 291332 995348
rect 291396 995346 291443 995348
rect 291745 995346 291811 995349
rect 301497 995346 301563 995349
rect 291396 995344 291488 995346
rect 291438 995288 291488 995344
rect 291396 995286 291488 995288
rect 291745 995344 301563 995346
rect 291745 995288 291750 995344
rect 291806 995288 301502 995344
rect 301558 995288 301563 995344
rect 291745 995286 301563 995288
rect 291396 995284 291443 995286
rect 291377 995283 291443 995284
rect 291745 995283 291811 995286
rect 301497 995283 301563 995286
rect 301681 995346 301747 995349
rect 304441 995346 304507 995349
rect 301681 995344 304507 995346
rect 301681 995288 301686 995344
rect 301742 995288 304446 995344
rect 304502 995288 304507 995344
rect 301681 995286 304507 995288
rect 306330 995346 306390 995830
rect 307201 995346 307267 995349
rect 306330 995344 307267 995346
rect 306330 995288 307206 995344
rect 307262 995288 307267 995344
rect 306330 995286 307267 995288
rect 301681 995283 301747 995286
rect 304441 995283 304507 995286
rect 307201 995283 307267 995286
rect 239903 995208 248154 995210
rect 239903 995152 239908 995208
rect 239964 995152 248154 995208
rect 239903 995150 248154 995152
rect 239903 995147 239969 995150
rect 173157 995072 209882 995074
rect 173157 995016 173162 995072
rect 173218 995016 209882 995072
rect 173157 995014 209882 995016
rect 248321 995074 248387 995077
rect 251817 995074 251883 995077
rect 248321 995072 251883 995074
rect 248321 995016 248326 995072
rect 248382 995016 251822 995072
rect 251878 995016 251883 995072
rect 248321 995014 251883 995016
rect 173157 995011 173223 995014
rect 248321 995011 248387 995014
rect 251817 995011 251883 995014
rect 280797 995074 280863 995077
rect 312862 995074 312922 996132
rect 383285 996026 383351 996029
rect 383285 996024 386706 996026
rect 383285 995968 383290 996024
rect 383346 995968 386706 996024
rect 383285 995966 386706 995968
rect 383285 995963 383351 995966
rect 385033 995756 385099 995757
rect 384982 995692 384988 995756
rect 385052 995754 385099 995756
rect 386646 995754 386706 995966
rect 388621 995754 388687 995757
rect 416129 995754 416195 995757
rect 385052 995752 385144 995754
rect 385094 995696 385144 995752
rect 385052 995694 385144 995696
rect 386646 995752 388687 995754
rect 386646 995696 388626 995752
rect 388682 995696 388687 995752
rect 386646 995694 388687 995696
rect 385052 995692 385099 995694
rect 385033 995691 385099 995692
rect 388621 995691 388687 995694
rect 389130 995752 416195 995754
rect 389130 995696 416134 995752
rect 416190 995696 416195 995752
rect 389130 995694 416195 995696
rect 382917 995482 382983 995485
rect 387885 995482 387951 995485
rect 388161 995484 388227 995485
rect 382917 995480 387951 995482
rect 382917 995424 382922 995480
rect 382978 995424 387890 995480
rect 387946 995424 387951 995480
rect 382917 995422 387951 995424
rect 382917 995419 382983 995422
rect 387885 995419 387951 995422
rect 388110 995420 388116 995484
rect 388180 995482 388227 995484
rect 388180 995480 388272 995482
rect 388222 995424 388272 995480
rect 388180 995422 388272 995424
rect 388180 995420 388227 995422
rect 388161 995419 388227 995420
rect 389130 995346 389190 995694
rect 416129 995691 416195 995694
rect 399845 995482 399911 995485
rect 415393 995482 415459 995485
rect 399845 995480 415459 995482
rect 399845 995424 399850 995480
rect 399906 995424 415398 995480
rect 415454 995424 415459 995480
rect 399845 995422 415459 995424
rect 399845 995419 399911 995422
rect 415393 995419 415459 995422
rect 388302 995286 389190 995346
rect 380893 995210 380959 995213
rect 388302 995210 388362 995286
rect 380893 995208 388362 995210
rect 380893 995152 380898 995208
rect 380954 995152 388362 995208
rect 380893 995150 388362 995152
rect 380893 995147 380959 995150
rect 280797 995072 312922 995074
rect 280797 995016 280802 995072
rect 280858 995016 312922 995072
rect 280797 995014 312922 995016
rect 388437 995074 388503 995077
rect 430990 995074 431050 996132
rect 469857 996104 469862 996160
rect 469918 996104 489930 996160
rect 519537 996160 527190 996162
rect 469857 996102 489930 996104
rect 469857 996099 469923 996102
rect 454861 995890 454927 995893
rect 454861 995888 482202 995890
rect 454861 995832 454866 995888
rect 454922 995832 482202 995888
rect 454861 995830 482202 995832
rect 454861 995827 454927 995830
rect 482142 995754 482202 995830
rect 483749 995754 483815 995757
rect 485589 995756 485655 995757
rect 485589 995754 485636 995756
rect 482142 995752 483815 995754
rect 482142 995696 483754 995752
rect 483810 995696 483815 995752
rect 482142 995694 483815 995696
rect 485544 995752 485636 995754
rect 485544 995696 485594 995752
rect 485544 995694 485636 995696
rect 483749 995691 483815 995694
rect 485589 995692 485636 995694
rect 485700 995692 485706 995756
rect 485589 995691 485655 995692
rect 446397 995618 446463 995621
rect 474733 995618 474799 995621
rect 480713 995618 480779 995621
rect 481265 995620 481331 995621
rect 446397 995616 474799 995618
rect 446397 995560 446402 995616
rect 446458 995560 474738 995616
rect 474794 995560 474799 995616
rect 446397 995558 474799 995560
rect 446397 995555 446463 995558
rect 474733 995555 474799 995558
rect 474966 995616 480779 995618
rect 474966 995560 480718 995616
rect 480774 995560 480779 995616
rect 474966 995558 480779 995560
rect 471421 995346 471487 995349
rect 474966 995346 475026 995558
rect 480713 995555 480779 995558
rect 481214 995556 481220 995620
rect 481284 995618 481331 995620
rect 489870 995618 489930 996102
rect 503662 995828 503668 995892
rect 503732 995890 503738 995892
rect 506197 995890 506263 995893
rect 503732 995888 506263 995890
rect 503732 995832 506202 995888
rect 506258 995832 506263 995888
rect 503732 995830 506263 995832
rect 503732 995828 503738 995830
rect 506197 995827 506263 995830
rect 506430 995618 506490 996132
rect 481284 995616 481376 995618
rect 481326 995560 481376 995616
rect 481284 995558 481376 995560
rect 489870 995558 506490 995618
rect 481284 995556 481331 995558
rect 481265 995555 481331 995556
rect 476481 995348 476547 995349
rect 471421 995344 475026 995346
rect 471421 995288 471426 995344
rect 471482 995288 475026 995344
rect 471421 995286 475026 995288
rect 471421 995283 471487 995286
rect 476430 995284 476436 995348
rect 476500 995346 476547 995348
rect 476500 995344 476592 995346
rect 476542 995288 476592 995344
rect 476500 995286 476592 995288
rect 476500 995284 476547 995286
rect 476798 995284 476804 995348
rect 476868 995346 476874 995348
rect 507166 995346 507226 996132
rect 476868 995286 507226 995346
rect 476868 995284 476874 995286
rect 476481 995283 476547 995284
rect 388437 995072 431050 995074
rect 388437 995016 388442 995072
rect 388498 995016 431050 995072
rect 388437 995014 431050 995016
rect 472249 995074 472315 995077
rect 476941 995074 477007 995077
rect 472249 995072 477007 995074
rect 472249 995016 472254 995072
rect 472310 995016 476946 995072
rect 477002 995016 477007 995072
rect 472249 995014 477007 995016
rect 280797 995011 280863 995014
rect 388437 995011 388503 995014
rect 472249 995011 472315 995014
rect 476941 995011 477007 995014
rect 480713 995074 480779 995077
rect 508822 995074 508882 996132
rect 519537 996104 519542 996160
rect 519598 996104 527190 996160
rect 519537 996102 527190 996104
rect 519537 996099 519603 996102
rect 522481 995754 522547 995757
rect 526069 995754 526135 995757
rect 522481 995752 526135 995754
rect 522481 995696 522486 995752
rect 522542 995696 526074 995752
rect 526130 995696 526135 995752
rect 522481 995694 526135 995696
rect 522481 995691 522547 995694
rect 526069 995691 526135 995694
rect 523861 995482 523927 995485
rect 524781 995482 524847 995485
rect 523861 995480 524847 995482
rect 523861 995424 523866 995480
rect 523922 995424 524786 995480
rect 524842 995424 524847 995480
rect 523861 995422 524847 995424
rect 527130 995482 527190 996102
rect 527958 995754 528018 996374
rect 536790 996432 549503 996434
rect 536790 996376 549442 996432
rect 549498 996376 549503 996432
rect 536790 996374 549503 996376
rect 528553 995754 528619 995757
rect 529105 995756 529171 995757
rect 533521 995756 533587 995757
rect 527958 995752 528619 995754
rect 527958 995696 528558 995752
rect 528614 995696 528619 995752
rect 527958 995694 528619 995696
rect 528553 995691 528619 995694
rect 529054 995692 529060 995756
rect 529124 995754 529171 995756
rect 529124 995752 529216 995754
rect 529166 995696 529216 995752
rect 529124 995694 529216 995696
rect 529124 995692 529171 995694
rect 533470 995692 533476 995756
rect 533540 995754 533587 995756
rect 536557 995754 536623 995757
rect 536790 995754 536850 996374
rect 549437 996371 549503 996374
rect 590561 996434 590627 996437
rect 590561 996432 633450 996434
rect 590561 996376 590566 996432
rect 590622 996376 633450 996432
rect 590561 996374 633450 996376
rect 590561 996371 590627 996374
rect 625613 996026 625679 996029
rect 625613 996024 629586 996026
rect 625613 995968 625618 996024
rect 625674 995968 629586 996024
rect 625613 995966 629586 995968
rect 625613 995963 625679 995966
rect 533540 995752 533632 995754
rect 533582 995696 533632 995752
rect 533540 995694 533632 995696
rect 536557 995752 536850 995754
rect 536557 995696 536562 995752
rect 536618 995696 536850 995752
rect 536557 995694 536850 995696
rect 625797 995754 625863 995757
rect 627177 995754 627243 995757
rect 625797 995752 627243 995754
rect 625797 995696 625802 995752
rect 625858 995696 627182 995752
rect 627238 995696 627243 995752
rect 625797 995694 627243 995696
rect 533540 995692 533587 995694
rect 529105 995691 529171 995692
rect 533521 995691 533587 995692
rect 536557 995691 536623 995694
rect 625797 995691 625863 995694
rect 627177 995691 627243 995694
rect 629526 995621 629586 995966
rect 629753 995756 629819 995757
rect 630857 995756 630923 995757
rect 629702 995692 629708 995756
rect 629772 995754 629819 995756
rect 629772 995752 629864 995754
rect 629814 995696 629864 995752
rect 629772 995694 629864 995696
rect 629772 995692 629819 995694
rect 630806 995692 630812 995756
rect 630876 995754 630923 995756
rect 633390 995754 633450 996374
rect 634537 995754 634603 995757
rect 630876 995752 630968 995754
rect 630918 995696 630968 995752
rect 630876 995694 630968 995696
rect 633390 995752 634603 995754
rect 633390 995696 634542 995752
rect 634598 995696 634603 995752
rect 633390 995694 634603 995696
rect 630876 995692 630923 995694
rect 629753 995691 629819 995692
rect 630857 995691 630923 995692
rect 634537 995691 634603 995694
rect 637665 995754 637731 995757
rect 642081 995754 642147 995757
rect 637665 995752 642147 995754
rect 637665 995696 637670 995752
rect 637726 995696 642086 995752
rect 642142 995696 642147 995752
rect 637665 995694 642147 995696
rect 637665 995691 637731 995694
rect 642081 995691 642147 995694
rect 629526 995616 629635 995621
rect 629526 995560 629574 995616
rect 629630 995560 629635 995616
rect 629526 995558 629635 995560
rect 629569 995555 629635 995558
rect 532693 995482 532759 995485
rect 527130 995480 532759 995482
rect 527130 995424 532698 995480
rect 532754 995424 532759 995480
rect 527130 995422 532759 995424
rect 523861 995419 523927 995422
rect 524781 995419 524847 995422
rect 532693 995419 532759 995422
rect 617149 995346 617215 995349
rect 635825 995346 635891 995349
rect 617149 995344 635891 995346
rect 617149 995288 617154 995344
rect 617210 995288 635830 995344
rect 635886 995288 635891 995344
rect 617149 995286 635891 995288
rect 617149 995283 617215 995286
rect 635825 995283 635891 995286
rect 538121 995210 538187 995213
rect 538305 995210 538371 995213
rect 538121 995208 538371 995210
rect 538121 995152 538126 995208
rect 538182 995152 538310 995208
rect 538366 995152 538371 995208
rect 538121 995150 538371 995152
rect 538121 995147 538187 995150
rect 538305 995147 538371 995150
rect 480713 995072 508882 995074
rect 480713 995016 480718 995072
rect 480774 995016 508882 995072
rect 480713 995014 508882 995016
rect 509049 995074 509115 995077
rect 511073 995074 511139 995077
rect 509049 995072 511139 995074
rect 509049 995016 509054 995072
rect 509110 995016 511078 995072
rect 511134 995016 511139 995072
rect 509049 995014 511139 995016
rect 480713 995011 480779 995014
rect 509049 995011 509115 995014
rect 511073 995011 511139 995014
rect 517513 995074 517579 995077
rect 530025 995074 530091 995077
rect 517513 995072 530091 995074
rect 517513 995016 517518 995072
rect 517574 995016 530030 995072
rect 530086 995016 530091 995072
rect 517513 995014 530091 995016
rect 517513 995011 517579 995014
rect 530025 995011 530091 995014
rect 590561 995074 590627 995077
rect 660573 995074 660639 995077
rect 590561 995072 660639 995074
rect 590561 995016 590566 995072
rect 590622 995016 660578 995072
rect 660634 995016 660639 995072
rect 590561 995014 660639 995016
rect 590561 995011 590627 995014
rect 660573 995011 660639 995014
rect 81985 994802 82051 994805
rect 97257 994802 97323 994805
rect 81985 994800 97323 994802
rect 81985 994744 81990 994800
rect 82046 994744 97262 994800
rect 97318 994744 97323 994800
rect 81985 994742 97323 994744
rect 81985 994739 82051 994742
rect 97257 994739 97323 994742
rect 133413 994802 133479 994805
rect 138749 994802 138815 994805
rect 133413 994800 138815 994802
rect 133413 994744 133418 994800
rect 133474 994744 138754 994800
rect 138810 994744 138815 994800
rect 133413 994742 138815 994744
rect 133413 994739 133479 994742
rect 138749 994739 138815 994742
rect 138933 994802 138999 994805
rect 144177 994802 144243 994805
rect 138933 994800 144243 994802
rect 138933 994744 138938 994800
rect 138994 994744 144182 994800
rect 144238 994744 144243 994800
rect 138933 994742 144243 994744
rect 138933 994739 138999 994742
rect 144177 994739 144243 994742
rect 181437 994802 181503 994805
rect 207013 994802 207079 994805
rect 181437 994800 207079 994802
rect 181437 994744 181442 994800
rect 181498 994744 207018 994800
rect 207074 994744 207079 994800
rect 181437 994742 207079 994744
rect 181437 994739 181503 994742
rect 207013 994739 207079 994742
rect 231577 994802 231643 994805
rect 255773 994802 255839 994805
rect 231577 994800 255839 994802
rect 231577 994744 231582 994800
rect 231638 994744 255778 994800
rect 255834 994744 255839 994800
rect 231577 994742 255839 994744
rect 231577 994739 231643 994742
rect 255773 994739 255839 994742
rect 285949 994802 286015 994805
rect 309133 994802 309199 994805
rect 285949 994800 309199 994802
rect 285949 994744 285954 994800
rect 286010 994744 309138 994800
rect 309194 994744 309199 994800
rect 285949 994742 309199 994744
rect 285949 994739 286015 994742
rect 309133 994739 309199 994742
rect 374821 994802 374887 994805
rect 392117 994802 392183 994805
rect 374821 994800 392183 994802
rect 374821 994744 374826 994800
rect 374882 994744 392122 994800
rect 392178 994744 392183 994800
rect 374821 994742 392183 994744
rect 374821 994739 374887 994742
rect 392117 994739 392183 994742
rect 464337 994802 464403 994805
rect 481633 994802 481699 994805
rect 464337 994800 481699 994802
rect 464337 994744 464342 994800
rect 464398 994744 481638 994800
rect 481694 994744 481699 994800
rect 464337 994742 481699 994744
rect 464337 994739 464403 994742
rect 481633 994739 481699 994742
rect 518157 994802 518223 994805
rect 537385 994802 537451 994805
rect 518157 994800 537451 994802
rect 518157 994744 518162 994800
rect 518218 994744 537390 994800
rect 537446 994744 537451 994800
rect 518157 994742 537451 994744
rect 518157 994739 518223 994742
rect 537385 994739 537451 994742
rect 570229 994802 570295 994805
rect 635181 994802 635247 994805
rect 570229 994800 635247 994802
rect 570229 994744 570234 994800
rect 570290 994744 635186 994800
rect 635242 994744 635247 994800
rect 570229 994742 635247 994744
rect 570229 994739 570295 994742
rect 635181 994739 635247 994742
rect 85297 994530 85363 994533
rect 93577 994530 93643 994533
rect 100017 994530 100083 994533
rect 85297 994528 93643 994530
rect 85297 994472 85302 994528
rect 85358 994472 93582 994528
rect 93638 994472 93643 994528
rect 85297 994470 93643 994472
rect 85297 994467 85363 994470
rect 93577 994467 93643 994470
rect 93810 994528 100083 994530
rect 93810 994472 100022 994528
rect 100078 994472 100083 994528
rect 93810 994470 100083 994472
rect 84469 994258 84535 994261
rect 93810 994258 93870 994470
rect 100017 994467 100083 994470
rect 133137 994530 133203 994533
rect 140589 994530 140655 994533
rect 133137 994528 140655 994530
rect 133137 994472 133142 994528
rect 133198 994472 140594 994528
rect 140650 994472 140655 994528
rect 133137 994470 140655 994472
rect 133137 994467 133203 994470
rect 140589 994467 140655 994470
rect 140773 994530 140839 994533
rect 144545 994530 144611 994533
rect 140773 994528 144611 994530
rect 140773 994472 140778 994528
rect 140834 994472 144550 994528
rect 144606 994472 144611 994528
rect 140773 994470 144611 994472
rect 140773 994467 140839 994470
rect 144545 994467 144611 994470
rect 187601 994530 187667 994533
rect 203517 994530 203583 994533
rect 243261 994532 243327 994533
rect 243261 994530 243308 994532
rect 187601 994528 203583 994530
rect 187601 994472 187606 994528
rect 187662 994472 203522 994528
rect 203578 994472 203583 994528
rect 187601 994470 203583 994472
rect 243216 994528 243308 994530
rect 243216 994472 243266 994528
rect 243216 994470 243308 994472
rect 187601 994467 187667 994470
rect 203517 994467 203583 994470
rect 243261 994468 243308 994470
rect 243372 994468 243378 994532
rect 243537 994530 243603 994533
rect 259453 994530 259519 994533
rect 243537 994528 259519 994530
rect 243537 994472 243542 994528
rect 243598 994472 259458 994528
rect 259514 994472 259519 994528
rect 243537 994470 259519 994472
rect 243261 994467 243327 994468
rect 243537 994467 243603 994470
rect 259453 994467 259519 994470
rect 287145 994530 287211 994533
rect 304257 994530 304323 994533
rect 287145 994528 304323 994530
rect 287145 994472 287150 994528
rect 287206 994472 304262 994528
rect 304318 994472 304323 994528
rect 287145 994470 304323 994472
rect 287145 994467 287211 994470
rect 304257 994467 304323 994470
rect 383101 994530 383167 994533
rect 400857 994530 400923 994533
rect 383101 994528 400923 994530
rect 383101 994472 383106 994528
rect 383162 994472 400862 994528
rect 400918 994472 400923 994528
rect 383101 994470 400923 994472
rect 383101 994467 383167 994470
rect 400857 994467 400923 994470
rect 465717 994530 465783 994533
rect 478597 994530 478663 994533
rect 465717 994528 478663 994530
rect 465717 994472 465722 994528
rect 465778 994472 478602 994528
rect 478658 994472 478663 994528
rect 465717 994470 478663 994472
rect 465717 994467 465783 994470
rect 478597 994467 478663 994470
rect 517697 994530 517763 994533
rect 532509 994530 532575 994533
rect 517697 994528 532575 994530
rect 517697 994472 517702 994528
rect 517758 994472 532514 994528
rect 532570 994472 532575 994528
rect 517697 994470 532575 994472
rect 517697 994467 517763 994470
rect 532509 994467 532575 994470
rect 572897 994530 572963 994533
rect 631501 994530 631567 994533
rect 572897 994528 631567 994530
rect 572897 994472 572902 994528
rect 572958 994472 631506 994528
rect 631562 994472 631567 994528
rect 572897 994470 631567 994472
rect 572897 994467 572963 994470
rect 631501 994467 631567 994470
rect 84469 994256 93870 994258
rect 84469 994200 84474 994256
rect 84530 994200 93870 994256
rect 84469 994198 93870 994200
rect 135897 994258 135963 994261
rect 152457 994258 152523 994261
rect 135897 994256 152523 994258
rect 135897 994200 135902 994256
rect 135958 994200 152462 994256
rect 152518 994200 152523 994256
rect 135897 994198 152523 994200
rect 84469 994195 84535 994198
rect 135897 994195 135963 994198
rect 152457 994195 152523 994198
rect 190361 994258 190427 994261
rect 200941 994258 201007 994261
rect 190361 994256 201007 994258
rect 190361 994200 190366 994256
rect 190422 994200 200946 994256
rect 201002 994200 201007 994256
rect 190361 994198 201007 994200
rect 190361 994195 190427 994198
rect 200941 994195 201007 994198
rect 226374 994196 226380 994260
rect 226444 994258 226450 994260
rect 251449 994258 251515 994261
rect 226444 994256 251515 994258
rect 226444 994200 251454 994256
rect 251510 994200 251515 994256
rect 226444 994198 251515 994200
rect 226444 994196 226450 994198
rect 251449 994195 251515 994198
rect 278630 994196 278636 994260
rect 278700 994258 278706 994260
rect 316401 994258 316467 994261
rect 278700 994256 316467 994258
rect 278700 994200 316406 994256
rect 316462 994200 316467 994256
rect 278700 994198 316467 994200
rect 278700 994196 278706 994198
rect 316401 994195 316467 994198
rect 449157 994258 449223 994261
rect 477953 994258 478019 994261
rect 449157 994256 478019 994258
rect 449157 994200 449162 994256
rect 449218 994200 477958 994256
rect 478014 994200 478019 994256
rect 449157 994198 478019 994200
rect 449157 994195 449223 994198
rect 477953 994195 478019 994198
rect 520917 994258 520983 994261
rect 532141 994258 532207 994261
rect 520917 994256 532207 994258
rect 520917 994200 520922 994256
rect 520978 994200 532146 994256
rect 532202 994200 532207 994256
rect 520917 994198 532207 994200
rect 520917 994195 520983 994198
rect 532141 994195 532207 994198
rect 568205 994258 568271 994261
rect 627913 994258 627979 994261
rect 568205 994256 627979 994258
rect 568205 994200 568210 994256
rect 568266 994200 627918 994256
rect 627974 994200 627979 994256
rect 568205 994198 627979 994200
rect 568205 994195 568271 994198
rect 627913 994195 627979 994198
rect 138749 993986 138815 993989
rect 145557 993986 145623 993989
rect 138749 993984 145623 993986
rect 138749 993928 138754 993984
rect 138810 993928 145562 993984
rect 145618 993928 145623 993984
rect 138749 993926 145623 993928
rect 138749 993923 138815 993926
rect 145557 993923 145623 993926
rect 188797 993986 188863 993989
rect 200757 993986 200823 993989
rect 188797 993984 200823 993986
rect 188797 993928 188802 993984
rect 188858 993928 200762 993984
rect 200818 993928 200823 993984
rect 188797 993926 200823 993928
rect 188797 993923 188863 993926
rect 200757 993923 200823 993926
rect 234521 993986 234587 993989
rect 243537 993986 243603 993989
rect 249057 993986 249123 993989
rect 234521 993984 243603 993986
rect 234521 993928 234526 993984
rect 234582 993928 243542 993984
rect 243598 993928 243603 993984
rect 234521 993926 243603 993928
rect 234521 993923 234587 993926
rect 243537 993923 243603 993926
rect 248370 993984 249123 993986
rect 248370 993928 249062 993984
rect 249118 993928 249123 993984
rect 248370 993926 249123 993928
rect 140589 993714 140655 993717
rect 149697 993714 149763 993717
rect 140589 993712 149763 993714
rect 140589 993656 140594 993712
rect 140650 993656 149702 993712
rect 149758 993656 149763 993712
rect 140589 993654 149763 993656
rect 140589 993651 140655 993654
rect 149697 993651 149763 993654
rect 239581 993714 239647 993717
rect 248370 993714 248430 993926
rect 249057 993923 249123 993926
rect 295517 993986 295583 993989
rect 310513 993986 310579 993989
rect 295517 993984 310579 993986
rect 295517 993928 295522 993984
rect 295578 993928 310518 993984
rect 310574 993928 310579 993984
rect 295517 993926 310579 993928
rect 295517 993923 295583 993926
rect 310513 993923 310579 993926
rect 239581 993712 248430 993714
rect 239581 993656 239586 993712
rect 239642 993656 248430 993712
rect 239581 993654 248430 993656
rect 239581 993651 239647 993654
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 42149 967602 42215 967605
rect 42609 967602 42675 967605
rect 42149 967600 42675 967602
rect 42149 967544 42154 967600
rect 42210 967544 42614 967600
rect 42670 967544 42675 967600
rect 42149 967542 42675 967544
rect 42149 967539 42215 967542
rect 42609 967539 42675 967542
rect 41454 967132 41460 967196
rect 41524 967194 41530 967196
rect 41781 967194 41847 967197
rect 41524 967192 41847 967194
rect 41524 967136 41786 967192
rect 41842 967136 41847 967192
rect 41524 967134 41847 967136
rect 41524 967132 41530 967134
rect 41781 967131 41847 967134
rect 42149 967194 42215 967197
rect 43437 967194 43503 967197
rect 42149 967192 43503 967194
rect 42149 967136 42154 967192
rect 42210 967136 43442 967192
rect 43498 967136 43503 967192
rect 42149 967134 43503 967136
rect 42149 967131 42215 967134
rect 43437 967131 43503 967134
rect 673361 966650 673427 966653
rect 675109 966650 675175 966653
rect 673361 966648 675175 966650
rect 673361 966592 673366 966648
rect 673422 966592 675114 966648
rect 675170 966592 675175 966648
rect 673361 966590 675175 966592
rect 673361 966587 673427 966590
rect 675109 966587 675175 966590
rect 675661 966516 675727 966517
rect 675661 966512 675708 966516
rect 675772 966514 675778 966516
rect 675661 966456 675666 966512
rect 675661 966452 675708 966456
rect 675772 966454 675818 966514
rect 675772 966452 675778 966454
rect 675661 966451 675727 966452
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 42425 964746 42491 964749
rect 43437 964746 43503 964749
rect 42425 964744 43503 964746
rect 42425 964688 42430 964744
rect 42486 964688 43442 964744
rect 43498 964688 43503 964744
rect 42425 964686 43503 964688
rect 42425 964683 42491 964686
rect 43437 964683 43503 964686
rect 675293 964746 675359 964749
rect 676806 964746 676812 964748
rect 675293 964744 676812 964746
rect 675293 964688 675298 964744
rect 675354 964688 676812 964744
rect 675293 964686 676812 964688
rect 675293 964683 675359 964686
rect 676806 964684 676812 964686
rect 676876 964684 676882 964748
rect 42425 963930 42491 963933
rect 43253 963930 43319 963933
rect 42425 963928 43319 963930
rect 42425 963872 42430 963928
rect 42486 963872 43258 963928
rect 43314 963872 43319 963928
rect 42425 963870 43319 963872
rect 42425 963867 42491 963870
rect 43253 963867 43319 963870
rect 42425 963386 42491 963389
rect 43069 963386 43135 963389
rect 42425 963384 43135 963386
rect 42425 963328 42430 963384
rect 42486 963328 43074 963384
rect 43130 963328 43135 963384
rect 42425 963326 43135 963328
rect 42425 963323 42491 963326
rect 43069 963323 43135 963326
rect 675477 963388 675543 963389
rect 675477 963384 675524 963388
rect 675588 963386 675594 963388
rect 675477 963328 675482 963384
rect 675477 963324 675524 963328
rect 675588 963326 675634 963386
rect 675588 963324 675594 963326
rect 675477 963323 675543 963324
rect 42425 963114 42491 963117
rect 44265 963114 44331 963117
rect 42425 963112 44331 963114
rect 42425 963056 42430 963112
rect 42486 963056 44270 963112
rect 44326 963056 44331 963112
rect 42425 963054 44331 963056
rect 42425 963051 42491 963054
rect 44265 963051 44331 963054
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 674281 962842 674347 962845
rect 675477 962842 675543 962845
rect 674281 962840 675543 962842
rect 674281 962784 674286 962840
rect 674342 962784 675482 962840
rect 675538 962784 675543 962840
rect 674281 962782 675543 962784
rect 674281 962779 674347 962782
rect 675477 962779 675543 962782
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 673177 960802 673243 960805
rect 675109 960802 675175 960805
rect 673177 960800 675175 960802
rect 673177 960744 673182 960800
rect 673238 960744 675114 960800
rect 675170 960744 675175 960800
rect 673177 960742 675175 960744
rect 673177 960739 673243 960742
rect 675109 960739 675175 960742
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 674925 959170 674991 959173
rect 675518 959170 675524 959172
rect 674925 959168 675524 959170
rect 674925 959112 674930 959168
rect 674986 959112 675524 959168
rect 674925 959110 675524 959112
rect 674925 959107 674991 959110
rect 675518 959108 675524 959110
rect 675588 959108 675594 959172
rect 42425 958762 42491 958765
rect 44449 958762 44515 958765
rect 42425 958760 44515 958762
rect 42425 958704 42430 958760
rect 42486 958704 44454 958760
rect 44510 958704 44515 958760
rect 42425 958702 44515 958704
rect 42425 958699 42491 958702
rect 44449 958699 44515 958702
rect 674649 958762 674715 958765
rect 675201 958762 675267 958765
rect 674649 958760 675267 958762
rect 674649 958704 674654 958760
rect 674710 958704 675206 958760
rect 675262 958704 675267 958760
rect 674649 958702 675267 958704
rect 674649 958699 674715 958702
rect 675201 958699 675267 958702
rect 41781 957812 41847 957813
rect 41781 957808 41828 957812
rect 41892 957810 41898 957812
rect 661677 957810 661743 957813
rect 675293 957810 675359 957813
rect 41781 957752 41786 957808
rect 41781 957748 41828 957752
rect 41892 957750 41938 957810
rect 661677 957808 675359 957810
rect 661677 957752 661682 957808
rect 661738 957752 675298 957808
rect 675354 957752 675359 957808
rect 661677 957750 675359 957752
rect 41892 957748 41898 957750
rect 41781 957747 41847 957748
rect 661677 957747 661743 957750
rect 675293 957747 675359 957750
rect 675753 957810 675819 957813
rect 676622 957810 676628 957812
rect 675753 957808 676628 957810
rect 675753 957752 675758 957808
rect 675814 957752 676628 957808
rect 675753 957750 676628 957752
rect 675753 957747 675819 957750
rect 676622 957748 676628 957750
rect 676692 957748 676698 957812
rect 674097 957130 674163 957133
rect 675477 957130 675543 957133
rect 674097 957128 675543 957130
rect 674097 957072 674102 957128
rect 674158 957072 675482 957128
rect 675538 957072 675543 957128
rect 674097 957070 675543 957072
rect 674097 957067 674163 957070
rect 675477 957067 675543 957070
rect 675753 956450 675819 956453
rect 676990 956450 676996 956452
rect 675753 956448 676996 956450
rect 675753 956392 675758 956448
rect 675814 956392 676996 956448
rect 675753 956390 676996 956392
rect 675753 956387 675819 956390
rect 676990 956388 676996 956390
rect 677060 956388 677066 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 41781 954680 41847 954685
rect 41781 954624 41786 954680
rect 41842 954624 41847 954680
rect 41781 954619 41847 954624
rect 675201 954682 675267 954685
rect 675702 954682 675708 954684
rect 675201 954680 675708 954682
rect 675201 954624 675206 954680
rect 675262 954624 675708 954680
rect 675201 954622 675708 954624
rect 675201 954619 675267 954622
rect 675702 954620 675708 954622
rect 675772 954620 675778 954684
rect 41784 954413 41844 954619
rect 41781 954408 41847 954413
rect 41781 954352 41786 954408
rect 41842 954352 41847 954408
rect 41781 954347 41847 954352
rect 674833 953458 674899 953461
rect 675477 953458 675543 953461
rect 674833 953456 675543 953458
rect 674833 953400 674838 953456
rect 674894 953400 675482 953456
rect 675538 953400 675543 953456
rect 674833 953398 675543 953400
rect 674833 953395 674899 953398
rect 675477 953395 675543 953398
rect 35157 952914 35223 952917
rect 41822 952914 41828 952916
rect 35157 952912 41828 952914
rect 35157 952856 35162 952912
rect 35218 952856 41828 952912
rect 35157 952854 41828 952856
rect 35157 952851 35223 952854
rect 41822 952852 41828 952854
rect 41892 952852 41898 952916
rect 37917 952506 37983 952509
rect 41454 952506 41460 952508
rect 37917 952504 41460 952506
rect 37917 952448 37922 952504
rect 37978 952448 41460 952504
rect 37917 952446 41460 952448
rect 37917 952443 37983 952446
rect 41454 952444 41460 952446
rect 41524 952444 41530 952508
rect 39297 952234 39363 952237
rect 41638 952234 41644 952236
rect 39297 952232 41644 952234
rect 39297 952176 39302 952232
rect 39358 952176 41644 952232
rect 39297 952174 41644 952176
rect 39297 952171 39363 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 672993 952234 673059 952237
rect 675569 952234 675635 952237
rect 672993 952232 675635 952234
rect 672993 952176 672998 952232
rect 673054 952176 675574 952232
rect 675630 952176 675635 952232
rect 672993 952174 675635 952176
rect 672993 952171 673059 952174
rect 675569 952171 675635 952174
rect 40033 951690 40099 951693
rect 41270 951690 41276 951692
rect 40033 951688 41276 951690
rect 40033 951632 40038 951688
rect 40094 951632 41276 951688
rect 40033 951630 41276 951632
rect 40033 951627 40099 951630
rect 41270 951628 41276 951630
rect 41340 951628 41346 951692
rect 676806 950676 676812 950740
rect 676876 950738 676882 950740
rect 683297 950738 683363 950741
rect 676876 950736 683363 950738
rect 676876 950680 683302 950736
rect 683358 950680 683363 950736
rect 676876 950678 683363 950680
rect 676876 950676 676882 950678
rect 683297 950675 683363 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 676070 949452 676076 949516
rect 676140 949514 676146 949516
rect 679617 949514 679683 949517
rect 676140 949512 679683 949514
rect 676140 949456 679622 949512
rect 679678 949456 679683 949512
rect 676140 949454 679683 949456
rect 676140 949452 676146 949454
rect 679617 949451 679683 949454
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 672717 947338 672783 947341
rect 683113 947338 683179 947341
rect 672717 947336 683179 947338
rect 672717 947280 672722 947336
rect 672778 947280 683118 947336
rect 683174 947280 683179 947336
rect 672717 947278 683179 947280
rect 672717 947275 672783 947278
rect 683113 947275 683179 947278
rect 31753 946658 31819 946661
rect 46197 946658 46263 946661
rect 31753 946656 46263 946658
rect 31753 946600 31758 946656
rect 31814 946600 46202 946656
rect 46258 946600 46263 946656
rect 31753 946598 46263 946600
rect 31753 946595 31819 946598
rect 46197 946595 46263 946598
rect 39757 943804 39823 943805
rect 39757 943800 39804 943804
rect 39868 943802 39874 943804
rect 39757 943744 39762 943800
rect 39757 943740 39804 943744
rect 39868 943742 39914 943802
rect 39868 943740 39874 943742
rect 40718 943740 40724 943804
rect 40788 943802 40794 943804
rect 42006 943802 42012 943804
rect 40788 943742 42012 943802
rect 40788 943740 40794 943742
rect 42006 943740 42012 943742
rect 42076 943740 42082 943804
rect 39757 943739 39823 943740
rect 45553 943530 45619 943533
rect 41492 943528 45619 943530
rect 41492 943472 45558 943528
rect 45614 943472 45619 943528
rect 41492 943470 45619 943472
rect 45553 943467 45619 943470
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 28717 942714 28783 942717
rect 28717 942712 28796 942714
rect 28717 942656 28722 942712
rect 28778 942656 28796 942712
rect 28717 942654 28796 942656
rect 28717 942651 28783 942654
rect 51717 942306 51783 942309
rect 41492 942304 51783 942306
rect 41492 942248 51722 942304
rect 51778 942248 51783 942304
rect 41492 942246 51783 942248
rect 51717 942243 51783 942246
rect 35801 941898 35867 941901
rect 35788 941896 35867 941898
rect 35788 941840 35806 941896
rect 35862 941840 35867 941896
rect 35788 941838 35867 941840
rect 35801 941835 35867 941838
rect 663057 941762 663123 941765
rect 676213 941762 676279 941765
rect 663057 941760 676279 941762
rect 663057 941704 663062 941760
rect 663118 941704 676218 941760
rect 676274 941704 676279 941760
rect 663057 941702 676279 941704
rect 663057 941699 663123 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 44633 941082 44699 941085
rect 41492 941080 44699 941082
rect 41492 941024 44638 941080
rect 44694 941024 44699 941080
rect 41492 941022 44699 941024
rect 44633 941019 44699 941022
rect 42057 940674 42123 940677
rect 41492 940672 42123 940674
rect 41492 940616 42062 940672
rect 42118 940616 42123 940672
rect 41492 940614 42123 940616
rect 42057 940611 42123 940614
rect 35801 940266 35867 940269
rect 35788 940264 35867 940266
rect 35788 940208 35806 940264
rect 35862 940208 35867 940264
rect 35788 940206 35867 940208
rect 35801 940203 35867 940206
rect 48957 940130 49023 940133
rect 41830 940128 49023 940130
rect 41830 940072 48962 940128
rect 49018 940072 49023 940128
rect 41830 940070 49023 940072
rect 41830 939858 41890 940070
rect 48957 940067 49023 940070
rect 41492 939798 41890 939858
rect 42057 939858 42123 939861
rect 50337 939858 50403 939861
rect 42057 939856 50403 939858
rect 42057 939800 42062 939856
rect 42118 939800 50342 939856
rect 50398 939800 50403 939856
rect 42057 939798 50403 939800
rect 42057 939795 42123 939798
rect 50337 939795 50403 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683113 939722 683179 939725
rect 683070 939720 683179 939722
rect 683070 939664 683118 939720
rect 683174 939664 683179 939720
rect 683070 939659 683179 939664
rect 683070 939556 683130 939659
rect 41776 939450 41782 939452
rect 41492 939390 41782 939450
rect 41776 939388 41782 939390
rect 41846 939388 41852 939452
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 36537 939042 36603 939045
rect 36524 939040 36603 939042
rect 36524 938984 36542 939040
rect 36598 938984 36603 939040
rect 36524 938982 36603 938984
rect 36537 938979 36603 938982
rect 37917 938634 37983 938637
rect 37917 938632 37996 938634
rect 37917 938576 37922 938632
rect 37978 938576 37996 938632
rect 37917 938574 37996 938576
rect 37917 938571 37983 938574
rect 669957 938498 670023 938501
rect 676262 938498 676322 938740
rect 669957 938496 676322 938498
rect 669957 938440 669962 938496
rect 670018 938440 676322 938496
rect 669957 938438 676322 938440
rect 669957 938435 670023 938438
rect 33777 938226 33843 938229
rect 33764 938224 33843 938226
rect 33764 938168 33782 938224
rect 33838 938168 33843 938224
rect 33764 938166 33843 938168
rect 33777 938163 33843 938166
rect 671797 938090 671863 938093
rect 674598 938090 674604 938092
rect 671797 938088 674604 938090
rect 671797 938032 671802 938088
rect 671858 938032 674604 938088
rect 671797 938030 674604 938032
rect 671797 938027 671863 938030
rect 674598 938028 674604 938030
rect 674668 938028 674674 938092
rect 676262 938090 676322 938332
rect 674790 938030 676322 938090
rect 35157 937818 35223 937821
rect 671613 937818 671679 937821
rect 674790 937818 674850 938030
rect 35157 937816 35236 937818
rect 35157 937760 35162 937816
rect 35218 937760 35236 937816
rect 35157 937758 35236 937760
rect 671613 937816 674850 937818
rect 671613 937760 671618 937816
rect 671674 937760 674850 937816
rect 671613 937758 674850 937760
rect 35157 937755 35223 937758
rect 671613 937755 671679 937758
rect 676446 937685 676506 937924
rect 674966 937620 674972 937684
rect 675036 937682 675042 937684
rect 675036 937622 676322 937682
rect 676446 937680 676555 937685
rect 676446 937624 676494 937680
rect 676550 937624 676555 937680
rect 676446 937622 676555 937624
rect 675036 937620 675042 937622
rect 668577 937546 668643 937549
rect 668577 937544 674850 937546
rect 668577 937488 668582 937544
rect 668638 937488 674850 937544
rect 676262 937516 676322 937622
rect 676489 937619 676555 937622
rect 668577 937486 674850 937488
rect 668577 937483 668643 937486
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 660297 937274 660363 937277
rect 674790 937274 674850 937486
rect 660297 937272 674666 937274
rect 660297 937216 660302 937272
rect 660358 937216 674666 937272
rect 660297 937214 674666 937216
rect 674790 937214 676322 937274
rect 660297 937211 660363 937214
rect 42793 937002 42859 937005
rect 41492 937000 42859 937002
rect 41492 936944 42798 937000
rect 42854 936944 42859 937000
rect 41492 936942 42859 936944
rect 42793 936939 42859 936942
rect 674606 936866 674666 937214
rect 676262 937108 676322 937214
rect 676489 936866 676555 936869
rect 674606 936864 676555 936866
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 44449 936322 44515 936325
rect 41830 936320 44515 936322
rect 41830 936264 44454 936320
rect 44510 936264 44515 936320
rect 41830 936262 44515 936264
rect 41830 936186 41890 936262
rect 44449 936259 44515 936262
rect 41492 936126 41890 936186
rect 39757 935778 39823 935781
rect 64462 935778 64522 936836
rect 674606 936808 676494 936864
rect 676550 936808 676555 936864
rect 674606 936806 676555 936808
rect 676489 936803 676555 936806
rect 672441 936458 672507 936461
rect 676262 936458 676322 936700
rect 672441 936456 676322 936458
rect 672441 936400 672446 936456
rect 672502 936400 676322 936456
rect 672441 936398 676322 936400
rect 672441 936395 672507 936398
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 39757 935776 39836 935778
rect 39757 935720 39762 935776
rect 39818 935720 39836 935776
rect 39757 935718 39836 935720
rect 48270 935718 64522 935778
rect 672625 935778 672691 935781
rect 676262 935778 676322 935884
rect 672625 935776 676322 935778
rect 672625 935720 672630 935776
rect 672686 935720 676322 935776
rect 672625 935718 676322 935720
rect 39757 935715 39823 935718
rect 41781 935642 41847 935645
rect 48270 935642 48330 935718
rect 672625 935715 672691 935718
rect 679617 935642 679683 935645
rect 41781 935640 48330 935642
rect 41781 935584 41786 935640
rect 41842 935584 48330 935640
rect 41781 935582 48330 935584
rect 679574 935640 679683 935642
rect 679574 935584 679622 935640
rect 679678 935584 679683 935640
rect 41781 935579 41847 935582
rect 679574 935579 679683 935584
rect 679574 935476 679634 935579
rect 43437 935370 43503 935373
rect 41492 935368 43503 935370
rect 41492 935312 43442 935368
rect 43498 935312 43503 935368
rect 41492 935310 43503 935312
rect 43437 935307 43503 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43069 934962 43135 934965
rect 41492 934960 43135 934962
rect 41492 934904 43074 934960
rect 43130 934904 43135 934960
rect 41492 934902 43135 934904
rect 43069 934899 43135 934902
rect 675293 934690 675359 934693
rect 675293 934688 676292 934690
rect 675293 934632 675298 934688
rect 675354 934632 676292 934688
rect 675293 934630 676292 934632
rect 675293 934627 675359 934630
rect 40033 934554 40099 934557
rect 40020 934552 40099 934554
rect 40020 934496 40038 934552
rect 40094 934496 40099 934552
rect 40020 934494 40099 934496
rect 40033 934491 40099 934494
rect 44265 934146 44331 934149
rect 41492 934144 44331 934146
rect 41492 934088 44270 934144
rect 44326 934088 44331 934144
rect 41492 934086 44331 934088
rect 44265 934083 44331 934086
rect 675109 934146 675175 934149
rect 676262 934146 676322 934252
rect 675109 934144 676322 934146
rect 675109 934088 675114 934144
rect 675170 934088 676322 934144
rect 675109 934086 676322 934088
rect 675109 934083 675175 934086
rect 674465 933874 674531 933877
rect 674465 933872 676292 933874
rect 674465 933816 674470 933872
rect 674526 933816 676292 933872
rect 674465 933814 676292 933816
rect 674465 933811 674531 933814
rect 43253 933738 43319 933741
rect 41492 933736 43319 933738
rect 41492 933680 43258 933736
rect 43314 933680 43319 933736
rect 41492 933678 43319 933680
rect 43253 933675 43319 933678
rect 43621 933330 43687 933333
rect 41492 933328 43687 933330
rect 41492 933272 43626 933328
rect 43682 933272 43687 933328
rect 41492 933270 43687 933272
rect 43621 933267 43687 933270
rect 673085 933194 673151 933197
rect 676262 933194 676322 933436
rect 673085 933192 676322 933194
rect 673085 933136 673090 933192
rect 673146 933136 676322 933192
rect 673085 933134 676322 933136
rect 673085 933131 673151 933134
rect 42333 932922 42399 932925
rect 41492 932920 42399 932922
rect 41492 932864 42338 932920
rect 42394 932864 42399 932920
rect 41492 932862 42399 932864
rect 42333 932859 42399 932862
rect 673361 932922 673427 932925
rect 676262 932922 676322 933028
rect 673361 932920 676322 932922
rect 673361 932864 673366 932920
rect 673422 932864 676322 932920
rect 673361 932862 676322 932864
rect 673361 932859 673427 932862
rect 674281 932650 674347 932653
rect 674281 932648 676292 932650
rect 674281 932592 674286 932648
rect 674342 932592 676292 932648
rect 674281 932590 676292 932592
rect 674281 932587 674347 932590
rect 683297 932378 683363 932381
rect 683254 932376 683363 932378
rect 683254 932320 683302 932376
rect 683358 932320 683363 932376
rect 683254 932315 683363 932320
rect 683254 932212 683314 932315
rect 43805 932106 43871 932109
rect 41492 932104 43871 932106
rect 41492 932048 43810 932104
rect 43866 932048 43871 932104
rect 41492 932046 43871 932048
rect 43805 932043 43871 932046
rect 676990 931908 676996 931972
rect 677060 931908 677066 931972
rect 676998 931804 677058 931908
rect 676622 931500 676628 931564
rect 676692 931500 676698 931564
rect 676630 931396 676690 931500
rect 673177 930746 673243 930749
rect 676262 930746 676322 930988
rect 673177 930744 676322 930746
rect 673177 930688 673182 930744
rect 673238 930688 676322 930744
rect 673177 930686 676322 930688
rect 673177 930683 673243 930686
rect 674649 930474 674715 930477
rect 676262 930474 676322 930580
rect 674649 930472 676322 930474
rect 674649 930416 674654 930472
rect 674710 930416 676322 930472
rect 674649 930414 676322 930416
rect 674649 930411 674715 930414
rect 674097 930202 674163 930205
rect 674097 930200 676292 930202
rect 674097 930144 674102 930200
rect 674158 930144 676292 930200
rect 674097 930142 676292 930144
rect 674097 930139 674163 930142
rect 670693 929522 670759 929525
rect 676262 929522 676322 929764
rect 670693 929520 676322 929522
rect 670693 929464 670698 929520
rect 670754 929464 676322 929520
rect 670693 929462 676322 929464
rect 670693 929459 670759 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 673361 928298 673427 928301
rect 676262 928298 676322 928540
rect 673361 928296 676322 928298
rect 673361 928240 673366 928296
rect 673422 928240 676322 928296
rect 673361 928238 676322 928240
rect 673361 928235 673427 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 41597 911978 41663 911981
rect 42006 911978 42012 911980
rect 41597 911976 42012 911978
rect 41597 911920 41602 911976
rect 41658 911920 42012 911976
rect 41597 911918 42012 911920
rect 41597 911915 41663 911918
rect 42006 911916 42012 911918
rect 42076 911916 42082 911980
rect 41413 911706 41479 911709
rect 42190 911706 42196 911708
rect 41413 911704 42196 911706
rect 41413 911648 41418 911704
rect 41474 911648 42196 911704
rect 41413 911646 42196 911648
rect 41413 911643 41479 911646
rect 42190 911644 42196 911646
rect 42260 911644 42266 911708
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 44081 892802 44147 892805
rect 55857 892802 55923 892805
rect 44081 892800 55923 892802
rect 44081 892744 44086 892800
rect 44142 892744 55862 892800
rect 55918 892744 55923 892800
rect 44081 892742 55923 892744
rect 44081 892739 44147 892742
rect 55857 892739 55923 892742
rect 42931 892530 42997 892533
rect 54477 892530 54543 892533
rect 42931 892528 54543 892530
rect 42931 892472 42936 892528
rect 42992 892472 54482 892528
rect 54538 892472 54543 892528
rect 42931 892470 54543 892472
rect 42931 892467 42997 892470
rect 54477 892467 54543 892470
rect 43069 892258 43135 892261
rect 53281 892258 53347 892261
rect 43069 892256 53347 892258
rect 43069 892200 43074 892256
rect 43130 892200 53286 892256
rect 53342 892200 53347 892256
rect 43069 892198 53347 892200
rect 43069 892195 43135 892198
rect 53281 892195 53347 892198
rect 44081 891986 44147 891989
rect 47577 891986 47643 891989
rect 44081 891984 47643 891986
rect 44081 891928 44086 891984
rect 44142 891928 47582 891984
rect 47638 891928 47643 891984
rect 44081 891926 47643 891928
rect 44081 891923 44147 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 669221 879202 669287 879205
rect 675017 879202 675083 879205
rect 669221 879200 675083 879202
rect 669221 879144 669226 879200
rect 669282 879144 675022 879200
rect 675078 879144 675083 879200
rect 669221 879142 675083 879144
rect 669221 879139 669287 879142
rect 675017 879139 675083 879142
rect 668761 877706 668827 877709
rect 675477 877706 675543 877709
rect 668761 877704 675543 877706
rect 668761 877648 668766 877704
rect 668822 877648 675482 877704
rect 675538 877648 675543 877704
rect 668761 877646 675543 877648
rect 668761 877643 668827 877646
rect 675477 877643 675543 877646
rect 675017 877298 675083 877301
rect 675385 877298 675451 877301
rect 675017 877296 675451 877298
rect 675017 877240 675022 877296
rect 675078 877240 675390 877296
rect 675446 877240 675451 877296
rect 675017 877238 675451 877240
rect 675017 877235 675083 877238
rect 675385 877235 675451 877238
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 670509 874034 670575 874037
rect 675477 874034 675543 874037
rect 670509 874032 675543 874034
rect 670509 873976 670514 874032
rect 670570 873976 675482 874032
rect 675538 873976 675543 874032
rect 670509 873974 675543 873976
rect 670509 873971 670575 873974
rect 675477 873971 675543 873974
rect 675661 874034 675727 874037
rect 675886 874034 675892 874036
rect 675661 874032 675892 874034
rect 675661 873976 675666 874032
rect 675722 873976 675892 874032
rect 675661 873974 675892 873976
rect 675661 873971 675727 873974
rect 675886 873972 675892 873974
rect 675956 873972 675962 874036
rect 669589 872266 669655 872269
rect 675109 872266 675175 872269
rect 675569 872266 675635 872269
rect 669589 872264 675175 872266
rect 669589 872208 669594 872264
rect 669650 872208 675114 872264
rect 675170 872208 675175 872264
rect 669589 872206 675175 872208
rect 669589 872203 669655 872206
rect 675109 872203 675175 872206
rect 675526 872264 675635 872266
rect 675526 872208 675574 872264
rect 675630 872208 675635 872264
rect 675526 872203 675635 872208
rect 675526 871994 675586 872203
rect 676806 871994 676812 871996
rect 675526 871934 676812 871994
rect 676806 871932 676812 871934
rect 676876 871932 676882 871996
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 673862 869484 673868 869548
rect 673932 869546 673938 869548
rect 675109 869546 675175 869549
rect 673932 869544 675175 869546
rect 673932 869488 675114 869544
rect 675170 869488 675175 869544
rect 673932 869486 675175 869488
rect 673932 869484 673938 869486
rect 675109 869483 675175 869486
rect 664437 868730 664503 868733
rect 675293 868730 675359 868733
rect 664437 868728 675359 868730
rect 664437 868672 664442 868728
rect 664498 868672 675298 868728
rect 675354 868672 675359 868728
rect 664437 868670 675359 868672
rect 664437 868667 664503 868670
rect 675293 868667 675359 868670
rect 673085 868458 673151 868461
rect 675477 868458 675543 868461
rect 673085 868456 675543 868458
rect 673085 868400 673090 868456
rect 673146 868400 675482 868456
rect 675538 868400 675543 868456
rect 673085 868398 675543 868400
rect 673085 868395 673151 868398
rect 675477 868395 675543 868398
rect 674005 868050 674071 868053
rect 675109 868050 675175 868053
rect 674005 868048 675175 868050
rect 674005 867992 674010 868048
rect 674066 867992 675114 868048
rect 675170 867992 675175 868048
rect 674005 867990 675175 867992
rect 674005 867987 674071 867990
rect 675109 867987 675175 867990
rect 671153 867234 671219 867237
rect 675477 867234 675543 867237
rect 671153 867232 675543 867234
rect 671153 867176 671158 867232
rect 671214 867176 675482 867232
rect 675538 867176 675543 867232
rect 671153 867174 675543 867176
rect 671153 867171 671219 867174
rect 675477 867171 675543 867174
rect 667841 866690 667907 866693
rect 674925 866690 674991 866693
rect 667841 866688 674991 866690
rect 667841 866632 667846 866688
rect 667902 866632 674930 866688
rect 674986 866632 674991 866688
rect 667841 866630 674991 866632
rect 667841 866627 667907 866630
rect 674925 866627 674991 866630
rect 674649 864786 674715 864789
rect 675201 864786 675267 864789
rect 674649 864784 675267 864786
rect 674649 864728 674654 864784
rect 674710 864728 675206 864784
rect 675262 864728 675267 864784
rect 674649 864726 675267 864728
rect 674649 864723 674715 864726
rect 675201 864723 675267 864726
rect 62757 858666 62823 858669
rect 62757 858664 64492 858666
rect 62757 858608 62762 858664
rect 62818 858608 64492 858664
rect 62757 858606 64492 858608
rect 62757 858603 62823 858606
rect 652385 856354 652451 856357
rect 650164 856352 652451 856354
rect 650164 856296 652390 856352
rect 652446 856296 652451 856352
rect 650164 856294 652451 856296
rect 652385 856291 652451 856294
rect 674465 854316 674531 854317
rect 674414 854314 674420 854316
rect 674374 854254 674420 854314
rect 674484 854312 674531 854316
rect 674526 854256 674531 854312
rect 674414 854252 674420 854254
rect 674484 854252 674531 854256
rect 674465 854251 674531 854252
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651833 843026 651899 843029
rect 650164 843024 651899 843026
rect 650164 842968 651838 843024
rect 651894 842968 651899 843024
rect 650164 842966 651899 842968
rect 651833 842963 651899 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 35801 816506 35867 816509
rect 651465 816506 651531 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 35801 816443 35867 816446
rect 651465 816443 651531 816446
rect 44449 816098 44515 816101
rect 41492 816096 44515 816098
rect 41492 816040 44454 816096
rect 44510 816040 44515 816096
rect 41492 816038 44515 816040
rect 44449 816035 44515 816038
rect 44633 815690 44699 815693
rect 41492 815688 44699 815690
rect 41492 815632 44638 815688
rect 44694 815632 44699 815688
rect 41492 815630 44699 815632
rect 44633 815627 44699 815630
rect 45001 815282 45067 815285
rect 41492 815280 45067 815282
rect 41492 815224 45006 815280
rect 45062 815224 45067 815280
rect 41492 815222 45067 815224
rect 45001 815219 45067 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 44633 814466 44699 814469
rect 41492 814464 44699 814466
rect 41492 814408 44638 814464
rect 44694 814408 44699 814464
rect 41492 814406 44699 814408
rect 44633 814403 44699 814406
rect 39982 814234 39988 814298
rect 40052 814234 40058 814298
rect 39990 814028 40050 814234
rect 44817 813650 44883 813653
rect 41492 813648 44883 813650
rect 41492 813592 44822 813648
rect 44878 813592 44883 813648
rect 41492 813590 44883 813592
rect 44817 813587 44883 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 41321 812834 41387 812837
rect 41308 812832 41387 812834
rect 41308 812776 41326 812832
rect 41382 812776 41387 812832
rect 41308 812774 41387 812776
rect 41321 812771 41387 812774
rect 40953 812426 41019 812429
rect 40940 812424 41019 812426
rect 40940 812368 40958 812424
rect 41014 812368 41019 812424
rect 40940 812366 41019 812368
rect 40953 812363 41019 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 35157 811610 35223 811613
rect 35157 811608 35236 811610
rect 35157 811552 35162 811608
rect 35218 811552 35236 811608
rect 35157 811550 35236 811552
rect 35157 811547 35223 811550
rect 35893 811202 35959 811205
rect 35893 811200 35972 811202
rect 35893 811144 35898 811200
rect 35954 811144 35972 811200
rect 35893 811142 35972 811144
rect 35893 811139 35959 811142
rect 43069 810794 43135 810797
rect 41492 810792 43135 810794
rect 41492 810736 43074 810792
rect 43130 810736 43135 810792
rect 41492 810734 43135 810736
rect 43069 810731 43135 810734
rect 44265 810386 44331 810389
rect 41492 810384 44331 810386
rect 41492 810328 44270 810384
rect 44326 810328 44331 810384
rect 41492 810326 44331 810328
rect 44265 810323 44331 810326
rect 42793 809978 42859 809981
rect 41492 809976 42859 809978
rect 41492 809920 42798 809976
rect 42854 809920 42859 809976
rect 41492 809918 42859 809920
rect 42793 809915 42859 809918
rect 43437 809570 43503 809573
rect 41492 809568 43503 809570
rect 41492 809512 43442 809568
rect 43498 809512 43503 809568
rect 41492 809510 43503 809512
rect 43437 809507 43503 809510
rect 41965 809162 42031 809165
rect 41492 809160 42031 809162
rect 41492 809104 41970 809160
rect 42026 809104 42031 809160
rect 41492 809102 42031 809104
rect 41965 809099 42031 809102
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 40769 808346 40835 808349
rect 40756 808344 40835 808346
rect 40756 808288 40774 808344
rect 40830 808288 40835 808344
rect 40756 808286 40835 808288
rect 40769 808283 40835 808286
rect 45185 807938 45251 807941
rect 41492 807936 45251 807938
rect 41492 807880 45190 807936
rect 45246 807880 45251 807936
rect 41492 807878 45251 807880
rect 45185 807875 45251 807878
rect 43253 807530 43319 807533
rect 41308 807528 43319 807530
rect 41308 807472 43258 807528
rect 43314 807472 43319 807528
rect 41308 807470 43319 807472
rect 43253 807467 43319 807470
rect 41462 806714 41522 807092
rect 42149 806714 42215 806717
rect 41462 806712 42215 806714
rect 41462 806684 42154 806712
rect 41492 806656 42154 806684
rect 42210 806656 42215 806712
rect 41492 806654 42215 806656
rect 42149 806651 42215 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43989 806306 44055 806309
rect 41492 806304 44055 806306
rect 41492 806248 43994 806304
rect 44050 806248 44055 806304
rect 41492 806246 44055 806248
rect 43989 806243 44055 806246
rect 40902 805428 40908 805492
rect 40972 805490 40978 805492
rect 41965 805490 42031 805493
rect 40972 805488 42031 805490
rect 40972 805432 41970 805488
rect 42026 805432 42031 805488
rect 40972 805430 42031 805432
rect 40972 805428 40978 805430
rect 41965 805427 42031 805430
rect 40585 805356 40651 805357
rect 40534 805354 40540 805356
rect 40494 805294 40540 805354
rect 40604 805352 40651 805356
rect 40646 805296 40651 805352
rect 40534 805292 40540 805294
rect 40604 805292 40651 805296
rect 40585 805291 40651 805292
rect 40769 805084 40835 805085
rect 40718 805082 40724 805084
rect 40678 805022 40724 805082
rect 40788 805080 40835 805084
rect 40830 805024 40835 805080
rect 40718 805020 40724 805022
rect 40788 805020 40835 805024
rect 40769 805019 40835 805020
rect 41137 804810 41203 804813
rect 42006 804810 42012 804812
rect 41137 804808 42012 804810
rect 41137 804752 41142 804808
rect 41198 804752 42012 804808
rect 41137 804750 42012 804752
rect 41137 804747 41203 804750
rect 42006 804748 42012 804750
rect 42076 804748 42082 804812
rect 40953 804538 41019 804541
rect 41638 804538 41644 804540
rect 40953 804536 41644 804538
rect 40953 804480 40958 804536
rect 41014 804480 41644 804536
rect 40953 804478 41644 804480
rect 40953 804475 41019 804478
rect 41638 804476 41644 804478
rect 41708 804476 41714 804540
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41689 802498 41755 802501
rect 42517 802498 42583 802501
rect 41689 802496 42583 802498
rect 41689 802440 41694 802496
rect 41750 802440 42522 802496
rect 42578 802440 42583 802496
rect 41689 802438 42583 802440
rect 41689 802435 41755 802438
rect 42517 802435 42583 802438
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 53097 799370 53163 799373
rect 51030 799368 53163 799370
rect 51030 799312 53102 799368
rect 53158 799312 53163 799368
rect 51030 799310 53163 799312
rect 42517 799234 42583 799237
rect 51030 799234 51090 799310
rect 53097 799307 53163 799310
rect 42517 799232 51090 799234
rect 42517 799176 42522 799232
rect 42578 799176 51090 799232
rect 42517 799174 51090 799176
rect 42517 799171 42583 799174
rect 42425 796786 42491 796789
rect 45185 796786 45251 796789
rect 42425 796784 45251 796786
rect 42425 796728 42430 796784
rect 42486 796728 45190 796784
rect 45246 796728 45251 796784
rect 42425 796726 45251 796728
rect 42425 796723 42491 796726
rect 45185 796723 45251 796726
rect 42149 796242 42215 796245
rect 43437 796242 43503 796245
rect 42149 796240 43503 796242
rect 42149 796184 42154 796240
rect 42210 796184 43442 796240
rect 43498 796184 43503 796240
rect 42149 796182 43503 796184
rect 42149 796179 42215 796182
rect 43437 796179 43503 796182
rect 40718 794956 40724 795020
rect 40788 795018 40794 795020
rect 40788 794958 42442 795018
rect 40788 794956 40794 794958
rect 42382 794341 42442 794958
rect 42382 794336 42491 794341
rect 42382 794280 42430 794336
rect 42486 794280 42491 794336
rect 42382 794278 42491 794280
rect 42425 794275 42491 794278
rect 40902 794140 40908 794204
rect 40972 794202 40978 794204
rect 41781 794202 41847 794205
rect 40972 794200 41847 794202
rect 40972 794144 41786 794200
rect 41842 794144 41847 794200
rect 40972 794142 41847 794144
rect 40972 794140 40978 794142
rect 41781 794139 41847 794142
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 42885 790802 42951 790805
rect 44265 790802 44331 790805
rect 42885 790800 44331 790802
rect 42885 790744 42890 790800
rect 42946 790744 44270 790800
rect 44326 790744 44331 790800
rect 42885 790742 44331 790744
rect 42885 790739 42951 790742
rect 44265 790739 44331 790742
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 669773 789442 669839 789445
rect 675201 789442 675267 789445
rect 669773 789440 675267 789442
rect 669773 789384 669778 789440
rect 669834 789384 675206 789440
rect 675262 789384 675267 789440
rect 669773 789382 675267 789384
rect 669773 789379 669839 789382
rect 675201 789379 675267 789382
rect 41638 788972 41644 789036
rect 41708 789034 41714 789036
rect 41708 788974 42074 789034
rect 41708 788972 41714 788974
rect 42014 788762 42074 788974
rect 42517 788762 42583 788765
rect 42014 788760 42583 788762
rect 42014 788704 42522 788760
rect 42578 788704 42583 788760
rect 42014 788702 42583 788704
rect 42517 788699 42583 788702
rect 41781 788628 41847 788629
rect 41781 788624 41828 788628
rect 41892 788626 41898 788628
rect 42701 788626 42767 788629
rect 62757 788626 62823 788629
rect 41781 788568 41786 788624
rect 41781 788564 41828 788568
rect 41892 788566 41938 788626
rect 42701 788624 62823 788626
rect 42701 788568 42706 788624
rect 42762 788568 62762 788624
rect 62818 788568 62823 788624
rect 42701 788566 62823 788568
rect 41892 788564 41898 788566
rect 41781 788563 41847 788564
rect 42701 788563 42767 788566
rect 62757 788563 62823 788566
rect 42425 788354 42491 788357
rect 43069 788354 43135 788357
rect 42425 788352 43135 788354
rect 42425 788296 42430 788352
rect 42486 788296 43074 788352
rect 43130 788296 43135 788352
rect 42425 788294 43135 788296
rect 42425 788291 42491 788294
rect 43069 788291 43135 788294
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 674465 788082 674531 788085
rect 675385 788082 675451 788085
rect 674465 788080 675451 788082
rect 674465 788024 674470 788080
rect 674526 788024 675390 788080
rect 675446 788024 675451 788080
rect 674465 788022 675451 788024
rect 674465 788019 674531 788022
rect 675385 788019 675451 788022
rect 674833 787268 674899 787269
rect 674782 787204 674788 787268
rect 674852 787266 674899 787268
rect 674852 787264 674944 787266
rect 674894 787208 674944 787264
rect 674852 787206 674944 787208
rect 674852 787204 674899 787206
rect 674833 787203 674899 787204
rect 674966 786660 674972 786724
rect 675036 786722 675042 786724
rect 675385 786722 675451 786725
rect 675036 786720 675451 786722
rect 675036 786664 675390 786720
rect 675446 786664 675451 786720
rect 675036 786662 675451 786664
rect 675036 786660 675042 786662
rect 675385 786659 675451 786662
rect 672625 784274 672691 784277
rect 675477 784274 675543 784277
rect 672625 784272 675543 784274
rect 672625 784216 672630 784272
rect 672686 784216 675482 784272
rect 675538 784216 675543 784272
rect 672625 784214 675543 784216
rect 672625 784211 672691 784214
rect 675477 784211 675543 784214
rect 668945 783866 669011 783869
rect 675477 783866 675543 783869
rect 668945 783864 675543 783866
rect 668945 783808 668950 783864
rect 669006 783808 675482 783864
rect 675538 783808 675543 783864
rect 668945 783806 675543 783808
rect 668945 783803 669011 783806
rect 675477 783803 675543 783806
rect 674925 783324 674991 783325
rect 674925 783322 674972 783324
rect 674880 783320 674972 783322
rect 674880 783264 674930 783320
rect 674880 783262 674972 783264
rect 674925 783260 674972 783262
rect 675036 783260 675042 783324
rect 674925 783259 674991 783260
rect 674281 783050 674347 783053
rect 675385 783050 675451 783053
rect 674281 783048 675451 783050
rect 674281 782992 674286 783048
rect 674342 782992 675390 783048
rect 675446 782992 675451 783048
rect 674281 782990 675451 782992
rect 674281 782987 674347 782990
rect 675385 782987 675451 782990
rect 674782 782716 674788 782780
rect 674852 782778 674858 782780
rect 675109 782778 675175 782781
rect 674852 782776 675175 782778
rect 674852 782720 675114 782776
rect 675170 782720 675175 782776
rect 674852 782718 675175 782720
rect 674852 782716 674858 782718
rect 675109 782715 675175 782718
rect 668209 782506 668275 782509
rect 675293 782506 675359 782509
rect 668209 782504 675359 782506
rect 668209 782448 668214 782504
rect 668270 782448 675298 782504
rect 675354 782448 675359 782504
rect 668209 782446 675359 782448
rect 668209 782443 668275 782446
rect 675293 782443 675359 782446
rect 675109 780738 675175 780741
rect 675109 780736 676230 780738
rect 675109 780680 675114 780736
rect 675170 780680 676230 780736
rect 675109 780678 676230 780680
rect 675109 780675 675175 780678
rect 676170 780602 676230 780678
rect 676990 780602 676996 780604
rect 676170 780542 676996 780602
rect 676990 780540 676996 780542
rect 677060 780540 677066 780604
rect 62757 780466 62823 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 62757 780403 62823 780406
rect 670325 780058 670391 780061
rect 675477 780058 675543 780061
rect 670325 780056 675543 780058
rect 670325 780000 670330 780056
rect 670386 780000 675482 780056
rect 675538 780000 675543 780056
rect 670325 779998 675543 780000
rect 670325 779995 670391 779998
rect 675477 779995 675543 779998
rect 673729 779242 673795 779245
rect 675293 779242 675359 779245
rect 673729 779240 675359 779242
rect 673729 779184 673734 779240
rect 673790 779184 675298 779240
rect 675354 779184 675359 779240
rect 673729 779182 675359 779184
rect 673729 779179 673795 779182
rect 675293 779179 675359 779182
rect 660297 778970 660363 778973
rect 670141 778970 670207 778973
rect 660297 778968 670207 778970
rect 660297 778912 660302 778968
rect 660358 778912 670146 778968
rect 670202 778912 670207 778968
rect 660297 778910 670207 778912
rect 660297 778907 660363 778910
rect 670141 778907 670207 778910
rect 674189 778698 674255 778701
rect 675477 778698 675543 778701
rect 674189 778696 675543 778698
rect 674189 778640 674194 778696
rect 674250 778640 675482 778696
rect 675538 778640 675543 778696
rect 674189 778638 675543 778640
rect 674189 778635 674255 778638
rect 675477 778635 675543 778638
rect 666461 778426 666527 778429
rect 670969 778426 671035 778429
rect 666461 778424 671035 778426
rect 666461 778368 666466 778424
rect 666522 778368 670974 778424
rect 671030 778368 671035 778424
rect 666461 778366 671035 778368
rect 666461 778363 666527 778366
rect 670969 778363 671035 778366
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 670141 777066 670207 777069
rect 675385 777066 675451 777069
rect 670141 777064 675451 777066
rect 670141 777008 670146 777064
rect 670202 777008 675390 777064
rect 675446 777008 675451 777064
rect 670141 777006 675451 777008
rect 670141 777003 670207 777006
rect 675385 777003 675451 777006
rect 652385 776658 652451 776661
rect 650164 776656 652451 776658
rect 650164 776600 652390 776656
rect 652446 776600 652451 776656
rect 650164 776598 652451 776600
rect 652385 776595 652451 776598
rect 670969 776522 671035 776525
rect 675477 776522 675543 776525
rect 670969 776520 675543 776522
rect 670969 776464 670974 776520
rect 671030 776464 675482 776520
rect 675538 776464 675543 776520
rect 670969 776462 675543 776464
rect 670969 776459 671035 776462
rect 675477 776459 675543 776462
rect 670141 775026 670207 775029
rect 675477 775026 675543 775029
rect 670141 775024 675543 775026
rect 670141 774968 670146 775024
rect 670202 774968 675482 775024
rect 675538 774968 675543 775024
rect 670141 774966 675543 774968
rect 670141 774963 670207 774966
rect 675477 774963 675543 774966
rect 41462 774346 41522 774452
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 41462 773938 41522 774044
rect 41462 773878 45570 773938
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 44449 773258 44515 773261
rect 41492 773256 44515 773258
rect 41492 773200 44454 773256
rect 44510 773200 44515 773256
rect 41492 773198 44515 773200
rect 44449 773195 44515 773198
rect 44449 772850 44515 772853
rect 41492 772848 44515 772850
rect 41492 772792 44454 772848
rect 44510 772792 44515 772848
rect 41492 772790 44515 772792
rect 45510 772850 45570 773878
rect 672901 773802 672967 773805
rect 675477 773802 675543 773805
rect 672901 773800 675543 773802
rect 672901 773744 672906 773800
rect 672962 773744 675482 773800
rect 675538 773744 675543 773800
rect 672901 773742 675543 773744
rect 672901 773739 672967 773742
rect 675477 773739 675543 773742
rect 55857 772850 55923 772853
rect 45510 772848 55923 772850
rect 45510 772792 55862 772848
rect 55918 772792 55923 772848
rect 45510 772790 55923 772792
rect 44449 772787 44515 772790
rect 55857 772787 55923 772790
rect 675886 772652 675892 772716
rect 675956 772714 675962 772716
rect 682377 772714 682443 772717
rect 675956 772712 682443 772714
rect 675956 772656 682382 772712
rect 682438 772656 682443 772712
rect 675956 772654 682443 772656
rect 675956 772652 675962 772654
rect 682377 772651 682443 772654
rect 45001 772442 45067 772445
rect 41492 772440 45067 772442
rect 41492 772384 45006 772440
rect 45062 772384 45067 772440
rect 41492 772382 45067 772384
rect 45001 772379 45067 772382
rect 44265 772034 44331 772037
rect 41492 772032 44331 772034
rect 41492 771976 44270 772032
rect 44326 771976 44331 772032
rect 41492 771974 44331 771976
rect 44265 771971 44331 771974
rect 674741 772034 674807 772037
rect 683205 772034 683271 772037
rect 674741 772032 683271 772034
rect 674741 771976 674746 772032
rect 674802 771976 683210 772032
rect 683266 771976 683271 772032
rect 674741 771974 683271 771976
rect 674741 771971 674807 771974
rect 683205 771971 683271 771974
rect 44633 771626 44699 771629
rect 41492 771624 44699 771626
rect 41492 771568 44638 771624
rect 44694 771568 44699 771624
rect 41492 771566 44699 771568
rect 44633 771563 44699 771566
rect 44817 771218 44883 771221
rect 41492 771216 44883 771218
rect 41492 771160 44822 771216
rect 44878 771160 44883 771216
rect 41492 771158 44883 771160
rect 44817 771155 44883 771158
rect 44633 770810 44699 770813
rect 41492 770808 44699 770810
rect 41492 770752 44638 770808
rect 44694 770752 44699 770808
rect 41492 770750 44699 770752
rect 44633 770747 44699 770750
rect 673913 770674 673979 770677
rect 683389 770674 683455 770677
rect 673913 770672 683455 770674
rect 673913 770616 673918 770672
rect 673974 770616 683394 770672
rect 683450 770616 683455 770672
rect 673913 770614 683455 770616
rect 673913 770611 673979 770614
rect 683389 770611 683455 770614
rect 44633 770402 44699 770405
rect 41492 770400 44699 770402
rect 41492 770344 44638 770400
rect 44694 770344 44699 770400
rect 41492 770342 44699 770344
rect 44633 770339 44699 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 676070 768708 676076 768772
rect 676140 768770 676146 768772
rect 680997 768770 681063 768773
rect 676140 768768 681063 768770
rect 676140 768712 681002 768768
rect 681058 768712 681063 768768
rect 676140 768710 681063 768712
rect 676140 768708 676146 768710
rect 680997 768707 681063 768710
rect 30974 768229 31034 768332
rect 30974 768224 31083 768229
rect 30974 768168 31022 768224
rect 31078 768168 31083 768224
rect 30974 768166 31083 768168
rect 31017 768163 31083 768166
rect 35574 767821 35634 767924
rect 35525 767816 35634 767821
rect 35801 767818 35867 767821
rect 35525 767760 35530 767816
rect 35586 767760 35634 767816
rect 35525 767758 35634 767760
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35525 767755 35591 767758
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 45093 766730 45159 766733
rect 41492 766728 45159 766730
rect 41492 766672 45098 766728
rect 45154 766672 45159 766728
rect 41492 766670 45159 766672
rect 45093 766667 45159 766670
rect 675201 766594 675267 766597
rect 675886 766594 675892 766596
rect 675201 766592 675892 766594
rect 675201 766536 675206 766592
rect 675262 766536 675892 766592
rect 675201 766534 675892 766536
rect 675201 766531 675267 766534
rect 675886 766532 675892 766534
rect 675956 766532 675962 766596
rect 42885 766322 42951 766325
rect 41492 766320 42951 766322
rect 41492 766264 42890 766320
rect 42946 766264 42951 766320
rect 41492 766262 42951 766264
rect 42885 766259 42951 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 41321 765778 41387 765781
rect 42701 765778 42767 765781
rect 41321 765776 42767 765778
rect 41321 765720 41326 765776
rect 41382 765720 42706 765776
rect 42762 765720 42767 765776
rect 41321 765718 42767 765720
rect 41321 765715 41387 765718
rect 42701 765715 42767 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 674833 765098 674899 765101
rect 676070 765098 676076 765100
rect 674833 765096 676076 765098
rect 40726 764964 40786 765068
rect 674833 765040 674838 765096
rect 674894 765040 676076 765096
rect 674833 765038 676076 765040
rect 674833 765035 674899 765038
rect 676070 765036 676076 765038
rect 676140 765036 676146 765100
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 45277 764826 45343 764829
rect 41462 764824 45343 764826
rect 41462 764768 45282 764824
rect 45338 764768 45343 764824
rect 41462 764766 45343 764768
rect 41462 764660 41522 764766
rect 45277 764763 45343 764766
rect 40033 764554 40099 764557
rect 41638 764554 41644 764556
rect 40033 764552 41644 764554
rect 40033 764496 40038 764552
rect 40094 764496 41644 764552
rect 40033 764494 41644 764496
rect 40033 764491 40099 764494
rect 41638 764492 41644 764494
rect 41708 764492 41714 764556
rect 46013 764282 46079 764285
rect 41492 764280 46079 764282
rect 41492 764224 46018 764280
rect 46074 764224 46079 764280
rect 41492 764222 46079 764224
rect 46013 764219 46079 764222
rect 37046 763333 37106 763844
rect 37046 763328 37155 763333
rect 651465 763330 651531 763333
rect 37046 763272 37094 763328
rect 37150 763272 37155 763328
rect 37046 763270 37155 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 37089 763267 37155 763270
rect 651465 763267 651531 763270
rect 43069 763058 43135 763061
rect 41492 763056 43135 763058
rect 41492 763000 43074 763056
rect 43130 763000 43135 763056
rect 41492 762998 43135 763000
rect 43069 762995 43135 762998
rect 671337 763058 671403 763061
rect 676029 763058 676095 763061
rect 671337 763056 676095 763058
rect 671337 763000 671342 763056
rect 671398 763000 676034 763056
rect 676090 763000 676095 763056
rect 671337 762998 676095 763000
rect 671337 762995 671403 762998
rect 676029 762995 676095 762998
rect 676949 761836 677015 761837
rect 676949 761832 676996 761836
rect 677060 761834 677066 761836
rect 676581 761792 676647 761793
rect 676581 761788 676628 761792
rect 676692 761790 676698 761792
rect 676581 761732 676586 761788
rect 676581 761728 676628 761732
rect 676692 761730 676738 761790
rect 676949 761776 676954 761832
rect 676949 761772 676996 761776
rect 677060 761774 677106 761834
rect 677060 761772 677066 761774
rect 676949 761771 677015 761772
rect 676692 761728 676698 761730
rect 676581 761727 676647 761728
rect 665817 761562 665883 761565
rect 665817 761560 676292 761562
rect 665817 761504 665822 761560
rect 665878 761504 676292 761560
rect 665817 761502 676292 761504
rect 665817 761499 665883 761502
rect 669270 761094 676292 761154
rect 663057 760474 663123 760477
rect 669270 760474 669330 761094
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 663057 760472 669330 760474
rect 663057 760416 663062 760472
rect 663118 760416 669330 760472
rect 663057 760414 669330 760416
rect 663057 760411 663123 760414
rect 671613 760338 671679 760341
rect 671613 760336 676292 760338
rect 671613 760280 671618 760336
rect 671674 760280 676292 760336
rect 671613 760278 676292 760280
rect 671613 760275 671679 760278
rect 671613 759930 671679 759933
rect 671613 759928 676292 759930
rect 671613 759872 671618 759928
rect 671674 759872 676292 759928
rect 671613 759870 676292 759872
rect 671613 759867 671679 759870
rect 671797 759522 671863 759525
rect 671797 759520 676292 759522
rect 671797 759464 671802 759520
rect 671858 759464 676292 759520
rect 671797 759462 676292 759464
rect 671797 759459 671863 759462
rect 672717 759114 672783 759117
rect 672717 759112 676292 759114
rect 672717 759056 672722 759112
rect 672778 759056 676292 759112
rect 672717 759054 676292 759056
rect 672717 759051 672783 759054
rect 41689 758842 41755 758845
rect 42241 758842 42307 758845
rect 41689 758840 42307 758842
rect 41689 758784 41694 758840
rect 41750 758784 42246 758840
rect 42302 758784 42307 758840
rect 41689 758782 42307 758784
rect 41689 758779 41755 758782
rect 42241 758779 42307 758782
rect 672349 758706 672415 758709
rect 672349 758704 676292 758706
rect 672349 758648 672354 758704
rect 672410 758648 676292 758704
rect 672349 758646 676292 758648
rect 672349 758643 672415 758646
rect 41689 758298 41755 758301
rect 42425 758298 42491 758301
rect 41689 758296 42491 758298
rect 41689 758240 41694 758296
rect 41750 758240 42430 758296
rect 42486 758240 42491 758296
rect 41689 758238 42491 758240
rect 41689 758235 41755 758238
rect 42425 758235 42491 758238
rect 671797 758298 671863 758301
rect 671797 758296 676292 758298
rect 671797 758240 671802 758296
rect 671858 758240 676292 758296
rect 671797 758238 676292 758240
rect 671797 758235 671863 758238
rect 39297 758026 39363 758029
rect 42241 758026 42307 758029
rect 39297 758024 42307 758026
rect 39297 757968 39302 758024
rect 39358 757968 42246 758024
rect 42302 757968 42307 758024
rect 39297 757966 42307 757968
rect 39297 757963 39363 757966
rect 42241 757963 42307 757966
rect 672165 757890 672231 757893
rect 672165 757888 676292 757890
rect 672165 757832 672170 757888
rect 672226 757832 676292 757888
rect 672165 757830 676292 757832
rect 672165 757827 672231 757830
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 670877 757482 670943 757485
rect 670877 757480 676292 757482
rect 670877 757424 670882 757480
rect 670938 757424 676292 757480
rect 670877 757422 676292 757424
rect 670877 757419 670943 757422
rect 39113 757346 39179 757349
rect 40350 757346 40356 757348
rect 39113 757344 40356 757346
rect 39113 757288 39118 757344
rect 39174 757288 40356 757344
rect 39113 757286 40356 757288
rect 39113 757283 39179 757286
rect 40350 757284 40356 757286
rect 40420 757284 40426 757348
rect 41781 757074 41847 757077
rect 680997 757074 681063 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 680997 757072 681076 757074
rect 680997 757016 681002 757072
rect 681058 757016 681076 757072
rect 680997 757014 681076 757016
rect 680997 757011 681063 757014
rect 41830 756669 41890 757011
rect 41830 756664 41939 756669
rect 41830 756608 41878 756664
rect 41934 756608 41939 756664
rect 41830 756606 41939 756608
rect 41873 756603 41939 756606
rect 683205 756666 683271 756669
rect 683205 756664 683284 756666
rect 683205 756608 683210 756664
rect 683266 756608 683284 756664
rect 683205 756606 683284 756608
rect 683205 756603 683271 756606
rect 42006 756332 42012 756396
rect 42076 756394 42082 756396
rect 46197 756394 46263 756397
rect 42076 756392 46263 756394
rect 42076 756336 46202 756392
rect 46258 756336 46263 756392
rect 42076 756334 46263 756336
rect 42076 756332 42082 756334
rect 46197 756331 46263 756334
rect 676170 756198 676292 756258
rect 676170 756122 676230 756198
rect 676078 756062 676230 756122
rect 668761 755986 668827 755989
rect 676078 755986 676138 756062
rect 668761 755984 676138 755986
rect 668761 755928 668766 755984
rect 668822 755928 676138 755984
rect 668761 755926 676138 755928
rect 668761 755923 668827 755926
rect 682377 755850 682443 755853
rect 682364 755848 682443 755850
rect 682364 755792 682382 755848
rect 682438 755792 682443 755848
rect 682364 755790 682443 755792
rect 682377 755787 682443 755790
rect 669589 755442 669655 755445
rect 669589 755440 676292 755442
rect 669589 755384 669594 755440
rect 669650 755384 676292 755440
rect 669589 755382 676292 755384
rect 669589 755379 669655 755382
rect 676949 755034 677015 755037
rect 676949 755032 677028 755034
rect 676949 754976 676954 755032
rect 677010 754976 677028 755032
rect 676949 754974 677028 754976
rect 676949 754971 677015 754974
rect 673862 754700 673868 754764
rect 673932 754762 673938 754764
rect 675845 754762 675911 754765
rect 673932 754760 675911 754762
rect 673932 754704 675850 754760
rect 675906 754704 675911 754760
rect 673932 754702 675911 754704
rect 673932 754700 673938 754702
rect 675845 754699 675911 754702
rect 676032 754566 676292 754626
rect 40350 754428 40356 754492
rect 40420 754490 40426 754492
rect 42425 754490 42491 754493
rect 676032 754490 676092 754566
rect 40420 754488 42491 754490
rect 40420 754432 42430 754488
rect 42486 754432 42491 754488
rect 40420 754430 42491 754432
rect 40420 754428 40426 754430
rect 42425 754427 42491 754430
rect 669270 754430 676092 754490
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 41965 754084 42031 754085
rect 41965 754080 42012 754084
rect 42076 754082 42082 754084
rect 41965 754024 41970 754080
rect 41965 754020 42012 754024
rect 42076 754022 42122 754082
rect 42076 754020 42082 754022
rect 41965 754019 42031 754020
rect 42241 753946 42307 753949
rect 42885 753946 42951 753949
rect 42241 753944 42951 753946
rect 42241 753888 42246 753944
rect 42302 753888 42890 753944
rect 42946 753888 42951 753944
rect 42241 753886 42951 753888
rect 42241 753883 42307 753886
rect 42885 753883 42951 753886
rect 669270 753541 669330 754430
rect 670509 754218 670575 754221
rect 670509 754216 676292 754218
rect 670509 754160 670514 754216
rect 670570 754160 676292 754216
rect 670509 754158 676292 754160
rect 670509 754155 670575 754158
rect 674414 753748 674420 753812
rect 674484 753810 674490 753812
rect 674484 753750 676292 753810
rect 674484 753748 674490 753750
rect 42885 753538 42951 753541
rect 45277 753538 45343 753541
rect 42885 753536 45343 753538
rect 42885 753480 42890 753536
rect 42946 753480 45282 753536
rect 45338 753480 45343 753536
rect 42885 753478 45343 753480
rect 42885 753475 42951 753478
rect 45277 753475 45343 753478
rect 669221 753536 669330 753541
rect 669221 753480 669226 753536
rect 669282 753480 669330 753536
rect 669221 753478 669330 753480
rect 669221 753475 669287 753478
rect 671153 753402 671219 753405
rect 671153 753400 676292 753402
rect 671153 753344 671158 753400
rect 671214 753344 676292 753400
rect 671153 753342 676292 753344
rect 671153 753339 671219 753342
rect 683389 752994 683455 752997
rect 683389 752992 683468 752994
rect 683389 752936 683394 752992
rect 683450 752936 683468 752992
rect 683389 752934 683468 752936
rect 683389 752931 683455 752934
rect 676029 752586 676095 752589
rect 676029 752584 676292 752586
rect 676029 752528 676034 752584
rect 676090 752528 676292 752584
rect 676029 752526 676292 752528
rect 676029 752523 676095 752526
rect 40718 752116 40724 752180
rect 40788 752178 40794 752180
rect 42241 752178 42307 752181
rect 683113 752178 683179 752181
rect 40788 752176 42307 752178
rect 40788 752120 42246 752176
rect 42302 752120 42307 752176
rect 40788 752118 42307 752120
rect 683100 752176 683179 752178
rect 683100 752120 683118 752176
rect 683174 752120 683179 752176
rect 683100 752118 683179 752120
rect 40788 752116 40794 752118
rect 42241 752115 42307 752118
rect 683113 752115 683179 752118
rect 42057 751770 42123 751773
rect 42885 751770 42951 751773
rect 42057 751768 42951 751770
rect 42057 751712 42062 751768
rect 42118 751712 42890 751768
rect 42946 751712 42951 751768
rect 42057 751710 42951 751712
rect 42057 751707 42123 751710
rect 42885 751707 42951 751710
rect 673085 751770 673151 751773
rect 673085 751768 676292 751770
rect 673085 751712 673090 751768
rect 673146 751712 676292 751768
rect 673085 751710 676292 751712
rect 673085 751707 673151 751710
rect 671061 751362 671127 751365
rect 671061 751360 676292 751362
rect 671061 751304 671066 751360
rect 671122 751304 676292 751360
rect 671061 751302 676292 751304
rect 671061 751299 671127 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 669270 750924 676660 750954
rect 669270 750894 676690 750924
rect 667841 750818 667907 750821
rect 669270 750818 669330 750894
rect 667841 750816 669330 750818
rect 667841 750760 667846 750816
rect 667902 750760 669330 750816
rect 667841 750758 669330 750760
rect 667841 750755 667907 750758
rect 676630 750516 676690 750894
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 671429 750138 671495 750141
rect 671429 750136 676292 750138
rect 671429 750080 671434 750136
rect 671490 750080 676292 750136
rect 671429 750078 676292 750080
rect 671429 750075 671495 750078
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 42425 749322 42491 749325
rect 45093 749322 45159 749325
rect 42425 749320 45159 749322
rect 42425 749264 42430 749320
rect 42486 749264 45098 749320
rect 45154 749264 45159 749320
rect 42425 749262 45159 749264
rect 42425 749259 42491 749262
rect 45093 749259 45159 749262
rect 41638 745044 41644 745108
rect 41708 745106 41714 745108
rect 42425 745106 42491 745109
rect 41708 745104 42491 745106
rect 41708 745048 42430 745104
rect 42486 745048 42491 745104
rect 41708 745046 42491 745048
rect 41708 745044 41714 745046
rect 42425 745043 42491 745046
rect 41822 744772 41828 744836
rect 41892 744834 41898 744836
rect 42241 744834 42307 744837
rect 41892 744832 42307 744834
rect 41892 744776 42246 744832
rect 42302 744776 42307 744832
rect 41892 744774 42307 744776
rect 41892 744772 41898 744774
rect 42241 744771 42307 744774
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 672257 743474 672323 743477
rect 674925 743474 674991 743477
rect 672257 743472 674991 743474
rect 672257 743416 672262 743472
rect 672318 743416 674930 743472
rect 674986 743416 674991 743472
rect 672257 743414 674991 743416
rect 672257 743411 672323 743414
rect 674925 743411 674991 743414
rect 667841 743202 667907 743205
rect 675109 743202 675175 743205
rect 667841 743200 675175 743202
rect 667841 743144 667846 743200
rect 667902 743144 675114 743200
rect 675170 743144 675175 743200
rect 667841 743142 675175 743144
rect 667841 743139 667907 743142
rect 675109 743139 675175 743142
rect 42701 743066 42767 743069
rect 62757 743066 62823 743069
rect 42701 743064 62823 743066
rect 42701 743008 42706 743064
rect 42762 743008 62762 743064
rect 62818 743008 62823 743064
rect 42701 743006 62823 743008
rect 42701 743003 42767 743006
rect 62757 743003 62823 743006
rect 666277 742522 666343 742525
rect 675017 742522 675083 742525
rect 666277 742520 675083 742522
rect 666277 742464 666282 742520
rect 666338 742464 675022 742520
rect 675078 742464 675083 742520
rect 666277 742462 675083 742464
rect 666277 742459 666343 742462
rect 675017 742459 675083 742462
rect 669405 741842 669471 741845
rect 674833 741842 674899 741845
rect 669405 741840 674899 741842
rect 669405 741784 669410 741840
rect 669466 741784 674838 741840
rect 674894 741784 674899 741840
rect 669405 741782 674899 741784
rect 669405 741779 669471 741782
rect 674833 741779 674899 741782
rect 674414 741508 674420 741572
rect 674484 741570 674490 741572
rect 675109 741570 675175 741573
rect 674484 741568 675175 741570
rect 674484 741512 675114 741568
rect 675170 741512 675175 741568
rect 674484 741510 675175 741512
rect 674484 741508 674490 741510
rect 675109 741507 675175 741510
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 672073 741162 672139 741165
rect 674925 741162 674991 741165
rect 672073 741160 674991 741162
rect 672073 741104 672078 741160
rect 672134 741104 674930 741160
rect 674986 741104 674991 741160
rect 672073 741102 674991 741104
rect 672073 741099 672139 741102
rect 674925 741099 674991 741102
rect 669589 738578 669655 738581
rect 675293 738578 675359 738581
rect 669589 738576 675359 738578
rect 669589 738520 669594 738576
rect 669650 738520 675298 738576
rect 675354 738520 675359 738576
rect 669589 738518 675359 738520
rect 669589 738515 669655 738518
rect 675293 738515 675359 738518
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675477 738170 675543 738173
rect 674668 738168 675543 738170
rect 674668 738112 675482 738168
rect 675538 738112 675543 738168
rect 674668 738110 675543 738112
rect 674668 738108 674674 738110
rect 675477 738107 675543 738110
rect 671245 737082 671311 737085
rect 675109 737082 675175 737085
rect 671245 737080 675175 737082
rect 671245 737024 671250 737080
rect 671306 737024 675114 737080
rect 675170 737024 675175 737080
rect 671245 737022 675175 737024
rect 671245 737019 671311 737022
rect 675109 737019 675175 737022
rect 652017 736810 652083 736813
rect 650164 736808 652083 736810
rect 650164 736752 652022 736808
rect 652078 736752 652083 736808
rect 650164 736750 652083 736752
rect 652017 736747 652083 736750
rect 668393 734770 668459 734773
rect 674925 734770 674991 734773
rect 668393 734768 674991 734770
rect 668393 734712 668398 734768
rect 668454 734712 674930 734768
rect 674986 734712 674991 734768
rect 668393 734710 674991 734712
rect 668393 734707 668459 734710
rect 674925 734707 674991 734710
rect 669129 734498 669195 734501
rect 675109 734498 675175 734501
rect 669129 734496 675175 734498
rect 669129 734440 669134 734496
rect 669190 734440 675114 734496
rect 675170 734440 675175 734496
rect 669129 734438 675175 734440
rect 669129 734435 669195 734438
rect 675109 734435 675175 734438
rect 670693 734092 670759 734093
rect 670693 734090 670740 734092
rect 670648 734088 670740 734090
rect 670648 734032 670698 734088
rect 670648 734030 670740 734032
rect 670693 734028 670740 734030
rect 670804 734028 670810 734092
rect 670693 734027 670759 734028
rect 673085 733682 673151 733685
rect 675109 733682 675175 733685
rect 673085 733680 675175 733682
rect 673085 733624 673090 733680
rect 673146 733624 675114 733680
rect 675170 733624 675175 733680
rect 673085 733622 675175 733624
rect 673085 733619 673151 733622
rect 675109 733619 675175 733622
rect 668393 733138 668459 733141
rect 674649 733138 674715 733141
rect 668393 733136 674715 733138
rect 668393 733080 668398 733136
rect 668454 733080 674654 733136
rect 674710 733080 674715 733136
rect 668393 733078 674715 733080
rect 668393 733075 668459 733078
rect 674649 733075 674715 733078
rect 674230 732804 674236 732868
rect 674300 732866 674306 732868
rect 675109 732866 675175 732869
rect 674300 732864 675175 732866
rect 674300 732808 675114 732864
rect 675170 732808 675175 732864
rect 674300 732806 675175 732808
rect 674300 732804 674306 732806
rect 675109 732803 675175 732806
rect 668761 731506 668827 731509
rect 674649 731506 674715 731509
rect 668761 731504 674715 731506
rect 668761 731448 668766 731504
rect 668822 731448 674654 731504
rect 674710 731448 674715 731504
rect 668761 731446 674715 731448
rect 668761 731443 668827 731446
rect 674649 731443 674715 731446
rect 41492 731310 51090 731370
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 44449 730146 44515 730149
rect 41492 730144 44515 730146
rect 41492 730088 44454 730144
rect 44510 730088 44515 730144
rect 41492 730086 44515 730088
rect 51030 730146 51090 731310
rect 671981 730554 672047 730557
rect 675109 730554 675175 730557
rect 671981 730552 675175 730554
rect 671981 730496 671986 730552
rect 672042 730496 675114 730552
rect 675170 730496 675175 730552
rect 671981 730494 675175 730496
rect 671981 730491 672047 730494
rect 675109 730491 675175 730494
rect 53097 730146 53163 730149
rect 51030 730144 53163 730146
rect 51030 730088 53102 730144
rect 53158 730088 53163 730144
rect 51030 730086 53163 730088
rect 44449 730083 44515 730086
rect 53097 730083 53163 730086
rect 45001 729738 45067 729741
rect 41492 729736 45067 729738
rect 41492 729680 45006 729736
rect 45062 729680 45067 729736
rect 41492 729678 45067 729680
rect 45001 729675 45067 729678
rect 44265 729330 44331 729333
rect 41492 729328 44331 729330
rect 41492 729272 44270 729328
rect 44326 729272 44331 729328
rect 41492 729270 44331 729272
rect 44265 729267 44331 729270
rect 44449 728922 44515 728925
rect 41492 728920 44515 728922
rect 41492 728864 44454 728920
rect 44510 728864 44515 728920
rect 41492 728862 44515 728864
rect 44449 728859 44515 728862
rect 675886 728724 675892 728788
rect 675956 728786 675962 728788
rect 676806 728786 676812 728788
rect 675956 728726 676812 728786
rect 675956 728724 675962 728726
rect 676806 728724 676812 728726
rect 676876 728724 676882 728788
rect 44817 728514 44883 728517
rect 41492 728512 44883 728514
rect 41492 728456 44822 728512
rect 44878 728456 44883 728512
rect 41492 728454 44883 728456
rect 44817 728451 44883 728454
rect 670693 728516 670759 728517
rect 670693 728512 670740 728516
rect 670804 728514 670810 728516
rect 670693 728456 670698 728512
rect 670693 728452 670740 728456
rect 670804 728454 670850 728514
rect 670804 728452 670810 728454
rect 670693 728451 670759 728452
rect 671429 728378 671495 728381
rect 673361 728378 673427 728381
rect 671429 728376 673427 728378
rect 671429 728320 671434 728376
rect 671490 728320 673366 728376
rect 673422 728320 673427 728376
rect 671429 728318 673427 728320
rect 671429 728315 671495 728318
rect 673361 728315 673427 728318
rect 62757 728242 62823 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 62757 728179 62823 728182
rect 44265 728106 44331 728109
rect 41492 728104 44331 728106
rect 41492 728048 44270 728104
rect 44326 728048 44331 728104
rect 41492 728046 44331 728048
rect 44265 728043 44331 728046
rect 671061 728106 671127 728109
rect 673361 728106 673427 728109
rect 671061 728104 673427 728106
rect 671061 728048 671066 728104
rect 671122 728048 673366 728104
rect 673422 728048 673427 728104
rect 671061 728046 673427 728048
rect 671061 728043 671127 728046
rect 673361 728043 673427 728046
rect 674281 727970 674347 727973
rect 683757 727970 683823 727973
rect 674281 727968 683823 727970
rect 674281 727912 674286 727968
rect 674342 727912 683762 727968
rect 683818 727912 683823 727968
rect 674281 727910 683823 727912
rect 674281 727907 674347 727910
rect 683757 727907 683823 727910
rect 44633 727698 44699 727701
rect 41492 727696 44699 727698
rect 41492 727640 44638 727696
rect 44694 727640 44699 727696
rect 41492 727638 44699 727640
rect 44633 727635 44699 727638
rect 44633 727426 44699 727429
rect 41830 727424 44699 727426
rect 41830 727368 44638 727424
rect 44694 727368 44699 727424
rect 41830 727366 44699 727368
rect 41830 727290 41890 727366
rect 44633 727363 44699 727366
rect 41492 727230 41890 727290
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 674097 726882 674163 726885
rect 674097 726880 677610 726882
rect 674097 726824 674102 726880
rect 674158 726824 677610 726880
rect 674097 726822 677610 726824
rect 674097 726819 674163 726822
rect 677550 726746 677610 726822
rect 683205 726746 683271 726749
rect 677550 726744 683271 726746
rect 677550 726688 683210 726744
rect 683266 726688 683271 726744
rect 677550 726686 683271 726688
rect 683205 726683 683271 726686
rect 674741 726610 674807 726613
rect 674741 726608 674850 726610
rect 674741 726552 674746 726608
rect 674802 726552 674850 726608
rect 674741 726547 674850 726552
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 674790 726474 674850 726547
rect 683389 726474 683455 726477
rect 674790 726472 683455 726474
rect 674790 726416 683394 726472
rect 683450 726416 683455 726472
rect 674790 726414 683455 726416
rect 41321 726411 41387 726414
rect 683389 726411 683455 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 682377 725794 682443 725797
rect 676140 725792 682443 725794
rect 676140 725736 682382 725792
rect 682438 725736 682443 725792
rect 676140 725734 682443 725736
rect 676140 725732 676146 725734
rect 682377 725731 682443 725734
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 33777 725250 33843 725253
rect 33764 725248 33843 725250
rect 33764 725192 33782 725248
rect 33838 725192 33843 725248
rect 33764 725190 33843 725192
rect 33777 725187 33843 725190
rect 673729 725114 673795 725117
rect 683573 725114 683639 725117
rect 673729 725112 683639 725114
rect 673729 725056 673734 725112
rect 673790 725056 683578 725112
rect 683634 725056 683639 725112
rect 673729 725054 683639 725056
rect 673729 725051 673795 725054
rect 683573 725051 683639 725054
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 40677 724434 40743 724437
rect 40677 724432 40756 724434
rect 40677 724376 40682 724432
rect 40738 724376 40756 724432
rect 40677 724374 40756 724376
rect 40677 724371 40743 724374
rect 33041 724026 33107 724029
rect 33028 724024 33107 724026
rect 33028 723968 33046 724024
rect 33102 723968 33107 724024
rect 33028 723966 33107 723968
rect 33041 723963 33107 723966
rect 45185 723618 45251 723621
rect 41492 723616 45251 723618
rect 41492 723560 45190 723616
rect 45246 723560 45251 723616
rect 41492 723558 45251 723560
rect 45185 723555 45251 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 31661 723210 31727 723213
rect 31661 723208 31740 723210
rect 31661 723152 31666 723208
rect 31722 723152 31740 723208
rect 31661 723150 31740 723152
rect 31661 723147 31727 723150
rect 44817 722802 44883 722805
rect 41492 722800 44883 722802
rect 41492 722744 44822 722800
rect 44878 722744 44883 722800
rect 41492 722742 44883 722744
rect 44817 722739 44883 722742
rect 41873 722394 41939 722397
rect 41492 722392 41939 722394
rect 41492 722336 41878 722392
rect 41934 722336 41939 722392
rect 41492 722334 41939 722336
rect 41873 722331 41939 722334
rect 40726 721772 40786 721956
rect 40350 721708 40356 721772
rect 40420 721708 40426 721772
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 40358 721548 40418 721708
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 46933 721170 46999 721173
rect 41492 721168 46999 721170
rect 41492 721112 46938 721168
rect 46994 721112 46999 721168
rect 41492 721110 46999 721112
rect 46933 721107 46999 721110
rect 42149 720354 42215 720357
rect 41492 720352 42215 720354
rect 41492 720296 42154 720352
rect 42210 720296 42215 720352
rect 41492 720294 42215 720296
rect 42149 720291 42215 720294
rect 47853 719946 47919 719949
rect 41492 719944 47919 719946
rect 41492 719888 47858 719944
rect 47914 719888 47919 719944
rect 41492 719886 47919 719888
rect 47853 719883 47919 719886
rect 41689 719674 41755 719677
rect 42517 719674 42583 719677
rect 41689 719672 42583 719674
rect 41689 719616 41694 719672
rect 41750 719616 42522 719672
rect 42578 719616 42583 719672
rect 41689 719614 42583 719616
rect 41689 719611 41755 719614
rect 42517 719611 42583 719614
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41873 718586 41939 718589
rect 40604 718584 41939 718586
rect 40604 718528 41878 718584
rect 41934 718528 41939 718584
rect 40604 718526 41939 718528
rect 40604 718524 40610 718526
rect 41873 718523 41939 718526
rect 40350 716756 40356 716820
rect 40420 716818 40426 716820
rect 40902 716818 40908 716820
rect 40420 716758 40908 716818
rect 40420 716756 40426 716758
rect 40902 716756 40908 716758
rect 40972 716756 40978 716820
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 659610 716078 676292 716138
rect 658917 716002 658983 716005
rect 659610 716002 659670 716078
rect 658917 716000 659670 716002
rect 658917 715944 658922 716000
rect 658978 715944 659670 716000
rect 658917 715942 659670 715944
rect 658917 715939 658983 715942
rect 41137 715866 41203 715869
rect 41689 715866 41755 715869
rect 42701 715866 42767 715869
rect 41137 715864 41430 715866
rect 41137 715808 41142 715864
rect 41198 715808 41430 715864
rect 41137 715806 41430 715808
rect 41137 715803 41203 715806
rect 41370 715594 41430 715806
rect 41689 715864 42767 715866
rect 41689 715808 41694 715864
rect 41750 715808 42706 715864
rect 42762 715808 42767 715864
rect 41689 715806 42767 715808
rect 41689 715803 41755 715806
rect 42701 715803 42767 715806
rect 669957 715730 670023 715733
rect 669957 715728 676292 715730
rect 669957 715672 669962 715728
rect 670018 715672 676292 715728
rect 669957 715670 676292 715672
rect 669957 715667 670023 715670
rect 42885 715594 42951 715597
rect 41370 715592 42951 715594
rect 41370 715536 42890 715592
rect 42946 715536 42951 715592
rect 41370 715534 42951 715536
rect 42885 715531 42951 715534
rect 62113 715322 62179 715325
rect 671613 715322 671679 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 671613 715320 676292 715322
rect 671613 715264 671618 715320
rect 671674 715264 676292 715320
rect 671613 715262 676292 715264
rect 62113 715259 62179 715262
rect 671613 715259 671679 715262
rect 671613 714914 671679 714917
rect 671613 714912 676292 714914
rect 671613 714856 671618 714912
rect 671674 714856 676292 714912
rect 671613 714854 676292 714856
rect 671613 714851 671679 714854
rect 40677 714778 40743 714781
rect 41822 714778 41828 714780
rect 40677 714776 41828 714778
rect 40677 714720 40682 714776
rect 40738 714720 41828 714776
rect 40677 714718 41828 714720
rect 40677 714715 40743 714718
rect 41822 714716 41828 714718
rect 41892 714716 41898 714780
rect 41965 714644 42031 714645
rect 41965 714640 42012 714644
rect 42076 714642 42082 714644
rect 41965 714584 41970 714640
rect 41965 714580 42012 714584
rect 42076 714582 42122 714642
rect 42076 714580 42082 714582
rect 41965 714579 42031 714580
rect 672717 714506 672783 714509
rect 672717 714504 676292 714506
rect 672717 714448 672722 714504
rect 672778 714448 676292 714504
rect 672717 714446 676292 714448
rect 672717 714443 672783 714446
rect 671429 714098 671495 714101
rect 671429 714096 676292 714098
rect 671429 714040 671434 714096
rect 671490 714040 676292 714096
rect 671429 714038 676292 714040
rect 671429 714035 671495 714038
rect 671797 713690 671863 713693
rect 671797 713688 676292 713690
rect 671797 713632 671802 713688
rect 671858 713632 676292 713688
rect 671797 713630 676292 713632
rect 671797 713627 671863 713630
rect 670877 713282 670943 713285
rect 670877 713280 676292 713282
rect 670877 713224 670882 713280
rect 670938 713224 676292 713280
rect 670877 713222 676292 713224
rect 670877 713219 670943 713222
rect 671061 712874 671127 712877
rect 671061 712872 676292 712874
rect 671061 712816 671066 712872
rect 671122 712816 676292 712872
rect 671061 712814 676292 712816
rect 671061 712811 671127 712814
rect 671061 712466 671127 712469
rect 671061 712464 676292 712466
rect 671061 712408 671066 712464
rect 671122 712408 676292 712464
rect 671061 712406 676292 712408
rect 671061 712403 671127 712406
rect 47577 712194 47643 712197
rect 42198 712192 47643 712194
rect 42198 712136 47582 712192
rect 47638 712136 47643 712192
rect 42198 712134 47643 712136
rect 42198 711109 42258 712134
rect 47577 712131 47643 712134
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 666461 711650 666527 711653
rect 666461 711648 676292 711650
rect 666461 711592 666466 711648
rect 666522 711592 676292 711648
rect 666461 711590 676292 711592
rect 666461 711587 666527 711590
rect 683389 711242 683455 711245
rect 683389 711240 683468 711242
rect 683389 711184 683394 711240
rect 683450 711184 683468 711240
rect 683389 711182 683468 711184
rect 683389 711179 683455 711182
rect 42198 711104 42307 711109
rect 42198 711048 42246 711104
rect 42302 711048 42307 711104
rect 42198 711046 42307 711048
rect 42241 711043 42307 711046
rect 682377 710834 682443 710837
rect 682364 710832 682443 710834
rect 682364 710776 682382 710832
rect 682438 710776 682443 710832
rect 682364 710774 682443 710776
rect 682377 710771 682443 710774
rect 668209 710426 668275 710429
rect 668209 710424 676292 710426
rect 668209 710368 668214 710424
rect 668270 710368 676292 710424
rect 668209 710366 676292 710368
rect 668209 710363 668275 710366
rect 651465 710290 651531 710293
rect 650164 710288 651531 710290
rect 650164 710232 651470 710288
rect 651526 710232 651531 710288
rect 650164 710230 651531 710232
rect 651465 710227 651531 710230
rect 672901 710018 672967 710021
rect 672901 710016 676292 710018
rect 672901 709960 672906 710016
rect 672962 709960 676292 710016
rect 672901 709958 676292 709960
rect 672901 709955 672967 709958
rect 41965 709884 42031 709885
rect 41965 709880 42012 709884
rect 42076 709882 42082 709884
rect 41965 709824 41970 709880
rect 41965 709820 42012 709824
rect 42076 709822 42122 709882
rect 42076 709820 42082 709822
rect 41965 709819 42031 709820
rect 669773 709610 669839 709613
rect 669773 709608 676292 709610
rect 669773 709552 669778 709608
rect 669834 709552 676292 709608
rect 669773 709550 676292 709552
rect 669773 709547 669839 709550
rect 44817 709474 44883 709477
rect 42198 709472 44883 709474
rect 42198 709416 44822 709472
rect 44878 709416 44883 709472
rect 42198 709414 44883 709416
rect 42198 709205 42258 709414
rect 44817 709411 44883 709414
rect 42198 709200 42307 709205
rect 42198 709144 42246 709200
rect 42302 709144 42307 709200
rect 42198 709142 42307 709144
rect 42241 709139 42307 709142
rect 672533 709202 672599 709205
rect 672533 709200 676292 709202
rect 672533 709144 672538 709200
rect 672594 709144 676292 709200
rect 672533 709142 676292 709144
rect 672533 709139 672599 709142
rect 668945 708794 669011 708797
rect 668945 708792 676292 708794
rect 668945 708736 668950 708792
rect 669006 708736 676292 708792
rect 668945 708734 676292 708736
rect 668945 708731 669011 708734
rect 40902 708460 40908 708524
rect 40972 708522 40978 708524
rect 41781 708522 41847 708525
rect 40972 708520 41847 708522
rect 40972 708464 41786 708520
rect 41842 708464 41847 708520
rect 40972 708462 41847 708464
rect 40972 708460 40978 708462
rect 41781 708459 41847 708462
rect 673545 708386 673611 708389
rect 673545 708384 676292 708386
rect 673545 708328 673550 708384
rect 673606 708328 676292 708384
rect 673545 708326 676292 708328
rect 673545 708323 673611 708326
rect 683573 707978 683639 707981
rect 683573 707976 683652 707978
rect 683573 707920 683578 707976
rect 683634 707920 683652 707976
rect 683573 707918 683652 707920
rect 683573 707915 683639 707918
rect 683757 707570 683823 707573
rect 683757 707568 683836 707570
rect 683757 707512 683762 707568
rect 683818 707512 683836 707568
rect 683757 707510 683836 707512
rect 683757 707507 683823 707510
rect 670325 707162 670391 707165
rect 670325 707160 676292 707162
rect 670325 707104 670330 707160
rect 670386 707104 676292 707160
rect 670325 707102 676292 707104
rect 670325 707099 670391 707102
rect 40718 706692 40724 706756
rect 40788 706754 40794 706756
rect 41781 706754 41847 706757
rect 40788 706752 41847 706754
rect 40788 706696 41786 706752
rect 41842 706696 41847 706752
rect 40788 706694 41847 706696
rect 40788 706692 40794 706694
rect 41781 706691 41847 706694
rect 42149 706754 42215 706757
rect 42701 706754 42767 706757
rect 42149 706752 42767 706754
rect 42149 706696 42154 706752
rect 42210 706696 42706 706752
rect 42762 706696 42767 706752
rect 42149 706694 42767 706696
rect 42149 706691 42215 706694
rect 42701 706691 42767 706694
rect 683205 706754 683271 706757
rect 683205 706752 683284 706754
rect 683205 706696 683210 706752
rect 683266 706696 683284 706752
rect 683205 706694 683284 706696
rect 683205 706691 683271 706694
rect 674373 706346 674439 706349
rect 674373 706344 676292 706346
rect 674373 706288 674378 706344
rect 674434 706288 676292 706344
rect 674373 706286 676292 706288
rect 674373 706283 674439 706286
rect 670141 705938 670207 705941
rect 670141 705936 676292 705938
rect 670141 705880 670146 705936
rect 670202 705908 676292 705936
rect 670202 705880 676322 705908
rect 670141 705878 676322 705880
rect 670141 705875 670207 705878
rect 42241 705530 42307 705533
rect 45185 705530 45251 705533
rect 42241 705528 45251 705530
rect 42241 705472 42246 705528
rect 42302 705472 45190 705528
rect 45246 705472 45251 705528
rect 676262 705500 676322 705878
rect 42241 705470 45251 705472
rect 42241 705467 42307 705470
rect 45185 705467 45251 705470
rect 673310 705060 673316 705124
rect 673380 705122 673386 705124
rect 673380 705062 676292 705122
rect 673380 705060 673386 705062
rect 40534 704244 40540 704308
rect 40604 704306 40610 704308
rect 41781 704306 41847 704309
rect 40604 704304 41847 704306
rect 40604 704248 41786 704304
rect 41842 704248 41847 704304
rect 40604 704246 41847 704248
rect 40604 704244 40610 704246
rect 41781 704243 41847 704246
rect 42057 703082 42123 703085
rect 42701 703082 42767 703085
rect 42057 703080 42767 703082
rect 42057 703024 42062 703080
rect 42118 703024 42706 703080
rect 42762 703024 42767 703080
rect 42057 703022 42767 703024
rect 42057 703019 42123 703022
rect 42701 703019 42767 703022
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42333 701858 42399 701861
rect 41892 701856 42399 701858
rect 41892 701800 42338 701856
rect 42394 701800 42399 701856
rect 41892 701798 42399 701800
rect 41892 701796 41898 701798
rect 42333 701795 42399 701798
rect 41638 701524 41644 701588
rect 41708 701586 41714 701588
rect 42609 701586 42675 701589
rect 41708 701584 42675 701586
rect 41708 701528 42614 701584
rect 42670 701528 42675 701584
rect 41708 701526 42675 701528
rect 41708 701524 41714 701526
rect 42609 701523 42675 701526
rect 669221 701178 669287 701181
rect 675109 701178 675175 701181
rect 669221 701176 675175 701178
rect 669221 701120 669226 701176
rect 669282 701120 675114 701176
rect 675170 701120 675175 701176
rect 669221 701118 675175 701120
rect 669221 701115 669287 701118
rect 675109 701115 675175 701118
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 666461 699818 666527 699821
rect 674833 699818 674899 699821
rect 666461 699816 674899 699818
rect 666461 699760 666466 699816
rect 666522 699760 674838 699816
rect 674894 699760 674899 699816
rect 666461 699758 674899 699760
rect 666461 699755 666527 699758
rect 674833 699755 674899 699758
rect 41689 697914 41755 697917
rect 62757 697914 62823 697917
rect 41689 697912 62823 697914
rect 41689 697856 41694 697912
rect 41750 697856 62762 697912
rect 62818 697856 62823 697912
rect 41689 697854 62823 697856
rect 41689 697851 41755 697854
rect 62757 697851 62823 697854
rect 674557 697234 674623 697237
rect 675109 697234 675175 697237
rect 674557 697232 675175 697234
rect 674557 697176 674562 697232
rect 674618 697176 675114 697232
rect 675170 697176 675175 697232
rect 674557 697174 675175 697176
rect 674557 697171 674623 697174
rect 675109 697171 675175 697174
rect 651465 696962 651531 696965
rect 650164 696960 651531 696962
rect 650164 696904 651470 696960
rect 651526 696904 651531 696960
rect 650164 696902 651531 696904
rect 651465 696899 651531 696902
rect 669773 696962 669839 696965
rect 674741 696962 674807 696965
rect 669773 696960 674807 696962
rect 669773 696904 669778 696960
rect 669834 696904 674746 696960
rect 674802 696904 674807 696960
rect 669773 696902 674807 696904
rect 669773 696899 669839 696902
rect 674741 696899 674807 696902
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676990 694106 676996 694108
rect 675894 694046 676996 694106
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 674005 693154 674071 693157
rect 675477 693154 675543 693157
rect 674005 693152 675543 693154
rect 674005 693096 674010 693152
rect 674066 693096 675482 693152
rect 675538 693096 675543 693152
rect 674005 693094 675543 693096
rect 674005 693091 674071 693094
rect 675477 693091 675543 693094
rect 674189 692882 674255 692885
rect 675109 692882 675175 692885
rect 674189 692880 675175 692882
rect 674189 692824 674194 692880
rect 674250 692824 675114 692880
rect 675170 692824 675175 692880
rect 674189 692822 675175 692824
rect 674189 692819 674255 692822
rect 675109 692819 675175 692822
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 670417 690434 670483 690437
rect 675109 690434 675175 690437
rect 670417 690432 675175 690434
rect 670417 690376 670422 690432
rect 670478 690376 675114 690432
rect 675170 690376 675175 690432
rect 670417 690374 675175 690376
rect 670417 690371 670483 690374
rect 675109 690371 675175 690374
rect 673453 690162 673519 690165
rect 675385 690162 675451 690165
rect 673453 690160 675451 690162
rect 673453 690104 673458 690160
rect 673514 690104 675390 690160
rect 675446 690104 675451 690160
rect 673453 690102 675451 690104
rect 673453 690099 673519 690102
rect 675385 690099 675451 690102
rect 674557 689754 674623 689757
rect 674782 689754 674788 689756
rect 674557 689752 674788 689754
rect 674557 689696 674562 689752
rect 674618 689696 674788 689752
rect 674557 689694 674788 689696
rect 674557 689691 674623 689694
rect 674782 689692 674788 689694
rect 674852 689692 674858 689756
rect 663057 689346 663123 689349
rect 674925 689346 674991 689349
rect 663057 689344 674991 689346
rect 663057 689288 663062 689344
rect 663118 689288 674930 689344
rect 674986 689288 674991 689344
rect 663057 689286 674991 689288
rect 663057 689283 663123 689286
rect 674925 689283 674991 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 673269 689074 673335 689077
rect 675109 689074 675175 689077
rect 673269 689072 675175 689074
rect 673269 689016 673274 689072
rect 673330 689016 675114 689072
rect 675170 689016 675175 689072
rect 673269 689014 675175 689016
rect 673269 689011 673335 689014
rect 675109 689011 675175 689014
rect 674741 688804 674807 688805
rect 674741 688802 674788 688804
rect 674696 688800 674788 688802
rect 674696 688744 674746 688800
rect 674696 688742 674788 688744
rect 674741 688740 674788 688742
rect 674852 688740 674858 688804
rect 674741 688739 674807 688740
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 41321 687714 41387 687717
rect 41308 687712 41387 687714
rect 41308 687656 41326 687712
rect 41382 687656 41387 687712
rect 41308 687654 41387 687656
rect 41321 687651 41387 687654
rect 671797 687442 671863 687445
rect 675109 687442 675175 687445
rect 671797 687440 675175 687442
rect 671797 687384 671802 687440
rect 671858 687384 675114 687440
rect 675170 687384 675175 687440
rect 671797 687382 675175 687384
rect 671797 687379 671863 687382
rect 675109 687379 675175 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 45001 686898 45067 686901
rect 41492 686896 45067 686898
rect 41492 686840 45006 686896
rect 45062 686840 45067 686896
rect 41492 686838 45067 686840
rect 45001 686835 45067 686838
rect 44817 686490 44883 686493
rect 41492 686488 44883 686490
rect 41492 686432 44822 686488
rect 44878 686432 44883 686488
rect 41492 686430 44883 686432
rect 44817 686427 44883 686430
rect 668025 686218 668091 686221
rect 675109 686218 675175 686221
rect 668025 686216 675175 686218
rect 668025 686160 668030 686216
rect 668086 686160 675114 686216
rect 675170 686160 675175 686216
rect 668025 686158 675175 686160
rect 668025 686155 668091 686158
rect 675109 686155 675175 686158
rect 44449 686082 44515 686085
rect 41492 686080 44515 686082
rect 41492 686024 44454 686080
rect 44510 686024 44515 686080
rect 41492 686022 44515 686024
rect 44449 686019 44515 686022
rect 672441 685946 672507 685949
rect 674925 685946 674991 685949
rect 672441 685944 674991 685946
rect 672441 685888 672446 685944
rect 672502 685888 674930 685944
rect 674986 685888 674991 685944
rect 672441 685886 674991 685888
rect 672441 685883 672507 685886
rect 674925 685883 674991 685886
rect 45001 685674 45067 685677
rect 41492 685672 45067 685674
rect 41492 685616 45006 685672
rect 45062 685616 45067 685672
rect 41492 685614 45067 685616
rect 45001 685611 45067 685614
rect 670233 685402 670299 685405
rect 675109 685402 675175 685405
rect 670233 685400 675175 685402
rect 670233 685344 670238 685400
rect 670294 685344 675114 685400
rect 675170 685344 675175 685400
rect 670233 685342 675175 685344
rect 670233 685339 670299 685342
rect 675109 685339 675175 685342
rect 44265 685266 44331 685269
rect 41492 685264 44331 685266
rect 41492 685208 44270 685264
rect 44326 685208 44331 685264
rect 41492 685206 44331 685208
rect 44265 685203 44331 685206
rect 44357 684858 44423 684861
rect 41492 684856 44423 684858
rect 41492 684800 44362 684856
rect 44418 684800 44423 684856
rect 41492 684798 44423 684800
rect 44357 684795 44423 684798
rect 44633 684450 44699 684453
rect 41492 684448 44699 684450
rect 41492 684392 44638 684448
rect 44694 684392 44699 684448
rect 41492 684390 44699 684392
rect 44633 684387 44699 684390
rect 45369 684042 45435 684045
rect 41492 684040 45435 684042
rect 41492 683984 45374 684040
rect 45430 683984 45435 684040
rect 41492 683982 45435 683984
rect 45369 683979 45435 683982
rect 42190 683634 42196 683636
rect 41492 683574 42196 683634
rect 42190 683572 42196 683574
rect 42260 683572 42266 683636
rect 651649 683634 651715 683637
rect 650164 683632 651715 683634
rect 650164 683576 651654 683632
rect 651710 683576 651715 683632
rect 650164 683574 651715 683576
rect 651649 683571 651715 683574
rect 41321 683226 41387 683229
rect 41308 683224 41387 683226
rect 41308 683168 41326 683224
rect 41382 683168 41387 683224
rect 41308 683166 41387 683168
rect 41321 683163 41387 683166
rect 42006 682818 42012 682820
rect 41492 682758 42012 682818
rect 42006 682756 42012 682758
rect 42076 682756 42082 682820
rect 41321 682410 41387 682413
rect 41308 682408 41387 682410
rect 41308 682352 41326 682408
rect 41382 682352 41387 682408
rect 41308 682350 41387 682352
rect 41321 682347 41387 682350
rect 674414 682348 674420 682412
rect 674484 682410 674490 682412
rect 683205 682410 683271 682413
rect 674484 682408 683271 682410
rect 674484 682352 683210 682408
rect 683266 682352 683271 682408
rect 674484 682350 683271 682352
rect 674484 682348 674490 682350
rect 683205 682347 683271 682350
rect 40033 682002 40099 682005
rect 40020 682000 40099 682002
rect 40020 681944 40038 682000
rect 40094 681944 40099 682000
rect 40020 681942 40099 681944
rect 40033 681939 40099 681942
rect 41689 681866 41755 681869
rect 42609 681866 42675 681869
rect 41689 681864 42675 681866
rect 41689 681808 41694 681864
rect 41750 681808 42614 681864
rect 42670 681808 42675 681864
rect 41689 681806 42675 681808
rect 41689 681803 41755 681806
rect 42609 681803 42675 681806
rect 36721 681594 36787 681597
rect 36708 681592 36787 681594
rect 36708 681536 36726 681592
rect 36782 681536 36787 681592
rect 36708 681534 36787 681536
rect 36721 681531 36787 681534
rect 36537 681186 36603 681189
rect 36524 681184 36603 681186
rect 36524 681128 36542 681184
rect 36598 681128 36603 681184
rect 36524 681126 36603 681128
rect 36537 681123 36603 681126
rect 674230 680988 674236 681052
rect 674300 681050 674306 681052
rect 683389 681050 683455 681053
rect 674300 681048 683455 681050
rect 674300 680992 683394 681048
rect 683450 680992 683455 681048
rect 674300 680990 683455 680992
rect 674300 680988 674306 680990
rect 683389 680987 683455 680990
rect 35157 680778 35223 680781
rect 35157 680776 35236 680778
rect 35157 680720 35162 680776
rect 35218 680720 35236 680776
rect 35157 680718 35236 680720
rect 35157 680715 35223 680718
rect 44541 680370 44607 680373
rect 41492 680368 44607 680370
rect 41492 680312 44546 680368
rect 44602 680312 44607 680368
rect 41492 680310 44607 680312
rect 44541 680307 44607 680310
rect 42793 679962 42859 679965
rect 41492 679960 42859 679962
rect 41492 679904 42798 679960
rect 42854 679904 42859 679960
rect 41492 679902 42859 679904
rect 42793 679899 42859 679902
rect 44173 679554 44239 679557
rect 41492 679552 44239 679554
rect 41492 679496 44178 679552
rect 44234 679496 44239 679552
rect 41492 679494 44239 679496
rect 44173 679491 44239 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40902 678928 40908 678992
rect 40972 678928 40978 678992
rect 40910 678708 40970 678928
rect 41822 678330 41828 678332
rect 41492 678270 41828 678330
rect 41822 678268 41828 678270
rect 41892 678268 41898 678332
rect 45645 677922 45711 677925
rect 41492 677920 45711 677922
rect 41492 677864 45650 677920
rect 45706 677864 45711 677920
rect 41492 677862 45711 677864
rect 45645 677859 45711 677862
rect 41822 677588 41828 677652
rect 41892 677650 41898 677652
rect 42190 677650 42196 677652
rect 41892 677590 42196 677650
rect 41892 677588 41898 677590
rect 42190 677588 42196 677590
rect 42260 677588 42266 677652
rect 39990 677109 40050 677484
rect 41689 677378 41755 677381
rect 42701 677378 42767 677381
rect 41689 677376 42767 677378
rect 41689 677320 41694 677376
rect 41750 677320 42706 677376
rect 42762 677320 42767 677376
rect 41689 677318 42767 677320
rect 41689 677315 41755 677318
rect 42701 677315 42767 677318
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 47669 676698 47735 676701
rect 41492 676696 47735 676698
rect 41492 676640 47674 676696
rect 47730 676640 47735 676696
rect 41492 676638 47735 676640
rect 47669 676635 47735 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 661677 673162 661743 673165
rect 676489 673162 676555 673165
rect 661677 673160 676555 673162
rect 661677 673104 661682 673160
rect 661738 673104 676494 673160
rect 676550 673104 676555 673160
rect 661677 673102 676555 673104
rect 661677 673099 661743 673102
rect 676489 673099 676555 673102
rect 40125 671258 40191 671261
rect 40350 671258 40356 671260
rect 40125 671256 40356 671258
rect 40125 671200 40130 671256
rect 40186 671200 40356 671256
rect 40125 671198 40356 671200
rect 40125 671195 40191 671198
rect 40350 671196 40356 671198
rect 40420 671196 40426 671260
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 676489 671122 676555 671125
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 676446 671120 676555 671122
rect 676446 671064 676494 671120
rect 676550 671064 676555 671120
rect 667197 671059 667263 671062
rect 676446 671059 676555 671064
rect 36537 670986 36603 670989
rect 41822 670986 41828 670988
rect 36537 670984 41828 670986
rect 36537 670928 36542 670984
rect 36598 670928 41828 670984
rect 36537 670926 41828 670928
rect 36537 670923 36603 670926
rect 41822 670924 41828 670926
rect 41892 670924 41898 670988
rect 676446 670956 676506 671059
rect 651465 670442 651531 670445
rect 650164 670440 651531 670442
rect 650164 670384 651470 670440
rect 651526 670384 651531 670440
rect 650164 670382 651531 670384
rect 651465 670379 651531 670382
rect 668577 670442 668643 670445
rect 676262 670442 676322 670548
rect 668577 670440 676322 670442
rect 668577 670384 668582 670440
rect 668638 670384 676322 670440
rect 668577 670382 676322 670384
rect 668577 670379 668643 670382
rect 671613 670170 671679 670173
rect 671613 670168 676292 670170
rect 671613 670112 671618 670168
rect 671674 670112 676292 670168
rect 671613 670110 676292 670112
rect 671613 670107 671679 670110
rect 671429 669898 671495 669901
rect 676489 669898 676555 669901
rect 671429 669896 676555 669898
rect 671429 669840 671434 669896
rect 671490 669840 676494 669896
rect 676550 669840 676555 669896
rect 671429 669838 676555 669840
rect 671429 669835 671495 669838
rect 676489 669835 676555 669838
rect 671613 669490 671679 669493
rect 676262 669490 676322 669732
rect 676489 669490 676555 669493
rect 671613 669488 676322 669490
rect 671613 669432 671618 669488
rect 671674 669432 676322 669488
rect 671613 669430 676322 669432
rect 676446 669488 676555 669490
rect 676446 669432 676494 669488
rect 676550 669432 676555 669488
rect 671613 669427 671679 669430
rect 676446 669427 676555 669432
rect 42190 669292 42196 669356
rect 42260 669354 42266 669356
rect 48957 669354 49023 669357
rect 42260 669352 49023 669354
rect 42260 669296 48962 669352
rect 49018 669296 49023 669352
rect 676446 669324 676506 669427
rect 42260 669294 49023 669296
rect 42260 669292 42266 669294
rect 48957 669291 49023 669294
rect 671429 668674 671495 668677
rect 676262 668674 676322 668916
rect 671429 668672 676322 668674
rect 671429 668616 671434 668672
rect 671490 668616 676322 668672
rect 671429 668614 676322 668616
rect 671429 668611 671495 668614
rect 670877 668266 670943 668269
rect 676262 668266 676322 668508
rect 670877 668264 676322 668266
rect 670877 668208 670882 668264
rect 670938 668208 676322 668264
rect 670877 668206 676322 668208
rect 670877 668203 670943 668206
rect 670877 667994 670943 667997
rect 676262 667994 676322 668100
rect 670877 667992 676322 667994
rect 670877 667936 670882 667992
rect 670938 667936 676322 667992
rect 670877 667934 676322 667936
rect 670877 667931 670943 667934
rect 42241 667860 42307 667861
rect 42190 667796 42196 667860
rect 42260 667858 42307 667860
rect 42260 667856 42352 667858
rect 42302 667800 42352 667856
rect 42260 667798 42352 667800
rect 42260 667796 42307 667798
rect 42241 667795 42307 667796
rect 40350 667524 40356 667588
rect 40420 667586 40426 667588
rect 42425 667586 42491 667589
rect 40420 667584 42491 667586
rect 40420 667528 42430 667584
rect 42486 667528 42491 667584
rect 40420 667526 42491 667528
rect 40420 667524 40426 667526
rect 42425 667523 42491 667526
rect 674833 667450 674899 667453
rect 676262 667450 676322 667692
rect 674833 667448 676322 667450
rect 674833 667392 674838 667448
rect 674894 667392 676322 667448
rect 674833 667390 676322 667392
rect 674833 667387 674899 667390
rect 42241 667178 42307 667181
rect 42885 667178 42951 667181
rect 42241 667176 42951 667178
rect 42241 667120 42246 667176
rect 42302 667120 42890 667176
rect 42946 667120 42951 667176
rect 42241 667118 42951 667120
rect 42241 667115 42307 667118
rect 42885 667115 42951 667118
rect 40902 666980 40908 667044
rect 40972 667042 40978 667044
rect 42006 667042 42012 667044
rect 40972 666982 42012 667042
rect 40972 666980 40978 666982
rect 42006 666980 42012 666982
rect 42076 666980 42082 667044
rect 672625 667042 672691 667045
rect 676262 667042 676322 667284
rect 672625 667040 676322 667042
rect 672625 666984 672630 667040
rect 672686 666984 676322 667040
rect 672625 666982 676322 666984
rect 683205 667042 683271 667045
rect 683205 667040 683314 667042
rect 683205 666984 683210 667040
rect 683266 666984 683314 667040
rect 672625 666979 672691 666982
rect 683205 666979 683314 666984
rect 683254 666876 683314 666979
rect 44173 666634 44239 666637
rect 42198 666632 44239 666634
rect 42198 666576 44178 666632
rect 44234 666576 44239 666632
rect 42198 666574 44239 666576
rect 42198 666093 42258 666574
rect 44173 666571 44239 666574
rect 671061 666634 671127 666637
rect 674833 666634 674899 666637
rect 671061 666632 674899 666634
rect 671061 666576 671066 666632
rect 671122 666576 674838 666632
rect 674894 666576 674899 666632
rect 671061 666574 674899 666576
rect 671061 666571 671127 666574
rect 674833 666571 674899 666574
rect 669589 666362 669655 666365
rect 674414 666362 674420 666364
rect 669589 666360 674420 666362
rect 669589 666304 669594 666360
rect 669650 666304 674420 666360
rect 669589 666302 674420 666304
rect 669589 666299 669655 666302
rect 674414 666300 674420 666302
rect 674484 666300 674490 666364
rect 676262 666226 676322 666468
rect 674790 666166 676322 666226
rect 42198 666088 42307 666093
rect 42198 666032 42246 666088
rect 42302 666032 42307 666088
rect 42198 666030 42307 666032
rect 42241 666027 42307 666030
rect 671981 666090 672047 666093
rect 674790 666090 674850 666166
rect 671981 666088 674850 666090
rect 671981 666032 671986 666088
rect 672042 666032 674850 666088
rect 671981 666030 674850 666032
rect 671981 666027 672047 666030
rect 672257 665818 672323 665821
rect 673494 665818 673500 665820
rect 672257 665816 673500 665818
rect 672257 665760 672262 665816
rect 672318 665760 673500 665816
rect 672257 665758 673500 665760
rect 672257 665755 672323 665758
rect 673494 665756 673500 665758
rect 673564 665756 673570 665820
rect 676262 665818 676322 666060
rect 673870 665758 676322 665818
rect 673678 665620 673684 665684
rect 673748 665682 673754 665684
rect 673870 665682 673930 665758
rect 673748 665622 673930 665682
rect 673748 665620 673754 665622
rect 666277 665546 666343 665549
rect 666277 665544 673470 665546
rect 666277 665488 666282 665544
rect 666338 665488 673470 665544
rect 666277 665486 673470 665488
rect 666277 665483 666343 665486
rect 40718 665348 40724 665412
rect 40788 665410 40794 665412
rect 41781 665410 41847 665413
rect 40788 665408 41847 665410
rect 40788 665352 41786 665408
rect 41842 665352 41847 665408
rect 40788 665350 41847 665352
rect 673410 665410 673470 665486
rect 676262 665410 676322 665652
rect 673410 665350 676322 665410
rect 40788 665348 40794 665350
rect 41781 665347 41847 665350
rect 667841 665274 667907 665277
rect 667841 665272 673378 665274
rect 667841 665216 667846 665272
rect 667902 665216 673378 665272
rect 667841 665214 673378 665216
rect 667841 665211 667907 665214
rect 673318 665138 673378 665214
rect 673678 665138 673684 665140
rect 673318 665078 673684 665138
rect 673678 665076 673684 665078
rect 673748 665076 673754 665140
rect 674414 665076 674420 665140
rect 674484 665138 674490 665140
rect 676262 665138 676322 665244
rect 674484 665078 676322 665138
rect 674484 665076 674490 665078
rect 668761 664594 668827 664597
rect 676262 664594 676322 664836
rect 668761 664592 676322 664594
rect 668761 664536 668766 664592
rect 668822 664536 676322 664592
rect 668761 664534 676322 664536
rect 668761 664531 668827 664534
rect 673678 664260 673684 664324
rect 673748 664322 673754 664324
rect 676262 664322 676322 664428
rect 673748 664262 676322 664322
rect 673748 664260 673754 664262
rect 41965 664052 42031 664053
rect 41965 664048 42012 664052
rect 42076 664050 42082 664052
rect 41965 663992 41970 664048
rect 41965 663988 42012 663992
rect 42076 663990 42122 664050
rect 42076 663988 42082 663990
rect 41965 663987 42031 663988
rect 672073 663914 672139 663917
rect 676262 663914 676322 664020
rect 672073 663912 676322 663914
rect 672073 663856 672078 663912
rect 672134 663856 676322 663912
rect 672073 663854 676322 663856
rect 672073 663851 672139 663854
rect 42149 663506 42215 663509
rect 42885 663506 42951 663509
rect 42149 663504 42951 663506
rect 42149 663448 42154 663504
rect 42210 663448 42890 663504
rect 42946 663448 42951 663504
rect 42149 663446 42951 663448
rect 42149 663443 42215 663446
rect 42885 663443 42951 663446
rect 669405 663370 669471 663373
rect 676262 663370 676322 663612
rect 669405 663368 676322 663370
rect 669405 663312 669410 663368
rect 669466 663312 676322 663368
rect 669405 663310 676322 663312
rect 683389 663370 683455 663373
rect 683389 663368 683498 663370
rect 683389 663312 683394 663368
rect 683450 663312 683498 663368
rect 669405 663307 669471 663310
rect 683389 663307 683498 663312
rect 683438 663204 683498 663307
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 42241 662962 42307 662965
rect 44541 662962 44607 662965
rect 42241 662960 44607 662962
rect 42241 662904 42246 662960
rect 42302 662904 44546 662960
rect 44602 662904 44607 662960
rect 42241 662902 44607 662904
rect 42241 662899 42307 662902
rect 44541 662899 44607 662902
rect 40534 662628 40540 662692
rect 40604 662690 40610 662692
rect 42241 662690 42307 662693
rect 40604 662688 42307 662690
rect 40604 662632 42246 662688
rect 42302 662632 42307 662688
rect 40604 662630 42307 662632
rect 40604 662628 40610 662630
rect 42241 662627 42307 662630
rect 669037 662554 669103 662557
rect 676262 662554 676322 662796
rect 669037 662552 676322 662554
rect 669037 662496 669042 662552
rect 669098 662496 676322 662552
rect 669037 662494 676322 662496
rect 669037 662491 669103 662494
rect 674598 662220 674604 662284
rect 674668 662282 674674 662284
rect 676262 662282 676322 662388
rect 674668 662222 676322 662282
rect 674668 662220 674674 662222
rect 674833 661874 674899 661877
rect 676262 661874 676322 661980
rect 674833 661872 676322 661874
rect 674833 661816 674838 661872
rect 674894 661816 676322 661872
rect 674833 661814 676322 661816
rect 674833 661811 674899 661814
rect 673085 661602 673151 661605
rect 673085 661600 676292 661602
rect 673085 661544 673090 661600
rect 673146 661544 676292 661600
rect 673085 661542 676292 661544
rect 673085 661539 673151 661542
rect 671245 661330 671311 661333
rect 674833 661330 674899 661333
rect 671245 661328 674899 661330
rect 671245 661272 671250 661328
rect 671306 661272 674838 661328
rect 674894 661272 674899 661328
rect 671245 661270 674899 661272
rect 671245 661267 671311 661270
rect 674833 661267 674899 661270
rect 667841 661058 667907 661061
rect 676262 661058 676322 661164
rect 667841 661056 676322 661058
rect 667841 661000 667846 661056
rect 667902 661000 676322 661056
rect 667841 660998 676322 661000
rect 667841 660995 667907 660998
rect 675293 660242 675359 660245
rect 676262 660242 676322 660756
rect 675293 660240 676322 660242
rect 675293 660184 675298 660240
rect 675354 660184 676322 660240
rect 675293 660182 676322 660184
rect 675293 660179 675359 660182
rect 670601 659970 670667 659973
rect 670601 659968 676292 659970
rect 670601 659912 670606 659968
rect 670662 659912 676292 659968
rect 670601 659910 676292 659912
rect 670601 659907 670667 659910
rect 668393 659698 668459 659701
rect 675293 659698 675359 659701
rect 668393 659696 675359 659698
rect 668393 659640 668398 659696
rect 668454 659640 675298 659696
rect 675354 659640 675359 659696
rect 668393 659638 675359 659640
rect 668393 659635 668459 659638
rect 675293 659635 675359 659638
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42609 658610 42675 658613
rect 41708 658608 42675 658610
rect 41708 658552 42614 658608
rect 42670 658552 42675 658608
rect 41708 658550 42675 658552
rect 41708 658548 41714 658550
rect 42609 658547 42675 658550
rect 41822 658276 41828 658340
rect 41892 658338 41898 658340
rect 42425 658338 42491 658341
rect 41892 658336 42491 658338
rect 41892 658280 42430 658336
rect 42486 658280 42491 658336
rect 41892 658278 42491 658280
rect 41892 658276 41898 658278
rect 42425 658275 42491 658278
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 651465 657114 651531 657117
rect 650164 657112 651531 657114
rect 650164 657056 651470 657112
rect 651526 657056 651531 657112
rect 650164 657054 651531 657056
rect 651465 657051 651531 657054
rect 671981 654258 672047 654261
rect 675201 654258 675267 654261
rect 671981 654256 675267 654258
rect 671981 654200 671986 654256
rect 672042 654200 675206 654256
rect 675262 654200 675267 654256
rect 671981 654198 675267 654200
rect 671981 654195 672047 654198
rect 675201 654195 675267 654198
rect 675385 652900 675451 652901
rect 675334 652898 675340 652900
rect 675294 652838 675340 652898
rect 675404 652896 675451 652900
rect 675446 652840 675451 652896
rect 675334 652836 675340 652838
rect 675404 652836 675451 652840
rect 675385 652835 675451 652836
rect 675477 651540 675543 651541
rect 675477 651536 675524 651540
rect 675588 651538 675594 651540
rect 675477 651480 675482 651536
rect 675477 651476 675524 651480
rect 675588 651478 675634 651538
rect 675588 651476 675594 651478
rect 675477 651475 675543 651476
rect 674281 650314 674347 650317
rect 674238 650312 674347 650314
rect 674238 650256 674286 650312
rect 674342 650256 674347 650312
rect 674238 650251 674347 650256
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674238 649637 674298 650251
rect 674189 649632 674298 649637
rect 674189 649576 674194 649632
rect 674250 649576 674298 649632
rect 674189 649574 674298 649576
rect 674189 649571 674255 649574
rect 674230 648892 674236 648956
rect 674300 648954 674306 648956
rect 675385 648954 675451 648957
rect 674300 648952 675451 648954
rect 674300 648896 675390 648952
rect 675446 648896 675451 648952
rect 674300 648894 675451 648896
rect 674300 648892 674306 648894
rect 675385 648891 675451 648894
rect 673085 648682 673151 648685
rect 675109 648682 675175 648685
rect 673085 648680 675175 648682
rect 673085 648624 673090 648680
rect 673146 648624 675114 648680
rect 675170 648624 675175 648680
rect 673085 648622 675175 648624
rect 673085 648619 673151 648622
rect 675109 648619 675175 648622
rect 672809 647866 672875 647869
rect 675385 647866 675451 647869
rect 672809 647864 675451 647866
rect 672809 647808 672814 647864
rect 672870 647808 675390 647864
rect 675446 647808 675451 647864
rect 672809 647806 675451 647808
rect 672809 647803 672875 647806
rect 675385 647803 675451 647806
rect 668209 647322 668275 647325
rect 675109 647322 675175 647325
rect 668209 647320 675175 647322
rect 668209 647264 668214 647320
rect 668270 647264 675114 647320
rect 675170 647264 675175 647320
rect 668209 647262 675175 647264
rect 668209 647259 668275 647262
rect 675109 647259 675175 647262
rect 35801 646778 35867 646781
rect 35801 646776 35910 646778
rect 35801 646720 35806 646776
rect 35862 646720 35910 646776
rect 35801 646715 35910 646720
rect 35850 646642 35910 646715
rect 51717 646642 51783 646645
rect 35850 646640 51783 646642
rect 35850 646584 51722 646640
rect 51778 646584 51783 646640
rect 35850 646582 51783 646584
rect 51717 646579 51783 646582
rect 674189 645146 674255 645149
rect 674598 645146 674604 645148
rect 674189 645144 674604 645146
rect 674189 645088 674194 645144
rect 674250 645088 674604 645144
rect 674189 645086 674604 645088
rect 674189 645083 674255 645086
rect 674598 645084 674604 645086
rect 674668 645084 674674 645148
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 675753 644738 675819 644741
rect 676806 644738 676812 644740
rect 675753 644736 676812 644738
rect 675753 644680 675758 644736
rect 675814 644680 676812 644736
rect 675753 644678 676812 644680
rect 675753 644675 675819 644678
rect 676806 644676 676812 644678
rect 676876 644676 676882 644740
rect 35758 644504 35818 644675
rect 673821 644602 673887 644605
rect 675109 644602 675175 644605
rect 673821 644600 675175 644602
rect 673821 644544 673826 644600
rect 673882 644544 675114 644600
rect 675170 644544 675175 644600
rect 673821 644542 675175 644544
rect 673821 644539 673887 644542
rect 675109 644539 675175 644542
rect 41462 643922 41522 644096
rect 675109 643922 675175 643925
rect 41462 643862 45570 643922
rect 41462 643650 41522 643688
rect 44817 643650 44883 643653
rect 41462 643648 44883 643650
rect 41462 643592 44822 643648
rect 44878 643592 44883 643648
rect 41462 643590 44883 643592
rect 44817 643587 44883 643590
rect 44633 643378 44699 643381
rect 41462 643376 44699 643378
rect 41462 643320 44638 643376
rect 44694 643320 44699 643376
rect 41462 643318 44699 643320
rect 41462 643280 41522 643318
rect 44633 643315 44699 643318
rect 45510 643242 45570 643862
rect 663750 643920 675175 643922
rect 663750 643864 675114 643920
rect 675170 643864 675175 643920
rect 663750 643862 675175 643864
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 661677 643786 661743 643789
rect 663750 643786 663810 643862
rect 675109 643859 675175 643862
rect 661677 643784 663810 643786
rect 661677 643728 661682 643784
rect 661738 643728 663810 643784
rect 661677 643726 663810 643728
rect 661677 643723 661743 643726
rect 671889 643514 671955 643517
rect 675385 643514 675451 643517
rect 671889 643512 675451 643514
rect 671889 643456 671894 643512
rect 671950 643456 675390 643512
rect 675446 643456 675451 643512
rect 671889 643454 675451 643456
rect 671889 643451 671955 643454
rect 675385 643451 675451 643454
rect 55857 643242 55923 643245
rect 45510 643240 55923 643242
rect 45510 643184 55862 643240
rect 55918 643184 55923 643240
rect 45510 643182 55923 643184
rect 55857 643179 55923 643182
rect 45001 643106 45067 643109
rect 41462 643104 45067 643106
rect 41462 643048 45006 643104
rect 45062 643048 45067 643104
rect 41462 643046 45067 643048
rect 41462 642872 41522 643046
rect 45001 643043 45067 643046
rect 44817 642562 44883 642565
rect 41462 642560 44883 642562
rect 41462 642504 44822 642560
rect 44878 642504 44883 642560
rect 41462 642502 44883 642504
rect 41462 642464 41522 642502
rect 44817 642499 44883 642502
rect 44357 642290 44423 642293
rect 41462 642288 44423 642290
rect 41462 642232 44362 642288
rect 44418 642232 44423 642288
rect 41462 642230 44423 642232
rect 41462 642056 41522 642230
rect 44357 642227 44423 642230
rect 673637 641746 673703 641749
rect 675293 641746 675359 641749
rect 673637 641744 675359 641746
rect 673637 641688 673642 641744
rect 673698 641688 675298 641744
rect 675354 641688 675359 641744
rect 673637 641686 675359 641688
rect 673637 641683 673703 641686
rect 675293 641683 675359 641686
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 45369 641474 45435 641477
rect 41462 641472 45435 641474
rect 41462 641416 45374 641472
rect 45430 641416 45435 641472
rect 41462 641414 45435 641416
rect 41462 641240 41522 641414
rect 45369 641411 45435 641414
rect 41781 641202 41847 641205
rect 45185 641202 45251 641205
rect 41781 641200 45251 641202
rect 41781 641144 41786 641200
rect 41842 641144 45190 641200
rect 45246 641144 45251 641200
rect 41781 641142 45251 641144
rect 41781 641139 41847 641142
rect 45185 641139 45251 641142
rect 45001 640930 45067 640933
rect 41462 640928 45067 640930
rect 41462 640872 45006 640928
rect 45062 640872 45067 640928
rect 41462 640870 45067 640872
rect 41462 640832 41522 640870
rect 45001 640867 45067 640870
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 675150 640460 675156 640524
rect 675220 640522 675226 640524
rect 675385 640522 675451 640525
rect 675220 640520 675451 640522
rect 675220 640464 675390 640520
rect 675446 640464 675451 640520
rect 675220 640462 675451 640464
rect 675220 640460 675226 640462
rect 675385 640459 675451 640462
rect 35574 639845 35634 640016
rect 35574 639840 35683 639845
rect 35574 639784 35622 639840
rect 35678 639784 35683 639840
rect 35574 639782 35683 639784
rect 35617 639779 35683 639782
rect 35758 639437 35818 639608
rect 35758 639432 35867 639437
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35758 639374 35867 639376
rect 35801 639371 35867 639374
rect 41822 639230 41828 639232
rect 41492 639170 41828 639230
rect 41822 639168 41828 639170
rect 41892 639168 41898 639232
rect 35758 638621 35818 638792
rect 668945 638754 669011 638757
rect 675477 638754 675543 638757
rect 668945 638752 675543 638754
rect 668945 638696 668950 638752
rect 669006 638696 675482 638752
rect 675538 638696 675543 638752
rect 668945 638694 675543 638696
rect 668945 638691 669011 638694
rect 675477 638691 675543 638694
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 40033 638618 40099 638621
rect 41638 638618 41644 638620
rect 40033 638616 41644 638618
rect 40033 638560 40038 638616
rect 40094 638560 41644 638616
rect 40033 638558 41644 638560
rect 40033 638555 40099 638558
rect 41638 638556 41644 638558
rect 41708 638556 41714 638620
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 41781 638210 41847 638213
rect 47209 638210 47275 638213
rect 41781 638208 47275 638210
rect 41781 638152 41786 638208
rect 41842 638152 47214 638208
rect 47270 638152 47275 638208
rect 41781 638150 47275 638152
rect 32397 638147 32463 638150
rect 41781 638147 41847 638150
rect 47209 638147 47275 638150
rect 675334 638012 675340 638076
rect 675404 638074 675410 638076
rect 675753 638074 675819 638077
rect 675404 638072 675819 638074
rect 675404 638016 675758 638072
rect 675814 638016 675819 638072
rect 675404 638014 675819 638016
rect 675404 638012 675410 638014
rect 675753 638011 675819 638014
rect 41462 637802 41522 637976
rect 45829 637802 45895 637805
rect 675569 637804 675635 637805
rect 41462 637800 45895 637802
rect 41462 637744 45834 637800
rect 45890 637744 45895 637800
rect 41462 637742 45895 637744
rect 45829 637739 45895 637742
rect 675518 637740 675524 637804
rect 675588 637802 675635 637804
rect 675588 637800 675680 637802
rect 675630 637744 675680 637800
rect 675588 637742 675680 637744
rect 675588 637740 675635 637742
rect 675569 637739 675635 637740
rect 675201 637668 675267 637669
rect 675150 637604 675156 637668
rect 675220 637666 675267 637668
rect 675220 637664 675312 637666
rect 675262 637608 675312 637664
rect 675220 637606 675312 637608
rect 675220 637604 675267 637606
rect 675201 637603 675267 637604
rect 41781 637598 41847 637601
rect 41492 637596 41847 637598
rect 41492 637540 41786 637596
rect 41842 637540 41847 637596
rect 41492 637538 41847 637540
rect 41781 637535 41847 637538
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 46381 636986 46447 636989
rect 41462 636984 46447 636986
rect 41462 636928 46386 636984
rect 46442 636928 46447 636984
rect 41462 636926 46447 636928
rect 46381 636923 46447 636926
rect 673453 636850 673519 636853
rect 683389 636850 683455 636853
rect 673453 636848 683455 636850
rect 673453 636792 673458 636848
rect 673514 636792 683394 636848
rect 683450 636792 683455 636848
rect 673453 636790 683455 636792
rect 673453 636787 673519 636790
rect 683389 636787 683455 636790
rect 35758 636581 35818 636752
rect 35758 636576 35867 636581
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35758 636518 35867 636520
rect 35801 636515 35867 636518
rect 47393 636442 47459 636445
rect 41462 636440 47459 636442
rect 41462 636384 47398 636440
rect 47454 636384 47459 636440
rect 41462 636382 47459 636384
rect 41462 636344 41522 636382
rect 47393 636379 47459 636382
rect 41462 635762 41522 635936
rect 42793 635762 42859 635765
rect 41462 635760 42859 635762
rect 41462 635704 42798 635760
rect 42854 635704 42859 635760
rect 41462 635702 42859 635704
rect 42793 635699 42859 635702
rect 674189 635762 674255 635765
rect 683573 635762 683639 635765
rect 674189 635760 683639 635762
rect 674189 635704 674194 635760
rect 674250 635704 683578 635760
rect 683634 635704 683639 635760
rect 674189 635702 683639 635704
rect 674189 635699 674255 635702
rect 683573 635699 683639 635702
rect 41462 635354 41522 635528
rect 672625 635490 672691 635493
rect 683757 635490 683823 635493
rect 672625 635488 683823 635490
rect 672625 635432 672630 635488
rect 672686 635432 683762 635488
rect 683818 635432 683823 635488
rect 672625 635430 683823 635432
rect 672625 635427 672691 635430
rect 683757 635427 683823 635430
rect 44173 635354 44239 635357
rect 41462 635352 44239 635354
rect 41462 635296 44178 635352
rect 44234 635296 44239 635352
rect 41462 635294 44239 635296
rect 44173 635291 44239 635294
rect 40542 634948 40602 635120
rect 40534 634884 40540 634948
rect 40604 634884 40610 634948
rect 41462 634538 41522 634712
rect 44357 634538 44423 634541
rect 41462 634536 44423 634538
rect 41462 634480 44362 634536
rect 44418 634480 44423 634536
rect 41462 634478 44423 634480
rect 44357 634475 44423 634478
rect 41462 633858 41522 634304
rect 42241 633858 42307 633861
rect 41462 633856 42307 633858
rect 41462 633800 42246 633856
rect 42302 633800 42307 633856
rect 41462 633798 42307 633800
rect 42241 633795 42307 633798
rect 41462 633450 41522 633488
rect 43437 633450 43503 633453
rect 41462 633448 43503 633450
rect 41462 633392 43442 633448
rect 43498 633392 43503 633448
rect 41462 633390 43503 633392
rect 43437 633387 43503 633390
rect 675150 632980 675156 633044
rect 675220 633042 675226 633044
rect 675569 633042 675635 633045
rect 675220 633040 675635 633042
rect 675220 632984 675574 633040
rect 675630 632984 675635 633040
rect 675220 632982 675635 632984
rect 675220 632980 675226 632982
rect 675569 632979 675635 632982
rect 675753 631410 675819 631413
rect 676070 631410 676076 631412
rect 675753 631408 676076 631410
rect 675753 631352 675758 631408
rect 675814 631352 676076 631408
rect 675753 631350 676076 631352
rect 675753 631347 675819 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 651465 630594 651531 630597
rect 650164 630592 651531 630594
rect 650164 630536 651470 630592
rect 651526 630536 651531 630592
rect 650164 630534 651531 630536
rect 651465 630531 651531 630534
rect 674925 629778 674991 629781
rect 675518 629778 675524 629780
rect 674925 629776 675524 629778
rect 674925 629720 674930 629776
rect 674986 629720 675524 629776
rect 674925 629718 675524 629720
rect 674925 629715 674991 629718
rect 675518 629716 675524 629718
rect 675588 629716 675594 629780
rect 652017 627874 652083 627877
rect 675845 627874 675911 627877
rect 652017 627872 675911 627874
rect 652017 627816 652022 627872
rect 652078 627816 675850 627872
rect 675906 627816 675911 627872
rect 652017 627814 675911 627816
rect 652017 627811 652083 627814
rect 675845 627811 675911 627814
rect 42006 626588 42012 626652
rect 42076 626650 42082 626652
rect 50337 626650 50403 626653
rect 42076 626648 50403 626650
rect 42076 626592 50342 626648
rect 50398 626592 50403 626648
rect 42076 626590 50403 626592
rect 42076 626588 42082 626590
rect 50337 626587 50403 626590
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 669270 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 671613 625154 671679 625157
rect 671613 625152 676292 625154
rect 671613 625096 671618 625152
rect 671674 625096 676292 625152
rect 671613 625094 676292 625096
rect 671613 625091 671679 625094
rect 42241 625020 42307 625021
rect 42190 625018 42196 625020
rect 42150 624958 42196 625018
rect 42260 625016 42307 625020
rect 42302 624960 42307 625016
rect 42190 624956 42196 624958
rect 42260 624956 42307 624960
rect 42241 624955 42307 624956
rect 671061 624746 671127 624749
rect 671061 624744 676292 624746
rect 671061 624688 671066 624744
rect 671122 624688 676292 624744
rect 671061 624686 676292 624688
rect 671061 624683 671127 624686
rect 42057 624476 42123 624477
rect 42006 624412 42012 624476
rect 42076 624474 42123 624476
rect 42076 624472 42168 624474
rect 42118 624416 42168 624472
rect 42076 624414 42168 624416
rect 42076 624412 42123 624414
rect 42057 624411 42123 624412
rect 671245 624338 671311 624341
rect 671245 624336 676292 624338
rect 671245 624280 671250 624336
rect 671306 624280 676292 624336
rect 671245 624278 676292 624280
rect 671245 624275 671311 624278
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 672257 623930 672323 623933
rect 672257 623928 676292 623930
rect 672257 623872 672262 623928
rect 672318 623872 676292 623928
rect 672257 623870 676292 623872
rect 672257 623867 672323 623870
rect 670877 623522 670943 623525
rect 670877 623520 676292 623522
rect 670877 623464 670882 623520
rect 670938 623464 676292 623520
rect 670877 623462 676292 623464
rect 670877 623459 670943 623462
rect 674465 623250 674531 623253
rect 683113 623250 683179 623253
rect 674465 623248 683179 623250
rect 674465 623192 674470 623248
rect 674526 623192 683118 623248
rect 683174 623192 683179 623248
rect 674465 623190 683179 623192
rect 674465 623187 674531 623190
rect 683113 623187 683179 623190
rect 670877 622842 670943 622845
rect 676262 622842 676322 623084
rect 670877 622840 676322 622842
rect 670877 622784 670882 622840
rect 670938 622784 676322 622840
rect 670877 622782 676322 622784
rect 683757 622842 683823 622845
rect 683757 622840 683866 622842
rect 683757 622784 683762 622840
rect 683818 622784 683866 622840
rect 670877 622779 670943 622782
rect 683757 622779 683866 622784
rect 683806 622676 683866 622779
rect 671613 622434 671679 622437
rect 671613 622432 674666 622434
rect 671613 622376 671618 622432
rect 671674 622376 674666 622432
rect 671613 622374 674666 622376
rect 671613 622371 671679 622374
rect 674606 622298 674666 622374
rect 674606 622238 676292 622298
rect 40534 622100 40540 622164
rect 40604 622162 40610 622164
rect 41781 622162 41847 622165
rect 674465 622162 674531 622165
rect 40604 622160 41847 622162
rect 40604 622104 41786 622160
rect 41842 622104 41847 622160
rect 40604 622102 41847 622104
rect 40604 622100 40610 622102
rect 41781 622099 41847 622102
rect 669270 622160 674531 622162
rect 669270 622104 674470 622160
rect 674526 622104 674531 622160
rect 669270 622102 674531 622104
rect 669270 622029 669330 622102
rect 674465 622099 674531 622102
rect 669221 622024 669330 622029
rect 669221 621968 669226 622024
rect 669282 621968 669330 622024
rect 669221 621966 669330 621968
rect 669221 621963 669287 621966
rect 672625 621890 672691 621893
rect 672625 621888 676292 621890
rect 672625 621832 672630 621888
rect 672686 621832 676292 621888
rect 672625 621830 676292 621832
rect 672625 621827 672691 621830
rect 668025 621754 668091 621757
rect 668025 621752 669330 621754
rect 668025 621696 668030 621752
rect 668086 621696 669330 621752
rect 668025 621694 669330 621696
rect 668025 621691 668091 621694
rect 42149 621618 42215 621621
rect 47393 621618 47459 621621
rect 42149 621616 47459 621618
rect 42149 621560 42154 621616
rect 42210 621560 47398 621616
rect 47454 621560 47459 621616
rect 42149 621558 47459 621560
rect 669270 621618 669330 621694
rect 669270 621558 676322 621618
rect 42149 621555 42215 621558
rect 47393 621555 47459 621558
rect 676262 621452 676322 621558
rect 666461 621210 666527 621213
rect 672625 621210 672691 621213
rect 666461 621208 672691 621210
rect 666461 621152 666466 621208
rect 666522 621152 672630 621208
rect 672686 621152 672691 621208
rect 666461 621150 672691 621152
rect 666461 621147 666527 621150
rect 672625 621147 672691 621150
rect 675158 621150 676322 621210
rect 674465 620938 674531 620941
rect 675158 620938 675218 621150
rect 676262 621044 676322 621150
rect 674465 620936 675218 620938
rect 674465 620880 674470 620936
rect 674526 620880 675218 620936
rect 674465 620878 675218 620880
rect 674465 620875 674531 620878
rect 42057 620802 42123 620805
rect 44173 620802 44239 620805
rect 42057 620800 44239 620802
rect 42057 620744 42062 620800
rect 42118 620744 44178 620800
rect 44234 620744 44239 620800
rect 42057 620742 44239 620744
rect 42057 620739 42123 620742
rect 44173 620739 44239 620742
rect 669773 620666 669839 620669
rect 669773 620664 676292 620666
rect 669773 620608 669778 620664
rect 669834 620608 676292 620664
rect 669773 620606 676292 620608
rect 669773 620603 669839 620606
rect 41965 620258 42031 620261
rect 42190 620258 42196 620260
rect 41965 620256 42196 620258
rect 41965 620200 41970 620256
rect 42026 620200 42196 620256
rect 41965 620198 42196 620200
rect 41965 620195 42031 620198
rect 42190 620196 42196 620198
rect 42260 620196 42266 620260
rect 670417 620258 670483 620261
rect 670417 620256 676292 620258
rect 670417 620200 670422 620256
rect 670478 620200 676292 620256
rect 670417 620198 676292 620200
rect 670417 620195 670483 620198
rect 672441 619850 672507 619853
rect 672441 619848 676292 619850
rect 672441 619792 672446 619848
rect 672502 619792 676292 619848
rect 672441 619790 676292 619792
rect 672441 619787 672507 619790
rect 674281 619442 674347 619445
rect 674281 619440 676292 619442
rect 674281 619384 674286 619440
rect 674342 619384 676292 619440
rect 674281 619382 676292 619384
rect 674281 619379 674347 619382
rect 42425 619306 42491 619309
rect 46381 619306 46447 619309
rect 42425 619304 46447 619306
rect 42425 619248 42430 619304
rect 42486 619248 46386 619304
rect 46442 619248 46447 619304
rect 42425 619246 46447 619248
rect 42425 619243 42491 619246
rect 46381 619243 46447 619246
rect 676990 619108 676996 619172
rect 677060 619108 677066 619172
rect 42609 619034 42675 619037
rect 47209 619034 47275 619037
rect 42609 619032 47275 619034
rect 42609 618976 42614 619032
rect 42670 618976 47214 619032
rect 47270 618976 47275 619032
rect 676998 619004 677058 619108
rect 42609 618974 47275 618976
rect 42609 618971 42675 618974
rect 47209 618971 47275 618974
rect 683573 618762 683639 618765
rect 683573 618760 683682 618762
rect 683573 618704 683578 618760
rect 683634 618704 683682 618760
rect 683573 618699 683682 618704
rect 683622 618596 683682 618699
rect 671429 618218 671495 618221
rect 671429 618216 676292 618218
rect 671429 618160 671434 618216
rect 671490 618160 676292 618216
rect 671429 618158 676292 618160
rect 671429 618155 671495 618158
rect 683113 617946 683179 617949
rect 682886 617944 683179 617946
rect 682886 617888 683118 617944
rect 683174 617888 683179 617944
rect 682886 617886 683179 617888
rect 682886 617780 682946 617886
rect 683113 617883 683179 617886
rect 674005 617402 674071 617405
rect 674005 617400 676292 617402
rect 674005 617344 674010 617400
rect 674066 617344 676292 617400
rect 674005 617342 676292 617344
rect 674005 617339 674071 617342
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683389 617130 683455 617133
rect 683389 617128 683498 617130
rect 683389 617072 683394 617128
rect 683450 617072 683498 617128
rect 683389 617067 683498 617072
rect 683438 616964 683498 617067
rect 673269 616586 673335 616589
rect 673269 616584 676292 616586
rect 673269 616528 673274 616584
rect 673330 616528 676292 616584
rect 673269 616526 676292 616528
rect 673269 616523 673335 616526
rect 669773 616178 669839 616181
rect 669773 616176 676292 616178
rect 669773 616120 669778 616176
rect 669834 616120 676292 616176
rect 669773 616118 676292 616120
rect 669773 616115 669839 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 42241 616042 42307 616045
rect 41524 616040 42307 616042
rect 41524 615984 42246 616040
rect 42302 615984 42307 616040
rect 41524 615982 42307 615984
rect 41524 615980 41530 615982
rect 42241 615979 42307 615982
rect 41781 615772 41847 615773
rect 41781 615768 41828 615772
rect 41892 615770 41898 615772
rect 670233 615770 670299 615773
rect 41781 615712 41786 615768
rect 41781 615708 41828 615712
rect 41892 615710 41938 615770
rect 670233 615768 676292 615770
rect 670233 615712 670238 615768
rect 670294 615740 676292 615768
rect 670294 615712 676322 615740
rect 670233 615710 676322 615712
rect 41892 615708 41898 615710
rect 41781 615707 41847 615708
rect 670233 615707 670299 615710
rect 42885 615634 42951 615637
rect 45829 615634 45895 615637
rect 42885 615632 45895 615634
rect 42885 615576 42890 615632
rect 42946 615576 45834 615632
rect 45890 615576 45895 615632
rect 42885 615574 45895 615576
rect 42885 615571 42951 615574
rect 45829 615571 45895 615574
rect 676262 615332 676322 615710
rect 670417 614954 670483 614957
rect 670417 614952 676292 614954
rect 670417 614896 670422 614952
rect 670478 614896 676292 614952
rect 670417 614894 676292 614896
rect 670417 614891 670483 614894
rect 44173 614138 44239 614141
rect 47761 614138 47827 614141
rect 44173 614136 47827 614138
rect 44173 614080 44178 614136
rect 44234 614080 47766 614136
rect 47822 614080 47827 614136
rect 44173 614078 47827 614080
rect 44173 614075 44239 614078
rect 47761 614075 47827 614078
rect 41781 612780 41847 612781
rect 41781 612776 41828 612780
rect 41892 612778 41898 612780
rect 41781 612720 41786 612776
rect 41781 612716 41828 612720
rect 41892 612718 41938 612778
rect 41892 612716 41898 612718
rect 41781 612715 41847 612716
rect 43069 612370 43135 612373
rect 43713 612370 43779 612373
rect 43069 612368 43779 612370
rect 43069 612312 43074 612368
rect 43130 612312 43718 612368
rect 43774 612312 43779 612368
rect 43069 612310 43779 612312
rect 43069 612307 43135 612310
rect 43713 612307 43779 612310
rect 44265 611010 44331 611013
rect 45645 611010 45711 611013
rect 44265 611008 45711 611010
rect 44265 610952 44270 611008
rect 44326 610952 45650 611008
rect 45706 610952 45711 611008
rect 44265 610950 45711 610952
rect 44265 610947 44331 610950
rect 45645 610947 45711 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 666461 608834 666527 608837
rect 674833 608834 674899 608837
rect 666461 608832 674899 608834
rect 666461 608776 666466 608832
rect 666522 608776 674838 608832
rect 674894 608776 674899 608832
rect 666461 608774 674899 608776
rect 666461 608771 666527 608774
rect 674833 608771 674899 608774
rect 669221 608562 669287 608565
rect 675017 608562 675083 608565
rect 669221 608560 675083 608562
rect 669221 608504 669226 608560
rect 669282 608504 675022 608560
rect 675078 608504 675083 608560
rect 669221 608502 675083 608504
rect 669221 608499 669287 608502
rect 675017 608499 675083 608502
rect 668393 608018 668459 608021
rect 675477 608018 675543 608021
rect 668393 608016 675543 608018
rect 668393 607960 668398 608016
rect 668454 607960 675482 608016
rect 675538 607960 675543 608016
rect 668393 607958 675543 607960
rect 668393 607955 668459 607958
rect 675477 607955 675543 607958
rect 675017 607746 675083 607749
rect 675477 607746 675543 607749
rect 675017 607744 675543 607746
rect 675017 607688 675022 607744
rect 675078 607688 675482 607744
rect 675538 607688 675543 607744
rect 675017 607686 675543 607688
rect 675017 607683 675083 607686
rect 675477 607683 675543 607686
rect 674833 607202 674899 607205
rect 675477 607202 675543 607205
rect 674833 607200 675543 607202
rect 674833 607144 674838 607200
rect 674894 607144 675482 607200
rect 675538 607144 675543 607200
rect 674833 607142 675543 607144
rect 674833 607139 674899 607142
rect 675477 607139 675543 607142
rect 674649 604618 674715 604621
rect 675477 604618 675543 604621
rect 674649 604616 675543 604618
rect 674649 604560 674654 604616
rect 674710 604560 675482 604616
rect 675538 604560 675543 604616
rect 674649 604558 675543 604560
rect 674649 604555 674715 604558
rect 675477 604555 675543 604558
rect 673361 604346 673427 604349
rect 675477 604346 675543 604349
rect 673361 604344 675543 604346
rect 673361 604288 673366 604344
rect 673422 604288 675482 604344
rect 675538 604288 675543 604344
rect 673361 604286 675543 604288
rect 673361 604283 673427 604286
rect 675477 604283 675543 604286
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 674005 603530 674071 603533
rect 675477 603530 675543 603533
rect 674005 603528 675543 603530
rect 674005 603472 674010 603528
rect 674066 603472 675482 603528
rect 675538 603472 675543 603528
rect 674005 603470 675543 603472
rect 674005 603467 674071 603470
rect 675477 603467 675543 603470
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675477 602986 675543 602989
rect 674484 602984 675543 602986
rect 674484 602928 675482 602984
rect 675538 602928 675543 602984
rect 674484 602926 675543 602928
rect 674484 602924 674490 602926
rect 675477 602923 675543 602926
rect 674833 602306 674899 602309
rect 675385 602306 675451 602309
rect 674833 602304 675451 602306
rect 674833 602248 674838 602304
rect 674894 602248 675390 602304
rect 675446 602248 675451 602304
rect 674833 602246 675451 602248
rect 674833 602243 674899 602246
rect 675385 602243 675451 602246
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 50337 601354 50403 601357
rect 41492 601352 50403 601354
rect 41492 601296 50342 601352
rect 50398 601296 50403 601352
rect 41492 601294 50403 601296
rect 50337 601291 50403 601294
rect 46197 600946 46263 600949
rect 41492 600944 46263 600946
rect 41492 600888 46202 600944
rect 46258 600888 46263 600944
rect 41492 600886 46263 600888
rect 46197 600883 46263 600886
rect 670233 600674 670299 600677
rect 675109 600674 675175 600677
rect 670233 600672 675175 600674
rect 670233 600616 670238 600672
rect 670294 600616 675114 600672
rect 675170 600616 675175 600672
rect 670233 600614 675175 600616
rect 670233 600611 670299 600614
rect 675109 600611 675175 600614
rect 44633 600538 44699 600541
rect 41492 600536 44699 600538
rect 41492 600480 44638 600536
rect 44694 600480 44699 600536
rect 41492 600478 44699 600480
rect 44633 600475 44699 600478
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 674281 600130 674347 600133
rect 675109 600130 675175 600133
rect 674281 600128 675175 600130
rect 674281 600072 674286 600128
rect 674342 600072 675114 600128
rect 675170 600072 675175 600128
rect 674281 600070 675175 600072
rect 674281 600067 674347 600070
rect 675109 600067 675175 600070
rect 44817 599722 44883 599725
rect 41492 599720 44883 599722
rect 41492 599664 44822 599720
rect 44878 599664 44883 599720
rect 41492 599662 44883 599664
rect 44817 599659 44883 599662
rect 660297 599586 660363 599589
rect 675109 599586 675175 599589
rect 660297 599584 675175 599586
rect 660297 599528 660302 599584
rect 660358 599528 675114 599584
rect 675170 599528 675175 599584
rect 660297 599526 675175 599528
rect 660297 599523 660363 599526
rect 675109 599523 675175 599526
rect 44817 599314 44883 599317
rect 41492 599312 44883 599314
rect 41492 599256 44822 599312
rect 44878 599256 44883 599312
rect 41492 599254 44883 599256
rect 44817 599251 44883 599254
rect 674465 599042 674531 599045
rect 675293 599042 675359 599045
rect 674465 599040 675359 599042
rect 674465 598984 674470 599040
rect 674526 598984 675298 599040
rect 675354 598984 675359 599040
rect 674465 598982 675359 598984
rect 674465 598979 674531 598982
rect 675293 598979 675359 598982
rect 45185 598906 45251 598909
rect 41492 598904 45251 598906
rect 41492 598848 45190 598904
rect 45246 598848 45251 598904
rect 41492 598846 45251 598848
rect 45185 598843 45251 598846
rect 45185 598498 45251 598501
rect 41492 598496 45251 598498
rect 41492 598440 45190 598496
rect 45246 598440 45251 598496
rect 41492 598438 45251 598440
rect 45185 598435 45251 598438
rect 673453 598498 673519 598501
rect 675477 598498 675543 598501
rect 673453 598496 675543 598498
rect 673453 598440 673458 598496
rect 673514 598440 675482 598496
rect 675538 598440 675543 598496
rect 673453 598438 675543 598440
rect 673453 598435 673519 598438
rect 675477 598435 675543 598438
rect 45001 598090 45067 598093
rect 41492 598088 45067 598090
rect 41492 598032 45006 598088
rect 45062 598032 45067 598088
rect 41492 598030 45067 598032
rect 45001 598027 45067 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41492 597622 42994 597682
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 42934 597005 42994 597622
rect 672625 597410 672691 597413
rect 675385 597410 675451 597413
rect 672625 597408 675451 597410
rect 672625 597352 672630 597408
rect 672686 597352 675390 597408
rect 675446 597352 675451 597408
rect 672625 597350 675451 597352
rect 672625 597347 672691 597350
rect 675385 597347 675451 597350
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 42425 596866 42491 596869
rect 41492 596864 42491 596866
rect 41492 596808 42430 596864
rect 42486 596808 42491 596864
rect 41492 596806 42491 596808
rect 42425 596803 42491 596806
rect 674925 596730 674991 596733
rect 675702 596730 675708 596732
rect 674925 596728 675708 596730
rect 674925 596672 674930 596728
rect 674986 596672 675708 596728
rect 674925 596670 675708 596672
rect 674925 596667 674991 596670
rect 675702 596668 675708 596670
rect 675772 596668 675778 596732
rect 41822 596458 41828 596460
rect 41492 596398 41828 596458
rect 41822 596396 41828 596398
rect 41892 596396 41898 596460
rect 41229 596050 41295 596053
rect 41229 596048 41308 596050
rect 41229 595992 41234 596048
rect 41290 595992 41308 596048
rect 41229 595990 41308 595992
rect 41229 595987 41295 595990
rect 33777 595642 33843 595645
rect 33764 595640 33843 595642
rect 33764 595584 33782 595640
rect 33838 595584 33843 595640
rect 33764 595582 33843 595584
rect 33777 595579 33843 595582
rect 36537 595234 36603 595237
rect 36524 595232 36603 595234
rect 36524 595176 36542 595232
rect 36598 595176 36603 595232
rect 36524 595174 36603 595176
rect 36537 595171 36603 595174
rect 32397 594826 32463 594829
rect 671061 594826 671127 594829
rect 675293 594826 675359 594829
rect 32397 594824 32476 594826
rect 32397 594768 32402 594824
rect 32458 594768 32476 594824
rect 32397 594766 32476 594768
rect 671061 594824 675359 594826
rect 671061 594768 671066 594824
rect 671122 594768 675298 594824
rect 675354 594768 675359 594824
rect 671061 594766 675359 594768
rect 32397 594763 32463 594766
rect 671061 594763 671127 594766
rect 675293 594763 675359 594766
rect 37917 594418 37983 594421
rect 674925 594418 674991 594421
rect 37917 594416 37996 594418
rect 37917 594360 37922 594416
rect 37978 594360 37996 594416
rect 37917 594358 37996 594360
rect 674925 594416 676230 594418
rect 674925 594360 674930 594416
rect 674986 594360 676230 594416
rect 674925 594358 676230 594360
rect 37917 594355 37983 594358
rect 674925 594355 674991 594358
rect 676170 594146 676230 594358
rect 676990 594146 676996 594148
rect 676170 594086 676996 594146
rect 676990 594084 676996 594086
rect 677060 594084 677066 594148
rect 42793 594010 42859 594013
rect 41492 594008 42859 594010
rect 41492 593952 42798 594008
rect 42854 593952 42859 594008
rect 41492 593950 42859 593952
rect 42793 593947 42859 593950
rect 675017 593874 675083 593877
rect 675518 593874 675524 593876
rect 675017 593872 675524 593874
rect 675017 593816 675022 593872
rect 675078 593816 675524 593872
rect 675017 593814 675524 593816
rect 675017 593811 675083 593814
rect 675518 593812 675524 593814
rect 675588 593812 675594 593876
rect 40677 593602 40743 593605
rect 668761 593602 668827 593605
rect 675385 593602 675451 593605
rect 40677 593600 40756 593602
rect 40677 593544 40682 593600
rect 40738 593544 40756 593600
rect 40677 593542 40756 593544
rect 668761 593600 675451 593602
rect 668761 593544 668766 593600
rect 668822 593544 675390 593600
rect 675446 593544 675451 593600
rect 668761 593542 675451 593544
rect 40677 593539 40743 593542
rect 668761 593539 668827 593542
rect 675385 593539 675451 593542
rect 42057 593194 42123 593197
rect 41492 593192 42123 593194
rect 41492 593136 42062 593192
rect 42118 593136 42123 593192
rect 41492 593134 42123 593136
rect 42057 593131 42123 593134
rect 673637 593194 673703 593197
rect 673637 593192 676138 593194
rect 673637 593136 673642 593192
rect 673698 593136 676138 593192
rect 673637 593134 676138 593136
rect 673637 593131 673703 593134
rect 675150 592860 675156 592924
rect 675220 592922 675226 592924
rect 675845 592922 675911 592925
rect 675220 592920 675911 592922
rect 675220 592864 675850 592920
rect 675906 592864 675911 592920
rect 675220 592862 675911 592864
rect 676078 592922 676138 593134
rect 683481 592922 683547 592925
rect 676078 592920 683547 592922
rect 676078 592864 683486 592920
rect 683542 592864 683547 592920
rect 676078 592862 683547 592864
rect 675220 592860 675226 592862
rect 675845 592859 675911 592862
rect 683481 592859 683547 592862
rect 41873 592786 41939 592789
rect 41492 592784 41939 592786
rect 41492 592728 41878 592784
rect 41934 592728 41939 592784
rect 41492 592726 41939 592728
rect 41873 592723 41939 592726
rect 674230 592588 674236 592652
rect 674300 592650 674306 592652
rect 683297 592650 683363 592653
rect 674300 592648 683363 592650
rect 674300 592592 683302 592648
rect 683358 592592 683363 592648
rect 674300 592590 683363 592592
rect 674300 592588 674306 592590
rect 683297 592587 683363 592590
rect 41822 592378 41828 592380
rect 41492 592318 41828 592378
rect 41822 592316 41828 592318
rect 41892 592316 41898 592380
rect 675702 592316 675708 592380
rect 675772 592378 675778 592380
rect 676029 592378 676095 592381
rect 675772 592376 676095 592378
rect 675772 592320 676034 592376
rect 676090 592320 676095 592376
rect 675772 592318 676095 592320
rect 675772 592316 675778 592318
rect 676029 592315 676095 592318
rect 44449 591970 44515 591973
rect 41492 591968 44515 591970
rect 41492 591912 44454 591968
rect 44510 591912 44515 591968
rect 41492 591910 44515 591912
rect 44449 591907 44515 591910
rect 43846 591562 43852 591564
rect 41492 591502 43852 591562
rect 43846 591500 43852 591502
rect 43916 591500 43922 591564
rect 673821 591290 673887 591293
rect 683113 591290 683179 591293
rect 673821 591288 683179 591290
rect 673821 591232 673826 591288
rect 673882 591232 683118 591288
rect 683174 591232 683179 591288
rect 673821 591230 683179 591232
rect 673821 591227 673887 591230
rect 683113 591227 683179 591230
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 652385 590746 652451 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 652451 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 652390 590744
rect 652446 590688 652451 590744
rect 650164 590686 652451 590688
rect 39941 590683 40007 590686
rect 652385 590683 652451 590686
rect 676070 590548 676076 590612
rect 676140 590610 676146 590612
rect 680997 590610 681063 590613
rect 676140 590608 681063 590610
rect 676140 590552 681002 590608
rect 681058 590552 681063 590608
rect 676140 590550 681063 590552
rect 676140 590548 676146 590550
rect 680997 590547 681063 590550
rect 43437 590338 43503 590341
rect 41492 590336 43503 590338
rect 41492 590280 43442 590336
rect 43498 590280 43503 590336
rect 41492 590278 43503 590280
rect 43437 590275 43503 590278
rect 40493 589660 40559 589661
rect 40493 589656 40540 589660
rect 40604 589658 40610 589660
rect 40493 589600 40498 589656
rect 40493 589596 40540 589600
rect 40604 589598 40650 589658
rect 40604 589596 40610 589598
rect 41270 589596 41276 589660
rect 41340 589658 41346 589660
rect 41822 589658 41828 589660
rect 41340 589598 41828 589658
rect 41340 589596 41346 589598
rect 41822 589596 41828 589598
rect 41892 589596 41898 589660
rect 40493 589595 40559 589596
rect 40902 589324 40908 589388
rect 40972 589386 40978 589388
rect 42057 589386 42123 589389
rect 40972 589384 42123 589386
rect 40972 589328 42062 589384
rect 42118 589328 42123 589384
rect 40972 589326 42123 589328
rect 40972 589324 40978 589326
rect 42057 589323 42123 589326
rect 39941 585986 40007 585989
rect 40350 585986 40356 585988
rect 39941 585984 40356 585986
rect 39941 585928 39946 585984
rect 40002 585928 40356 585984
rect 39941 585926 40356 585928
rect 39941 585923 40007 585926
rect 40350 585924 40356 585926
rect 40420 585924 40426 585988
rect 41505 585986 41571 585989
rect 42701 585986 42767 585989
rect 41505 585984 42767 585986
rect 41505 585928 41510 585984
rect 41566 585928 42706 585984
rect 42762 585928 42767 585984
rect 41505 585926 42767 585928
rect 41505 585923 41571 585926
rect 42701 585923 42767 585926
rect 32397 585714 32463 585717
rect 41822 585714 41828 585716
rect 32397 585712 41828 585714
rect 32397 585656 32402 585712
rect 32458 585656 41828 585712
rect 32397 585654 41828 585656
rect 32397 585651 32463 585654
rect 41822 585652 41828 585654
rect 41892 585652 41898 585716
rect 39665 585306 39731 585309
rect 42374 585306 42380 585308
rect 39665 585304 42380 585306
rect 39665 585248 39670 585304
rect 39726 585248 42380 585304
rect 39665 585246 42380 585248
rect 39665 585243 39731 585246
rect 42374 585244 42380 585246
rect 42444 585244 42450 585308
rect 40217 585034 40283 585037
rect 42241 585034 42307 585037
rect 40217 585032 42307 585034
rect 40217 584976 40222 585032
rect 40278 584976 42246 585032
rect 42302 584976 42307 585032
rect 40217 584974 42307 584976
rect 40217 584971 40283 584974
rect 42241 584971 42307 584974
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40677 584626 40743 584629
rect 41086 584626 41092 584628
rect 40677 584624 41092 584626
rect 40677 584568 40682 584624
rect 40738 584568 41092 584624
rect 40677 584566 41092 584568
rect 40677 584563 40743 584566
rect 41086 584564 41092 584566
rect 41156 584564 41162 584628
rect 41413 584626 41479 584629
rect 42006 584626 42012 584628
rect 41413 584624 42012 584626
rect 41413 584568 41418 584624
rect 41474 584568 42012 584624
rect 41413 584566 42012 584568
rect 41413 584563 41479 584566
rect 42006 584564 42012 584566
rect 42076 584564 42082 584628
rect 40350 582524 40356 582588
rect 40420 582586 40426 582588
rect 41781 582586 41847 582589
rect 40420 582584 41847 582586
rect 40420 582528 41786 582584
rect 41842 582528 41847 582584
rect 40420 582526 41847 582528
rect 40420 582524 40426 582526
rect 41781 582523 41847 582526
rect 47577 582450 47643 582453
rect 42566 582448 47643 582450
rect 42566 582392 47582 582448
rect 47638 582392 47643 582448
rect 42566 582390 47643 582392
rect 42152 582330 42626 582390
rect 47577 582387 47643 582390
rect 42152 581634 42212 582330
rect 42152 581574 42258 581634
rect 42198 581501 42258 581574
rect 42198 581496 42307 581501
rect 42198 581440 42246 581496
rect 42302 581440 42307 581496
rect 42198 581438 42307 581440
rect 42241 581435 42307 581438
rect 661861 581090 661927 581093
rect 661861 581088 676292 581090
rect 661861 581032 661866 581088
rect 661922 581032 676292 581088
rect 661861 581030 676292 581032
rect 661861 581027 661927 581030
rect 673821 580818 673887 580821
rect 673821 580816 676322 580818
rect 673821 580760 673826 580816
rect 673882 580760 676322 580816
rect 673821 580758 676322 580760
rect 673821 580755 673887 580758
rect 40902 580620 40908 580684
rect 40972 580682 40978 580684
rect 42425 580682 42491 580685
rect 40972 580680 42491 580682
rect 40972 580624 42430 580680
rect 42486 580624 42491 580680
rect 676262 580652 676322 580758
rect 40972 580622 42491 580624
rect 40972 580620 40978 580622
rect 42425 580619 42491 580622
rect 671429 580546 671495 580549
rect 674833 580546 674899 580549
rect 671429 580544 674899 580546
rect 671429 580488 671434 580544
rect 671490 580488 674838 580544
rect 674894 580488 674899 580544
rect 671429 580486 674899 580488
rect 671429 580483 671495 580486
rect 674833 580483 674899 580486
rect 41086 580212 41092 580276
rect 41156 580274 41162 580276
rect 41781 580274 41847 580277
rect 41156 580272 41847 580274
rect 41156 580216 41786 580272
rect 41842 580216 41847 580272
rect 41156 580214 41847 580216
rect 41156 580212 41162 580214
rect 41781 580211 41847 580214
rect 42057 580138 42123 580141
rect 42014 580136 42123 580138
rect 42014 580080 42062 580136
rect 42118 580080 42123 580136
rect 42014 580075 42123 580080
rect 669957 580138 670023 580141
rect 676262 580138 676322 580244
rect 669957 580136 676322 580138
rect 669957 580080 669962 580136
rect 670018 580080 676322 580136
rect 669957 580078 676322 580080
rect 669957 580075 670023 580078
rect 40718 579940 40724 580004
rect 40788 580002 40794 580004
rect 42014 580002 42074 580075
rect 40788 579942 42074 580002
rect 40788 579940 40794 579942
rect 674833 579866 674899 579869
rect 674833 579864 676292 579866
rect 674833 579808 674838 579864
rect 674894 579808 676292 579864
rect 674833 579806 676292 579808
rect 674833 579803 674899 579806
rect 664437 579730 664503 579733
rect 673821 579730 673887 579733
rect 664437 579728 673887 579730
rect 664437 579672 664442 579728
rect 664498 579672 673826 579728
rect 673882 579672 673887 579728
rect 664437 579670 673887 579672
rect 664437 579667 664503 579670
rect 673821 579667 673887 579670
rect 674833 579458 674899 579461
rect 674833 579456 676292 579458
rect 674833 579400 674838 579456
rect 674894 579400 676292 579456
rect 674833 579398 676292 579400
rect 674833 579395 674899 579398
rect 672993 579186 673059 579189
rect 672993 579184 676322 579186
rect 672993 579128 672998 579184
rect 673054 579128 676322 579184
rect 672993 579126 676322 579128
rect 672993 579123 673059 579126
rect 676262 579020 676322 579126
rect 42057 578914 42123 578917
rect 44449 578914 44515 578917
rect 42057 578912 44515 578914
rect 42057 578856 42062 578912
rect 42118 578856 44454 578912
rect 44510 578856 44515 578912
rect 42057 578854 44515 578856
rect 42057 578851 42123 578854
rect 44449 578851 44515 578854
rect 671337 578914 671403 578917
rect 674833 578914 674899 578917
rect 671337 578912 674899 578914
rect 671337 578856 671342 578912
rect 671398 578856 674838 578912
rect 674894 578856 674899 578912
rect 671337 578854 674899 578856
rect 671337 578851 671403 578854
rect 674833 578851 674899 578854
rect 672441 578642 672507 578645
rect 672441 578640 676292 578642
rect 672441 578584 672446 578640
rect 672502 578584 676292 578640
rect 672441 578582 676292 578584
rect 672441 578579 672507 578582
rect 42241 578368 42307 578373
rect 675477 578370 675543 578373
rect 42241 578312 42246 578368
rect 42302 578312 42307 578368
rect 42241 578307 42307 578312
rect 674606 578368 675543 578370
rect 674606 578312 675482 578368
rect 675538 578312 675543 578368
rect 674606 578310 675543 578312
rect 42244 577829 42304 578307
rect 671521 578098 671587 578101
rect 674606 578098 674666 578310
rect 675477 578307 675543 578310
rect 676262 578098 676322 578204
rect 671521 578096 674666 578098
rect 671521 578040 671526 578096
rect 671582 578040 674666 578096
rect 671521 578038 674666 578040
rect 674790 578038 676322 578098
rect 671521 578035 671587 578038
rect 42241 577824 42307 577829
rect 42241 577768 42246 577824
rect 42302 577768 42307 577824
rect 42241 577763 42307 577768
rect 670877 577690 670943 577693
rect 674790 577690 674850 578038
rect 670877 577688 674850 577690
rect 670877 577632 670882 577688
rect 670938 577632 674850 577688
rect 670877 577630 674850 577632
rect 675293 577690 675359 577693
rect 676262 577690 676322 577796
rect 675293 577688 676322 577690
rect 675293 577632 675298 577688
rect 675354 577632 676322 577688
rect 675293 577630 676322 577632
rect 670877 577627 670943 577630
rect 675293 577627 675359 577630
rect 651465 577418 651531 577421
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 651465 577355 651531 577358
rect 671705 577282 671771 577285
rect 676262 577282 676322 577388
rect 671705 577280 676322 577282
rect 671705 577224 671710 577280
rect 671766 577224 676322 577280
rect 671705 577222 676322 577224
rect 671705 577219 671771 577222
rect 675477 577010 675543 577013
rect 675477 577008 676292 577010
rect 675477 576952 675482 577008
rect 675538 576952 676292 577008
rect 675477 576950 676292 576952
rect 675477 576947 675543 576950
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 42241 576874 42307 576877
rect 40604 576872 42307 576874
rect 40604 576816 42246 576872
rect 42302 576816 42307 576872
rect 40604 576814 42307 576816
rect 40604 576812 40610 576814
rect 42241 576811 42307 576814
rect 671337 576874 671403 576877
rect 675293 576874 675359 576877
rect 671337 576872 675359 576874
rect 671337 576816 671342 576872
rect 671398 576816 675298 576872
rect 675354 576816 675359 576872
rect 671337 576814 675359 576816
rect 671337 576811 671403 576814
rect 675293 576811 675359 576814
rect 41965 576602 42031 576605
rect 42190 576602 42196 576604
rect 41965 576600 42196 576602
rect 41965 576544 41970 576600
rect 42026 576544 42196 576600
rect 41965 576542 42196 576544
rect 41965 576539 42031 576542
rect 42190 576540 42196 576542
rect 42260 576540 42266 576604
rect 675845 576602 675911 576605
rect 675845 576600 676292 576602
rect 675845 576544 675850 576600
rect 675906 576544 676292 576600
rect 675845 576542 676292 576544
rect 675845 576539 675911 576542
rect 676990 576404 676996 576468
rect 677060 576404 677066 576468
rect 676998 576164 677058 576404
rect 680997 576058 681063 576061
rect 680997 576056 681106 576058
rect 680997 576000 681002 576056
rect 681058 576000 681106 576056
rect 680997 575995 681106 576000
rect 681046 575756 681106 575995
rect 674925 575378 674991 575381
rect 674925 575376 676292 575378
rect 674925 575320 674930 575376
rect 674986 575320 676292 575376
rect 674925 575318 676292 575320
rect 674925 575315 674991 575318
rect 668209 574834 668275 574837
rect 676262 574834 676322 574940
rect 668209 574832 676322 574834
rect 668209 574776 668214 574832
rect 668270 574776 676322 574832
rect 668209 574774 676322 574776
rect 668209 574771 668275 574774
rect 668945 574426 669011 574429
rect 676262 574426 676322 574532
rect 668945 574424 676322 574426
rect 668945 574368 668950 574424
rect 669006 574368 676322 574424
rect 668945 574366 676322 574368
rect 668945 574363 669011 574366
rect 42149 574154 42215 574157
rect 42885 574154 42951 574157
rect 42149 574152 42951 574154
rect 42149 574096 42154 574152
rect 42210 574096 42890 574152
rect 42946 574096 42951 574152
rect 42149 574094 42951 574096
rect 42149 574091 42215 574094
rect 42885 574091 42951 574094
rect 671981 574154 672047 574157
rect 671981 574152 676292 574154
rect 671981 574096 671986 574152
rect 672042 574096 676292 574152
rect 671981 574094 676292 574096
rect 671981 574091 672047 574094
rect 683297 574018 683363 574021
rect 683254 574016 683363 574018
rect 683254 573960 683302 574016
rect 683358 573960 683363 574016
rect 683254 573955 683363 573960
rect 683254 573716 683314 573955
rect 41965 573204 42031 573205
rect 41965 573200 42012 573204
rect 42076 573202 42082 573204
rect 673085 573202 673151 573205
rect 676262 573202 676322 573308
rect 683481 573202 683547 573205
rect 41965 573144 41970 573200
rect 41965 573140 42012 573144
rect 42076 573142 42122 573202
rect 673085 573200 676322 573202
rect 673085 573144 673090 573200
rect 673146 573144 676322 573200
rect 673085 573142 676322 573144
rect 683438 573200 683547 573202
rect 683438 573144 683486 573200
rect 683542 573144 683547 573200
rect 42076 573140 42082 573142
rect 41965 573139 42031 573140
rect 673085 573139 673151 573142
rect 683438 573139 683547 573144
rect 683438 572900 683498 573139
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 676814 572492 676874 572732
rect 672809 571978 672875 571981
rect 676262 571978 676322 572084
rect 683113 571978 683179 571981
rect 672809 571976 676322 571978
rect 672809 571920 672814 571976
rect 672870 571920 676322 571976
rect 672809 571918 676322 571920
rect 683070 571976 683179 571978
rect 683070 571920 683118 571976
rect 683174 571920 683179 571976
rect 672809 571915 672875 571918
rect 683070 571915 683179 571920
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 41454 571644 41460 571708
rect 41524 571706 41530 571708
rect 42425 571706 42491 571709
rect 41524 571704 42491 571706
rect 41524 571648 42430 571704
rect 42486 571648 42491 571704
rect 683070 571676 683130 571915
rect 41524 571646 42491 571648
rect 41524 571644 41530 571646
rect 42425 571643 42491 571646
rect 41822 571372 41828 571436
rect 41892 571434 41898 571436
rect 42241 571434 42307 571437
rect 41892 571432 42307 571434
rect 41892 571376 42246 571432
rect 42302 571376 42307 571432
rect 41892 571374 42307 571376
rect 41892 571372 41898 571374
rect 42241 571371 42307 571374
rect 671797 571162 671863 571165
rect 676262 571162 676322 571268
rect 671797 571160 676322 571162
rect 671797 571104 671802 571160
rect 671858 571104 676322 571160
rect 671797 571102 676322 571104
rect 671797 571099 671863 571102
rect 41638 570964 41644 571028
rect 41708 571026 41714 571028
rect 42057 571026 42123 571029
rect 41708 571024 42123 571026
rect 41708 570968 42062 571024
rect 42118 570968 42123 571024
rect 41708 570966 42123 570968
rect 41708 570964 41714 570966
rect 42057 570963 42123 570966
rect 676262 570754 676322 570860
rect 682377 570754 682443 570757
rect 674790 570694 676322 570754
rect 682334 570752 682443 570754
rect 682334 570696 682382 570752
rect 682438 570696 682443 570752
rect 671705 570346 671771 570349
rect 674790 570346 674850 570694
rect 671705 570344 674850 570346
rect 671705 570288 671710 570344
rect 671766 570288 674850 570344
rect 671705 570286 674850 570288
rect 682334 570691 682443 570696
rect 671705 570283 671771 570286
rect 682334 570044 682394 570691
rect 671981 569530 672047 569533
rect 676262 569530 676322 569636
rect 671981 569528 676322 569530
rect 671981 569472 671986 569528
rect 672042 569472 676322 569528
rect 671981 569470 676322 569472
rect 671981 569467 672047 569470
rect 62113 569258 62179 569261
rect 51030 569256 62179 569258
rect 51030 569200 62118 569256
rect 62174 569200 62179 569256
rect 51030 569198 62179 569200
rect 42241 569122 42307 569125
rect 51030 569122 51090 569198
rect 62113 569195 62179 569198
rect 42241 569120 51090 569122
rect 42241 569064 42246 569120
rect 42302 569064 51090 569120
rect 42241 569062 51090 569064
rect 42241 569059 42307 569062
rect 669037 564498 669103 564501
rect 675293 564498 675359 564501
rect 669037 564496 675359 564498
rect 669037 564440 669042 564496
rect 669098 564440 675298 564496
rect 675354 564440 675359 564496
rect 669037 564438 675359 564440
rect 669037 564435 669103 564438
rect 675293 564435 675359 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675477 562732 675543 562733
rect 675477 562728 675524 562732
rect 675588 562730 675594 562732
rect 675477 562672 675482 562728
rect 675477 562668 675524 562672
rect 675588 562670 675634 562730
rect 675588 562668 675594 562670
rect 675477 562667 675543 562668
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 674833 559738 674899 559741
rect 675293 559738 675359 559741
rect 674833 559736 675359 559738
rect 674833 559680 674838 559736
rect 674894 559680 675298 559736
rect 675354 559680 675359 559736
rect 674833 559678 675359 559680
rect 674833 559675 674899 559678
rect 675293 559675 675359 559678
rect 672257 559466 672323 559469
rect 675385 559466 675451 559469
rect 672257 559464 675451 559466
rect 672257 559408 672262 559464
rect 672318 559408 675390 559464
rect 675446 559408 675451 559464
rect 672257 559406 675451 559408
rect 672257 559403 672323 559406
rect 675385 559403 675451 559406
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 42057 558514 42123 558517
rect 41492 558512 42123 558514
rect 41492 558456 42062 558512
rect 42118 558456 42123 558512
rect 41492 558454 42123 558456
rect 42057 558451 42123 558454
rect 673821 558378 673887 558381
rect 675385 558378 675451 558381
rect 673821 558376 675451 558378
rect 673821 558320 673826 558376
rect 673882 558320 675390 558376
rect 675446 558320 675451 558376
rect 673821 558318 675451 558320
rect 673821 558315 673887 558318
rect 675385 558315 675451 558318
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 48957 557834 49023 557837
rect 41830 557832 49023 557834
rect 41830 557776 48962 557832
rect 49018 557776 49023 557832
rect 41830 557774 49023 557776
rect 41830 557698 41890 557774
rect 48957 557771 49023 557774
rect 41492 557638 41890 557698
rect 675753 557698 675819 557701
rect 676254 557698 676260 557700
rect 675753 557696 676260 557698
rect 675753 557640 675758 557696
rect 675814 557640 676260 557696
rect 675753 557638 676260 557640
rect 675753 557635 675819 557638
rect 676254 557636 676260 557638
rect 676324 557636 676330 557700
rect 42057 557562 42123 557565
rect 51717 557562 51783 557565
rect 42057 557560 51783 557562
rect 42057 557504 42062 557560
rect 42118 557504 51722 557560
rect 51778 557504 51783 557560
rect 42057 557502 51783 557504
rect 42057 557499 42123 557502
rect 51717 557499 51783 557502
rect 668209 557562 668275 557565
rect 674925 557562 674991 557565
rect 668209 557560 674991 557562
rect 668209 557504 668214 557560
rect 668270 557504 674930 557560
rect 674986 557504 674991 557560
rect 668209 557502 674991 557504
rect 668209 557499 668275 557502
rect 674925 557499 674991 557502
rect 44633 557290 44699 557293
rect 41492 557288 44699 557290
rect 41492 557232 44638 557288
rect 44694 557232 44699 557288
rect 41492 557230 44699 557232
rect 44633 557227 44699 557230
rect 45553 556882 45619 556885
rect 41492 556880 45619 556882
rect 41492 556824 45558 556880
rect 45614 556824 45619 556880
rect 41492 556822 45619 556824
rect 45553 556819 45619 556822
rect 44817 556474 44883 556477
rect 41492 556472 44883 556474
rect 41492 556416 44822 556472
rect 44878 556416 44883 556472
rect 41492 556414 44883 556416
rect 44817 556411 44883 556414
rect 44817 556066 44883 556069
rect 41492 556064 44883 556066
rect 41492 556008 44822 556064
rect 44878 556008 44883 556064
rect 41492 556006 44883 556008
rect 44817 556003 44883 556006
rect 674925 555794 674991 555797
rect 675477 555794 675543 555797
rect 674925 555792 675543 555794
rect 674925 555736 674930 555792
rect 674986 555736 675482 555792
rect 675538 555736 675543 555792
rect 674925 555734 675543 555736
rect 674925 555731 674991 555734
rect 675477 555731 675543 555734
rect 45001 555658 45067 555661
rect 41492 555656 45067 555658
rect 41492 555600 45006 555656
rect 45062 555600 45067 555656
rect 41492 555598 45067 555600
rect 45001 555595 45067 555598
rect 44357 555250 44423 555253
rect 41492 555248 44423 555250
rect 41492 555192 44362 555248
rect 44418 555192 44423 555248
rect 41492 555190 44423 555192
rect 44357 555187 44423 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 669589 554706 669655 554709
rect 675385 554706 675451 554709
rect 669589 554704 675451 554706
rect 669589 554648 669594 554704
rect 669650 554648 675390 554704
rect 675446 554648 675451 554704
rect 669589 554646 675451 554648
rect 669589 554643 669655 554646
rect 675385 554643 675451 554646
rect 44725 554434 44791 554437
rect 41492 554432 44791 554434
rect 41492 554376 44730 554432
rect 44786 554376 44791 554432
rect 41492 554374 44791 554376
rect 44725 554371 44791 554374
rect 35617 554026 35683 554029
rect 35604 554024 35683 554026
rect 35604 553968 35622 554024
rect 35678 553968 35683 554024
rect 35604 553966 35683 553968
rect 35617 553963 35683 553966
rect 659101 554026 659167 554029
rect 670049 554026 670115 554029
rect 659101 554024 670115 554026
rect 659101 553968 659106 554024
rect 659162 553968 670054 554024
rect 670110 553968 670115 554024
rect 659101 553966 670115 553968
rect 659101 553963 659167 553966
rect 670049 553963 670115 553966
rect 675753 554026 675819 554029
rect 676806 554026 676812 554028
rect 675753 554024 676812 554026
rect 675753 553968 675758 554024
rect 675814 553968 676812 554024
rect 675753 553966 676812 553968
rect 675753 553963 675819 553966
rect 676806 553964 676812 553966
rect 676876 553964 676882 554028
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 673085 553482 673151 553485
rect 675385 553482 675451 553485
rect 673085 553480 675451 553482
rect 673085 553424 673090 553480
rect 673146 553424 675390 553480
rect 675446 553424 675451 553480
rect 673085 553422 675451 553424
rect 673085 553419 673151 553422
rect 675385 553419 675451 553422
rect 40861 553210 40927 553213
rect 41781 553212 41847 553213
rect 40861 553208 40940 553210
rect 40861 553152 40866 553208
rect 40922 553152 40940 553208
rect 40861 553150 40940 553152
rect 41781 553208 41828 553212
rect 41892 553210 41898 553212
rect 41781 553152 41786 553208
rect 40861 553147 40927 553150
rect 41781 553148 41828 553152
rect 41892 553150 41938 553210
rect 41892 553148 41898 553150
rect 41781 553147 41847 553148
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 43161 552394 43227 552397
rect 41492 552392 43227 552394
rect 41492 552336 43166 552392
rect 43222 552336 43227 552392
rect 41492 552334 43227 552336
rect 43161 552331 43227 552334
rect 670877 552122 670943 552125
rect 675385 552122 675451 552125
rect 670877 552120 675451 552122
rect 670877 552064 670882 552120
rect 670938 552064 675390 552120
rect 675446 552064 675451 552120
rect 670877 552062 675451 552064
rect 670877 552059 670943 552062
rect 675385 552059 675451 552062
rect 33777 551986 33843 551989
rect 33764 551984 33843 551986
rect 33764 551928 33782 551984
rect 33838 551928 33843 551984
rect 33764 551926 33843 551928
rect 33777 551923 33843 551926
rect 45093 551578 45159 551581
rect 41492 551576 45159 551578
rect 41492 551520 45098 551576
rect 45154 551520 45159 551576
rect 41492 551518 45159 551520
rect 45093 551515 45159 551518
rect 670049 551578 670115 551581
rect 675385 551578 675451 551581
rect 670049 551576 675451 551578
rect 670049 551520 670054 551576
rect 670110 551520 675390 551576
rect 675446 551520 675451 551576
rect 670049 551518 675451 551520
rect 670049 551515 670115 551518
rect 675385 551515 675451 551518
rect 41229 551170 41295 551173
rect 41229 551168 41308 551170
rect 41229 551112 41234 551168
rect 41290 551112 41308 551168
rect 41229 551110 41308 551112
rect 41229 551107 41295 551110
rect 651465 550898 651531 550901
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 651465 550835 651531 550838
rect 44541 550762 44607 550765
rect 41492 550760 44607 550762
rect 41492 550704 44546 550760
rect 44602 550704 44607 550760
rect 41492 550702 44607 550704
rect 44541 550699 44607 550702
rect 675017 550490 675083 550493
rect 675886 550490 675892 550492
rect 675017 550488 675892 550490
rect 675017 550432 675022 550488
rect 675078 550432 675892 550488
rect 675017 550430 675892 550432
rect 675017 550427 675083 550430
rect 675886 550428 675892 550430
rect 675956 550428 675962 550492
rect 42057 550354 42123 550357
rect 41492 550352 42123 550354
rect 41492 550296 42062 550352
rect 42118 550296 42123 550352
rect 41492 550294 42123 550296
rect 42057 550291 42123 550294
rect 675753 550218 675819 550221
rect 676990 550218 676996 550220
rect 675753 550216 676996 550218
rect 675753 550160 675758 550216
rect 675814 550160 676996 550216
rect 675753 550158 676996 550160
rect 675753 550155 675819 550158
rect 676990 550156 676996 550158
rect 677060 550156 677066 550220
rect 41873 549946 41939 549949
rect 41492 549944 41939 549946
rect 41492 549888 41878 549944
rect 41934 549888 41939 549944
rect 41492 549886 41939 549888
rect 41873 549883 41939 549886
rect 41229 549538 41295 549541
rect 41229 549536 41308 549538
rect 41229 549480 41234 549536
rect 41290 549480 41308 549536
rect 41229 549478 41308 549480
rect 41229 549475 41295 549478
rect 41689 549402 41755 549405
rect 42977 549402 43043 549405
rect 41689 549400 43043 549402
rect 41689 549344 41694 549400
rect 41750 549344 42982 549400
rect 43038 549344 43043 549400
rect 41689 549342 43043 549344
rect 41689 549339 41755 549342
rect 42977 549339 43043 549342
rect 45277 549130 45343 549133
rect 41492 549128 45343 549130
rect 41492 549072 45282 549128
rect 45338 549072 45343 549128
rect 41492 549070 45343 549072
rect 45277 549067 45343 549070
rect 44173 548722 44239 548725
rect 41492 548720 44239 548722
rect 41492 548664 44178 548720
rect 44234 548664 44239 548720
rect 41492 548662 44239 548664
rect 44173 548659 44239 548662
rect 673637 548450 673703 548453
rect 675477 548450 675543 548453
rect 673637 548448 675543 548450
rect 673637 548392 673642 548448
rect 673698 548392 675482 548448
rect 675538 548392 675543 548448
rect 673637 548390 675543 548392
rect 673637 548387 673703 548390
rect 675477 548387 675543 548390
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 28766 547498 28826 547890
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 675937 547636 676003 547637
rect 675886 547634 675892 547636
rect 675846 547574 675892 547634
rect 675956 547632 676003 547636
rect 675998 547576 676003 547632
rect 675886 547572 675892 547574
rect 675956 547572 676003 547576
rect 676254 547572 676260 547636
rect 676324 547634 676330 547636
rect 677409 547634 677475 547637
rect 676324 547632 677475 547634
rect 676324 547576 677414 547632
rect 677470 547576 677475 547632
rect 676324 547574 677475 547576
rect 676324 547572 676330 547574
rect 675937 547571 676003 547572
rect 677409 547571 677475 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 43805 547090 43871 547093
rect 41492 547088 43871 547090
rect 41492 547032 43810 547088
rect 43866 547032 43871 547088
rect 41492 547030 43871 547032
rect 43805 547027 43871 547030
rect 674005 547090 674071 547093
rect 683389 547090 683455 547093
rect 674005 547088 683455 547090
rect 674005 547032 674010 547088
rect 674066 547032 683394 547088
rect 683450 547032 683455 547088
rect 674005 547030 683455 547032
rect 674005 547027 674071 547030
rect 683389 547027 683455 547030
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40718 545668 40724 545732
rect 40788 545730 40794 545732
rect 42057 545730 42123 545733
rect 40788 545728 42123 545730
rect 40788 545672 42062 545728
rect 42118 545672 42123 545728
rect 40788 545670 42123 545672
rect 40788 545668 40794 545670
rect 42057 545667 42123 545670
rect 674281 545730 674347 545733
rect 683205 545730 683271 545733
rect 674281 545728 683271 545730
rect 674281 545672 674286 545728
rect 674342 545672 683210 545728
rect 683266 545672 683271 545728
rect 674281 545670 683271 545672
rect 674281 545667 674347 545670
rect 683205 545667 683271 545670
rect 40534 545396 40540 545460
rect 40604 545458 40610 545460
rect 41873 545458 41939 545461
rect 40604 545456 41939 545458
rect 40604 545400 41878 545456
rect 41934 545400 41939 545456
rect 40604 545398 41939 545400
rect 40604 545396 40610 545398
rect 41873 545395 41939 545398
rect 675293 544916 675359 544917
rect 675293 544914 675340 544916
rect 675248 544912 675340 544914
rect 675248 544856 675298 544912
rect 675248 544854 675340 544856
rect 675293 544852 675340 544854
rect 675404 544852 675410 544916
rect 675293 544851 675359 544852
rect 674833 544506 674899 544509
rect 675518 544506 675524 544508
rect 674833 544504 675524 544506
rect 674833 544448 674838 544504
rect 674894 544448 675524 544504
rect 674833 544446 675524 544448
rect 674833 544443 674899 544446
rect 675518 544444 675524 544446
rect 675588 544444 675594 544508
rect 674833 543962 674899 543965
rect 675477 543962 675543 543965
rect 674833 543960 675543 543962
rect 674833 543904 674838 543960
rect 674894 543904 675482 543960
rect 675538 543904 675543 543960
rect 674833 543902 675543 543904
rect 674833 543899 674899 543902
rect 675477 543899 675543 543902
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 663057 538794 663123 538797
rect 676029 538794 676095 538797
rect 663057 538792 676095 538794
rect 663057 538736 663062 538792
rect 663118 538736 676034 538792
rect 676090 538736 676095 538792
rect 663057 538734 676095 538736
rect 663057 538731 663123 538734
rect 676029 538731 676095 538734
rect 40718 538188 40724 538252
rect 40788 538250 40794 538252
rect 42241 538250 42307 538253
rect 40788 538248 42307 538250
rect 40788 538192 42246 538248
rect 42302 538192 42307 538248
rect 40788 538190 42307 538192
rect 40788 538188 40794 538190
rect 42241 538187 42307 538190
rect 42057 537978 42123 537981
rect 42609 537978 42675 537981
rect 42057 537976 42675 537978
rect 42057 537920 42062 537976
rect 42118 537920 42614 537976
rect 42670 537920 42675 537976
rect 42057 537918 42675 537920
rect 42057 537915 42123 537918
rect 42609 537915 42675 537918
rect 651465 537570 651531 537573
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 651465 537507 651531 537510
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 668577 535875 668643 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 42149 535258 42215 535261
rect 44173 535258 44239 535261
rect 42149 535256 44239 535258
rect 42149 535200 42154 535256
rect 42210 535200 44178 535256
rect 44234 535200 44239 535256
rect 42149 535198 44239 535200
rect 42149 535195 42215 535198
rect 44173 535195 44239 535198
rect 676262 535122 676322 535296
rect 669270 535062 676322 535122
rect 40534 534924 40540 534988
rect 40604 534986 40610 534988
rect 41781 534986 41847 534989
rect 40604 534984 41847 534986
rect 40604 534928 41786 534984
rect 41842 534928 41847 534984
rect 40604 534926 41847 534928
rect 40604 534924 40610 534926
rect 41781 534923 41847 534926
rect 42149 534442 42215 534445
rect 45277 534442 45343 534445
rect 42149 534440 45343 534442
rect 42149 534384 42154 534440
rect 42210 534384 45282 534440
rect 45338 534384 45343 534440
rect 42149 534382 45343 534384
rect 42149 534379 42215 534382
rect 45277 534379 45343 534382
rect 667197 534442 667263 534445
rect 669270 534442 669330 535062
rect 671245 534850 671311 534853
rect 676262 534850 676322 534888
rect 671245 534848 676322 534850
rect 671245 534792 671250 534848
rect 671306 534792 676322 534848
rect 671245 534790 676322 534792
rect 671245 534787 671311 534790
rect 672441 534578 672507 534581
rect 675753 534578 675819 534581
rect 672441 534576 675819 534578
rect 672441 534520 672446 534576
rect 672502 534520 675758 534576
rect 675814 534520 675819 534576
rect 672441 534518 675819 534520
rect 672441 534515 672507 534518
rect 675753 534515 675819 534518
rect 667197 534440 669330 534442
rect 667197 534384 667202 534440
rect 667258 534384 669330 534440
rect 667197 534382 669330 534384
rect 667197 534379 667263 534382
rect 672809 534306 672875 534309
rect 676262 534306 676322 534480
rect 672809 534304 676322 534306
rect 672809 534248 672814 534304
rect 672870 534248 676322 534304
rect 672809 534246 676322 534248
rect 672809 534243 672875 534246
rect 675753 534102 675819 534105
rect 675753 534100 676292 534102
rect 675753 534044 675758 534100
rect 675814 534044 676292 534100
rect 675753 534042 676292 534044
rect 675753 534039 675819 534042
rect 42149 533898 42215 533901
rect 43161 533898 43227 533901
rect 42149 533896 43227 533898
rect 42149 533840 42154 533896
rect 42210 533840 43166 533896
rect 43222 533840 43227 533896
rect 42149 533838 43227 533840
rect 42149 533835 42215 533838
rect 43161 533835 43227 533838
rect 674414 533836 674420 533900
rect 674484 533898 674490 533900
rect 683573 533898 683639 533901
rect 674484 533896 683639 533898
rect 674484 533840 683578 533896
rect 683634 533840 683639 533896
rect 674484 533838 683639 533840
rect 674484 533836 674490 533838
rect 683573 533835 683639 533838
rect 675753 533694 675819 533697
rect 675753 533692 676292 533694
rect 675753 533636 675758 533692
rect 675814 533636 676292 533692
rect 675753 533634 676292 533636
rect 675753 533631 675819 533634
rect 671429 533490 671495 533493
rect 671429 533488 676322 533490
rect 671429 533432 671434 533488
rect 671490 533432 676322 533488
rect 671429 533430 676322 533432
rect 671429 533427 671495 533430
rect 676262 533256 676322 533430
rect 42241 533218 42307 533221
rect 42977 533218 43043 533221
rect 42241 533216 43043 533218
rect 42241 533160 42246 533216
rect 42302 533160 42982 533216
rect 43038 533160 43043 533216
rect 42241 533158 43043 533160
rect 42241 533155 42307 533158
rect 42977 533155 43043 533158
rect 674189 533218 674255 533221
rect 675753 533218 675819 533221
rect 674189 533216 675819 533218
rect 674189 533160 674194 533216
rect 674250 533160 675758 533216
rect 675814 533160 675819 533216
rect 674189 533158 675819 533160
rect 674189 533155 674255 533158
rect 675753 533155 675819 533158
rect 674005 532946 674071 532949
rect 674005 532944 676322 532946
rect 674005 532888 674010 532944
rect 674066 532888 676322 532944
rect 674005 532886 676322 532888
rect 674005 532883 674071 532886
rect 676262 532848 676322 532886
rect 42517 532810 42583 532813
rect 44541 532810 44607 532813
rect 42517 532808 44607 532810
rect 42517 532752 42522 532808
rect 42578 532752 44546 532808
rect 44602 532752 44607 532808
rect 42517 532750 44607 532752
rect 42517 532747 42583 532750
rect 44541 532747 44607 532750
rect 62113 532810 62179 532813
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 62113 532747 62179 532750
rect 671521 532674 671587 532677
rect 671521 532672 676322 532674
rect 671521 532616 671526 532672
rect 671582 532616 676322 532672
rect 671521 532614 676322 532616
rect 671521 532611 671587 532614
rect 676262 532440 676322 532614
rect 676262 531994 676322 532032
rect 676170 531934 676322 531994
rect 672441 531858 672507 531861
rect 676170 531858 676230 531934
rect 672441 531856 676230 531858
rect 672441 531800 672446 531856
rect 672502 531800 676230 531856
rect 672441 531798 676230 531800
rect 672441 531795 672507 531798
rect 666461 531450 666527 531453
rect 676262 531450 676322 531624
rect 666461 531448 676322 531450
rect 666461 531392 666466 531448
rect 666522 531392 676322 531448
rect 666461 531390 676322 531392
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 666461 531387 666527 531390
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 41454 530572 41460 530636
rect 41524 530634 41530 530636
rect 42517 530634 42583 530637
rect 41524 530632 42583 530634
rect 41524 530576 42522 530632
rect 42578 530576 42583 530632
rect 41524 530574 42583 530576
rect 41524 530572 41530 530574
rect 42517 530571 42583 530574
rect 668393 530634 668459 530637
rect 676262 530634 676322 530808
rect 668393 530632 676322 530634
rect 668393 530576 668398 530632
rect 668454 530576 676322 530632
rect 668393 530574 676322 530576
rect 668393 530571 668459 530574
rect 674649 530362 674715 530365
rect 676262 530362 676322 530400
rect 674649 530360 676322 530362
rect 674649 530304 674654 530360
rect 674710 530304 676322 530360
rect 674649 530302 676322 530304
rect 674649 530299 674715 530302
rect 42149 530090 42215 530093
rect 42701 530090 42767 530093
rect 42149 530088 42767 530090
rect 42149 530032 42154 530088
rect 42210 530032 42706 530088
rect 42762 530032 42767 530088
rect 42149 530030 42767 530032
rect 42149 530027 42215 530030
rect 42701 530027 42767 530030
rect 670233 530090 670299 530093
rect 670233 530088 676322 530090
rect 670233 530032 670238 530088
rect 670294 530032 676322 530088
rect 670233 530030 676322 530032
rect 670233 530027 670299 530030
rect 676262 529992 676322 530030
rect 42609 529682 42675 529685
rect 45093 529682 45159 529685
rect 42609 529680 45159 529682
rect 42609 529624 42614 529680
rect 42670 529624 45098 529680
rect 45154 529624 45159 529680
rect 42609 529622 45159 529624
rect 42609 529619 42675 529622
rect 45093 529619 45159 529622
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 671521 529410 671587 529413
rect 676262 529410 676322 529584
rect 671521 529408 676322 529410
rect 671521 529352 671526 529408
rect 671582 529352 676322 529408
rect 671521 529350 676322 529352
rect 671521 529347 671587 529350
rect 41638 529076 41644 529140
rect 41708 529138 41714 529140
rect 42885 529138 42951 529141
rect 41708 529136 42951 529138
rect 41708 529080 42890 529136
rect 42946 529080 42951 529136
rect 41708 529078 42951 529080
rect 41708 529076 41714 529078
rect 42885 529075 42951 529078
rect 669221 529002 669287 529005
rect 676262 529002 676322 529176
rect 669221 529000 676322 529002
rect 669221 528944 669226 529000
rect 669282 528944 676322 529000
rect 669221 528942 676322 528944
rect 669221 528939 669287 528942
rect 673269 528730 673335 528733
rect 676262 528730 676322 528768
rect 673269 528728 676322 528730
rect 673269 528672 673274 528728
rect 673330 528672 676322 528728
rect 673269 528670 676322 528672
rect 673269 528667 673335 528670
rect 668761 528594 668827 528597
rect 671521 528594 671587 528597
rect 668761 528592 671587 528594
rect 668761 528536 668766 528592
rect 668822 528536 671526 528592
rect 671582 528536 671587 528592
rect 668761 528534 671587 528536
rect 668761 528531 668827 528534
rect 671521 528531 671587 528534
rect 683389 528594 683455 528597
rect 683389 528592 683498 528594
rect 683389 528536 683394 528592
rect 683450 528536 683498 528592
rect 683389 528531 683498 528536
rect 683438 528360 683498 528531
rect 672625 528186 672691 528189
rect 672625 528184 676322 528186
rect 672625 528128 672630 528184
rect 672686 528128 676322 528184
rect 672625 528126 676322 528128
rect 672625 528123 672691 528126
rect 676262 527952 676322 528126
rect 674465 527778 674531 527781
rect 674465 527776 676322 527778
rect 674465 527720 674470 527776
rect 674526 527720 676322 527776
rect 674465 527718 676322 527720
rect 674465 527715 674531 527718
rect 676262 527544 676322 527718
rect 683573 527370 683639 527373
rect 683573 527368 683682 527370
rect 683573 527312 683578 527368
rect 683634 527312 683682 527368
rect 683573 527307 683682 527312
rect 683622 527136 683682 527307
rect 683205 526962 683271 526965
rect 683205 526960 683314 526962
rect 683205 526904 683210 526960
rect 683266 526904 683314 526960
rect 683205 526899 683314 526904
rect 683254 526728 683314 526899
rect 673453 526554 673519 526557
rect 673453 526552 676322 526554
rect 673453 526496 673458 526552
rect 673514 526496 676322 526552
rect 673453 526494 676322 526496
rect 673453 526491 673519 526494
rect 676262 526320 676322 526494
rect 676814 525741 676874 525912
rect 671061 525738 671127 525741
rect 671061 525736 676322 525738
rect 671061 525680 671066 525736
rect 671122 525680 676322 525736
rect 671061 525678 676322 525680
rect 676814 525736 676923 525741
rect 676814 525680 676862 525736
rect 676918 525680 676923 525736
rect 676814 525678 676923 525680
rect 671061 525675 671127 525678
rect 676262 525096 676322 525678
rect 676857 525675 676923 525678
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 675477 513770 675543 513773
rect 676029 513770 676095 513773
rect 675477 513768 676095 513770
rect 675477 513712 675482 513768
rect 675538 513712 676034 513768
rect 676090 513712 676095 513768
rect 675477 513710 676095 513712
rect 675477 513707 675543 513710
rect 676029 513707 676095 513710
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683573 503706 683639 503709
rect 677060 503704 683639 503706
rect 677060 503648 683578 503704
rect 683634 503648 683639 503704
rect 677060 503646 683639 503648
rect 677060 503644 677066 503646
rect 683573 503643 683639 503646
rect 676806 503372 676812 503436
rect 676876 503434 676882 503436
rect 683389 503434 683455 503437
rect 676876 503432 683455 503434
rect 676876 503376 683394 503432
rect 683450 503376 683455 503432
rect 676876 503374 683455 503376
rect 676876 503372 676882 503374
rect 683389 503371 683455 503374
rect 675109 502618 675175 502621
rect 675845 502618 675911 502621
rect 675109 502616 675911 502618
rect 675109 502560 675114 502616
rect 675170 502560 675850 502616
rect 675906 502560 675911 502616
rect 675109 502558 675911 502560
rect 675109 502555 675175 502558
rect 675845 502555 675911 502558
rect 671705 500986 671771 500989
rect 676397 500986 676463 500989
rect 671705 500984 676463 500986
rect 671705 500928 671710 500984
rect 671766 500928 676402 500984
rect 676458 500928 676463 500984
rect 671705 500926 676463 500928
rect 671705 500923 671771 500926
rect 676397 500923 676463 500926
rect 652569 497722 652635 497725
rect 650164 497720 652635 497722
rect 650164 497664 652574 497720
rect 652630 497664 652635 497720
rect 650164 497662 652635 497664
rect 652569 497659 652635 497662
rect 666001 494050 666067 494053
rect 675845 494050 675911 494053
rect 666001 494048 675911 494050
rect 666001 493992 666006 494048
rect 666062 493992 675850 494048
rect 675906 493992 675911 494048
rect 666001 493990 675911 493992
rect 666001 493987 666067 493990
rect 675845 493987 675911 493990
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 663750 492086 676292 492146
rect 658917 492010 658983 492013
rect 663750 492010 663810 492086
rect 658917 492008 663810 492010
rect 658917 491952 658922 492008
rect 658978 491952 663810 492008
rect 658917 491950 663810 491952
rect 658917 491947 658983 491950
rect 664621 491738 664687 491741
rect 664621 491736 676292 491738
rect 664621 491680 664626 491736
rect 664682 491680 676292 491736
rect 664621 491678 676292 491680
rect 664621 491675 664687 491678
rect 683113 491330 683179 491333
rect 683100 491328 683179 491330
rect 683100 491272 683118 491328
rect 683174 491272 683179 491328
rect 683100 491270 683179 491272
rect 683113 491267 683179 491270
rect 672901 490922 672967 490925
rect 672901 490920 676292 490922
rect 672901 490864 672906 490920
rect 672962 490864 676292 490920
rect 672901 490862 676292 490864
rect 672901 490859 672967 490862
rect 676029 490514 676095 490517
rect 676029 490512 676292 490514
rect 676029 490456 676034 490512
rect 676090 490456 676292 490512
rect 676029 490454 676292 490456
rect 676029 490451 676095 490454
rect 674189 490106 674255 490109
rect 674189 490104 676292 490106
rect 674189 490048 674194 490104
rect 674250 490048 676292 490104
rect 674189 490046 676292 490048
rect 674189 490043 674255 490046
rect 672901 489698 672967 489701
rect 672901 489696 676292 489698
rect 672901 489640 672906 489696
rect 672962 489640 676292 489696
rect 672901 489638 676292 489640
rect 672901 489635 672967 489638
rect 672717 489290 672783 489293
rect 672717 489288 676292 489290
rect 672717 489232 672722 489288
rect 672778 489232 676292 489288
rect 672717 489230 676292 489232
rect 672717 489227 672783 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 672441 488474 672507 488477
rect 672441 488472 676292 488474
rect 672441 488416 672446 488472
rect 672502 488416 676292 488472
rect 672441 488414 676292 488416
rect 672441 488411 672507 488414
rect 672441 488066 672507 488069
rect 672441 488064 676292 488066
rect 672441 488008 672446 488064
rect 672502 488008 676292 488064
rect 672441 488006 676292 488008
rect 672441 488003 672507 488006
rect 679617 487658 679683 487661
rect 679604 487656 679683 487658
rect 679604 487600 679622 487656
rect 679678 487600 679683 487656
rect 679604 487598 679683 487600
rect 679617 487595 679683 487598
rect 683573 487250 683639 487253
rect 683573 487248 683652 487250
rect 683573 487192 683578 487248
rect 683634 487192 683652 487248
rect 683573 487190 683652 487192
rect 683573 487187 683639 487190
rect 680997 486842 681063 486845
rect 680997 486840 681076 486842
rect 680997 486784 681002 486840
rect 681058 486784 681076 486840
rect 680997 486782 681076 486784
rect 680997 486779 681063 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 668209 486026 668275 486029
rect 668209 486024 676292 486026
rect 668209 485968 668214 486024
rect 668270 485968 676292 486024
rect 668209 485966 676292 485968
rect 668209 485963 668275 485966
rect 673637 485618 673703 485621
rect 673637 485616 676292 485618
rect 673637 485560 673642 485616
rect 673698 485560 676292 485616
rect 673637 485558 676292 485560
rect 673637 485555 673703 485558
rect 669270 485150 676292 485210
rect 669037 485074 669103 485077
rect 669270 485074 669330 485150
rect 669037 485072 669330 485074
rect 669037 485016 669042 485072
rect 669098 485016 669330 485072
rect 669037 485014 669330 485016
rect 669037 485011 669103 485014
rect 672165 484802 672231 484805
rect 672165 484800 676292 484802
rect 672165 484744 672170 484800
rect 672226 484744 676292 484800
rect 672165 484742 676292 484744
rect 672165 484739 672231 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 673821 484394 673887 484397
rect 673821 484392 676292 484394
rect 673821 484336 673826 484392
rect 673882 484336 676292 484392
rect 673821 484334 676292 484336
rect 673821 484331 673887 484334
rect 670877 483986 670943 483989
rect 670877 483984 676292 483986
rect 670877 483928 670882 483984
rect 670938 483928 676292 483984
rect 670877 483926 676292 483928
rect 670877 483923 670943 483926
rect 683389 483578 683455 483581
rect 683389 483576 683468 483578
rect 683389 483520 683394 483576
rect 683450 483520 683468 483576
rect 683389 483518 683468 483520
rect 683389 483515 683455 483518
rect 677409 483170 677475 483173
rect 677396 483168 677475 483170
rect 677396 483112 677414 483168
rect 677470 483112 677475 483168
rect 677396 483110 677475 483112
rect 677409 483107 677475 483110
rect 674925 483034 674991 483037
rect 675845 483034 675911 483037
rect 674925 483032 675911 483034
rect 674925 482976 674930 483032
rect 674986 482976 675850 483032
rect 675906 482976 675911 483032
rect 674925 482974 675911 482976
rect 674925 482971 674991 482974
rect 675845 482971 675911 482974
rect 669589 482762 669655 482765
rect 669589 482760 676292 482762
rect 669589 482704 669594 482760
rect 669650 482704 676292 482760
rect 669589 482702 676292 482704
rect 669589 482699 669655 482702
rect 673085 482354 673151 482357
rect 673085 482352 676292 482354
rect 673085 482296 673090 482352
rect 673146 482296 676292 482352
rect 673085 482294 676292 482296
rect 673085 482291 673151 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675661 480722 675727 480725
rect 675661 480720 676292 480722
rect 675661 480664 675666 480720
rect 675722 480664 676292 480720
rect 675661 480662 676292 480664
rect 675661 480659 675727 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 674598 475356 674604 475420
rect 674668 475418 674674 475420
rect 677133 475418 677199 475421
rect 674668 475416 677199 475418
rect 674668 475360 677138 475416
rect 677194 475360 677199 475416
rect 674668 475358 677199 475360
rect 674668 475356 674674 475358
rect 677133 475355 677199 475358
rect 673269 474876 673335 474877
rect 673269 474874 673316 474876
rect 673224 474872 673316 474874
rect 673224 474816 673274 474872
rect 673224 474814 673316 474816
rect 673269 474812 673316 474814
rect 673380 474812 673386 474876
rect 673269 474811 673335 474812
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 674833 456378 674899 456381
rect 675845 456378 675911 456381
rect 674833 456376 675911 456378
rect 674833 456320 674838 456376
rect 674894 456320 675850 456376
rect 675906 456320 675911 456376
rect 674833 456318 675911 456320
rect 674833 456315 674899 456318
rect 675845 456315 675911 456318
rect 667841 456106 667907 456109
rect 673453 456106 673519 456109
rect 667841 456104 673519 456106
rect 667841 456048 667846 456104
rect 667902 456048 673458 456104
rect 673514 456048 673519 456104
rect 667841 456046 673519 456048
rect 667841 456043 667907 456046
rect 673453 456043 673519 456046
rect 673821 456106 673887 456109
rect 675845 456106 675911 456109
rect 673821 456104 675911 456106
rect 673821 456048 673826 456104
rect 673882 456048 675850 456104
rect 675906 456048 675911 456104
rect 673821 456046 675911 456048
rect 673821 456043 673887 456046
rect 675845 456043 675911 456046
rect 670601 455834 670667 455837
rect 673729 455834 673795 455837
rect 670601 455832 673795 455834
rect 670601 455776 670606 455832
rect 670662 455776 673734 455832
rect 673790 455776 673795 455832
rect 670601 455774 673795 455776
rect 670601 455771 670667 455774
rect 673729 455771 673795 455774
rect 670417 455426 670483 455429
rect 673499 455426 673565 455429
rect 670417 455424 673565 455426
rect 670417 455368 670422 455424
rect 670478 455368 673504 455424
rect 673560 455368 673565 455424
rect 670417 455366 673565 455368
rect 670417 455363 670483 455366
rect 673499 455363 673565 455366
rect 669773 455154 669839 455157
rect 673381 455154 673447 455157
rect 669773 455152 673447 455154
rect 669773 455096 669778 455152
rect 669834 455096 673386 455152
rect 673442 455096 673447 455152
rect 669773 455094 673447 455096
rect 669773 455091 669839 455094
rect 673381 455091 673447 455094
rect 673545 455154 673611 455157
rect 676673 455154 676739 455157
rect 673545 455152 676739 455154
rect 673545 455096 673550 455152
rect 673606 455096 676678 455152
rect 676734 455096 676739 455152
rect 673545 455094 676739 455096
rect 673545 455091 673611 455094
rect 676673 455091 676739 455094
rect 673039 454882 673105 454885
rect 675477 454882 675543 454885
rect 673039 454880 675543 454882
rect 673039 454824 673044 454880
rect 673100 454824 675482 454880
rect 675538 454824 675543 454880
rect 673039 454822 675543 454824
rect 673039 454819 673105 454822
rect 675477 454819 675543 454822
rect 62113 454610 62179 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 62113 454547 62179 454550
rect 672809 454474 672875 454477
rect 675661 454474 675727 454477
rect 672809 454472 675727 454474
rect 672809 454416 672814 454472
rect 672870 454416 675666 454472
rect 675722 454416 675727 454472
rect 672809 454414 675727 454416
rect 672809 454411 672875 454414
rect 675661 454411 675727 454414
rect 672947 454202 673013 454205
rect 675937 454202 676003 454205
rect 672947 454200 676003 454202
rect 672947 454144 672952 454200
rect 673008 454144 675942 454200
rect 675998 454144 676003 454200
rect 672947 454142 676003 454144
rect 672947 454139 673013 454142
rect 675937 454139 676003 454142
rect 672257 453930 672323 453933
rect 674833 453930 674899 453933
rect 672257 453928 674899 453930
rect 672257 453872 672262 453928
rect 672318 453872 674838 453928
rect 674894 453872 674899 453928
rect 672257 453870 674899 453872
rect 672257 453867 672323 453870
rect 674833 453867 674899 453870
rect 675334 453732 675340 453796
rect 675404 453794 675410 453796
rect 676121 453794 676187 453797
rect 675404 453792 676187 453794
rect 675404 453736 676126 453792
rect 676182 453736 676187 453792
rect 675404 453734 676187 453736
rect 675404 453732 675410 453734
rect 676121 453731 676187 453734
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45553 429722 45619 429725
rect 41492 429720 45619 429722
rect 41492 429664 45558 429720
rect 45614 429664 45619 429720
rect 41492 429662 45619 429664
rect 45553 429659 45619 429662
rect 45185 429314 45251 429317
rect 41492 429312 45251 429314
rect 41492 429256 45190 429312
rect 45246 429256 45251 429312
rect 41492 429254 45251 429256
rect 45185 429251 45251 429254
rect 44909 428906 44975 428909
rect 41492 428904 44975 428906
rect 41492 428848 44914 428904
rect 44970 428848 44975 428904
rect 41492 428846 44975 428848
rect 44909 428843 44975 428846
rect 45001 428498 45067 428501
rect 41492 428496 45067 428498
rect 41492 428440 45006 428496
rect 45062 428440 45067 428496
rect 41492 428438 45067 428440
rect 45001 428435 45067 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44357 428090 44423 428093
rect 41492 428088 44423 428090
rect 41492 428032 44362 428088
rect 44418 428032 44423 428088
rect 41492 428030 44423 428032
rect 44357 428027 44423 428030
rect 44449 427682 44515 427685
rect 41492 427680 44515 427682
rect 41492 427624 44454 427680
rect 44510 427624 44515 427680
rect 41492 427622 44515 427624
rect 44449 427619 44515 427622
rect 44725 427274 44791 427277
rect 41492 427272 44791 427274
rect 41492 427216 44730 427272
rect 44786 427216 44791 427272
rect 41492 427214 44791 427216
rect 44725 427211 44791 427214
rect 44265 426866 44331 426869
rect 41492 426864 44331 426866
rect 41492 426808 44270 426864
rect 44326 426808 44331 426864
rect 41492 426806 44331 426808
rect 44265 426803 44331 426806
rect 46933 426458 46999 426461
rect 41492 426456 46999 426458
rect 41492 426400 46938 426456
rect 46994 426400 46999 426456
rect 41492 426398 46999 426400
rect 46933 426395 46999 426398
rect 40953 426050 41019 426053
rect 40940 426048 41019 426050
rect 40940 425992 40958 426048
rect 41014 425992 41019 426048
rect 40940 425990 41019 425992
rect 40953 425987 41019 425990
rect 40769 425642 40835 425645
rect 40756 425640 40835 425642
rect 40756 425584 40774 425640
rect 40830 425584 40835 425640
rect 40756 425582 40835 425584
rect 40769 425579 40835 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 36537 424418 36603 424421
rect 36524 424416 36603 424418
rect 36524 424360 36542 424416
rect 36598 424360 36603 424416
rect 36524 424358 36603 424360
rect 36537 424355 36603 424358
rect 41321 424010 41387 424013
rect 41308 424008 41387 424010
rect 41308 423952 41326 424008
rect 41382 423952 41387 424008
rect 41308 423950 41387 423952
rect 41321 423947 41387 423950
rect 47117 423602 47183 423605
rect 41492 423600 47183 423602
rect 41492 423544 47122 423600
rect 47178 423544 47183 423600
rect 41492 423542 47183 423544
rect 47117 423539 47183 423542
rect 41462 423168 41844 423228
rect 41462 423164 41522 423168
rect 41784 423061 41844 423168
rect 41781 423056 41847 423061
rect 41781 423000 41786 423056
rect 41842 423000 41847 423056
rect 41781 422995 41847 423000
rect 42149 422786 42215 422789
rect 41492 422784 42215 422786
rect 41492 422728 42154 422784
rect 42210 422728 42215 422784
rect 41492 422726 42215 422728
rect 42149 422723 42215 422726
rect 44633 422514 44699 422517
rect 41692 422512 44699 422514
rect 41692 422456 44638 422512
rect 44694 422456 44699 422512
rect 41692 422454 44699 422456
rect 41692 422412 41752 422454
rect 44633 422451 44699 422454
rect 41278 422352 41752 422412
rect 41278 422348 41338 422352
rect 41781 422242 41847 422245
rect 43069 422242 43135 422245
rect 41781 422240 43135 422242
rect 41781 422184 41786 422240
rect 41842 422184 43074 422240
rect 43130 422184 43135 422240
rect 41781 422182 43135 422184
rect 41781 422179 41847 422182
rect 43069 422179 43135 422182
rect 40493 421970 40559 421973
rect 40493 421968 40572 421970
rect 40493 421912 40498 421968
rect 40554 421912 40572 421968
rect 40493 421910 40572 421912
rect 40493 421907 40559 421910
rect 41781 421562 41847 421565
rect 41492 421560 41847 421562
rect 41492 421504 41786 421560
rect 41842 421504 41847 421560
rect 41492 421502 41847 421504
rect 41781 421499 41847 421502
rect 43253 421154 43319 421157
rect 41492 421152 43319 421154
rect 41492 421096 43258 421152
rect 43314 421096 43319 421152
rect 41492 421094 43319 421096
rect 43253 421091 43319 421094
rect 44817 420746 44883 420749
rect 41492 420744 44883 420746
rect 41492 420688 44822 420744
rect 44878 420688 44883 420744
rect 41492 420686 44883 420688
rect 44817 420683 44883 420686
rect 41462 419930 41522 420308
rect 42517 419930 42583 419933
rect 41462 419928 42583 419930
rect 41462 419900 42522 419928
rect 41492 419872 42522 419900
rect 42578 419872 42583 419928
rect 41492 419870 42583 419872
rect 42517 419867 42583 419870
rect 43989 419522 44055 419525
rect 41492 419520 44055 419522
rect 41492 419464 43994 419520
rect 44050 419464 44055 419520
rect 41492 419462 44055 419464
rect 43989 419459 44055 419462
rect 40769 418842 40835 418845
rect 41638 418842 41644 418844
rect 40769 418840 41644 418842
rect 40769 418784 40774 418840
rect 40830 418784 41644 418840
rect 40769 418782 41644 418784
rect 40769 418779 40835 418782
rect 41638 418780 41644 418782
rect 41708 418780 41714 418844
rect 40493 418708 40559 418709
rect 40493 418704 40540 418708
rect 40604 418706 40610 418708
rect 40493 418648 40498 418704
rect 40493 418644 40540 418648
rect 40604 418646 40650 418706
rect 40604 418644 40610 418646
rect 40493 418643 40559 418644
rect 40718 418508 40724 418572
rect 40788 418570 40794 418572
rect 42149 418570 42215 418573
rect 40788 418568 42215 418570
rect 40788 418512 42154 418568
rect 42210 418512 42215 418568
rect 40788 418510 42215 418512
rect 40788 418508 40794 418510
rect 42149 418507 42215 418510
rect 41781 418298 41847 418301
rect 45369 418298 45435 418301
rect 41781 418296 45435 418298
rect 41781 418240 41786 418296
rect 41842 418240 45374 418296
rect 45430 418240 45435 418296
rect 41781 418238 45435 418240
rect 41781 418235 41847 418238
rect 45369 418235 45435 418238
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 675334 410484 675340 410548
rect 675404 410546 675410 410548
rect 676029 410546 676095 410549
rect 675404 410544 676095 410546
rect 675404 410488 676034 410544
rect 676090 410488 676095 410544
rect 675404 410486 676095 410488
rect 675404 410484 675410 410486
rect 676029 410483 676095 410486
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 43253 407826 43319 407829
rect 42425 407824 43319 407826
rect 42425 407768 42430 407824
rect 42486 407768 43258 407824
rect 43314 407768 43319 407824
rect 42425 407766 43319 407768
rect 42425 407763 42491 407766
rect 43253 407763 43319 407766
rect 42425 407146 42491 407149
rect 44633 407146 44699 407149
rect 42425 407144 44699 407146
rect 42425 407088 42430 407144
rect 42486 407088 44638 407144
rect 44694 407088 44699 407144
rect 42425 407086 44699 407088
rect 42425 407083 42491 407086
rect 44633 407083 44699 407086
rect 42425 406874 42491 406877
rect 45369 406874 45435 406877
rect 42425 406872 45435 406874
rect 42425 406816 42430 406872
rect 42486 406816 45374 406872
rect 45430 406816 45435 406872
rect 42425 406814 45435 406816
rect 42425 406811 42491 406814
rect 45369 406811 45435 406814
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 660297 405650 660363 405653
rect 675845 405650 675911 405653
rect 660297 405648 675911 405650
rect 660297 405592 660302 405648
rect 660358 405592 675850 405648
rect 675906 405592 675911 405648
rect 660297 405590 675911 405592
rect 660297 405587 660363 405590
rect 675845 405587 675911 405590
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669957 403746 670023 403749
rect 676262 403746 676322 403852
rect 669957 403744 676322 403746
rect 669957 403688 669962 403744
rect 670018 403688 676322 403744
rect 669957 403686 676322 403688
rect 669957 403683 670023 403686
rect 675845 403474 675911 403477
rect 675845 403472 676292 403474
rect 675845 403416 675850 403472
rect 675906 403416 676292 403472
rect 675845 403414 676292 403416
rect 675845 403411 675911 403414
rect 683113 403338 683179 403341
rect 682886 403336 683179 403338
rect 682886 403280 683118 403336
rect 683174 403280 683179 403336
rect 682886 403278 683179 403280
rect 682886 403036 682946 403278
rect 683113 403275 683179 403278
rect 42333 402930 42399 402933
rect 43069 402930 43135 402933
rect 42333 402928 43135 402930
rect 42333 402872 42338 402928
rect 42394 402872 43074 402928
rect 43130 402872 43135 402928
rect 42333 402870 43135 402872
rect 42333 402867 42399 402870
rect 43069 402867 43135 402870
rect 676029 402658 676095 402661
rect 676029 402656 676292 402658
rect 676029 402600 676034 402656
rect 676090 402600 676292 402656
rect 676029 402598 676292 402600
rect 676029 402595 676095 402598
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674833 402250 674899 402253
rect 674833 402248 676292 402250
rect 674833 402192 674838 402248
rect 674894 402192 676292 402248
rect 674833 402190 676292 402192
rect 674833 402187 674899 402190
rect 672625 401978 672691 401981
rect 672625 401976 676322 401978
rect 672625 401920 672630 401976
rect 672686 401920 676322 401976
rect 672625 401918 676322 401920
rect 672625 401915 672691 401918
rect 41454 401780 41460 401844
rect 41524 401842 41530 401844
rect 41781 401842 41847 401845
rect 41524 401840 41847 401842
rect 41524 401784 41786 401840
rect 41842 401784 41847 401840
rect 676262 401812 676322 401918
rect 41524 401782 41847 401784
rect 41524 401780 41530 401782
rect 41781 401779 41847 401782
rect 672993 401706 673059 401709
rect 674833 401706 674899 401709
rect 672993 401704 674899 401706
rect 672993 401648 672998 401704
rect 673054 401648 674838 401704
rect 674894 401648 674899 401704
rect 672993 401646 674899 401648
rect 672993 401643 673059 401646
rect 674833 401643 674899 401646
rect 673177 401298 673243 401301
rect 676262 401298 676322 401404
rect 673177 401296 676322 401298
rect 673177 401240 673182 401296
rect 673238 401240 676322 401296
rect 673177 401238 676322 401240
rect 673177 401235 673243 401238
rect 676806 401236 676812 401300
rect 676876 401236 676882 401300
rect 676814 400996 676874 401236
rect 672257 400482 672323 400485
rect 676262 400482 676322 400588
rect 672257 400480 676322 400482
rect 672257 400424 672262 400480
rect 672318 400424 676322 400480
rect 672257 400422 676322 400424
rect 672257 400419 672323 400422
rect 42425 400210 42491 400213
rect 47117 400210 47183 400213
rect 42425 400208 47183 400210
rect 42425 400152 42430 400208
rect 42486 400152 47122 400208
rect 47178 400152 47183 400208
rect 42425 400150 47183 400152
rect 42425 400147 42491 400150
rect 47117 400147 47183 400150
rect 672441 400074 672507 400077
rect 676262 400074 676322 400180
rect 672441 400072 676322 400074
rect 672441 400016 672446 400072
rect 672502 400016 676322 400072
rect 672441 400014 676322 400016
rect 672441 400011 672507 400014
rect 42425 399802 42491 399805
rect 46933 399802 46999 399805
rect 42425 399800 46999 399802
rect 42425 399744 42430 399800
rect 42486 399744 46938 399800
rect 46994 399744 46999 399800
rect 42425 399742 46999 399744
rect 42425 399739 42491 399742
rect 46933 399739 46999 399742
rect 674649 399802 674715 399805
rect 674649 399800 676292 399802
rect 674649 399744 674654 399800
rect 674710 399744 676292 399800
rect 674649 399742 676292 399744
rect 674649 399739 674715 399742
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41781 398852 41847 398853
rect 41781 398848 41828 398852
rect 41892 398850 41898 398852
rect 41781 398792 41786 398848
rect 41781 398788 41828 398792
rect 41892 398790 41938 398850
rect 41892 398788 41898 398790
rect 675886 398788 675892 398852
rect 675956 398850 675962 398852
rect 676262 398850 676322 398956
rect 675956 398790 676322 398850
rect 675956 398788 675962 398790
rect 41781 398787 41847 398788
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 674281 397354 674347 397357
rect 674281 397352 676292 397354
rect 674281 397296 674286 397352
rect 674342 397296 676292 397352
rect 674281 397294 676292 397296
rect 674281 397291 674347 397294
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 673361 396674 673427 396677
rect 673361 396672 676322 396674
rect 673361 396616 673366 396672
rect 673422 396616 676322 396672
rect 673361 396614 676322 396616
rect 673361 396611 673427 396614
rect 676262 396508 676322 396614
rect 673913 396130 673979 396133
rect 673913 396128 676292 396130
rect 673913 396072 673918 396128
rect 673974 396072 676292 396128
rect 673913 396070 676292 396072
rect 673913 396067 673979 396070
rect 673729 395722 673795 395725
rect 673729 395720 676292 395722
rect 673729 395664 673734 395720
rect 673790 395664 676292 395720
rect 673729 395662 676292 395664
rect 673729 395659 673795 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 673545 394362 673611 394365
rect 676262 394362 676322 394468
rect 673545 394360 676322 394362
rect 673545 394304 673550 394360
rect 673606 394304 676322 394360
rect 673545 394302 676322 394304
rect 673545 394299 673611 394302
rect 674465 394090 674531 394093
rect 674465 394088 676292 394090
rect 674465 394032 674470 394088
rect 674526 394032 676292 394088
rect 674465 394030 676292 394032
rect 674465 394027 674531 394030
rect 674097 393682 674163 393685
rect 674097 393680 676292 393682
rect 674097 393624 674102 393680
rect 674158 393624 676292 393680
rect 674097 393622 676292 393624
rect 674097 393619 674163 393622
rect 676070 393076 676076 393140
rect 676140 393138 676146 393140
rect 676262 393138 676322 393244
rect 676140 393078 676322 393138
rect 676140 393076 676146 393078
rect 676262 392836 676322 393078
rect 672717 392594 672783 392597
rect 672717 392592 676322 392594
rect 672717 392536 672722 392592
rect 672778 392536 676322 392592
rect 672717 392534 676322 392536
rect 672717 392531 672783 392534
rect 676262 392428 676322 392534
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 41492 387638 51090 387698
rect 41492 387230 49250 387290
rect 41137 387154 41203 387157
rect 41094 387152 41203 387154
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387091 41203 387096
rect 41094 386852 41154 387091
rect 41873 387018 41939 387021
rect 48957 387018 49023 387021
rect 41873 387016 49023 387018
rect 41873 386960 41878 387016
rect 41934 386960 48962 387016
rect 49018 386960 49023 387016
rect 41873 386958 49023 386960
rect 41873 386955 41939 386958
rect 48957 386955 49023 386958
rect 41321 386746 41387 386749
rect 41278 386744 41387 386746
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386683 41387 386688
rect 41505 386746 41571 386749
rect 45185 386746 45251 386749
rect 41505 386744 45251 386746
rect 41505 386688 41510 386744
rect 41566 386688 45190 386744
rect 45246 386688 45251 386744
rect 41505 386686 45251 386688
rect 41505 386683 41571 386686
rect 45185 386683 45251 386686
rect 41278 386444 41338 386683
rect 49190 386474 49250 387230
rect 51030 386746 51090 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 51717 386746 51783 386749
rect 51030 386744 51783 386746
rect 51030 386688 51722 386744
rect 51778 386688 51783 386744
rect 51030 386686 51783 386688
rect 51717 386683 51783 386686
rect 51901 386474 51967 386477
rect 49190 386472 51967 386474
rect 49190 386416 51906 386472
rect 51962 386416 51967 386472
rect 49190 386414 51967 386416
rect 51901 386411 51967 386414
rect 45185 386066 45251 386069
rect 41492 386064 45251 386066
rect 41492 386008 45190 386064
rect 45246 386008 45251 386064
rect 41492 386006 45251 386008
rect 45185 386003 45251 386006
rect 45001 385658 45067 385661
rect 41492 385656 45067 385658
rect 41492 385600 45006 385656
rect 45062 385600 45067 385656
rect 41492 385598 45067 385600
rect 45001 385595 45067 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 672993 385250 673059 385253
rect 673545 385250 673611 385253
rect 672993 385248 673611 385250
rect 672993 385192 672998 385248
rect 673054 385192 673550 385248
rect 673606 385192 673611 385248
rect 672993 385190 673611 385192
rect 672993 385187 673059 385190
rect 673545 385187 673611 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 44449 384842 44515 384845
rect 41492 384840 44515 384842
rect 41492 384784 44454 384840
rect 44510 384784 44515 384840
rect 41492 384782 44515 384784
rect 44449 384779 44515 384782
rect 45185 384434 45251 384437
rect 41492 384432 45251 384434
rect 41492 384376 45190 384432
rect 45246 384376 45251 384432
rect 41492 384374 45251 384376
rect 45185 384371 45251 384374
rect 44265 384026 44331 384029
rect 41492 384024 44331 384026
rect 41492 383968 44270 384024
rect 44326 383968 44331 384024
rect 41492 383966 44331 383968
rect 44265 383963 44331 383966
rect 45369 383618 45435 383621
rect 41492 383616 45435 383618
rect 41492 383560 45374 383616
rect 45430 383560 45435 383616
rect 41492 383558 45435 383560
rect 45369 383555 45435 383558
rect 41094 383077 41154 383180
rect 41094 383072 41203 383077
rect 41094 383016 41142 383072
rect 41198 383016 41203 383072
rect 41094 383014 41203 383016
rect 41137 383011 41203 383014
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 41689 382258 41755 382261
rect 42793 382258 42859 382261
rect 41689 382256 42859 382258
rect 41689 382200 41694 382256
rect 41750 382200 42798 382256
rect 42854 382200 42859 382256
rect 41689 382198 42859 382200
rect 41689 382195 41755 382198
rect 42793 382195 42859 382198
rect 673361 382258 673427 382261
rect 675385 382258 675451 382261
rect 673361 382256 675451 382258
rect 673361 382200 673366 382256
rect 673422 382200 675390 382256
rect 675446 382200 675451 382256
rect 673361 382198 675451 382200
rect 673361 382195 673427 382198
rect 675385 382195 675451 382198
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 40726 381445 40786 381548
rect 40726 381440 40835 381445
rect 40726 381384 40774 381440
rect 40830 381384 40835 381440
rect 40726 381382 40835 381384
rect 40769 381379 40835 381382
rect 673913 381442 673979 381445
rect 675109 381442 675175 381445
rect 673913 381440 675175 381442
rect 673913 381384 673918 381440
rect 673974 381384 675114 381440
rect 675170 381384 675175 381440
rect 673913 381382 675175 381384
rect 673913 381379 673979 381382
rect 675109 381379 675175 381382
rect 41278 381037 41338 381140
rect 41278 381032 41387 381037
rect 41278 380976 41326 381032
rect 41382 380976 41387 381032
rect 41278 380974 41387 380976
rect 41321 380971 41387 380974
rect 46933 380762 46999 380765
rect 41492 380760 46999 380762
rect 41492 380704 46938 380760
rect 46994 380704 46999 380760
rect 41492 380702 46999 380704
rect 46933 380699 46999 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 45553 380354 45619 380357
rect 41492 380352 45619 380354
rect 41492 380296 45558 380352
rect 45614 380296 45619 380352
rect 41492 380294 45619 380296
rect 45553 380291 45619 380294
rect 44449 379946 44515 379949
rect 41492 379944 44515 379946
rect 41492 379888 44454 379944
rect 44510 379888 44515 379944
rect 41492 379886 44515 379888
rect 44449 379883 44515 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 41689 379402 41755 379405
rect 42977 379402 43043 379405
rect 41689 379400 43043 379402
rect 41689 379344 41694 379400
rect 41750 379344 42982 379400
rect 43038 379344 43043 379400
rect 41689 379342 43043 379344
rect 41689 379339 41755 379342
rect 42977 379339 43043 379342
rect 673085 379402 673151 379405
rect 675293 379402 675359 379405
rect 673085 379400 675359 379402
rect 673085 379344 673090 379400
rect 673146 379344 675298 379400
rect 675354 379344 675359 379400
rect 673085 379342 675359 379344
rect 673085 379339 673151 379342
rect 675293 379339 675359 379342
rect 47117 379130 47183 379133
rect 41492 379128 47183 379130
rect 41492 379072 47122 379128
rect 47178 379072 47183 379128
rect 41492 379070 47183 379072
rect 47117 379067 47183 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 40769 378586 40835 378589
rect 41822 378586 41828 378588
rect 40769 378584 41828 378586
rect 40769 378528 40774 378584
rect 40830 378528 41828 378584
rect 40769 378526 41828 378528
rect 40769 378523 40835 378526
rect 41822 378524 41828 378526
rect 41892 378524 41898 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 652017 378178 652083 378181
rect 650164 378176 652083 378178
rect 650164 378120 652022 378176
rect 652078 378120 652083 378176
rect 650164 378118 652083 378120
rect 652017 378115 652083 378118
rect 674281 378042 674347 378045
rect 674782 378042 674788 378044
rect 674281 378040 674788 378042
rect 674281 377984 674286 378040
rect 674342 377984 674788 378040
rect 674281 377982 674788 377984
rect 674281 377979 674347 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 41321 377770 41387 377773
rect 42333 377770 42399 377773
rect 41321 377768 42399 377770
rect 41321 377712 41326 377768
rect 41382 377712 42338 377768
rect 42394 377712 42399 377768
rect 41321 377710 42399 377712
rect 41321 377707 41387 377710
rect 42333 377707 42399 377710
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 35758 376549 35818 377060
rect 674465 376682 674531 376685
rect 675109 376682 675175 376685
rect 674465 376680 675175 376682
rect 674465 376624 674470 376680
rect 674526 376624 675114 376680
rect 675170 376624 675175 376680
rect 674465 376622 675175 376624
rect 674465 376619 674531 376622
rect 675109 376619 675175 376622
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 40033 376546 40099 376549
rect 41638 376546 41644 376548
rect 40033 376544 41644 376546
rect 40033 376488 40038 376544
rect 40094 376488 41644 376544
rect 40033 376486 41644 376488
rect 40033 376483 40099 376486
rect 41638 376484 41644 376486
rect 41708 376484 41714 376548
rect 62113 376274 62179 376277
rect 62113 376272 64492 376274
rect 28950 376141 29010 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 62113 376211 62179 376214
rect 28901 376136 29010 376141
rect 28901 376080 28906 376136
rect 28962 376080 29010 376136
rect 28901 376078 29010 376080
rect 28901 376075 28967 376078
rect 39481 375730 39547 375733
rect 40350 375730 40356 375732
rect 39481 375728 40356 375730
rect 39481 375672 39486 375728
rect 39542 375672 40356 375728
rect 39481 375670 40356 375672
rect 39481 375667 39547 375670
rect 40350 375668 40356 375670
rect 40420 375668 40426 375732
rect 673729 375458 673795 375461
rect 675109 375458 675175 375461
rect 673729 375456 675175 375458
rect 673729 375400 673734 375456
rect 673790 375400 675114 375456
rect 675170 375400 675175 375456
rect 673729 375398 675175 375400
rect 673729 375395 673795 375398
rect 675109 375395 675175 375398
rect 675293 375050 675359 375053
rect 675886 375050 675892 375052
rect 675293 375048 675892 375050
rect 675293 374992 675298 375048
rect 675354 374992 675892 375048
rect 675293 374990 675892 374992
rect 675293 374987 675359 374990
rect 675886 374988 675892 374990
rect 675956 374988 675962 375052
rect 675753 373010 675819 373013
rect 676070 373010 676076 373012
rect 675753 373008 676076 373010
rect 675753 372952 675758 373008
rect 675814 372952 676076 373008
rect 675753 372950 676076 372952
rect 675753 372947 675819 372950
rect 676070 372948 676076 372950
rect 676140 372948 676146 373012
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 41689 371922 41755 371925
rect 43345 371922 43411 371925
rect 41689 371920 43411 371922
rect 41689 371864 41694 371920
rect 41750 371864 43350 371920
rect 43406 371864 43411 371920
rect 41689 371862 43411 371864
rect 41689 371859 41755 371862
rect 43345 371859 43411 371862
rect 40350 368596 40356 368660
rect 40420 368658 40426 368660
rect 41781 368658 41847 368661
rect 40420 368656 41847 368658
rect 40420 368600 41786 368656
rect 41842 368600 41847 368656
rect 40420 368598 41847 368600
rect 40420 368596 40426 368598
rect 41781 368595 41847 368598
rect 42425 367026 42491 367029
rect 46197 367026 46263 367029
rect 42425 367024 46263 367026
rect 42425 366968 42430 367024
rect 42486 366968 46202 367024
rect 46258 366968 46263 367024
rect 42425 366966 46263 366968
rect 42425 366963 42491 366966
rect 46197 366963 46263 366966
rect 42425 365802 42491 365805
rect 42977 365802 43043 365805
rect 42425 365800 43043 365802
rect 42425 365744 42430 365800
rect 42486 365744 42982 365800
rect 43038 365744 43043 365800
rect 42425 365742 43043 365744
rect 42425 365739 42491 365742
rect 42977 365739 43043 365742
rect 651649 364850 651715 364853
rect 650164 364848 651715 364850
rect 650164 364792 651654 364848
rect 651710 364792 651715 364848
rect 650164 364790 651715 364792
rect 651649 364787 651715 364790
rect 40902 364244 40908 364308
rect 40972 364306 40978 364308
rect 41781 364306 41847 364309
rect 40972 364304 41847 364306
rect 40972 364248 41786 364304
rect 41842 364248 41847 364304
rect 40972 364246 41847 364248
rect 40972 364244 40978 364246
rect 41781 364243 41847 364246
rect 40718 363564 40724 363628
rect 40788 363626 40794 363628
rect 41781 363626 41847 363629
rect 40788 363624 41847 363626
rect 40788 363568 41786 363624
rect 41842 363568 41847 363624
rect 40788 363566 41847 363568
rect 40788 363564 40794 363566
rect 41781 363563 41847 363566
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 41781 362948 41847 362949
rect 41781 362944 41828 362948
rect 41892 362946 41898 362948
rect 41781 362888 41786 362944
rect 41781 362884 41828 362888
rect 41892 362886 41938 362946
rect 41892 362884 41898 362886
rect 41781 362883 41847 362884
rect 42425 361586 42491 361589
rect 47117 361586 47183 361589
rect 42425 361584 47183 361586
rect 42425 361528 42430 361584
rect 42486 361528 47122 361584
rect 47178 361528 47183 361584
rect 42425 361526 47183 361528
rect 42425 361523 42491 361526
rect 47117 361523 47183 361526
rect 670141 360906 670207 360909
rect 675845 360906 675911 360909
rect 670141 360904 675911 360906
rect 670141 360848 670146 360904
rect 670202 360848 675850 360904
rect 675906 360848 675911 360904
rect 670141 360846 675911 360848
rect 670141 360843 670207 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 42149 359954 42215 359957
rect 44449 359954 44515 359957
rect 42149 359952 44515 359954
rect 42149 359896 42154 359952
rect 42210 359896 44454 359952
rect 44510 359896 44515 359952
rect 42149 359894 44515 359896
rect 42149 359891 42215 359894
rect 44449 359891 44515 359894
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 665817 358730 665883 358733
rect 665817 358728 676292 358730
rect 665817 358672 665822 358728
rect 665878 358672 676292 358728
rect 665817 358670 676292 358672
rect 665817 358667 665883 358670
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 672993 357506 673059 357509
rect 672993 357504 676292 357506
rect 672993 357448 672998 357504
rect 673054 357448 676292 357504
rect 672993 357446 676292 357448
rect 672993 357443 673059 357446
rect 42425 357370 42491 357373
rect 45553 357370 45619 357373
rect 42425 357368 45619 357370
rect 42425 357312 42430 357368
rect 42486 357312 45558 357368
rect 45614 357312 45619 357368
rect 42425 357310 45619 357312
rect 42425 357307 42491 357310
rect 45553 357307 45619 357310
rect 673361 357098 673427 357101
rect 673361 357096 676292 357098
rect 673361 357040 673366 357096
rect 673422 357040 676292 357096
rect 673361 357038 676292 357040
rect 673361 357035 673427 357038
rect 44265 356690 44331 356693
rect 45645 356690 45711 356693
rect 44265 356688 45711 356690
rect 44265 356632 44270 356688
rect 44326 356632 45650 356688
rect 45706 356632 45711 356688
rect 44265 356630 45711 356632
rect 44265 356627 44331 356630
rect 45645 356627 45711 356630
rect 673177 356690 673243 356693
rect 673177 356688 676292 356690
rect 673177 356632 673182 356688
rect 673238 356632 676292 356688
rect 673177 356630 676292 356632
rect 673177 356627 673243 356630
rect 673913 356282 673979 356285
rect 673913 356280 676292 356282
rect 673913 356224 673918 356280
rect 673974 356224 676292 356280
rect 673913 356222 676292 356224
rect 673913 356219 673979 356222
rect 42425 356146 42491 356149
rect 46933 356146 46999 356149
rect 42425 356144 46999 356146
rect 42425 356088 42430 356144
rect 42486 356088 46938 356144
rect 46994 356088 46999 356144
rect 42425 356086 46999 356088
rect 42425 356083 42491 356086
rect 46933 356083 46999 356086
rect 43345 355874 43411 355877
rect 45921 355874 45987 355877
rect 43345 355872 45987 355874
rect 43345 355816 43350 355872
rect 43406 355816 45926 355872
rect 45982 355816 45987 355872
rect 43345 355814 45987 355816
rect 43345 355811 43411 355814
rect 45921 355811 45987 355814
rect 672257 355874 672323 355877
rect 672257 355872 676292 355874
rect 672257 355816 672262 355872
rect 672318 355816 676292 355872
rect 672257 355814 676292 355816
rect 672257 355811 672323 355814
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 673085 355466 673151 355469
rect 673085 355464 676292 355466
rect 673085 355408 673090 355464
rect 673146 355408 676292 355464
rect 673085 355406 676292 355408
rect 673085 355403 673151 355406
rect 674649 355058 674715 355061
rect 674649 355056 676292 355058
rect 674649 355000 674654 355056
rect 674710 355000 676292 355056
rect 674649 354998 676292 355000
rect 674649 354995 674715 354998
rect 672533 354650 672599 354653
rect 672533 354648 676292 354650
rect 672533 354592 672538 354648
rect 672594 354592 676292 354648
rect 672533 354590 676292 354592
rect 672533 354587 672599 354590
rect 43897 354244 43963 354245
rect 43846 354180 43852 354244
rect 43916 354242 43963 354244
rect 43916 354240 44008 354242
rect 43958 354184 44008 354240
rect 43916 354182 44008 354184
rect 43916 354180 43963 354182
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 43897 354179 43963 354180
rect 44214 353772 44220 353836
rect 44284 353834 44290 353836
rect 44725 353834 44791 353837
rect 44284 353832 44791 353834
rect 44284 353776 44730 353832
rect 44786 353776 44791 353832
rect 44284 353774 44791 353776
rect 44284 353772 44290 353774
rect 44725 353771 44791 353774
rect 676029 353834 676095 353837
rect 676029 353832 676292 353834
rect 676029 353776 676034 353832
rect 676090 353776 676292 353832
rect 676029 353774 676292 353776
rect 676029 353771 676095 353774
rect 674741 353426 674807 353429
rect 674741 353424 676292 353426
rect 674741 353368 674746 353424
rect 674802 353368 676292 353424
rect 674741 353366 676292 353368
rect 674741 353363 674807 353366
rect 675518 352956 675524 353020
rect 675588 353018 675594 353020
rect 675588 352958 676292 353018
rect 675588 352956 675594 352958
rect 673545 352610 673611 352613
rect 673545 352608 676292 352610
rect 673545 352552 673550 352608
rect 673606 352552 676292 352608
rect 673545 352550 676292 352552
rect 673545 352547 673611 352550
rect 674557 352202 674623 352205
rect 674557 352200 676292 352202
rect 674557 352144 674562 352200
rect 674618 352144 676292 352200
rect 674557 352142 676292 352144
rect 674557 352139 674623 352142
rect 675886 351868 675892 351932
rect 675956 351930 675962 351932
rect 675956 351870 676230 351930
rect 675956 351868 675962 351870
rect 676170 351794 676230 351870
rect 676170 351734 676292 351794
rect 651465 351658 651531 351661
rect 650164 351656 651531 351658
rect 650164 351600 651470 351656
rect 651526 351600 651531 351656
rect 650164 351598 651531 351600
rect 651465 351595 651531 351598
rect 672901 351386 672967 351389
rect 672901 351384 676292 351386
rect 672901 351328 672906 351384
rect 672962 351328 676292 351384
rect 672901 351326 676292 351328
rect 672901 351323 672967 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 673729 350570 673795 350573
rect 673729 350568 676292 350570
rect 673729 350512 673734 350568
rect 673790 350512 676292 350568
rect 673729 350510 676292 350512
rect 673729 350507 673795 350510
rect 62757 350298 62823 350301
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 62757 350235 62823 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 672165 349754 672231 349757
rect 672165 349752 676292 349754
rect 672165 349696 672170 349752
rect 672226 349696 676292 349752
rect 672165 349694 676292 349696
rect 672165 349691 672231 349694
rect 674373 349482 674439 349485
rect 674373 349480 676230 349482
rect 674373 349424 674378 349480
rect 674434 349424 676230 349480
rect 674373 349422 676230 349424
rect 674373 349419 674439 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 675937 349212 676003 349213
rect 675886 349210 675892 349212
rect 675846 349150 675892 349210
rect 675956 349208 676003 349212
rect 675998 349152 676003 349208
rect 675886 349148 675892 349150
rect 675956 349148 676003 349152
rect 675937 349147 676003 349148
rect 671981 348938 672047 348941
rect 671981 348936 676292 348938
rect 671981 348880 671986 348936
rect 672042 348880 676292 348936
rect 671981 348878 676292 348880
rect 671981 348875 672047 348878
rect 670141 348530 670207 348533
rect 670141 348528 676292 348530
rect 670141 348472 670146 348528
rect 670202 348472 676292 348528
rect 670141 348470 676292 348472
rect 670141 348467 670207 348470
rect 672349 347714 672415 347717
rect 683070 347714 683130 348092
rect 672349 347712 683130 347714
rect 672349 347656 672354 347712
rect 672410 347684 683130 347712
rect 672410 347656 683100 347684
rect 672349 347654 683100 347656
rect 672349 347651 672415 347654
rect 669957 347306 670023 347309
rect 669957 347304 676292 347306
rect 669957 347248 669962 347304
rect 670018 347248 676292 347304
rect 669957 347246 676292 347248
rect 669957 347243 670023 347246
rect 38285 346354 38351 346357
rect 49141 346354 49207 346357
rect 38285 346352 49207 346354
rect 38285 346296 38290 346352
rect 38346 346296 49146 346352
rect 49202 346296 49207 346352
rect 38285 346294 49207 346296
rect 38285 346291 38351 346294
rect 49141 346291 49207 346294
rect 28901 344314 28967 344317
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 28901 344312 29010 344314
rect 28901 344256 28906 344312
rect 28962 344256 29010 344312
rect 28901 344251 29010 344256
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 28950 344148 29010 344251
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 28582 343740 28642 343843
rect 45001 343362 45067 343365
rect 41492 343360 45067 343362
rect 41492 343304 45006 343360
rect 45062 343304 45067 343360
rect 41492 343302 45067 343304
rect 45001 343299 45067 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 44214 342682 44220 342684
rect 41462 342622 44220 342682
rect 41462 342516 41522 342622
rect 44214 342620 44220 342622
rect 44284 342620 44290 342684
rect 44398 342138 44404 342140
rect 41492 342078 44404 342138
rect 44398 342076 44404 342078
rect 44468 342076 44474 342140
rect 45277 341730 45343 341733
rect 41492 341728 45343 341730
rect 41492 341672 45282 341728
rect 45338 341672 45343 341728
rect 41492 341670 45343 341672
rect 45277 341667 45343 341670
rect 45277 341322 45343 341325
rect 41492 341320 45343 341322
rect 41492 341264 45282 341320
rect 45338 341264 45343 341320
rect 41492 341262 45343 341264
rect 45277 341259 45343 341262
rect 45461 340914 45527 340917
rect 41492 340912 45527 340914
rect 41492 340856 45466 340912
rect 45522 340856 45527 340912
rect 41492 340854 45527 340856
rect 45461 340851 45527 340854
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340234 675819 340237
rect 676622 340234 676628 340236
rect 675753 340232 676628 340234
rect 675753 340176 675758 340232
rect 675814 340176 676628 340232
rect 675753 340174 676628 340176
rect 675753 340171 675819 340174
rect 676622 340172 676628 340174
rect 676692 340172 676698 340236
rect 45829 340098 45895 340101
rect 41492 340096 45895 340098
rect 41492 340040 45834 340096
rect 45890 340040 45895 340096
rect 41492 340038 45895 340040
rect 45829 340035 45895 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 45645 339282 45711 339285
rect 41492 339280 45711 339282
rect 41492 339224 45650 339280
rect 45706 339224 45711 339280
rect 41492 339222 45711 339224
rect 45645 339219 45711 339222
rect 675385 339012 675451 339013
rect 675334 339010 675340 339012
rect 675294 338950 675340 339010
rect 675404 339008 675451 339012
rect 675446 338952 675451 339008
rect 675334 338948 675340 338950
rect 675404 338948 675451 338952
rect 675385 338947 675451 338948
rect 34470 338605 34530 338844
rect 34421 338600 34530 338605
rect 34421 338544 34426 338600
rect 34482 338544 34530 338600
rect 34421 338542 34530 338544
rect 34421 338539 34487 338542
rect 46013 338466 46079 338469
rect 41492 338464 46079 338466
rect 41492 338408 46018 338464
rect 46074 338408 46079 338464
rect 41492 338406 46079 338408
rect 46013 338403 46079 338406
rect 651465 338330 651531 338333
rect 650164 338328 651531 338330
rect 650164 338272 651470 338328
rect 651526 338272 651531 338328
rect 650164 338270 651531 338272
rect 651465 338267 651531 338270
rect 672901 338058 672967 338061
rect 675109 338058 675175 338061
rect 672901 338056 675175 338058
rect 41462 337788 41522 338028
rect 672901 338000 672906 338056
rect 672962 338000 675114 338056
rect 675170 338000 675175 338056
rect 672901 337998 675175 338000
rect 672901 337995 672967 337998
rect 675109 337995 675175 337998
rect 675569 337788 675635 337789
rect 41454 337724 41460 337788
rect 41524 337724 41530 337788
rect 675518 337786 675524 337788
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 41278 337514 41338 337620
rect 42926 337514 42932 337516
rect 41278 337454 42932 337514
rect 42926 337452 42932 337454
rect 42996 337452 43002 337516
rect 43110 337242 43116 337244
rect 41492 337182 43116 337242
rect 43110 337180 43116 337182
rect 43180 337180 43186 337244
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 40542 336564 40602 336804
rect 673545 336698 673611 336701
rect 675109 336698 675175 336701
rect 673545 336696 675175 336698
rect 673545 336640 673550 336696
rect 673606 336640 675114 336696
rect 675170 336640 675175 336696
rect 673545 336638 675175 336640
rect 673545 336635 673611 336638
rect 675109 336635 675175 336638
rect 675753 336698 675819 336701
rect 676438 336698 676444 336700
rect 675753 336696 676444 336698
rect 675753 336640 675758 336696
rect 675814 336640 676444 336696
rect 675753 336638 676444 336640
rect 675753 336635 675819 336638
rect 676438 336636 676444 336638
rect 676508 336636 676514 336700
rect 40534 336500 40540 336564
rect 40604 336500 40610 336564
rect 43294 336426 43300 336428
rect 41492 336366 43300 336426
rect 43294 336364 43300 336366
rect 43364 336364 43370 336428
rect 34421 336154 34487 336157
rect 41822 336154 41828 336156
rect 34421 336152 41828 336154
rect 34421 336096 34426 336152
rect 34482 336096 41828 336152
rect 34421 336094 41828 336096
rect 34421 336091 34487 336094
rect 41822 336092 41828 336094
rect 41892 336092 41898 336156
rect 41462 335746 41522 335988
rect 42742 335746 42748 335748
rect 41462 335686 42748 335746
rect 42742 335684 42748 335686
rect 42812 335684 42818 335748
rect 40726 335340 40786 335580
rect 40718 335276 40724 335340
rect 40788 335276 40794 335340
rect 41462 334930 41522 335172
rect 41462 334870 43914 334930
rect 41462 334658 41522 334764
rect 41462 334598 42258 334658
rect 42198 334386 42258 334598
rect 42742 334596 42748 334660
rect 42812 334658 42818 334660
rect 43069 334658 43135 334661
rect 42812 334656 43135 334658
rect 42812 334600 43074 334656
rect 43130 334600 43135 334656
rect 42812 334598 43135 334600
rect 42812 334596 42818 334598
rect 43069 334595 43135 334598
rect 43294 334596 43300 334660
rect 43364 334658 43370 334660
rect 43621 334658 43687 334661
rect 43364 334656 43687 334658
rect 43364 334600 43626 334656
rect 43682 334600 43687 334656
rect 43364 334598 43687 334600
rect 43854 334658 43914 334870
rect 44265 334658 44331 334661
rect 43854 334656 44331 334658
rect 43854 334600 44270 334656
rect 44326 334600 44331 334656
rect 43854 334598 44331 334600
rect 43364 334596 43370 334598
rect 43621 334595 43687 334598
rect 44265 334595 44331 334598
rect 42793 334386 42859 334389
rect 42198 334384 42859 334386
rect 41462 334114 41522 334356
rect 42198 334328 42798 334384
rect 42854 334328 42859 334384
rect 42198 334326 42859 334328
rect 42793 334323 42859 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 672165 333978 672231 333981
rect 675293 333978 675359 333981
rect 672165 333976 675359 333978
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 672165 333920 672170 333976
rect 672226 333920 675298 333976
rect 675354 333920 675359 333976
rect 672165 333918 675359 333920
rect 672165 333915 672231 333918
rect 675293 333915 675359 333918
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 674373 332754 674439 332757
rect 675109 332754 675175 332757
rect 674373 332752 675175 332754
rect 674373 332696 674378 332752
rect 674434 332696 675114 332752
rect 675170 332696 675175 332752
rect 674373 332694 675175 332696
rect 674373 332691 674439 332694
rect 675109 332691 675175 332694
rect 671981 332346 672047 332349
rect 675109 332346 675175 332349
rect 671981 332344 675175 332346
rect 671981 332288 671986 332344
rect 672042 332288 675114 332344
rect 675170 332288 675175 332344
rect 671981 332286 675175 332288
rect 671981 332283 672047 332286
rect 675109 332283 675175 332286
rect 675753 332346 675819 332349
rect 676254 332346 676260 332348
rect 675753 332344 676260 332346
rect 675753 332288 675758 332344
rect 675814 332288 676260 332344
rect 675753 332286 676260 332288
rect 675753 332283 675819 332286
rect 676254 332284 676260 332286
rect 676324 332284 676330 332348
rect 673729 331122 673795 331125
rect 675109 331122 675175 331125
rect 673729 331120 675175 331122
rect 673729 331064 673734 331120
rect 673790 331064 675114 331120
rect 675170 331064 675175 331120
rect 673729 331062 675175 331064
rect 673729 331059 673795 331062
rect 675109 331059 675175 331062
rect 37917 328402 37983 328405
rect 41638 328402 41644 328404
rect 37917 328400 41644 328402
rect 37917 328344 37922 328400
rect 37978 328344 41644 328400
rect 37917 328342 41644 328344
rect 37917 328339 37983 328342
rect 41638 328340 41644 328342
rect 41708 328340 41714 328404
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 672349 327586 672415 327589
rect 675109 327586 675175 327589
rect 672349 327584 675175 327586
rect 672349 327528 672354 327584
rect 672410 327528 675114 327584
rect 675170 327528 675175 327584
rect 672349 327526 675175 327528
rect 672349 327523 672415 327526
rect 675109 327523 675175 327526
rect 41454 326708 41460 326772
rect 41524 326770 41530 326772
rect 41781 326770 41847 326773
rect 41524 326768 41847 326770
rect 41524 326712 41786 326768
rect 41842 326712 41847 326768
rect 41524 326710 41847 326712
rect 41524 326708 41530 326710
rect 41781 326707 41847 326710
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41454 324804 41460 324868
rect 41524 324866 41530 324868
rect 41781 324866 41847 324869
rect 41524 324864 41847 324866
rect 41524 324808 41786 324864
rect 41842 324808 41847 324864
rect 41524 324806 41847 324808
rect 41524 324804 41530 324806
rect 41781 324803 41847 324806
rect 43437 323098 43503 323101
rect 43437 323096 45570 323098
rect 43437 323040 43442 323096
rect 43498 323040 45570 323096
rect 43437 323038 45570 323040
rect 43437 323035 43503 323038
rect 45510 322962 45570 323038
rect 64462 322962 64522 324156
rect 45510 322902 64522 322962
rect 42057 322826 42123 322829
rect 43621 322826 43687 322829
rect 42057 322824 43687 322826
rect 42057 322768 42062 322824
rect 42118 322768 43626 322824
rect 43682 322768 43687 322824
rect 42057 322766 43687 322768
rect 42057 322763 42123 322766
rect 43621 322763 43687 322766
rect 42425 321466 42491 321469
rect 53097 321466 53163 321469
rect 42425 321464 53163 321466
rect 42425 321408 42430 321464
rect 42486 321408 53102 321464
rect 53158 321408 53163 321464
rect 42425 321406 53163 321408
rect 42425 321403 42491 321406
rect 53097 321403 53163 321406
rect 42425 320106 42491 320109
rect 44265 320106 44331 320109
rect 42425 320104 44331 320106
rect 42425 320048 42430 320104
rect 42486 320048 44270 320104
rect 44326 320048 44331 320104
rect 42425 320046 44331 320048
rect 42425 320043 42491 320046
rect 44265 320043 44331 320046
rect 42425 319426 42491 319429
rect 46013 319426 46079 319429
rect 42425 319424 46079 319426
rect 42425 319368 42430 319424
rect 42486 319368 46018 319424
rect 46074 319368 46079 319424
rect 42425 319366 46079 319368
rect 42425 319363 42491 319366
rect 46013 319363 46079 319366
rect 40718 317460 40724 317524
rect 40788 317522 40794 317524
rect 42241 317522 42307 317525
rect 40788 317520 42307 317522
rect 40788 317464 42246 317520
rect 42302 317464 42307 317520
rect 40788 317462 42307 317464
rect 40788 317460 40794 317462
rect 42241 317459 42307 317462
rect 40534 316644 40540 316708
rect 40604 316706 40610 316708
rect 41781 316706 41847 316709
rect 40604 316704 41847 316706
rect 40604 316648 41786 316704
rect 41842 316648 41847 316704
rect 40604 316646 41847 316648
rect 40604 316644 40610 316646
rect 41781 316643 41847 316646
rect 42149 316026 42215 316029
rect 43110 316026 43116 316028
rect 42149 316024 43116 316026
rect 42149 315968 42154 316024
rect 42210 315968 43116 316024
rect 42149 315966 43116 315968
rect 42149 315963 42215 315966
rect 43110 315964 43116 315966
rect 43180 315964 43186 316028
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 663057 315482 663123 315485
rect 676029 315482 676095 315485
rect 663057 315480 676095 315482
rect 663057 315424 663062 315480
rect 663118 315424 676034 315480
rect 676090 315424 676095 315480
rect 663057 315422 676095 315424
rect 663057 315419 663123 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 45829 313714 45895 313717
rect 42149 313712 45895 313714
rect 42149 313656 42154 313712
rect 42210 313656 45834 313712
rect 45890 313656 45895 313712
rect 42149 313654 45895 313656
rect 42149 313651 42215 313654
rect 45829 313651 45895 313654
rect 667197 313714 667263 313717
rect 667197 313712 676292 313714
rect 667197 313656 667202 313712
rect 667258 313656 676292 313712
rect 667197 313654 676292 313656
rect 667197 313651 667263 313654
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 669270 312838 676292 312898
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 42149 312354 42215 312357
rect 45645 312354 45711 312357
rect 42149 312352 45711 312354
rect 42149 312296 42154 312352
rect 42210 312296 45650 312352
rect 45706 312296 45711 312352
rect 42149 312294 45711 312296
rect 42149 312291 42215 312294
rect 45645 312291 45711 312294
rect 668577 311946 668643 311949
rect 669270 311946 669330 312838
rect 673269 312490 673335 312493
rect 673269 312488 676292 312490
rect 673269 312432 673274 312488
rect 673330 312432 676292 312488
rect 673269 312430 676292 312432
rect 673269 312427 673335 312430
rect 672901 312082 672967 312085
rect 672901 312080 676292 312082
rect 672901 312024 672906 312080
rect 672962 312024 676292 312080
rect 672901 312022 676292 312024
rect 672901 312019 672967 312022
rect 668577 311944 669330 311946
rect 668577 311888 668582 311944
rect 668638 311888 669330 311944
rect 668577 311886 669330 311888
rect 668577 311883 668643 311886
rect 651465 311810 651531 311813
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 651465 311747 651531 311750
rect 673913 311674 673979 311677
rect 673913 311672 676292 311674
rect 673913 311616 673918 311672
rect 673974 311616 676292 311672
rect 673913 311614 676292 311616
rect 673913 311611 673979 311614
rect 44173 311538 44239 311541
rect 44582 311538 44588 311540
rect 44173 311536 44588 311538
rect 44173 311480 44178 311536
rect 44234 311480 44588 311536
rect 44173 311478 44588 311480
rect 44173 311475 44239 311478
rect 44582 311476 44588 311478
rect 44652 311476 44658 311540
rect 44357 311268 44423 311269
rect 44357 311264 44404 311268
rect 44468 311266 44474 311268
rect 673085 311266 673151 311269
rect 44357 311208 44362 311264
rect 44357 311204 44404 311208
rect 44468 311206 44514 311266
rect 673085 311264 676292 311266
rect 673085 311208 673090 311264
rect 673146 311208 676292 311264
rect 673085 311206 676292 311208
rect 44468 311204 44474 311206
rect 44357 311203 44423 311204
rect 673085 311203 673151 311206
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 62113 311067 62179 311070
rect 673269 310858 673335 310861
rect 673269 310856 676292 310858
rect 673269 310800 673274 310856
rect 673330 310800 676292 310856
rect 673269 310798 676292 310800
rect 673269 310795 673335 310798
rect 673821 310450 673887 310453
rect 673821 310448 676292 310450
rect 673821 310392 673826 310448
rect 673882 310392 676292 310448
rect 673821 310390 676292 310392
rect 673821 310387 673887 310390
rect 672533 310042 672599 310045
rect 672533 310040 676292 310042
rect 672533 309984 672538 310040
rect 672594 309984 676292 310040
rect 672533 309982 676292 309984
rect 672533 309979 672599 309982
rect 674649 309634 674715 309637
rect 674649 309632 676292 309634
rect 674649 309576 674654 309632
rect 674710 309576 676292 309632
rect 674649 309574 676292 309576
rect 674649 309571 674715 309574
rect 675017 309226 675083 309229
rect 675017 309224 676292 309226
rect 675017 309168 675022 309224
rect 675078 309168 676292 309224
rect 675017 309166 676292 309168
rect 675017 309163 675083 309166
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 676029 308002 676095 308005
rect 676029 308000 676292 308002
rect 676029 307944 676034 308000
rect 676090 307944 676292 308000
rect 676029 307942 676292 307944
rect 676029 307939 676095 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 675886 306716 675892 306780
rect 675956 306778 675962 306780
rect 675956 306718 676292 306778
rect 675956 306716 675962 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 676489 305962 676555 305965
rect 676476 305960 676555 305962
rect 676476 305904 676494 305960
rect 676550 305904 676555 305960
rect 676476 305902 676555 305904
rect 676489 305899 676555 305902
rect 674465 305554 674531 305557
rect 674465 305552 676292 305554
rect 674465 305496 674470 305552
rect 674526 305496 676292 305552
rect 674465 305494 676292 305496
rect 674465 305491 674531 305494
rect 676673 305146 676739 305149
rect 676660 305144 676739 305146
rect 676660 305088 676678 305144
rect 676734 305088 676739 305144
rect 676660 305086 676739 305088
rect 676673 305083 676739 305086
rect 674741 304738 674807 304741
rect 674741 304736 676292 304738
rect 674741 304680 674746 304736
rect 674802 304680 676292 304736
rect 674741 304678 676292 304680
rect 674741 304675 674807 304678
rect 673361 304330 673427 304333
rect 673361 304328 676292 304330
rect 673361 304272 673366 304328
rect 673422 304272 676292 304328
rect 673361 304270 676292 304272
rect 673361 304267 673427 304270
rect 674238 303998 676230 304058
rect 674238 303925 674298 303998
rect 674189 303920 674298 303925
rect 674189 303864 674194 303920
rect 674250 303864 674298 303920
rect 674189 303862 674298 303864
rect 676170 303922 676230 303998
rect 676170 303862 676292 303922
rect 674189 303859 674255 303862
rect 675201 303786 675267 303789
rect 676029 303786 676095 303789
rect 675201 303784 676095 303786
rect 675201 303728 675206 303784
rect 675262 303728 676034 303784
rect 676090 303728 676095 303784
rect 675201 303726 676095 303728
rect 675201 303723 675267 303726
rect 676029 303723 676095 303726
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 41781 303106 41847 303109
rect 46381 303106 46447 303109
rect 41781 303104 46447 303106
rect 41781 303048 41786 303104
rect 41842 303048 46386 303104
rect 46442 303048 46447 303104
rect 41781 303046 46447 303048
rect 41781 303043 41847 303046
rect 46381 303043 46447 303046
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 669221 302290 669287 302293
rect 669221 302288 676292 302290
rect 669221 302232 669226 302288
rect 669282 302232 676292 302288
rect 669221 302230 676292 302232
rect 669221 302227 669287 302230
rect 674833 302018 674899 302021
rect 675201 302018 675267 302021
rect 674833 302016 675267 302018
rect 674833 301960 674838 302016
rect 674894 301960 675206 302016
rect 675262 301960 675267 302016
rect 674833 301958 675267 301960
rect 674833 301955 674899 301958
rect 675201 301955 675267 301958
rect 676489 301612 676555 301613
rect 676438 301610 676444 301612
rect 676398 301550 676444 301610
rect 676508 301608 676555 301612
rect 676550 301552 676555 301608
rect 676438 301548 676444 301550
rect 676508 301548 676555 301552
rect 676489 301547 676555 301548
rect 672441 301474 672507 301477
rect 676029 301474 676095 301477
rect 676673 301476 676739 301477
rect 672441 301472 676095 301474
rect 672441 301416 672446 301472
rect 672502 301416 676034 301472
rect 676090 301416 676095 301472
rect 672441 301414 676095 301416
rect 672441 301411 672507 301414
rect 676029 301411 676095 301414
rect 676622 301412 676628 301476
rect 676692 301474 676739 301476
rect 676692 301472 676784 301474
rect 676734 301416 676784 301472
rect 676692 301414 676784 301416
rect 676692 301412 676739 301414
rect 676673 301411 676739 301412
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44357 300114 44423 300117
rect 41492 300112 44423 300114
rect 41492 300056 44362 300112
rect 44418 300056 44423 300112
rect 41492 300054 44423 300056
rect 44357 300051 44423 300054
rect 42885 299706 42951 299709
rect 41492 299704 42951 299706
rect 41492 299648 42890 299704
rect 42946 299648 42951 299704
rect 41492 299646 42951 299648
rect 42885 299643 42951 299646
rect 44173 299298 44239 299301
rect 41492 299296 44239 299298
rect 41492 299240 44178 299296
rect 44234 299240 44239 299296
rect 41492 299238 44239 299240
rect 44173 299235 44239 299238
rect 43253 298890 43319 298893
rect 41492 298888 43319 298890
rect 41492 298832 43258 298888
rect 43314 298832 43319 298888
rect 41492 298830 43319 298832
rect 43253 298827 43319 298830
rect 45461 298482 45527 298485
rect 652201 298482 652267 298485
rect 41492 298480 45527 298482
rect 41492 298424 45466 298480
rect 45522 298424 45527 298480
rect 41492 298422 45527 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 45461 298419 45527 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 44173 298074 44239 298077
rect 41492 298072 44239 298074
rect 41492 298016 44178 298072
rect 44234 298016 44239 298072
rect 41492 298014 44239 298016
rect 44173 298011 44239 298014
rect 675702 298012 675708 298076
rect 675772 298074 675778 298076
rect 678237 298074 678303 298077
rect 675772 298072 678303 298074
rect 675772 298016 678242 298072
rect 678298 298016 678303 298072
rect 675772 298014 678303 298016
rect 675772 298012 675778 298014
rect 678237 298011 678303 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 45001 297258 45067 297261
rect 41492 297256 45067 297258
rect 41492 297200 45006 297256
rect 45062 297200 45067 297256
rect 41492 297198 45067 297200
rect 45001 297195 45067 297198
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 675385 296578 675451 296581
rect 676029 296578 676095 296581
rect 675385 296576 676095 296578
rect 675385 296520 675390 296576
rect 675446 296520 676034 296576
rect 676090 296520 676095 296576
rect 675385 296518 676095 296520
rect 675385 296515 675451 296518
rect 676029 296515 676095 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 41321 296034 41387 296037
rect 41308 296032 41387 296034
rect 41308 295976 41326 296032
rect 41382 295976 41387 296032
rect 41308 295974 41387 295976
rect 41321 295971 41387 295974
rect 674833 295898 674899 295901
rect 675477 295898 675543 295901
rect 674833 295896 675543 295898
rect 674833 295840 674838 295896
rect 674894 295840 675482 295896
rect 675538 295840 675543 295896
rect 674833 295838 675543 295840
rect 674833 295835 674899 295838
rect 675477 295835 675543 295838
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 43069 295218 43135 295221
rect 41492 295216 43135 295218
rect 41492 295160 43074 295216
rect 43130 295160 43135 295216
rect 41492 295158 43135 295160
rect 43069 295155 43135 295158
rect 675753 295218 675819 295221
rect 676254 295218 676260 295220
rect 675753 295216 676260 295218
rect 675753 295160 675758 295216
rect 675814 295160 676260 295216
rect 675753 295158 676260 295160
rect 675753 295155 675819 295158
rect 676254 295156 676260 295158
rect 676324 295156 676330 295220
rect 32397 294810 32463 294813
rect 32397 294808 32476 294810
rect 32397 294752 32402 294808
rect 32458 294752 32476 294808
rect 32397 294750 32476 294752
rect 32397 294747 32463 294750
rect 674925 294538 674991 294541
rect 675477 294538 675543 294541
rect 674925 294536 675543 294538
rect 674925 294480 674930 294536
rect 674986 294480 675482 294536
rect 675538 294480 675543 294536
rect 674925 294478 675543 294480
rect 674925 294475 674991 294478
rect 675477 294475 675543 294478
rect 44357 294402 44423 294405
rect 41492 294400 44423 294402
rect 41492 294344 44362 294400
rect 44418 294344 44423 294400
rect 41492 294342 44423 294344
rect 44357 294339 44423 294342
rect 43621 293994 43687 293997
rect 41492 293992 43687 293994
rect 41492 293936 43626 293992
rect 43682 293936 43687 293992
rect 41492 293934 43687 293936
rect 43621 293931 43687 293934
rect 44633 293586 44699 293589
rect 41492 293584 44699 293586
rect 41492 293528 44638 293584
rect 44694 293528 44699 293584
rect 41492 293526 44699 293528
rect 44633 293523 44699 293526
rect 43989 293178 44055 293181
rect 41492 293176 44055 293178
rect 41492 293120 43994 293176
rect 44050 293120 44055 293176
rect 41492 293118 44055 293120
rect 43989 293115 44055 293118
rect 675017 292770 675083 292773
rect 675477 292770 675543 292773
rect 675017 292768 675543 292770
rect 40910 292592 40970 292740
rect 675017 292712 675022 292768
rect 675078 292712 675482 292768
rect 675538 292712 675543 292768
rect 675017 292710 675543 292712
rect 675017 292707 675083 292710
rect 675477 292707 675543 292710
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40542 292332 40602 292528
rect 41781 292500 41847 292501
rect 41781 292496 41828 292500
rect 41892 292498 41898 292500
rect 41781 292440 41786 292496
rect 41781 292436 41828 292440
rect 41892 292438 41938 292498
rect 41892 292436 41898 292438
rect 41781 292435 41847 292436
rect 43805 291954 43871 291957
rect 41492 291952 43871 291954
rect 41492 291896 43810 291952
rect 43866 291896 43871 291952
rect 41492 291894 43871 291896
rect 43805 291891 43871 291894
rect 45185 291682 45251 291685
rect 41830 291680 45251 291682
rect 41830 291624 45190 291680
rect 45246 291624 45251 291680
rect 41830 291622 45251 291624
rect 41830 291546 41890 291622
rect 45185 291619 45251 291622
rect 41492 291486 41890 291546
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 41492 291078 51090 291138
rect 46197 290730 46263 290733
rect 41492 290728 46263 290730
rect 41492 290672 46202 290728
rect 46258 290672 46263 290728
rect 41492 290670 46263 290672
rect 46197 290667 46263 290670
rect 41781 290460 41847 290461
rect 41781 290456 41828 290460
rect 41892 290458 41898 290460
rect 41781 290400 41786 290456
rect 41781 290396 41828 290400
rect 41892 290398 41938 290458
rect 41892 290396 41898 290398
rect 41781 290395 41847 290396
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 49141 289914 49207 289917
rect 41492 289912 49207 289914
rect 41492 289856 49146 289912
rect 49202 289856 49207 289912
rect 41492 289854 49207 289856
rect 51030 289914 51090 291078
rect 674741 291002 674807 291005
rect 675385 291002 675451 291005
rect 674741 291000 675451 291002
rect 674741 290944 674746 291000
rect 674802 290944 675390 291000
rect 675446 290944 675451 291000
rect 674741 290942 675451 290944
rect 674741 290939 674807 290942
rect 675385 290939 675451 290942
rect 51717 289914 51783 289917
rect 51030 289912 51783 289914
rect 51030 289856 51722 289912
rect 51778 289856 51783 289912
rect 51030 289854 51783 289856
rect 49141 289851 49207 289854
rect 51717 289851 51783 289854
rect 673361 287874 673427 287877
rect 675109 287874 675175 287877
rect 673361 287872 675175 287874
rect 673361 287816 673366 287872
rect 673422 287816 675114 287872
rect 675170 287816 675175 287872
rect 673361 287814 675175 287816
rect 673361 287811 673427 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676622 287058 676628 287060
rect 675753 287056 676628 287058
rect 675753 287000 675758 287056
rect 675814 287000 676628 287056
rect 675753 286998 676628 287000
rect 675753 286995 675819 286998
rect 676622 286996 676628 286998
rect 676692 286996 676698 287060
rect 674281 286514 674347 286517
rect 675385 286514 675451 286517
rect 674281 286512 675451 286514
rect 674281 286456 674286 286512
rect 674342 286456 675390 286512
rect 675446 286456 675451 286512
rect 674281 286454 675451 286456
rect 674281 286451 674347 286454
rect 675385 286451 675451 286454
rect 674465 285562 674531 285565
rect 675477 285562 675543 285565
rect 674465 285560 675543 285562
rect 674465 285504 674470 285560
rect 674526 285504 675482 285560
rect 675538 285504 675543 285560
rect 674465 285502 675543 285504
rect 674465 285499 674531 285502
rect 675477 285499 675543 285502
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62941 285154 63007 285157
rect 62941 285152 64492 285154
rect 62941 285096 62946 285152
rect 63002 285096 64492 285152
rect 62941 285094 64492 285096
rect 62941 285091 63007 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 42149 279850 42215 279853
rect 43989 279850 44055 279853
rect 42149 279848 44055 279850
rect 42149 279792 42154 279848
rect 42210 279792 43994 279848
rect 44050 279792 44055 279848
rect 42149 279790 44055 279792
rect 42149 279787 42215 279790
rect 43989 279787 44055 279790
rect 42425 278762 42491 278765
rect 55857 278762 55923 278765
rect 42425 278760 55923 278762
rect 42425 278704 42430 278760
rect 42486 278704 55862 278760
rect 55918 278704 55923 278760
rect 42425 278702 55923 278704
rect 42425 278699 42491 278702
rect 55857 278699 55923 278702
rect 40718 278428 40724 278492
rect 40788 278490 40794 278492
rect 42333 278490 42399 278493
rect 40788 278488 42399 278490
rect 40788 278432 42338 278488
rect 42394 278432 42399 278488
rect 40788 278430 42399 278432
rect 40788 278428 40794 278430
rect 42333 278427 42399 278430
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 41781 277946 41847 277949
rect 40972 277944 41847 277946
rect 40972 277888 41786 277944
rect 41842 277888 41847 277944
rect 40972 277886 41847 277888
rect 40972 277884 40978 277886
rect 41781 277883 41847 277886
rect 42149 277946 42215 277949
rect 45185 277946 45251 277949
rect 42149 277944 45251 277946
rect 42149 277888 42154 277944
rect 42210 277888 45190 277944
rect 45246 277888 45251 277944
rect 42149 277886 45251 277888
rect 42149 277883 42215 277886
rect 45185 277883 45251 277886
rect 42057 277130 42123 277133
rect 43805 277130 43871 277133
rect 42057 277128 43871 277130
rect 42057 277072 42062 277128
rect 42118 277072 43810 277128
rect 43866 277072 43871 277128
rect 42057 277070 43871 277072
rect 42057 277067 42123 277070
rect 43805 277067 43871 277070
rect 42057 276586 42123 276589
rect 43069 276586 43135 276589
rect 42057 276584 43135 276586
rect 42057 276528 42062 276584
rect 42118 276528 43074 276584
rect 43130 276528 43135 276584
rect 42057 276526 43135 276528
rect 42057 276523 42123 276526
rect 43069 276523 43135 276526
rect 525517 275770 525583 275773
rect 527725 275770 527791 275773
rect 525517 275768 527791 275770
rect 525517 275712 525522 275768
rect 525578 275712 527730 275768
rect 527786 275712 527791 275768
rect 525517 275710 527791 275712
rect 525517 275707 525583 275710
rect 527725 275707 527791 275710
rect 535269 275362 535335 275365
rect 538857 275362 538923 275365
rect 535269 275360 538923 275362
rect 535269 275304 535274 275360
rect 535330 275304 538862 275360
rect 538918 275304 538923 275360
rect 535269 275302 538923 275304
rect 535269 275299 535335 275302
rect 538857 275299 538923 275302
rect 538213 275090 538279 275093
rect 544193 275090 544259 275093
rect 538213 275088 544259 275090
rect 538213 275032 538218 275088
rect 538274 275032 544198 275088
rect 544254 275032 544259 275088
rect 538213 275030 544259 275032
rect 538213 275027 538279 275030
rect 544193 275027 544259 275030
rect 530761 274954 530827 274957
rect 534165 274954 534231 274957
rect 530761 274952 534231 274954
rect 530761 274896 530766 274952
rect 530822 274896 534170 274952
rect 534226 274896 534231 274952
rect 530761 274894 534231 274896
rect 530761 274891 530827 274894
rect 534165 274891 534231 274894
rect 544377 274954 544443 274957
rect 546033 274954 546099 274957
rect 544377 274952 546099 274954
rect 544377 274896 544382 274952
rect 544438 274896 546038 274952
rect 546094 274896 546099 274952
rect 544377 274894 546099 274896
rect 544377 274891 544443 274894
rect 546033 274891 546099 274894
rect 538213 274682 538279 274685
rect 543181 274682 543247 274685
rect 538213 274680 543247 274682
rect 538213 274624 538218 274680
rect 538274 274624 543186 274680
rect 543242 274624 543247 274680
rect 538213 274622 543247 274624
rect 538213 274619 538279 274622
rect 543181 274619 543247 274622
rect 528507 274410 528573 274413
rect 537937 274410 538003 274413
rect 528507 274408 538003 274410
rect 528507 274352 528512 274408
rect 528568 274352 537942 274408
rect 537998 274352 538003 274408
rect 528507 274350 538003 274352
rect 528507 274347 528573 274350
rect 537937 274347 538003 274350
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 528093 274138 528159 274141
rect 528645 274138 528711 274141
rect 528093 274136 528711 274138
rect 528093 274080 528098 274136
rect 528154 274080 528650 274136
rect 528706 274080 528711 274136
rect 528093 274078 528711 274080
rect 528093 274075 528159 274078
rect 528645 274075 528711 274078
rect 538121 274138 538187 274141
rect 538305 274138 538371 274141
rect 538121 274136 538371 274138
rect 538121 274080 538126 274136
rect 538182 274080 538310 274136
rect 538366 274080 538371 274136
rect 538121 274078 538371 274080
rect 538121 274075 538187 274078
rect 538305 274075 538371 274078
rect 513189 274002 513255 274005
rect 514109 274002 514175 274005
rect 513189 274000 514175 274002
rect 513189 273944 513194 274000
rect 513250 273944 514114 274000
rect 514170 273944 514175 274000
rect 513189 273942 514175 273944
rect 513189 273939 513255 273942
rect 514109 273939 514175 273942
rect 521101 274002 521167 274005
rect 524045 274002 524111 274005
rect 521101 274000 524111 274002
rect 521101 273944 521106 274000
rect 521162 273944 524050 274000
rect 524106 273944 524111 274000
rect 521101 273942 524111 273944
rect 521101 273939 521167 273942
rect 524045 273939 524111 273942
rect 538857 273866 538923 273869
rect 635641 273866 635707 273869
rect 538857 273864 635707 273866
rect 538857 273808 538862 273864
rect 538918 273808 635646 273864
rect 635702 273808 635707 273864
rect 538857 273806 635707 273808
rect 538857 273803 538923 273806
rect 635641 273803 635707 273806
rect 42057 273458 42123 273461
rect 44633 273458 44699 273461
rect 42057 273456 44699 273458
rect 42057 273400 42062 273456
rect 42118 273400 44638 273456
rect 44694 273400 44699 273456
rect 42057 273398 44699 273400
rect 42057 273395 42123 273398
rect 44633 273395 44699 273398
rect 42057 273050 42123 273053
rect 43621 273050 43687 273053
rect 42057 273048 43687 273050
rect 42057 272992 42062 273048
rect 42118 272992 43626 273048
rect 43682 272992 43687 273048
rect 42057 272990 43687 272992
rect 42057 272987 42123 272990
rect 43621 272987 43687 272990
rect 527909 272914 527975 272917
rect 528645 272914 528711 272917
rect 527909 272912 528711 272914
rect 527909 272856 527914 272912
rect 527970 272856 528650 272912
rect 528706 272856 528711 272912
rect 527909 272854 528711 272856
rect 527909 272851 527975 272854
rect 528645 272851 528711 272854
rect 538213 272778 538279 272781
rect 545113 272778 545179 272781
rect 538213 272776 545179 272778
rect 538213 272720 538218 272776
rect 538274 272720 545118 272776
rect 545174 272720 545179 272776
rect 538213 272718 545179 272720
rect 538213 272715 538279 272718
rect 545113 272715 545179 272718
rect 521469 272506 521535 272509
rect 528369 272506 528435 272509
rect 521469 272504 528435 272506
rect 521469 272448 521474 272504
rect 521530 272448 528374 272504
rect 528430 272448 528435 272504
rect 521469 272446 528435 272448
rect 521469 272443 521535 272446
rect 528369 272443 528435 272446
rect 528553 272506 528619 272509
rect 531681 272506 531747 272509
rect 528553 272504 531747 272506
rect 528553 272448 528558 272504
rect 528614 272448 531686 272504
rect 531742 272448 531747 272504
rect 528553 272446 531747 272448
rect 528553 272443 528619 272446
rect 531681 272443 531747 272446
rect 540697 272506 540763 272509
rect 626441 272506 626507 272509
rect 540697 272504 626507 272506
rect 540697 272448 540702 272504
rect 540758 272448 626446 272504
rect 626502 272448 626507 272504
rect 540697 272446 626507 272448
rect 540697 272443 540763 272446
rect 626441 272443 626507 272446
rect 533705 272234 533771 272237
rect 538305 272234 538371 272237
rect 533705 272232 538371 272234
rect 533705 272176 533710 272232
rect 533766 272176 538310 272232
rect 538366 272176 538371 272232
rect 533705 272174 538371 272176
rect 533705 272171 533771 272174
rect 538305 272171 538371 272174
rect 519721 271690 519787 271693
rect 525885 271690 525951 271693
rect 519721 271688 525951 271690
rect 519721 271632 519726 271688
rect 519782 271632 525890 271688
rect 525946 271632 525951 271688
rect 519721 271630 525951 271632
rect 519721 271627 519787 271630
rect 525885 271627 525951 271630
rect 523493 271418 523559 271421
rect 525701 271418 525767 271421
rect 523493 271416 525767 271418
rect 523493 271360 523498 271416
rect 523554 271360 525706 271416
rect 525762 271360 525767 271416
rect 523493 271358 525767 271360
rect 523493 271355 523559 271358
rect 525701 271355 525767 271358
rect 529841 271418 529907 271421
rect 538029 271418 538095 271421
rect 529841 271416 538095 271418
rect 529841 271360 529846 271416
rect 529902 271360 538034 271416
rect 538090 271360 538095 271416
rect 529841 271358 538095 271360
rect 529841 271355 529907 271358
rect 538029 271355 538095 271358
rect 514293 271282 514359 271285
rect 518341 271282 518407 271285
rect 514293 271280 518407 271282
rect 514293 271224 514298 271280
rect 514354 271224 518346 271280
rect 518402 271224 518407 271280
rect 514293 271222 518407 271224
rect 514293 271219 514359 271222
rect 518341 271219 518407 271222
rect 524137 271146 524203 271149
rect 617977 271146 618043 271149
rect 524137 271144 618043 271146
rect 524137 271088 524142 271144
rect 524198 271088 617982 271144
rect 618038 271088 618043 271144
rect 524137 271086 618043 271088
rect 524137 271083 524203 271086
rect 617977 271083 618043 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 480253 270738 480319 270741
rect 483105 270738 483171 270741
rect 480253 270736 483171 270738
rect 480253 270680 480258 270736
rect 480314 270680 483110 270736
rect 483166 270680 483171 270736
rect 480253 270678 483171 270680
rect 480253 270675 480319 270678
rect 483105 270675 483171 270678
rect 504909 270602 504975 270605
rect 507853 270602 507919 270605
rect 504909 270600 507919 270602
rect 504909 270544 504914 270600
rect 504970 270544 507858 270600
rect 507914 270544 507919 270600
rect 504909 270542 507919 270544
rect 504909 270539 504975 270542
rect 507853 270539 507919 270542
rect 536097 270602 536163 270605
rect 537845 270602 537911 270605
rect 536097 270600 537911 270602
rect 536097 270544 536102 270600
rect 536158 270544 537850 270600
rect 537906 270544 537911 270600
rect 536097 270542 537911 270544
rect 536097 270539 536163 270542
rect 537845 270539 537911 270542
rect 538029 270602 538095 270605
rect 539593 270602 539659 270605
rect 538029 270600 539659 270602
rect 538029 270544 538034 270600
rect 538090 270544 539598 270600
rect 539654 270544 539659 270600
rect 538029 270542 539659 270544
rect 538029 270539 538095 270542
rect 539593 270539 539659 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 42425 270466 42491 270469
rect 44357 270466 44423 270469
rect 42425 270464 44423 270466
rect 42425 270408 42430 270464
rect 42486 270408 44362 270464
rect 44418 270408 44423 270464
rect 42425 270406 44423 270408
rect 42425 270403 42491 270406
rect 44357 270403 44423 270406
rect 494237 270330 494303 270333
rect 574921 270330 574987 270333
rect 494237 270328 574987 270330
rect 494237 270272 494242 270328
rect 494298 270272 574926 270328
rect 574982 270272 574987 270328
rect 494237 270270 574987 270272
rect 494237 270267 494303 270270
rect 574921 270267 574987 270270
rect 482277 270058 482343 270061
rect 484577 270058 484643 270061
rect 532785 270058 532851 270061
rect 482277 270056 484643 270058
rect 482277 270000 482282 270056
rect 482338 270000 484582 270056
rect 484638 270000 484643 270056
rect 482277 269998 484643 270000
rect 482277 269995 482343 269998
rect 484577 269995 484643 269998
rect 528510 270056 532851 270058
rect 528510 270000 532790 270056
rect 532846 270000 532851 270056
rect 528510 269998 532851 270000
rect 136541 269786 136607 269789
rect 139945 269786 140011 269789
rect 136541 269784 140011 269786
rect 136541 269728 136546 269784
rect 136602 269728 139950 269784
rect 140006 269728 140011 269784
rect 136541 269726 140011 269728
rect 136541 269723 136607 269726
rect 139945 269723 140011 269726
rect 475745 269786 475811 269789
rect 478873 269786 478939 269789
rect 475745 269784 478939 269786
rect 475745 269728 475750 269784
rect 475806 269728 478878 269784
rect 478934 269728 478939 269784
rect 475745 269726 478939 269728
rect 475745 269723 475811 269726
rect 478873 269723 478939 269726
rect 504725 269786 504791 269789
rect 528510 269786 528570 269998
rect 532785 269995 532851 269998
rect 533061 270058 533127 270061
rect 630673 270058 630739 270061
rect 533061 270056 630739 270058
rect 533061 270000 533066 270056
rect 533122 270000 630678 270056
rect 630734 270000 630739 270056
rect 533061 269998 630739 270000
rect 533061 269995 533127 269998
rect 630673 269995 630739 269998
rect 504725 269784 528570 269786
rect 504725 269728 504730 269784
rect 504786 269728 528570 269784
rect 504725 269726 528570 269728
rect 531313 269786 531379 269789
rect 534717 269786 534783 269789
rect 531313 269784 534783 269786
rect 531313 269728 531318 269784
rect 531374 269728 534722 269784
rect 534778 269728 534783 269784
rect 531313 269726 534783 269728
rect 504725 269723 504791 269726
rect 531313 269723 531379 269726
rect 534717 269723 534783 269726
rect 538029 269786 538095 269789
rect 637573 269786 637639 269789
rect 538029 269784 637639 269786
rect 538029 269728 538034 269784
rect 538090 269728 637578 269784
rect 637634 269728 637639 269784
rect 538029 269726 637639 269728
rect 538029 269723 538095 269726
rect 637573 269723 637639 269726
rect 671337 269786 671403 269789
rect 676029 269786 676095 269789
rect 671337 269784 676095 269786
rect 671337 269728 671342 269784
rect 671398 269728 676034 269784
rect 676090 269728 676095 269784
rect 671337 269726 676095 269728
rect 671337 269723 671403 269726
rect 676029 269723 676095 269726
rect 475377 269514 475443 269517
rect 476297 269514 476363 269517
rect 475377 269512 476363 269514
rect 475377 269456 475382 269512
rect 475438 269456 476302 269512
rect 476358 269456 476363 269512
rect 475377 269454 476363 269456
rect 475377 269451 475443 269454
rect 476297 269451 476363 269454
rect 484301 269514 484367 269517
rect 490005 269514 490071 269517
rect 484301 269512 490071 269514
rect 484301 269456 484306 269512
rect 484362 269456 490010 269512
rect 490066 269456 490071 269512
rect 484301 269454 490071 269456
rect 484301 269451 484367 269454
rect 490005 269451 490071 269454
rect 537845 269514 537911 269517
rect 538397 269514 538463 269517
rect 537845 269512 538463 269514
rect 537845 269456 537850 269512
rect 537906 269456 538402 269512
rect 538458 269456 538463 269512
rect 537845 269454 538463 269456
rect 537845 269451 537911 269454
rect 538397 269451 538463 269454
rect 479057 269378 479123 269381
rect 480345 269378 480411 269381
rect 479057 269376 480411 269378
rect 479057 269320 479062 269376
rect 479118 269320 480350 269376
rect 480406 269320 480411 269376
rect 479057 269318 480411 269320
rect 479057 269315 479123 269318
rect 480345 269315 480411 269318
rect 541433 269378 541499 269381
rect 543549 269378 543615 269381
rect 541433 269376 543615 269378
rect 541433 269320 541438 269376
rect 541494 269320 543554 269376
rect 543610 269320 543615 269376
rect 541433 269318 543615 269320
rect 541433 269315 541499 269318
rect 543549 269315 543615 269318
rect 468753 269242 468819 269245
rect 476021 269242 476087 269245
rect 468753 269240 476087 269242
rect 468753 269184 468758 269240
rect 468814 269184 476026 269240
rect 476082 269184 476087 269240
rect 468753 269182 476087 269184
rect 468753 269179 468819 269182
rect 476021 269179 476087 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 538213 269106 538279 269109
rect 544377 269106 544443 269109
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 538213 269104 544443 269106
rect 538213 269048 538218 269104
rect 538274 269048 544382 269104
rect 544438 269048 544443 269104
rect 538213 269046 544443 269048
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 538213 269043 538279 269046
rect 544377 269043 544443 269046
rect 527173 268562 527239 268565
rect 528921 268562 528987 268565
rect 676262 268562 676322 268668
rect 527173 268560 528987 268562
rect 527173 268504 527178 268560
rect 527234 268504 528926 268560
rect 528982 268504 528987 268560
rect 527173 268502 528987 268504
rect 527173 268499 527239 268502
rect 528921 268499 528987 268502
rect 663750 268502 676322 268562
rect 513833 268426 513899 268429
rect 514937 268426 515003 268429
rect 513833 268424 515003 268426
rect 513833 268368 513838 268424
rect 513894 268368 514942 268424
rect 514998 268368 515003 268424
rect 513833 268366 515003 268368
rect 513833 268363 513899 268366
rect 514937 268363 515003 268366
rect 543687 268426 543753 268429
rect 549437 268426 549503 268429
rect 543687 268424 549503 268426
rect 543687 268368 543692 268424
rect 543748 268368 549442 268424
rect 549498 268368 549503 268424
rect 543687 268366 549503 268368
rect 543687 268363 543753 268366
rect 549437 268363 549503 268366
rect 523493 268290 523559 268293
rect 527541 268290 527607 268293
rect 523493 268288 527607 268290
rect 523493 268232 523498 268288
rect 523554 268232 527546 268288
rect 527602 268232 527607 268288
rect 523493 268230 527607 268232
rect 523493 268227 523559 268230
rect 527541 268227 527607 268230
rect 528553 268290 528619 268293
rect 535637 268290 535703 268293
rect 528553 268288 535703 268290
rect 528553 268232 528558 268288
rect 528614 268232 535642 268288
rect 535698 268232 535703 268288
rect 528553 268230 535703 268232
rect 528553 268227 528619 268230
rect 535637 268227 535703 268230
rect 661677 268154 661743 268157
rect 663750 268154 663810 268502
rect 676029 268290 676095 268293
rect 676029 268288 676292 268290
rect 676029 268232 676034 268288
rect 676090 268232 676292 268288
rect 676029 268230 676292 268232
rect 676029 268227 676095 268230
rect 683113 268154 683179 268157
rect 661677 268152 663810 268154
rect 661677 268096 661682 268152
rect 661738 268096 663810 268152
rect 661677 268094 663810 268096
rect 682886 268152 683179 268154
rect 682886 268096 683118 268152
rect 683174 268096 683179 268152
rect 682886 268094 683179 268096
rect 661677 268091 661743 268094
rect 539225 268018 539291 268021
rect 543825 268018 543891 268021
rect 539225 268016 543891 268018
rect 539225 267960 539230 268016
rect 539286 267960 543830 268016
rect 543886 267960 543891 268016
rect 539225 267958 543891 267960
rect 539225 267955 539291 267958
rect 543825 267955 543891 267958
rect 544009 267882 544075 267885
rect 552657 267882 552723 267885
rect 544009 267880 552723 267882
rect 544009 267824 544014 267880
rect 544070 267824 552662 267880
rect 552718 267824 552723 267880
rect 682886 267852 682946 268094
rect 683113 268091 683179 268094
rect 544009 267822 552723 267824
rect 544009 267819 544075 267822
rect 552657 267819 552723 267822
rect 518893 267610 518959 267613
rect 521653 267610 521719 267613
rect 518893 267608 521719 267610
rect 518893 267552 518898 267608
rect 518954 267552 521658 267608
rect 521714 267552 521719 267608
rect 518893 267550 521719 267552
rect 518893 267547 518959 267550
rect 521653 267547 521719 267550
rect 528553 267610 528619 267613
rect 531865 267610 531931 267613
rect 528553 267608 531931 267610
rect 528553 267552 528558 267608
rect 528614 267552 531870 267608
rect 531926 267552 531931 267608
rect 528553 267550 531931 267552
rect 528553 267547 528619 267550
rect 531865 267547 531931 267550
rect 537569 267610 537635 267613
rect 538305 267610 538371 267613
rect 537569 267608 538371 267610
rect 537569 267552 537574 267608
rect 537630 267552 538310 267608
rect 538366 267552 538371 267608
rect 537569 267550 538371 267552
rect 537569 267547 537635 267550
rect 538305 267547 538371 267550
rect 539685 267610 539751 267613
rect 539685 267608 553410 267610
rect 539685 267552 539690 267608
rect 539746 267552 553410 267608
rect 539685 267550 553410 267552
rect 539685 267547 539751 267550
rect 504909 267474 504975 267477
rect 508037 267474 508103 267477
rect 504909 267472 508103 267474
rect 504909 267416 504914 267472
rect 504970 267416 508042 267472
rect 508098 267416 508103 267472
rect 504909 267414 508103 267416
rect 504909 267411 504975 267414
rect 508037 267411 508103 267414
rect 514661 267338 514727 267341
rect 518985 267338 519051 267341
rect 514661 267336 519051 267338
rect 514661 267280 514666 267336
rect 514722 267280 518990 267336
rect 519046 267280 519051 267336
rect 514661 267278 519051 267280
rect 514661 267275 514727 267278
rect 518985 267275 519051 267278
rect 522665 267338 522731 267341
rect 528645 267338 528711 267341
rect 522665 267336 528711 267338
rect 522665 267280 522670 267336
rect 522726 267280 528650 267336
rect 528706 267280 528711 267336
rect 522665 267278 528711 267280
rect 522665 267275 522731 267278
rect 528645 267275 528711 267278
rect 538213 267338 538279 267341
rect 543825 267338 543891 267341
rect 538213 267336 543891 267338
rect 538213 267280 538218 267336
rect 538274 267280 543830 267336
rect 543886 267280 543891 267336
rect 538213 267278 543891 267280
rect 553350 267338 553410 267550
rect 580257 267338 580323 267341
rect 553350 267336 580323 267338
rect 553350 267280 580262 267336
rect 580318 267280 580323 267336
rect 553350 267278 580323 267280
rect 538213 267275 538279 267278
rect 543825 267275 543891 267278
rect 580257 267275 580323 267278
rect 672901 267338 672967 267341
rect 676262 267338 676322 267444
rect 672901 267336 676322 267338
rect 672901 267280 672906 267336
rect 672962 267280 676322 267336
rect 672901 267278 676322 267280
rect 672901 267275 672967 267278
rect 40677 267066 40743 267069
rect 62757 267066 62823 267069
rect 40677 267064 62823 267066
rect 40677 267008 40682 267064
rect 40738 267008 62762 267064
rect 62818 267008 62823 267064
rect 40677 267006 62823 267008
rect 40677 267003 40743 267006
rect 62757 267003 62823 267006
rect 509233 267066 509299 267069
rect 517513 267066 517579 267069
rect 519169 267066 519235 267069
rect 509233 267064 517579 267066
rect 509233 267008 509238 267064
rect 509294 267008 517518 267064
rect 517574 267008 517579 267064
rect 509233 267006 517579 267008
rect 509233 267003 509299 267006
rect 517513 267003 517579 267006
rect 518022 267064 519235 267066
rect 518022 267008 519174 267064
rect 519230 267008 519235 267064
rect 518022 267006 519235 267008
rect 484853 266794 484919 266797
rect 487429 266794 487495 266797
rect 484853 266792 487495 266794
rect 484853 266736 484858 266792
rect 484914 266736 487434 266792
rect 487490 266736 487495 266792
rect 484853 266734 487495 266736
rect 484853 266731 484919 266734
rect 487429 266731 487495 266734
rect 517329 266794 517395 266797
rect 518022 266794 518082 267006
rect 519169 267003 519235 267006
rect 528461 267066 528527 267069
rect 528737 267066 528803 267069
rect 528461 267064 528570 267066
rect 528461 267008 528466 267064
rect 528522 267032 528570 267064
rect 528694 267064 528803 267066
rect 528694 267032 528742 267064
rect 528522 267008 528742 267032
rect 528798 267008 528803 267064
rect 528461 267003 528803 267008
rect 536373 267066 536439 267069
rect 538857 267066 538923 267069
rect 536373 267064 538923 267066
rect 536373 267008 536378 267064
rect 536434 267008 538862 267064
rect 538918 267008 538923 267064
rect 536373 267006 538923 267008
rect 536373 267003 536439 267006
rect 538857 267003 538923 267006
rect 542169 267066 542235 267069
rect 607857 267066 607923 267069
rect 542169 267064 607923 267066
rect 542169 267008 542174 267064
rect 542230 267008 607862 267064
rect 607918 267008 607923 267064
rect 542169 267006 607923 267008
rect 542169 267003 542235 267006
rect 607857 267003 607923 267006
rect 675017 267066 675083 267069
rect 675017 267064 676292 267066
rect 675017 267008 675022 267064
rect 675078 267008 676292 267064
rect 675017 267006 676292 267008
rect 675017 267003 675083 267006
rect 528510 266972 528754 267003
rect 517329 266792 518082 266794
rect 517329 266736 517334 266792
rect 517390 266736 518082 266792
rect 517329 266734 518082 266736
rect 518709 266794 518775 266797
rect 527449 266794 527515 266797
rect 518709 266792 527515 266794
rect 518709 266736 518714 266792
rect 518770 266736 527454 266792
rect 527510 266736 527515 266792
rect 518709 266734 527515 266736
rect 517329 266731 517395 266734
rect 518709 266731 518775 266734
rect 527449 266731 527515 266734
rect 540237 266794 540303 266797
rect 540881 266794 540947 266797
rect 540237 266792 540947 266794
rect 540237 266736 540242 266792
rect 540298 266736 540886 266792
rect 540942 266736 540947 266792
rect 540237 266734 540947 266736
rect 540237 266731 540303 266734
rect 540881 266731 540947 266734
rect 528737 266658 528803 266661
rect 537385 266658 537451 266661
rect 528737 266656 537451 266658
rect 528737 266600 528742 266656
rect 528798 266600 537390 266656
rect 537446 266600 537451 266656
rect 528737 266598 537451 266600
rect 528737 266595 528803 266598
rect 537385 266595 537451 266598
rect 673085 266522 673151 266525
rect 676262 266522 676322 266628
rect 673085 266520 676322 266522
rect 673085 266464 673090 266520
rect 673146 266464 676322 266520
rect 673085 266462 676322 266464
rect 673085 266459 673151 266462
rect 673085 266114 673151 266117
rect 676262 266114 676322 266220
rect 673085 266112 676322 266114
rect 673085 266056 673090 266112
rect 673146 266056 676322 266112
rect 673085 266054 676322 266056
rect 673085 266051 673151 266054
rect 673913 265842 673979 265845
rect 673913 265840 676292 265842
rect 673913 265784 673918 265840
rect 673974 265784 676292 265840
rect 673913 265782 676292 265784
rect 673913 265779 673979 265782
rect 675385 265434 675451 265437
rect 675385 265432 676292 265434
rect 675385 265376 675390 265432
rect 675446 265376 676292 265432
rect 675385 265374 676292 265376
rect 675385 265371 675451 265374
rect 674465 265026 674531 265029
rect 674465 265024 676292 265026
rect 674465 264968 674470 265024
rect 674526 264968 676292 265024
rect 674465 264966 676292 264968
rect 674465 264963 674531 264966
rect 674833 264482 674899 264485
rect 676262 264482 676322 264588
rect 674833 264480 676322 264482
rect 674833 264424 674838 264480
rect 674894 264424 676322 264480
rect 674833 264422 676322 264424
rect 674833 264419 674899 264422
rect 676446 264077 676506 264180
rect 671981 264074 672047 264077
rect 671981 264072 676322 264074
rect 671981 264016 671986 264072
rect 672042 264016 676322 264072
rect 671981 264014 676322 264016
rect 676446 264072 676555 264077
rect 676446 264016 676494 264072
rect 676550 264016 676555 264072
rect 676446 264014 676555 264016
rect 671981 264011 672047 264014
rect 672901 263802 672967 263805
rect 674833 263802 674899 263805
rect 672901 263800 674899 263802
rect 672901 263744 672906 263800
rect 672962 263744 674838 263800
rect 674894 263744 674899 263800
rect 676262 263772 676322 264014
rect 676489 264011 676555 264014
rect 672901 263742 674899 263744
rect 672901 263739 672967 263742
rect 674833 263739 674899 263742
rect 674966 263604 674972 263668
rect 675036 263666 675042 263668
rect 676489 263666 676555 263669
rect 675036 263664 676555 263666
rect 675036 263608 676494 263664
rect 676550 263608 676555 263664
rect 675036 263606 676555 263608
rect 675036 263604 675042 263606
rect 676489 263603 676555 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 674557 263122 674623 263125
rect 675385 263122 675451 263125
rect 674557 263120 675451 263122
rect 674557 263064 674562 263120
rect 674618 263064 675390 263120
rect 675446 263064 675451 263120
rect 674557 263062 675451 263064
rect 674557 263059 674623 263062
rect 675385 263059 675451 263062
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 676070 262380 676076 262444
rect 676140 262442 676146 262444
rect 676262 262442 676322 262548
rect 676140 262382 676322 262442
rect 676140 262380 676146 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671705 262170 671771 262173
rect 671705 262168 676292 262170
rect 671705 262112 671710 262168
rect 671766 262112 676292 262168
rect 671705 262110 676292 262112
rect 671705 262107 671771 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 678470 261221 678530 261324
rect 678421 261216 678530 261221
rect 678421 261160 678426 261216
rect 678482 261160 678530 261216
rect 678421 261158 678530 261160
rect 678421 261155 678487 261158
rect 674373 260946 674439 260949
rect 674373 260944 676292 260946
rect 674373 260888 674378 260944
rect 674434 260888 676292 260944
rect 674373 260886 676292 260888
rect 674373 260883 674439 260886
rect 673361 260538 673427 260541
rect 673361 260536 676292 260538
rect 673361 260480 673366 260536
rect 673422 260480 676292 260536
rect 673361 260478 676292 260480
rect 673361 260475 673427 260478
rect 35801 259994 35867 259997
rect 50337 259994 50403 259997
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 35801 259992 50403 259994
rect 35801 259936 35806 259992
rect 35862 259936 50342 259992
rect 50398 259936 50403 259992
rect 35801 259934 50403 259936
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 35801 259931 35867 259934
rect 50337 259931 50403 259934
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 671521 259722 671587 259725
rect 671521 259720 676292 259722
rect 671521 259664 671526 259720
rect 671582 259664 676292 259720
rect 671521 259662 676292 259664
rect 671521 259659 671587 259662
rect 673637 259314 673703 259317
rect 673637 259312 676292 259314
rect 673637 259256 673642 259312
rect 673698 259256 676292 259312
rect 673637 259254 676292 259256
rect 673637 259251 673703 259254
rect 671337 258906 671403 258909
rect 671337 258904 676292 258906
rect 671337 258848 671342 258904
rect 671398 258848 676292 258904
rect 671337 258846 676292 258848
rect 671337 258843 671403 258846
rect 673913 258498 673979 258501
rect 673913 258496 676292 258498
rect 673913 258440 673918 258496
rect 673974 258440 676292 258496
rect 673913 258438 676292 258440
rect 673913 258435 673979 258438
rect 35801 258362 35867 258365
rect 35758 258360 35867 258362
rect 35758 258304 35806 258360
rect 35862 258304 35867 258360
rect 35758 258299 35867 258304
rect 35758 258060 35818 258299
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 43437 257682 43503 257685
rect 41492 257680 43503 257682
rect 41492 257624 43442 257680
rect 43498 257624 43503 257680
rect 41492 257622 43503 257624
rect 43437 257619 43503 257622
rect 670601 257682 670667 257685
rect 676262 257682 676322 258060
rect 670601 257680 676322 257682
rect 670601 257624 670606 257680
rect 670662 257652 676322 257680
rect 670662 257624 676292 257652
rect 670601 257622 676292 257624
rect 670601 257619 670667 257622
rect 672257 257274 672323 257277
rect 672257 257272 676292 257274
rect 35758 257141 35818 257244
rect 672257 257216 672262 257272
rect 672318 257216 676292 257272
rect 672257 257214 676292 257216
rect 672257 257211 672323 257214
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 42885 256866 42951 256869
rect 41492 256864 42951 256866
rect 41492 256808 42890 256864
rect 42946 256808 42951 256864
rect 41492 256806 42951 256808
rect 42885 256803 42951 256806
rect 42793 256458 42859 256461
rect 41492 256456 42859 256458
rect 41492 256400 42798 256456
rect 42854 256400 42859 256456
rect 41492 256398 42859 256400
rect 42793 256395 42859 256398
rect 43253 256050 43319 256053
rect 41492 256048 43319 256050
rect 41492 255992 43258 256048
rect 43314 255992 43319 256048
rect 41492 255990 43319 255992
rect 43253 255987 43319 255990
rect 43621 255642 43687 255645
rect 553485 255642 553551 255645
rect 41492 255640 43687 255642
rect 41492 255584 43626 255640
rect 43682 255584 43687 255640
rect 41492 255582 43687 255584
rect 552460 255640 553551 255642
rect 552460 255584 553490 255640
rect 553546 255584 553551 255640
rect 552460 255582 553551 255584
rect 43621 255579 43687 255582
rect 553485 255579 553551 255582
rect 675385 255370 675451 255373
rect 676121 255370 676187 255373
rect 675385 255368 676187 255370
rect 675385 255312 675390 255368
rect 675446 255312 676126 255368
rect 676182 255312 676187 255368
rect 675385 255310 676187 255312
rect 675385 255307 675451 255310
rect 676121 255307 676187 255310
rect 44173 255234 44239 255237
rect 41492 255232 44239 255234
rect 41492 255176 44178 255232
rect 44234 255176 44239 255232
rect 41492 255174 44239 255176
rect 44173 255171 44239 255174
rect 42977 254826 43043 254829
rect 41492 254824 43043 254826
rect 41492 254768 42982 254824
rect 43038 254768 43043 254824
rect 41492 254766 43043 254768
rect 42977 254763 43043 254766
rect 45001 254418 45067 254421
rect 41492 254416 45067 254418
rect 41492 254360 45006 254416
rect 45062 254360 45067 254416
rect 41492 254358 45067 254360
rect 45001 254355 45067 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35390 253469 35450 253572
rect 35390 253464 35499 253469
rect 554405 253466 554471 253469
rect 35390 253408 35438 253464
rect 35494 253408 35499 253464
rect 35390 253406 35499 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35433 253403 35499 253406
rect 554405 253403 554471 253406
rect 35574 253061 35634 253164
rect 35574 253056 35683 253061
rect 35574 253000 35622 253056
rect 35678 253000 35683 253056
rect 35574 252998 35683 253000
rect 35617 252995 35683 252998
rect 35758 252653 35818 252756
rect 35758 252648 35867 252653
rect 35758 252592 35806 252648
rect 35862 252592 35867 252648
rect 35758 252590 35867 252592
rect 35801 252587 35867 252590
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 44633 251970 44699 251973
rect 41492 251968 44699 251970
rect 41492 251912 44638 251968
rect 44694 251912 44699 251968
rect 41492 251910 44699 251912
rect 44633 251907 44699 251910
rect 675109 251834 675175 251837
rect 676029 251834 676095 251837
rect 675109 251832 676095 251834
rect 675109 251776 675114 251832
rect 675170 251776 676034 251832
rect 676090 251776 676095 251832
rect 675109 251774 676095 251776
rect 675109 251771 675175 251774
rect 676029 251771 676095 251774
rect 40726 251428 40786 251532
rect 40718 251364 40724 251428
rect 40788 251364 40794 251428
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 43437 251154 43503 251157
rect 41492 251152 43503 251154
rect 41492 251096 43442 251152
rect 43498 251096 43503 251152
rect 41492 251094 43503 251096
rect 43437 251091 43503 251094
rect 45553 250746 45619 250749
rect 41492 250744 45619 250746
rect 41492 250688 45558 250744
rect 45614 250688 45619 250744
rect 41492 250686 45619 250688
rect 45553 250683 45619 250686
rect 45829 250338 45895 250341
rect 41492 250336 45895 250338
rect 41492 250280 45834 250336
rect 45890 250280 45895 250336
rect 41492 250278 45895 250280
rect 45829 250275 45895 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 674925 249930 674991 249933
rect 676070 249930 676076 249932
rect 674925 249928 676076 249930
rect 40542 249796 40602 249900
rect 674925 249872 674930 249928
rect 674986 249872 676076 249928
rect 674925 249870 676076 249872
rect 674925 249867 674991 249870
rect 676070 249868 676076 249870
rect 676140 249868 676146 249932
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675385 249658 675451 249661
rect 674852 249656 675451 249658
rect 674852 249600 675390 249656
rect 675446 249600 675451 249656
rect 674852 249598 675451 249600
rect 674852 249596 674858 249598
rect 675385 249595 675451 249598
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 43713 249114 43779 249117
rect 553853 249114 553919 249117
rect 41492 249112 43779 249114
rect 41492 249056 43718 249112
rect 43774 249056 43779 249112
rect 41492 249054 43779 249056
rect 552460 249112 553919 249114
rect 552460 249056 553858 249112
rect 553914 249056 553919 249112
rect 552460 249054 553919 249056
rect 43713 249051 43779 249054
rect 553853 249051 553919 249054
rect 44541 248706 44607 248709
rect 41492 248704 44607 248706
rect 41492 248648 44546 248704
rect 44602 248648 44607 248704
rect 41492 248646 44607 248648
rect 44541 248643 44607 248646
rect 44357 248298 44423 248301
rect 41492 248296 44423 248298
rect 41492 248240 44362 248296
rect 44418 248240 44423 248296
rect 41492 248238 44423 248240
rect 44357 248235 44423 248238
rect 41462 247754 41522 247860
rect 50521 247754 50587 247757
rect 41462 247752 50587 247754
rect 41462 247696 50526 247752
rect 50582 247696 50587 247752
rect 41462 247694 50587 247696
rect 50521 247691 50587 247694
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46933 247074 46999 247077
rect 41492 247072 46999 247074
rect 41492 247016 46938 247072
rect 46994 247016 46999 247072
rect 41492 247014 46999 247016
rect 46933 247011 46999 247014
rect 554405 246938 554471 246941
rect 552460 246936 554471 246938
rect 552460 246880 554410 246936
rect 554466 246880 554471 246936
rect 552460 246878 554471 246880
rect 554405 246875 554471 246878
rect 674281 246938 674347 246941
rect 675109 246938 675175 246941
rect 674281 246936 675175 246938
rect 674281 246880 674286 246936
rect 674342 246880 675114 246936
rect 675170 246880 675175 246936
rect 674281 246878 675175 246880
rect 674281 246875 674347 246878
rect 675109 246875 675175 246878
rect 41462 246530 41522 246636
rect 50337 246530 50403 246533
rect 41462 246528 50403 246530
rect 41462 246472 50342 246528
rect 50398 246472 50403 246528
rect 41462 246470 50403 246472
rect 50337 246467 50403 246470
rect 671521 245850 671587 245853
rect 675293 245850 675359 245853
rect 671521 245848 675359 245850
rect 671521 245792 671526 245848
rect 671582 245792 675298 245848
rect 675354 245792 675359 245848
rect 671521 245790 675359 245792
rect 671521 245787 671587 245790
rect 675293 245787 675359 245790
rect 671705 245578 671771 245581
rect 674782 245578 674788 245580
rect 671705 245576 674788 245578
rect 671705 245520 671710 245576
rect 671766 245520 674788 245576
rect 671705 245518 674788 245520
rect 671705 245515 671771 245518
rect 674782 245516 674788 245518
rect 674852 245516 674858 245580
rect 675886 245516 675892 245580
rect 675956 245578 675962 245580
rect 676806 245578 676812 245580
rect 675956 245518 676812 245578
rect 675956 245516 675962 245518
rect 676806 245516 676812 245518
rect 676876 245516 676882 245580
rect 673361 245306 673427 245309
rect 675334 245306 675340 245308
rect 673361 245304 675340 245306
rect 673361 245248 673366 245304
rect 673422 245248 675340 245304
rect 673361 245246 675340 245248
rect 673361 245243 673427 245246
rect 675334 245244 675340 245246
rect 675404 245244 675410 245308
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 40677 242858 40743 242861
rect 43253 242858 43319 242861
rect 40677 242856 43319 242858
rect 40677 242800 40682 242856
rect 40738 242800 43258 242856
rect 43314 242800 43319 242856
rect 40677 242798 43319 242800
rect 40677 242795 40743 242798
rect 43253 242795 43319 242798
rect 673637 242858 673703 242861
rect 675293 242858 675359 242861
rect 673637 242856 675359 242858
rect 673637 242800 673642 242856
rect 673698 242800 675298 242856
rect 675354 242800 675359 242856
rect 673637 242798 675359 242800
rect 673637 242795 673703 242798
rect 675293 242795 675359 242798
rect 553945 242586 554011 242589
rect 552460 242584 554011 242586
rect 552460 242528 553950 242584
rect 554006 242528 554011 242584
rect 552460 242526 554011 242528
rect 553945 242523 554011 242526
rect 675661 242314 675727 242317
rect 675886 242314 675892 242316
rect 675661 242312 675892 242314
rect 675661 242256 675666 242312
rect 675722 242256 675892 242312
rect 675661 242254 675892 242256
rect 675661 242251 675727 242254
rect 675886 242252 675892 242254
rect 675956 242252 675962 242316
rect 671337 241498 671403 241501
rect 675109 241498 675175 241501
rect 671337 241496 675175 241498
rect 671337 241440 671342 241496
rect 671398 241440 675114 241496
rect 675170 241440 675175 241496
rect 671337 241438 675175 241440
rect 671337 241435 671403 241438
rect 675109 241435 675175 241438
rect 553853 240410 553919 240413
rect 552460 240408 553919 240410
rect 552460 240352 553858 240408
rect 553914 240352 553919 240408
rect 552460 240350 553919 240352
rect 553853 240347 553919 240350
rect 675385 240276 675451 240277
rect 675334 240274 675340 240276
rect 675294 240214 675340 240274
rect 675404 240272 675451 240276
rect 675446 240216 675451 240272
rect 675334 240212 675340 240214
rect 675404 240212 675451 240216
rect 675385 240211 675451 240212
rect 40718 240076 40724 240140
rect 40788 240138 40794 240140
rect 41781 240138 41847 240141
rect 40788 240136 41847 240138
rect 40788 240080 41786 240136
rect 41842 240080 41847 240136
rect 40788 240078 41847 240080
rect 40788 240076 40794 240078
rect 41781 240075 41847 240078
rect 673085 240002 673151 240005
rect 673310 240002 673316 240004
rect 673085 240000 673316 240002
rect 673085 239944 673090 240000
rect 673146 239944 673316 240000
rect 673085 239942 673316 239944
rect 673085 239939 673151 239942
rect 673310 239940 673316 239942
rect 673380 239940 673386 240004
rect 42149 238506 42215 238509
rect 46933 238506 46999 238509
rect 42149 238504 46999 238506
rect 42149 238448 42154 238504
rect 42210 238448 46938 238504
rect 46994 238448 46999 238504
rect 42149 238446 46999 238448
rect 42149 238443 42215 238446
rect 46933 238443 46999 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 671889 238234 671955 238237
rect 675109 238234 675175 238237
rect 671889 238232 675175 238234
rect 671889 238176 671894 238232
rect 671950 238176 675114 238232
rect 675170 238176 675175 238232
rect 671889 238174 675175 238176
rect 671889 238171 671955 238174
rect 675109 238171 675175 238174
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42609 237418 42675 237421
rect 42076 237416 42675 237418
rect 42076 237360 42614 237416
rect 42670 237360 42675 237416
rect 42076 237358 42675 237360
rect 42076 237356 42082 237358
rect 42609 237355 42675 237358
rect 674782 237220 674788 237284
rect 674852 237282 674858 237284
rect 675109 237282 675175 237285
rect 674852 237280 675175 237282
rect 674852 237224 675114 237280
rect 675170 237224 675175 237280
rect 674852 237222 675175 237224
rect 674852 237220 674858 237222
rect 675109 237219 675175 237222
rect 673297 237146 673363 237149
rect 674046 237146 674052 237148
rect 673297 237144 674052 237146
rect 673297 237088 673302 237144
rect 673358 237088 674052 237144
rect 673297 237086 674052 237088
rect 673297 237083 673363 237086
rect 674046 237084 674052 237086
rect 674116 237084 674122 237148
rect 673521 236738 673587 236741
rect 669270 236736 673587 236738
rect 669270 236680 673526 236736
rect 673582 236680 673587 236736
rect 669270 236678 673587 236680
rect 666185 236194 666251 236197
rect 669270 236194 669330 236678
rect 673521 236675 673587 236678
rect 666185 236192 669330 236194
rect 666185 236136 666190 236192
rect 666246 236136 669330 236192
rect 666185 236134 669330 236136
rect 666185 236131 666251 236134
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 40534 235860 40540 235924
rect 40604 235922 40610 235924
rect 41781 235922 41847 235925
rect 40604 235920 41847 235922
rect 40604 235864 41786 235920
rect 41842 235864 41847 235920
rect 40604 235862 41847 235864
rect 40604 235860 40610 235862
rect 41781 235859 41847 235862
rect 42241 235922 42307 235925
rect 44357 235922 44423 235925
rect 42241 235920 44423 235922
rect 42241 235864 42246 235920
rect 42302 235864 44362 235920
rect 44418 235864 44423 235920
rect 42241 235862 44423 235864
rect 42241 235859 42307 235862
rect 44357 235859 44423 235862
rect 670601 235922 670667 235925
rect 674925 235922 674991 235925
rect 670601 235920 674991 235922
rect 670601 235864 670606 235920
rect 670662 235864 674930 235920
rect 674986 235864 674991 235920
rect 670601 235862 674991 235864
rect 670601 235859 670667 235862
rect 674925 235859 674991 235862
rect 673310 235180 673316 235244
rect 673380 235242 673386 235244
rect 676029 235242 676095 235245
rect 673380 235240 676095 235242
rect 673380 235184 676034 235240
rect 676090 235184 676095 235240
rect 673380 235182 676095 235184
rect 673380 235180 673386 235182
rect 676029 235179 676095 235182
rect 674465 234834 674531 234837
rect 675845 234834 675911 234837
rect 674465 234832 675911 234834
rect 674465 234776 674470 234832
rect 674526 234776 675850 234832
rect 675906 234776 675911 234832
rect 674465 234774 675911 234776
rect 674465 234771 674531 234774
rect 675845 234771 675911 234774
rect 42241 234562 42307 234565
rect 46013 234562 46079 234565
rect 42241 234560 46079 234562
rect 42241 234504 42246 234560
rect 42302 234504 46018 234560
rect 46074 234504 46079 234560
rect 42241 234502 46079 234504
rect 42241 234499 42307 234502
rect 46013 234499 46079 234502
rect 42241 234154 42307 234157
rect 44449 234154 44515 234157
rect 42241 234152 44515 234154
rect 42241 234096 42246 234152
rect 42302 234096 44454 234152
rect 44510 234096 44515 234152
rect 42241 234094 44515 234096
rect 42241 234091 42307 234094
rect 44449 234091 44515 234094
rect 663241 234154 663307 234157
rect 683205 234154 683271 234157
rect 663241 234152 683271 234154
rect 663241 234096 663246 234152
rect 663302 234096 683210 234152
rect 683266 234096 683271 234152
rect 663241 234094 683271 234096
rect 663241 234091 663307 234094
rect 683205 234091 683271 234094
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683665 233882 683731 233885
rect 658917 233880 683731 233882
rect 658917 233824 658922 233880
rect 658978 233824 683670 233880
rect 683726 233824 683731 233880
rect 658917 233822 683731 233824
rect 658917 233819 658983 233822
rect 683665 233819 683731 233822
rect 673269 233610 673335 233613
rect 675845 233610 675911 233613
rect 673269 233608 675911 233610
rect 673269 233552 673274 233608
rect 673330 233552 675850 233608
rect 675906 233552 675911 233608
rect 673269 233550 675911 233552
rect 673269 233547 673335 233550
rect 675845 233547 675911 233550
rect 42149 233338 42215 233341
rect 44633 233338 44699 233341
rect 42149 233336 44699 233338
rect 42149 233280 42154 233336
rect 42210 233280 44638 233336
rect 44694 233280 44699 233336
rect 42149 233278 44699 233280
rect 42149 233275 42215 233278
rect 44633 233275 44699 233278
rect 671286 233140 671292 233204
rect 671356 233202 671362 233204
rect 672257 233202 672323 233205
rect 671356 233200 672323 233202
rect 671356 233144 672262 233200
rect 672318 233144 672323 233200
rect 671356 233142 672323 233144
rect 671356 233140 671362 233142
rect 672257 233139 672323 233142
rect 670509 232658 670575 232661
rect 673729 232658 673795 232661
rect 670509 232656 673795 232658
rect 670509 232600 670514 232656
rect 670570 232600 673734 232656
rect 673790 232600 673795 232656
rect 670509 232598 673795 232600
rect 670509 232595 670575 232598
rect 673729 232595 673795 232598
rect 670325 232114 670391 232117
rect 673637 232114 673703 232117
rect 670325 232112 673703 232114
rect 670325 232056 670330 232112
rect 670386 232056 673642 232112
rect 673698 232056 673703 232112
rect 670325 232054 673703 232056
rect 670325 232051 670391 232054
rect 673637 232051 673703 232054
rect 675173 231842 675239 231845
rect 663750 231840 675239 231842
rect 663750 231784 675178 231840
rect 675234 231784 675239 231840
rect 663750 231782 675239 231784
rect 42241 231706 42307 231709
rect 43713 231706 43779 231709
rect 42241 231704 43779 231706
rect 42241 231648 42246 231704
rect 42302 231648 43718 231704
rect 43774 231648 43779 231704
rect 42241 231646 43779 231648
rect 42241 231643 42307 231646
rect 43713 231643 43779 231646
rect 663057 231706 663123 231709
rect 663750 231706 663810 231782
rect 675173 231779 675239 231782
rect 663057 231704 663810 231706
rect 663057 231648 663062 231704
rect 663118 231648 663810 231704
rect 663057 231646 663810 231648
rect 663057 231643 663123 231646
rect 669405 231570 669471 231573
rect 675063 231570 675129 231573
rect 669405 231568 675129 231570
rect 669405 231512 669410 231568
rect 669466 231512 675068 231568
rect 675124 231512 675129 231568
rect 669405 231510 675129 231512
rect 669405 231507 669471 231510
rect 675063 231507 675129 231510
rect 640241 231434 640307 231437
rect 669262 231434 669268 231436
rect 640241 231432 669268 231434
rect 640241 231376 640246 231432
rect 640302 231376 669268 231432
rect 640241 231374 669268 231376
rect 640241 231371 640307 231374
rect 669262 231372 669268 231374
rect 669332 231372 669338 231436
rect 665265 231162 665331 231165
rect 674725 231162 674791 231165
rect 665265 231160 674791 231162
rect 665265 231104 665270 231160
rect 665326 231104 674730 231160
rect 674786 231104 674791 231160
rect 665265 231102 674791 231104
rect 665265 231099 665331 231102
rect 674725 231099 674791 231102
rect 663241 230890 663307 230893
rect 674833 230890 674899 230893
rect 663241 230888 674899 230890
rect 663241 230832 663246 230888
rect 663302 230832 674838 230888
rect 674894 230832 674899 230888
rect 663241 230830 674899 230832
rect 663241 230827 663307 230830
rect 674833 230827 674899 230830
rect 664437 230618 664503 230621
rect 668209 230618 668275 230621
rect 664437 230616 668275 230618
rect 664437 230560 664442 230616
rect 664498 230560 668214 230616
rect 668270 230560 668275 230616
rect 664437 230558 668275 230560
rect 664437 230555 664503 230558
rect 668209 230555 668275 230558
rect 674511 230618 674577 230621
rect 676857 230618 676923 230621
rect 674511 230616 676923 230618
rect 674511 230560 674516 230616
rect 674572 230560 676862 230616
rect 676918 230560 676923 230616
rect 674511 230558 676923 230560
rect 674511 230555 674577 230558
rect 676857 230555 676923 230558
rect 668577 230482 668643 230485
rect 674389 230482 674455 230485
rect 668577 230480 674455 230482
rect 668577 230424 668582 230480
rect 668638 230424 674394 230480
rect 674450 230424 674455 230480
rect 668577 230422 674455 230424
rect 668577 230419 668643 230422
rect 674389 230419 674455 230422
rect 42149 230210 42215 230213
rect 45829 230210 45895 230213
rect 42149 230208 45895 230210
rect 42149 230152 42154 230208
rect 42210 230152 45834 230208
rect 45890 230152 45895 230208
rect 42149 230150 45895 230152
rect 42149 230147 42215 230150
rect 45829 230147 45895 230150
rect 639597 230210 639663 230213
rect 673453 230210 673519 230213
rect 639597 230208 673519 230210
rect 639597 230152 639602 230208
rect 639658 230152 673458 230208
rect 673514 230152 673519 230208
rect 639597 230150 673519 230152
rect 639597 230147 639663 230150
rect 673453 230147 673519 230150
rect 673729 230210 673795 230213
rect 676581 230210 676647 230213
rect 673729 230208 676647 230210
rect 673729 230152 673734 230208
rect 673790 230152 676586 230208
rect 676642 230152 676647 230208
rect 673729 230150 676647 230152
rect 673729 230147 673795 230150
rect 676581 230147 676647 230150
rect 42241 229938 42307 229941
rect 45553 229938 45619 229941
rect 42241 229936 45619 229938
rect 42241 229880 42246 229936
rect 42302 229880 45558 229936
rect 45614 229880 45619 229936
rect 42241 229878 45619 229880
rect 42241 229875 42307 229878
rect 45553 229875 45619 229878
rect 151353 229938 151419 229941
rect 152365 229938 152431 229941
rect 151353 229936 152431 229938
rect 151353 229880 151358 229936
rect 151414 229880 152370 229936
rect 152426 229880 152431 229936
rect 151353 229878 152431 229880
rect 151353 229875 151419 229878
rect 152365 229875 152431 229878
rect 674557 229938 674623 229941
rect 675109 229938 675175 229941
rect 674557 229936 675175 229938
rect 674557 229880 674562 229936
rect 674618 229880 675114 229936
rect 675170 229880 675175 229936
rect 674557 229878 675175 229880
rect 674557 229875 674623 229878
rect 675109 229875 675175 229878
rect 103605 229802 103671 229805
rect 145649 229802 145715 229805
rect 103605 229800 145715 229802
rect 103605 229744 103610 229800
rect 103666 229744 145654 229800
rect 145710 229744 145715 229800
rect 103605 229742 145715 229744
rect 103605 229739 103671 229742
rect 145649 229739 145715 229742
rect 637481 229802 637547 229805
rect 673729 229802 673795 229805
rect 637481 229800 673795 229802
rect 637481 229744 637486 229800
rect 637542 229744 673734 229800
rect 673790 229744 673795 229800
rect 637481 229742 673795 229744
rect 637481 229739 637547 229742
rect 673729 229739 673795 229742
rect 660941 229530 661007 229533
rect 673269 229530 673335 229533
rect 660941 229528 673335 229530
rect 660941 229472 660946 229528
rect 661002 229472 673274 229528
rect 673330 229472 673335 229528
rect 660941 229470 673335 229472
rect 660941 229467 661007 229470
rect 673269 229467 673335 229470
rect 146293 229258 146359 229261
rect 147949 229258 148015 229261
rect 146293 229256 148015 229258
rect 146293 229200 146298 229256
rect 146354 229200 147954 229256
rect 148010 229200 148015 229256
rect 146293 229198 148015 229200
rect 146293 229195 146359 229198
rect 147949 229195 148015 229198
rect 661677 229258 661743 229261
rect 668577 229258 668643 229261
rect 661677 229256 668643 229258
rect 661677 229200 661682 229256
rect 661738 229200 668582 229256
rect 668638 229200 668643 229256
rect 661677 229198 668643 229200
rect 661677 229195 661743 229198
rect 668577 229195 668643 229198
rect 673381 229258 673447 229261
rect 675109 229258 675175 229261
rect 673381 229256 675175 229258
rect 673381 229200 673386 229256
rect 673442 229200 675114 229256
rect 675170 229200 675175 229256
rect 673381 229198 675175 229200
rect 673381 229195 673447 229198
rect 675109 229195 675175 229198
rect 190545 229122 190611 229125
rect 192293 229122 192359 229125
rect 190545 229120 192359 229122
rect 190545 229064 190550 229120
rect 190606 229064 192298 229120
rect 192354 229064 192359 229120
rect 190545 229062 192359 229064
rect 190545 229059 190611 229062
rect 192293 229059 192359 229062
rect 157977 228986 158043 228989
rect 163865 228986 163931 228989
rect 157977 228984 163931 228986
rect 157977 228928 157982 228984
rect 158038 228928 163870 228984
rect 163926 228928 163931 228984
rect 157977 228926 163931 228928
rect 157977 228923 158043 228926
rect 163865 228923 163931 228926
rect 171133 228986 171199 228989
rect 172237 228986 172303 228989
rect 171133 228984 172303 228986
rect 171133 228928 171138 228984
rect 171194 228928 172242 228984
rect 172298 228928 172303 228984
rect 171133 228926 172303 228928
rect 171133 228923 171199 228926
rect 172237 228923 172303 228926
rect 172421 228986 172487 228989
rect 174077 228986 174143 228989
rect 172421 228984 174143 228986
rect 172421 228928 172426 228984
rect 172482 228928 174082 228984
rect 174138 228928 174143 228984
rect 172421 228926 174143 228928
rect 172421 228923 172487 228926
rect 174077 228923 174143 228926
rect 180609 228986 180675 228989
rect 181897 228986 181963 228989
rect 180609 228984 181963 228986
rect 180609 228928 180614 228984
rect 180670 228928 181902 228984
rect 181958 228928 181963 228984
rect 180609 228926 181963 228928
rect 180609 228923 180675 228926
rect 181897 228923 181963 228926
rect 672901 228986 672967 228989
rect 673310 228986 673316 228988
rect 672901 228984 673316 228986
rect 672901 228928 672906 228984
rect 672962 228928 673316 228984
rect 672901 228926 673316 228928
rect 672901 228923 672967 228926
rect 673310 228924 673316 228926
rect 673380 228924 673386 228988
rect 673545 228986 673611 228989
rect 673545 228984 675034 228986
rect 673545 228928 673550 228984
rect 673606 228928 675034 228984
rect 673545 228926 675034 228928
rect 673545 228923 673611 228926
rect 174261 228850 174327 228853
rect 175641 228850 175707 228853
rect 174261 228848 175707 228850
rect 174261 228792 174266 228848
rect 174322 228792 175646 228848
rect 175702 228792 175707 228848
rect 174261 228790 175707 228792
rect 174261 228787 174327 228790
rect 175641 228787 175707 228790
rect 669446 228788 669452 228852
rect 669516 228850 669522 228852
rect 672257 228850 672323 228853
rect 669516 228848 672323 228850
rect 669516 228792 672262 228848
rect 672318 228792 672323 228848
rect 669516 228790 672323 228792
rect 669516 228788 669522 228790
rect 672257 228787 672323 228790
rect 157425 228578 157491 228581
rect 158805 228578 158871 228581
rect 672901 228580 672967 228581
rect 672901 228578 672948 228580
rect 157425 228576 158871 228578
rect 157425 228520 157430 228576
rect 157486 228520 158810 228576
rect 158866 228520 158871 228576
rect 157425 228518 158871 228520
rect 672856 228576 672948 228578
rect 672856 228520 672906 228576
rect 672856 228518 672948 228520
rect 157425 228515 157491 228518
rect 158805 228515 158871 228518
rect 672901 228516 672948 228518
rect 673012 228516 673018 228580
rect 673381 228578 673447 228581
rect 674782 228578 674788 228580
rect 673381 228576 674788 228578
rect 673381 228520 673386 228576
rect 673442 228520 674788 228576
rect 673381 228518 674788 228520
rect 672901 228515 672967 228516
rect 673381 228515 673447 228518
rect 674782 228516 674788 228518
rect 674852 228516 674858 228580
rect 674974 228578 675034 228926
rect 677041 228578 677107 228581
rect 674974 228576 677107 228578
rect 674974 228520 677046 228576
rect 677102 228520 677107 228576
rect 674974 228518 677107 228520
rect 677041 228515 677107 228518
rect 166625 228442 166691 228445
rect 171593 228442 171659 228445
rect 166625 228440 171659 228442
rect 166625 228384 166630 228440
rect 166686 228384 171598 228440
rect 171654 228384 171659 228440
rect 166625 228382 171659 228384
rect 166625 228379 166691 228382
rect 171593 228379 171659 228382
rect 79961 228306 80027 228309
rect 160461 228306 160527 228309
rect 79961 228304 160527 228306
rect 79961 228248 79966 228304
rect 80022 228248 160466 228304
rect 160522 228248 160527 228304
rect 79961 228246 160527 228248
rect 79961 228243 80027 228246
rect 160461 228243 160527 228246
rect 134609 228034 134675 228037
rect 141141 228034 141207 228037
rect 134609 228032 141207 228034
rect 134609 227976 134614 228032
rect 134670 227976 141146 228032
rect 141202 227976 141207 228032
rect 134609 227974 141207 227976
rect 134609 227971 134675 227974
rect 141141 227971 141207 227974
rect 145925 228034 145991 228037
rect 150341 228034 150407 228037
rect 145925 228032 150407 228034
rect 145925 227976 145930 228032
rect 145986 227976 150346 228032
rect 150402 227976 150407 228032
rect 145925 227974 150407 227976
rect 145925 227971 145991 227974
rect 150341 227971 150407 227974
rect 155861 228034 155927 228037
rect 157793 228034 157859 228037
rect 155861 228032 157859 228034
rect 155861 227976 155866 228032
rect 155922 227976 157798 228032
rect 157854 227976 157859 228032
rect 155861 227974 157859 227976
rect 155861 227971 155927 227974
rect 157793 227971 157859 227974
rect 159633 227490 159699 227493
rect 166441 227490 166507 227493
rect 159633 227488 166507 227490
rect 159633 227432 159638 227488
rect 159694 227432 166446 227488
rect 166502 227432 166507 227488
rect 159633 227430 166507 227432
rect 159633 227427 159699 227430
rect 166441 227427 166507 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 151813 227354 151879 227357
rect 154665 227354 154731 227357
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 151813 227352 154731 227354
rect 151813 227296 151818 227352
rect 151874 227296 154670 227352
rect 154726 227296 154731 227352
rect 151813 227294 154731 227296
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 151813 227291 151879 227294
rect 154665 227291 154731 227294
rect 142153 227218 142219 227221
rect 143073 227218 143139 227221
rect 142153 227216 143139 227218
rect 142153 227160 142158 227216
rect 142214 227160 143078 227216
rect 143134 227160 143139 227216
rect 142153 227158 143139 227160
rect 142153 227155 142219 227158
rect 143073 227155 143139 227158
rect 670509 227218 670575 227221
rect 671102 227218 671108 227220
rect 670509 227216 671108 227218
rect 670509 227160 670514 227216
rect 670570 227160 671108 227216
rect 670509 227158 671108 227160
rect 670509 227155 670575 227158
rect 671102 227156 671108 227158
rect 671172 227156 671178 227220
rect 671889 227082 671955 227085
rect 674925 227082 674991 227085
rect 671889 227080 674991 227082
rect 671889 227024 671894 227080
rect 671950 227024 674930 227080
rect 674986 227024 674991 227080
rect 671889 227022 674991 227024
rect 671889 227019 671955 227022
rect 674925 227019 674991 227022
rect 73061 226946 73127 226949
rect 155309 226946 155375 226949
rect 73061 226944 155375 226946
rect 73061 226888 73066 226944
rect 73122 226888 155314 226944
rect 155370 226888 155375 226944
rect 73061 226886 155375 226888
rect 73061 226883 73127 226886
rect 155309 226883 155375 226886
rect 670509 226810 670575 226813
rect 671654 226810 671660 226812
rect 670509 226808 671660 226810
rect 670509 226752 670514 226808
rect 670570 226752 671660 226808
rect 670509 226750 671660 226752
rect 670509 226747 670575 226750
rect 671654 226748 671660 226750
rect 671724 226748 671730 226812
rect 672257 226810 672323 226813
rect 673126 226810 673132 226812
rect 672257 226808 673132 226810
rect 672257 226752 672262 226808
rect 672318 226752 673132 226808
rect 672257 226750 673132 226752
rect 672257 226747 672323 226750
rect 673126 226748 673132 226750
rect 673196 226748 673202 226812
rect 42149 226674 42215 226677
rect 43437 226674 43503 226677
rect 42149 226672 43503 226674
rect 42149 226616 42154 226672
rect 42210 226616 43442 226672
rect 43498 226616 43503 226672
rect 42149 226614 43503 226616
rect 42149 226611 42215 226614
rect 43437 226611 43503 226614
rect 150341 226674 150407 226677
rect 152273 226674 152339 226677
rect 671889 226676 671955 226677
rect 671838 226674 671844 226676
rect 150341 226672 152339 226674
rect 150341 226616 150346 226672
rect 150402 226616 152278 226672
rect 152334 226616 152339 226672
rect 150341 226614 152339 226616
rect 671798 226614 671844 226674
rect 671908 226672 671955 226676
rect 671950 226616 671955 226672
rect 150341 226611 150407 226614
rect 152273 226611 152339 226614
rect 671838 226612 671844 226614
rect 671908 226612 671955 226616
rect 671889 226611 671955 226612
rect 139301 226538 139367 226541
rect 142245 226538 142311 226541
rect 672027 226540 672093 226541
rect 139301 226536 142311 226538
rect 139301 226480 139306 226536
rect 139362 226480 142250 226536
rect 142306 226480 142311 226536
rect 139301 226478 142311 226480
rect 139301 226475 139367 226478
rect 142245 226475 142311 226478
rect 672022 226476 672028 226540
rect 672092 226538 672098 226540
rect 673177 226538 673243 226541
rect 675150 226538 675156 226540
rect 672092 226478 672184 226538
rect 673177 226536 675156 226538
rect 673177 226480 673182 226536
rect 673238 226480 675156 226536
rect 673177 226478 675156 226480
rect 672092 226476 672098 226478
rect 672027 226475 672093 226476
rect 673177 226475 673243 226478
rect 675150 226476 675156 226478
rect 675220 226476 675226 226540
rect 652753 226402 652819 226405
rect 671889 226402 671955 226405
rect 652753 226400 671955 226402
rect 652753 226344 652758 226400
rect 652814 226344 671894 226400
rect 671950 226344 671955 226400
rect 652753 226342 671955 226344
rect 652753 226339 652819 226342
rect 671889 226339 671955 226342
rect 673678 226204 673684 226268
rect 673748 226266 673754 226268
rect 674097 226266 674163 226269
rect 673748 226264 674163 226266
rect 673748 226208 674102 226264
rect 674158 226208 674163 226264
rect 673748 226206 674163 226208
rect 673748 226204 673754 226206
rect 674097 226203 674163 226206
rect 152917 226130 152983 226133
rect 157609 226130 157675 226133
rect 152917 226128 157675 226130
rect 152917 226072 152922 226128
rect 152978 226072 157614 226128
rect 157670 226072 157675 226128
rect 152917 226070 157675 226072
rect 152917 226067 152983 226070
rect 157609 226067 157675 226070
rect 176653 226130 176719 226133
rect 180793 226130 180859 226133
rect 176653 226128 180859 226130
rect 176653 226072 176658 226128
rect 176714 226072 180798 226128
rect 180854 226072 180859 226128
rect 176653 226070 180859 226072
rect 176653 226067 176719 226070
rect 180793 226067 180859 226070
rect 181069 226130 181135 226133
rect 186129 226130 186195 226133
rect 181069 226128 186195 226130
rect 181069 226072 181074 226128
rect 181130 226072 186134 226128
rect 186190 226072 186195 226128
rect 181069 226070 186195 226072
rect 181069 226067 181135 226070
rect 186129 226067 186195 226070
rect 670509 226130 670575 226133
rect 670509 226128 672090 226130
rect 670509 226072 670514 226128
rect 670570 226072 672090 226128
rect 670509 226070 672090 226072
rect 670509 226067 670575 226070
rect 170857 225994 170923 225997
rect 171225 225994 171291 225997
rect 170857 225992 171291 225994
rect 170857 225936 170862 225992
rect 170918 225936 171230 225992
rect 171286 225936 171291 225992
rect 170857 225934 171291 225936
rect 170857 225931 170923 225934
rect 171225 225931 171291 225934
rect 186405 225994 186471 225997
rect 188061 225994 188127 225997
rect 186405 225992 188127 225994
rect 186405 225936 186410 225992
rect 186466 225936 188066 225992
rect 188122 225936 188127 225992
rect 186405 225934 188127 225936
rect 672030 225994 672090 226070
rect 674097 225994 674163 225997
rect 672030 225992 674163 225994
rect 672030 225936 674102 225992
rect 674158 225936 674163 225992
rect 672030 225934 674163 225936
rect 186405 225931 186471 225934
rect 188061 225931 188127 225934
rect 674097 225931 674163 225934
rect 166809 225858 166875 225861
rect 169845 225858 169911 225861
rect 671337 225858 671403 225861
rect 166809 225856 169911 225858
rect 166809 225800 166814 225856
rect 166870 225800 169850 225856
rect 169906 225800 169911 225856
rect 166809 225798 169911 225800
rect 166809 225795 166875 225798
rect 169845 225795 169911 225798
rect 663750 225856 671403 225858
rect 663750 225800 671342 225856
rect 671398 225800 671403 225856
rect 663750 225798 671403 225800
rect 42425 225722 42491 225725
rect 43253 225722 43319 225725
rect 42425 225720 43319 225722
rect 42425 225664 42430 225720
rect 42486 225664 43258 225720
rect 43314 225664 43319 225720
rect 42425 225662 43319 225664
rect 42425 225659 42491 225662
rect 43253 225659 43319 225662
rect 171041 225722 171107 225725
rect 176929 225722 176995 225725
rect 171041 225720 176995 225722
rect 171041 225664 171046 225720
rect 171102 225664 176934 225720
rect 176990 225664 176995 225720
rect 171041 225662 176995 225664
rect 171041 225659 171107 225662
rect 176929 225659 176995 225662
rect 184841 225722 184907 225725
rect 186405 225722 186471 225725
rect 184841 225720 186471 225722
rect 184841 225664 184846 225720
rect 184902 225664 186410 225720
rect 186466 225664 186471 225720
rect 184841 225662 186471 225664
rect 184841 225659 184907 225662
rect 186405 225659 186471 225662
rect 142981 225586 143047 225589
rect 147397 225586 147463 225589
rect 142981 225584 147463 225586
rect 142981 225528 142986 225584
rect 143042 225528 147402 225584
rect 147458 225528 147463 225584
rect 142981 225526 147463 225528
rect 142981 225523 143047 225526
rect 147397 225523 147463 225526
rect 161565 225586 161631 225589
rect 166717 225586 166783 225589
rect 161565 225584 166783 225586
rect 161565 225528 161570 225584
rect 161626 225528 166722 225584
rect 166778 225528 166783 225584
rect 161565 225526 166783 225528
rect 161565 225523 161631 225526
rect 166717 225523 166783 225526
rect 650637 225586 650703 225589
rect 663750 225586 663810 225798
rect 671337 225795 671403 225798
rect 671813 225722 671879 225725
rect 672165 225722 672231 225725
rect 671813 225720 672231 225722
rect 671813 225664 671818 225720
rect 671874 225664 672170 225720
rect 672226 225664 672231 225720
rect 671813 225662 672231 225664
rect 671813 225659 671879 225662
rect 672165 225659 672231 225662
rect 672855 225722 672921 225725
rect 675661 225722 675727 225725
rect 672855 225720 675727 225722
rect 672855 225664 672860 225720
rect 672916 225664 675666 225720
rect 675722 225664 675727 225720
rect 672855 225662 675727 225664
rect 672855 225659 672921 225662
rect 675661 225659 675727 225662
rect 650637 225584 663810 225586
rect 650637 225528 650642 225584
rect 650698 225528 663810 225584
rect 650637 225526 663810 225528
rect 650637 225523 650703 225526
rect 186129 225450 186195 225453
rect 187049 225450 187115 225453
rect 186129 225448 187115 225450
rect 186129 225392 186134 225448
rect 186190 225392 187054 225448
rect 187110 225392 187115 225448
rect 186129 225390 187115 225392
rect 186129 225387 186195 225390
rect 187049 225387 187115 225390
rect 190545 225450 190611 225453
rect 194869 225450 194935 225453
rect 190545 225448 194935 225450
rect 190545 225392 190550 225448
rect 190606 225392 194874 225448
rect 194930 225392 194935 225448
rect 190545 225390 194935 225392
rect 190545 225387 190611 225390
rect 194869 225387 194935 225390
rect 671337 225450 671403 225453
rect 673637 225450 673703 225453
rect 671337 225448 673703 225450
rect 671337 225392 671342 225448
rect 671398 225392 673642 225448
rect 673698 225392 673703 225448
rect 671337 225390 673703 225392
rect 671337 225387 671403 225390
rect 673637 225387 673703 225390
rect 136357 225314 136423 225317
rect 142245 225314 142311 225317
rect 136357 225312 142311 225314
rect 136357 225256 136362 225312
rect 136418 225256 142250 225312
rect 142306 225256 142311 225312
rect 136357 225254 142311 225256
rect 136357 225251 136423 225254
rect 142245 225251 142311 225254
rect 176469 225314 176535 225317
rect 176745 225314 176811 225317
rect 176469 225312 176811 225314
rect 176469 225256 176474 225312
rect 176530 225256 176750 225312
rect 176806 225256 176811 225312
rect 176469 225254 176811 225256
rect 176469 225251 176535 225254
rect 176745 225251 176811 225254
rect 660205 225314 660271 225317
rect 667013 225314 667079 225317
rect 660205 225312 667079 225314
rect 660205 225256 660210 225312
rect 660266 225256 667018 225312
rect 667074 225256 667079 225312
rect 660205 225254 667079 225256
rect 660205 225251 660271 225254
rect 667013 225251 667079 225254
rect 185577 225178 185643 225181
rect 195513 225178 195579 225181
rect 185577 225176 195579 225178
rect 185577 225120 185582 225176
rect 185638 225120 195518 225176
rect 195574 225120 195579 225176
rect 185577 225118 195579 225120
rect 185577 225115 185643 225118
rect 195513 225115 195579 225118
rect 202597 225178 202663 225181
rect 205081 225178 205147 225181
rect 202597 225176 205147 225178
rect 202597 225120 202602 225176
rect 202658 225120 205086 225176
rect 205142 225120 205147 225176
rect 202597 225118 205147 225120
rect 202597 225115 202663 225118
rect 205081 225115 205147 225118
rect 671838 225116 671844 225180
rect 671908 225178 671914 225180
rect 674189 225178 674255 225181
rect 671908 225176 674255 225178
rect 671908 225120 674194 225176
rect 674250 225120 674255 225176
rect 671908 225118 674255 225120
rect 671908 225116 671914 225118
rect 674189 225115 674255 225118
rect 166533 225042 166599 225045
rect 171041 225042 171107 225045
rect 166533 225040 171107 225042
rect 166533 224984 166538 225040
rect 166594 224984 171046 225040
rect 171102 224984 171107 225040
rect 166533 224982 171107 224984
rect 166533 224979 166599 224982
rect 171041 224979 171107 224982
rect 655421 225042 655487 225045
rect 671245 225042 671311 225045
rect 655421 225040 671311 225042
rect 655421 224984 655426 225040
rect 655482 224984 671250 225040
rect 671306 224984 671311 225040
rect 655421 224982 671311 224984
rect 655421 224979 655487 224982
rect 671245 224979 671311 224982
rect 672901 224906 672967 224909
rect 673310 224906 673316 224908
rect 672901 224904 673316 224906
rect 672901 224848 672906 224904
rect 672962 224848 673316 224904
rect 672901 224846 673316 224848
rect 672901 224843 672967 224846
rect 673310 224844 673316 224846
rect 673380 224844 673386 224908
rect 671245 224770 671311 224773
rect 672073 224770 672139 224773
rect 671245 224768 672139 224770
rect 671245 224712 671250 224768
rect 671306 224712 672078 224768
rect 672134 224712 672139 224768
rect 671245 224710 672139 224712
rect 671245 224707 671311 224710
rect 672073 224707 672139 224710
rect 157333 224498 157399 224501
rect 162945 224498 163011 224501
rect 157333 224496 163011 224498
rect 157333 224440 157338 224496
rect 157394 224440 162950 224496
rect 163006 224440 163011 224496
rect 157333 224438 163011 224440
rect 157333 224435 157399 224438
rect 162945 224435 163011 224438
rect 658181 224498 658247 224501
rect 671889 224498 671955 224501
rect 675201 224498 675267 224501
rect 658181 224496 659670 224498
rect 658181 224440 658186 224496
rect 658242 224440 659670 224496
rect 658181 224438 659670 224440
rect 658181 224435 658247 224438
rect 152733 224362 152799 224365
rect 137970 224360 152799 224362
rect 137970 224304 152738 224360
rect 152794 224304 152799 224360
rect 137970 224302 152799 224304
rect 68921 224226 68987 224229
rect 137970 224226 138030 224302
rect 152733 224299 152799 224302
rect 68921 224224 138030 224226
rect 68921 224168 68926 224224
rect 68982 224168 138030 224224
rect 68921 224166 138030 224168
rect 170949 224226 171015 224229
rect 171409 224226 171475 224229
rect 170949 224224 171475 224226
rect 170949 224168 170954 224224
rect 171010 224168 171414 224224
rect 171470 224168 171475 224224
rect 170949 224166 171475 224168
rect 659610 224226 659670 224438
rect 671889 224496 675267 224498
rect 671889 224440 671894 224496
rect 671950 224440 675206 224496
rect 675262 224440 675267 224496
rect 671889 224438 675267 224440
rect 671889 224435 671955 224438
rect 675201 224435 675267 224438
rect 667013 224226 667079 224229
rect 659610 224224 667079 224226
rect 659610 224168 667018 224224
rect 667074 224168 667079 224224
rect 659610 224166 667079 224168
rect 68921 224163 68987 224166
rect 170949 224163 171015 224166
rect 171409 224163 171475 224166
rect 667013 224163 667079 224166
rect 671654 224164 671660 224228
rect 671724 224226 671730 224228
rect 675385 224226 675451 224229
rect 671724 224224 675451 224226
rect 671724 224168 675390 224224
rect 675446 224168 675451 224224
rect 671724 224166 675451 224168
rect 671724 224164 671730 224166
rect 675385 224163 675451 224166
rect 157425 224090 157491 224093
rect 154622 224088 157491 224090
rect 154622 224032 157430 224088
rect 157486 224032 157491 224088
rect 154622 224030 157491 224032
rect 154622 223991 154682 224030
rect 157425 224027 157491 224030
rect 154573 223986 154682 223991
rect 141417 223954 141483 223957
rect 145373 223954 145439 223957
rect 141417 223952 145439 223954
rect 141417 223896 141422 223952
rect 141478 223896 145378 223952
rect 145434 223896 145439 223952
rect 141417 223894 145439 223896
rect 141417 223891 141483 223894
rect 145373 223891 145439 223894
rect 146201 223954 146267 223957
rect 147673 223954 147739 223957
rect 146201 223952 147739 223954
rect 146201 223896 146206 223952
rect 146262 223896 147678 223952
rect 147734 223896 147739 223952
rect 154573 223930 154578 223986
rect 154634 223930 154682 223986
rect 154573 223928 154682 223930
rect 163957 223954 164023 223957
rect 170949 223954 171015 223957
rect 163957 223952 171015 223954
rect 154573 223925 154639 223928
rect 146201 223894 147739 223896
rect 146201 223891 146267 223894
rect 147673 223891 147739 223894
rect 163957 223896 163962 223952
rect 164018 223896 170954 223952
rect 171010 223896 171015 223952
rect 163957 223894 171015 223896
rect 163957 223891 164023 223894
rect 170949 223891 171015 223894
rect 658917 223954 658983 223957
rect 670601 223954 670667 223957
rect 658917 223952 670667 223954
rect 658917 223896 658922 223952
rect 658978 223896 670606 223952
rect 670662 223896 670667 223952
rect 658917 223894 670667 223896
rect 658917 223891 658983 223894
rect 670601 223891 670667 223894
rect 671102 223892 671108 223956
rect 671172 223954 671178 223956
rect 673453 223954 673519 223957
rect 671172 223952 673519 223954
rect 671172 223896 673458 223952
rect 673514 223896 673519 223952
rect 671172 223894 673519 223896
rect 671172 223892 671178 223894
rect 673453 223891 673519 223894
rect 151721 223818 151787 223821
rect 156873 223818 156939 223821
rect 679249 223818 679315 223821
rect 151721 223816 156939 223818
rect 151721 223760 151726 223816
rect 151782 223760 156878 223816
rect 156934 223760 156939 223816
rect 151721 223758 156939 223760
rect 151721 223755 151787 223758
rect 156873 223755 156939 223758
rect 679206 223816 679315 223818
rect 679206 223760 679254 223816
rect 679310 223760 679315 223816
rect 679206 223755 679315 223760
rect 656617 223682 656683 223685
rect 670509 223682 670575 223685
rect 656617 223680 670575 223682
rect 656617 223624 656622 223680
rect 656678 223624 670514 223680
rect 670570 223624 670575 223680
rect 656617 223622 670575 223624
rect 656617 223619 656683 223622
rect 670509 223619 670575 223622
rect 673494 223620 673500 223684
rect 673564 223682 673570 223684
rect 673913 223682 673979 223685
rect 673564 223680 673979 223682
rect 673564 223624 673918 223680
rect 673974 223624 673979 223680
rect 673564 223622 673979 223624
rect 673564 223620 673570 223622
rect 673913 223619 673979 223622
rect 679206 223516 679266 223755
rect 157241 223410 157307 223413
rect 157425 223410 157491 223413
rect 157241 223408 157491 223410
rect 157241 223352 157246 223408
rect 157302 223352 157430 223408
rect 157486 223352 157491 223408
rect 157241 223350 157491 223352
rect 157241 223347 157307 223350
rect 157425 223347 157491 223350
rect 158621 223410 158687 223413
rect 166441 223410 166507 223413
rect 158621 223408 166507 223410
rect 158621 223352 158626 223408
rect 158682 223352 166446 223408
rect 166502 223352 166507 223408
rect 158621 223350 166507 223352
rect 158621 223347 158687 223350
rect 166441 223347 166507 223350
rect 166257 223138 166323 223141
rect 170397 223138 170463 223141
rect 166257 223136 170463 223138
rect 166257 223080 166262 223136
rect 166318 223080 170402 223136
rect 170458 223080 170463 223136
rect 166257 223078 170463 223080
rect 166257 223075 166323 223078
rect 170397 223075 170463 223078
rect 651281 223138 651347 223141
rect 667841 223138 667907 223141
rect 683665 223138 683731 223141
rect 651281 223136 667907 223138
rect 651281 223080 651286 223136
rect 651342 223080 667846 223136
rect 667902 223080 667907 223136
rect 651281 223078 667907 223080
rect 683652 223136 683731 223138
rect 683652 223080 683670 223136
rect 683726 223080 683731 223136
rect 683652 223078 683731 223080
rect 651281 223075 651347 223078
rect 667841 223075 667907 223078
rect 683665 223075 683731 223078
rect 40677 222866 40743 222869
rect 62941 222866 63007 222869
rect 40677 222864 63007 222866
rect 40677 222808 40682 222864
rect 40738 222808 62946 222864
rect 63002 222808 63007 222864
rect 40677 222806 63007 222808
rect 40677 222803 40743 222806
rect 62941 222803 63007 222806
rect 123477 222866 123543 222869
rect 165613 222866 165679 222869
rect 123477 222864 165679 222866
rect 123477 222808 123482 222864
rect 123538 222808 165618 222864
rect 165674 222808 165679 222864
rect 123477 222806 165679 222808
rect 123477 222803 123543 222806
rect 165613 222803 165679 222806
rect 651833 222866 651899 222869
rect 666829 222866 666895 222869
rect 651833 222864 666895 222866
rect 651833 222808 651838 222864
rect 651894 222808 666834 222864
rect 666890 222808 666895 222864
rect 651833 222806 666895 222808
rect 651833 222803 651899 222806
rect 666829 222803 666895 222806
rect 683205 222730 683271 222733
rect 683205 222728 683284 222730
rect 683205 222672 683210 222728
rect 683266 222672 683284 222728
rect 683205 222670 683284 222672
rect 683205 222667 683271 222670
rect 166073 222594 166139 222597
rect 166993 222594 167059 222597
rect 166073 222592 167059 222594
rect 166073 222536 166078 222592
rect 166134 222536 166998 222592
rect 167054 222536 167059 222592
rect 166073 222534 167059 222536
rect 166073 222531 166139 222534
rect 166993 222531 167059 222534
rect 174813 222594 174879 222597
rect 175457 222594 175523 222597
rect 174813 222592 175523 222594
rect 174813 222536 174818 222592
rect 174874 222536 175462 222592
rect 175518 222536 175523 222592
rect 174813 222534 175523 222536
rect 174813 222531 174879 222534
rect 175457 222531 175523 222534
rect 570505 222594 570571 222597
rect 574829 222594 574895 222597
rect 570505 222592 574895 222594
rect 570505 222536 570510 222592
rect 570566 222536 574834 222592
rect 574890 222536 574895 222592
rect 570505 222534 574895 222536
rect 570505 222531 570571 222534
rect 574829 222531 574895 222534
rect 155309 222458 155375 222461
rect 157241 222458 157307 222461
rect 155309 222456 157307 222458
rect 155309 222400 155314 222456
rect 155370 222400 157246 222456
rect 157302 222400 157307 222456
rect 155309 222398 157307 222400
rect 155309 222395 155375 222398
rect 157241 222395 157307 222398
rect 203517 222458 203583 222461
rect 205081 222458 205147 222461
rect 203517 222456 205147 222458
rect 203517 222400 203522 222456
rect 203578 222400 205086 222456
rect 205142 222400 205147 222456
rect 203517 222398 205147 222400
rect 203517 222395 203583 222398
rect 205081 222395 205147 222398
rect 166809 222322 166875 222325
rect 168097 222322 168163 222325
rect 166809 222320 168163 222322
rect 166809 222264 166814 222320
rect 166870 222264 168102 222320
rect 168158 222264 168163 222320
rect 166809 222262 168163 222264
rect 166809 222259 166875 222262
rect 168097 222259 168163 222262
rect 562869 222322 562935 222325
rect 563329 222322 563395 222325
rect 562869 222320 563395 222322
rect 562869 222264 562874 222320
rect 562930 222264 563334 222320
rect 563390 222264 563395 222320
rect 562869 222262 563395 222264
rect 562869 222259 562935 222262
rect 563329 222259 563395 222262
rect 564893 222322 564959 222325
rect 567193 222322 567259 222325
rect 572437 222322 572503 222325
rect 564893 222320 572503 222322
rect 564893 222264 564898 222320
rect 564954 222264 567198 222320
rect 567254 222264 572442 222320
rect 572498 222264 572503 222320
rect 564893 222262 572503 222264
rect 564893 222259 564959 222262
rect 567193 222259 567259 222262
rect 572437 222259 572503 222262
rect 674741 222322 674807 222325
rect 674741 222320 676292 222322
rect 674741 222264 674746 222320
rect 674802 222264 676292 222320
rect 674741 222262 676292 222264
rect 674741 222259 674807 222262
rect 147305 222186 147371 222189
rect 152089 222186 152155 222189
rect 147305 222184 152155 222186
rect 147305 222128 147310 222184
rect 147366 222128 152094 222184
rect 152150 222128 152155 222184
rect 147305 222126 152155 222128
rect 147305 222123 147371 222126
rect 152089 222123 152155 222126
rect 171133 222186 171199 222189
rect 177573 222186 177639 222189
rect 171133 222184 177639 222186
rect 171133 222128 171138 222184
rect 171194 222128 177578 222184
rect 177634 222128 177639 222184
rect 171133 222126 177639 222128
rect 171133 222123 171199 222126
rect 177573 222123 177639 222126
rect 562317 222052 562383 222053
rect 562317 222050 562364 222052
rect 562272 222048 562364 222050
rect 562272 221992 562322 222048
rect 562272 221990 562364 221992
rect 562317 221988 562364 221990
rect 562428 221988 562434 222052
rect 562685 222050 562751 222053
rect 563513 222050 563579 222053
rect 562685 222048 563579 222050
rect 562685 221992 562690 222048
rect 562746 221992 563518 222048
rect 563574 221992 563579 222048
rect 562685 221990 563579 221992
rect 562317 221987 562383 221988
rect 562685 221987 562751 221990
rect 563513 221987 563579 221990
rect 564566 221988 564572 222052
rect 564636 222050 564642 222052
rect 565077 222050 565143 222053
rect 571057 222050 571123 222053
rect 564636 222048 571123 222050
rect 564636 221992 565082 222048
rect 565138 221992 571062 222048
rect 571118 221992 571123 222048
rect 564636 221990 571123 221992
rect 564636 221988 564642 221990
rect 565077 221987 565143 221990
rect 571057 221987 571123 221990
rect 572846 221988 572852 222052
rect 572916 222050 572922 222052
rect 576025 222050 576091 222053
rect 572916 222048 576091 222050
rect 572916 221992 576030 222048
rect 576086 221992 576091 222048
rect 572916 221990 576091 221992
rect 572916 221988 572922 221990
rect 576025 221987 576091 221990
rect 591941 222050 592007 222053
rect 599301 222050 599367 222053
rect 591941 222048 599367 222050
rect 591941 221992 591946 222048
rect 592002 221992 599306 222048
rect 599362 221992 599367 222048
rect 591941 221990 599367 221992
rect 591941 221987 592007 221990
rect 599301 221987 599367 221990
rect 665265 222050 665331 222053
rect 673453 222050 673519 222053
rect 665265 222048 673519 222050
rect 665265 221992 665270 222048
rect 665326 221992 673458 222048
rect 673514 221992 673519 222048
rect 665265 221990 673519 221992
rect 665265 221987 665331 221990
rect 673453 221987 673519 221990
rect 147489 221914 147555 221917
rect 149053 221914 149119 221917
rect 147489 221912 149119 221914
rect 147489 221856 147494 221912
rect 147550 221856 149058 221912
rect 149114 221856 149119 221912
rect 147489 221854 149119 221856
rect 147489 221851 147555 221854
rect 149053 221851 149119 221854
rect 170857 221914 170923 221917
rect 171409 221914 171475 221917
rect 170857 221912 171475 221914
rect 170857 221856 170862 221912
rect 170918 221856 171414 221912
rect 171470 221856 171475 221912
rect 170857 221854 171475 221856
rect 170857 221851 170923 221854
rect 171409 221851 171475 221854
rect 674649 221914 674715 221917
rect 674649 221912 676292 221914
rect 674649 221856 674654 221912
rect 674710 221856 676292 221912
rect 674649 221854 676292 221856
rect 674649 221851 674715 221854
rect 138565 221778 138631 221781
rect 146569 221778 146635 221781
rect 138565 221776 146635 221778
rect 138565 221720 138570 221776
rect 138626 221720 146574 221776
rect 146630 221720 146635 221776
rect 138565 221718 146635 221720
rect 138565 221715 138631 221718
rect 146569 221715 146635 221718
rect 519721 221778 519787 221781
rect 618253 221778 618319 221781
rect 519721 221776 618319 221778
rect 519721 221720 519726 221776
rect 519782 221720 618258 221776
rect 618314 221720 618319 221776
rect 519721 221718 618319 221720
rect 519721 221715 519787 221718
rect 618253 221715 618319 221718
rect 101857 221506 101923 221509
rect 178033 221506 178099 221509
rect 101857 221504 178099 221506
rect 101857 221448 101862 221504
rect 101918 221448 178038 221504
rect 178094 221448 178099 221504
rect 101857 221446 178099 221448
rect 101857 221443 101923 221446
rect 178033 221443 178099 221446
rect 517789 221506 517855 221509
rect 517973 221506 518039 221509
rect 616873 221506 616939 221509
rect 517789 221504 616939 221506
rect 517789 221448 517794 221504
rect 517850 221448 517978 221504
rect 518034 221448 616878 221504
rect 616934 221448 616939 221504
rect 517789 221446 616939 221448
rect 517789 221443 517855 221446
rect 517973 221443 518039 221446
rect 616873 221443 616939 221446
rect 657997 221506 658063 221509
rect 673637 221506 673703 221509
rect 657997 221504 673703 221506
rect 657997 221448 658002 221504
rect 658058 221448 673642 221504
rect 673698 221448 673703 221504
rect 657997 221446 673703 221448
rect 657997 221443 658063 221446
rect 673637 221443 673703 221446
rect 678421 221506 678487 221509
rect 678421 221504 678500 221506
rect 678421 221448 678426 221504
rect 678482 221448 678500 221504
rect 678421 221446 678500 221448
rect 678421 221443 678487 221446
rect 178309 221370 178375 221373
rect 185117 221370 185183 221373
rect 178309 221368 185183 221370
rect 178309 221312 178314 221368
rect 178370 221312 185122 221368
rect 185178 221312 185183 221368
rect 178309 221310 185183 221312
rect 178309 221307 178375 221310
rect 185117 221307 185183 221310
rect 142429 221234 142495 221237
rect 144177 221234 144243 221237
rect 142429 221232 144243 221234
rect 142429 221176 142434 221232
rect 142490 221176 144182 221232
rect 144238 221176 144243 221232
rect 142429 221174 144243 221176
rect 142429 221171 142495 221174
rect 144177 221171 144243 221174
rect 505921 221234 505987 221237
rect 597921 221234 597987 221237
rect 505921 221232 597987 221234
rect 505921 221176 505926 221232
rect 505982 221176 597926 221232
rect 597982 221176 597987 221232
rect 505921 221174 597987 221176
rect 505921 221171 505987 221174
rect 597921 221171 597987 221174
rect 659377 221234 659443 221237
rect 674925 221234 674991 221237
rect 659377 221232 674991 221234
rect 659377 221176 659382 221232
rect 659438 221176 674930 221232
rect 674986 221176 674991 221232
rect 659377 221174 674991 221176
rect 659377 221171 659443 221174
rect 674925 221171 674991 221174
rect 675158 221038 676292 221098
rect 487061 220962 487127 220965
rect 611445 220962 611511 220965
rect 487061 220960 611511 220962
rect 487061 220904 487066 220960
rect 487122 220904 611450 220960
rect 611506 220904 611511 220960
rect 487061 220902 611511 220904
rect 487061 220899 487127 220902
rect 611445 220899 611511 220902
rect 667841 220962 667907 220965
rect 675158 220962 675218 221038
rect 667841 220960 675218 220962
rect 667841 220904 667846 220960
rect 667902 220904 675218 220960
rect 667841 220902 675218 220904
rect 667841 220899 667907 220902
rect 141049 220826 141115 220829
rect 146385 220826 146451 220829
rect 141049 220824 146451 220826
rect 141049 220768 141054 220824
rect 141110 220768 146390 220824
rect 146446 220768 146451 220824
rect 141049 220766 146451 220768
rect 141049 220763 141115 220766
rect 146385 220763 146451 220766
rect 147213 220826 147279 220829
rect 148409 220826 148475 220829
rect 147213 220824 148475 220826
rect 147213 220768 147218 220824
rect 147274 220768 148414 220824
rect 148470 220768 148475 220824
rect 147213 220766 148475 220768
rect 147213 220763 147279 220766
rect 148409 220763 148475 220766
rect 150617 220826 150683 220829
rect 156137 220826 156203 220829
rect 150617 220824 156203 220826
rect 150617 220768 150622 220824
rect 150678 220768 156142 220824
rect 156198 220768 156203 220824
rect 150617 220766 156203 220768
rect 150617 220763 150683 220766
rect 156137 220763 156203 220766
rect 194869 220826 194935 220829
rect 196065 220826 196131 220829
rect 194869 220824 196131 220826
rect 194869 220768 194874 220824
rect 194930 220768 196070 220824
rect 196126 220768 196131 220824
rect 194869 220766 196131 220768
rect 194869 220763 194935 220766
rect 196065 220763 196131 220766
rect 548333 220690 548399 220693
rect 552381 220690 552447 220693
rect 554037 220690 554103 220693
rect 548333 220688 554103 220690
rect 548333 220632 548338 220688
rect 548394 220632 552386 220688
rect 552442 220632 554042 220688
rect 554098 220632 554103 220688
rect 548333 220630 554103 220632
rect 548333 220627 548399 220630
rect 552381 220627 552447 220630
rect 554037 220627 554103 220630
rect 563421 220690 563487 220693
rect 563421 220688 572362 220690
rect 563421 220632 563426 220688
rect 563482 220632 572362 220688
rect 563421 220630 572362 220632
rect 563421 220627 563487 220630
rect 153745 220554 153811 220557
rect 563237 220554 563303 220557
rect 137970 220552 153811 220554
rect 137970 220496 153750 220552
rect 153806 220496 153811 220552
rect 137970 220494 153811 220496
rect 72877 220418 72943 220421
rect 137970 220418 138030 220494
rect 153745 220491 153811 220494
rect 554224 220552 563303 220554
rect 554224 220496 563242 220552
rect 563298 220496 563303 220552
rect 554224 220494 563303 220496
rect 572302 220554 572362 220630
rect 572846 220628 572852 220692
rect 572916 220690 572922 220692
rect 575197 220690 575263 220693
rect 572916 220688 575263 220690
rect 572916 220632 575202 220688
rect 575258 220632 575263 220688
rect 572916 220630 575263 220632
rect 572916 220628 572922 220630
rect 575197 220627 575263 220630
rect 653029 220690 653095 220693
rect 671245 220690 671311 220693
rect 653029 220688 671311 220690
rect 653029 220632 653034 220688
rect 653090 220632 671250 220688
rect 671306 220632 671311 220688
rect 653029 220630 671311 220632
rect 653029 220627 653095 220630
rect 671245 220627 671311 220630
rect 678237 220690 678303 220693
rect 678237 220688 678316 220690
rect 678237 220632 678242 220688
rect 678298 220632 678316 220688
rect 678237 220630 678316 220632
rect 678237 220627 678303 220630
rect 572621 220554 572687 220557
rect 673821 220554 673887 220557
rect 572302 220552 572687 220554
rect 572302 220496 572626 220552
rect 572682 220496 572687 220552
rect 572302 220494 572687 220496
rect 72877 220416 138030 220418
rect 72877 220360 72882 220416
rect 72938 220360 138030 220416
rect 72877 220358 138030 220360
rect 157609 220418 157675 220421
rect 161565 220418 161631 220421
rect 157609 220416 161631 220418
rect 157609 220360 157614 220416
rect 157670 220360 161570 220416
rect 161626 220360 161631 220416
rect 157609 220358 161631 220360
rect 72877 220355 72943 220358
rect 157609 220355 157675 220358
rect 161565 220355 161631 220358
rect 532693 220418 532759 220421
rect 534165 220418 534231 220421
rect 532693 220416 534231 220418
rect 532693 220360 532698 220416
rect 532754 220360 534170 220416
rect 534226 220360 534231 220416
rect 532693 220358 534231 220360
rect 532693 220355 532759 220358
rect 534165 220355 534231 220358
rect 553669 220418 553735 220421
rect 554224 220418 554284 220494
rect 563237 220491 563303 220494
rect 572621 220491 572687 220494
rect 671478 220552 673887 220554
rect 671478 220496 673826 220552
rect 673882 220496 673887 220552
rect 671478 220494 673887 220496
rect 553669 220416 554284 220418
rect 553669 220360 553674 220416
rect 553730 220360 554284 220416
rect 553669 220358 554284 220360
rect 563789 220418 563855 220421
rect 578233 220420 578299 220421
rect 572110 220418 572116 220420
rect 563789 220416 572116 220418
rect 563789 220360 563794 220416
rect 563850 220360 572116 220416
rect 563789 220358 572116 220360
rect 553669 220355 553735 220358
rect 563789 220355 563855 220358
rect 572110 220356 572116 220358
rect 572180 220356 572186 220420
rect 578182 220418 578188 220420
rect 578142 220358 578188 220418
rect 578252 220416 578299 220420
rect 578294 220360 578299 220416
rect 578182 220356 578188 220358
rect 578252 220356 578299 220360
rect 578233 220355 578299 220356
rect 592033 220418 592099 220421
rect 599301 220418 599367 220421
rect 592033 220416 599367 220418
rect 592033 220360 592038 220416
rect 592094 220360 599306 220416
rect 599362 220360 599367 220416
rect 592033 220358 599367 220360
rect 592033 220355 592099 220358
rect 599301 220355 599367 220358
rect 643185 220418 643251 220421
rect 663425 220418 663491 220421
rect 643185 220416 663491 220418
rect 643185 220360 643190 220416
rect 643246 220360 663430 220416
rect 663486 220360 663491 220416
rect 643185 220358 663491 220360
rect 643185 220355 643251 220358
rect 663425 220355 663491 220358
rect 165153 220282 165219 220285
rect 167637 220282 167703 220285
rect 165153 220280 167703 220282
rect 165153 220224 165158 220280
rect 165214 220224 167642 220280
rect 167698 220224 167703 220280
rect 165153 220222 167703 220224
rect 165153 220219 165219 220222
rect 167637 220219 167703 220222
rect 543917 220282 543983 220285
rect 547137 220282 547203 220285
rect 543917 220280 547203 220282
rect 543917 220224 543922 220280
rect 543978 220224 547142 220280
rect 547198 220224 547203 220280
rect 543917 220222 547203 220224
rect 543917 220219 543983 220222
rect 547137 220219 547203 220222
rect 552841 220282 552907 220285
rect 554589 220282 554655 220285
rect 572805 220282 572871 220285
rect 573449 220282 573515 220285
rect 552841 220280 553594 220282
rect 552841 220224 552846 220280
rect 552902 220224 553594 220280
rect 552841 220222 553594 220224
rect 552841 220219 552907 220222
rect 70025 220146 70091 220149
rect 150801 220146 150867 220149
rect 70025 220144 150867 220146
rect 70025 220088 70030 220144
rect 70086 220088 150806 220144
rect 150862 220088 150867 220144
rect 70025 220086 150867 220088
rect 70025 220083 70091 220086
rect 150801 220083 150867 220086
rect 544929 220010 544995 220013
rect 553347 220010 553413 220013
rect 544929 220008 553413 220010
rect 544929 219952 544934 220008
rect 544990 219952 553352 220008
rect 553408 219952 553413 220008
rect 544929 219950 553413 219952
rect 553534 220010 553594 220222
rect 554589 220280 563162 220282
rect 554589 220224 554594 220280
rect 554650 220224 563162 220280
rect 554589 220222 563162 220224
rect 554589 220219 554655 220222
rect 563102 220146 563162 220222
rect 572302 220280 572871 220282
rect 572302 220224 572810 220280
rect 572866 220224 572871 220280
rect 572302 220222 572871 220224
rect 563605 220146 563671 220149
rect 564617 220146 564683 220149
rect 572302 220146 572362 220222
rect 572805 220219 572871 220222
rect 573038 220280 573515 220282
rect 573038 220224 573454 220280
rect 573510 220224 573515 220280
rect 573038 220222 573515 220224
rect 563102 220144 563671 220146
rect 563102 220088 563610 220144
rect 563666 220088 563671 220144
rect 563102 220086 563671 220088
rect 563605 220083 563671 220086
rect 563792 220144 564683 220146
rect 563792 220088 564622 220144
rect 564678 220088 564683 220144
rect 563792 220086 564683 220088
rect 553534 219950 563070 220010
rect 544929 219947 544995 219950
rect 553347 219947 553413 219950
rect 563010 219908 563070 219950
rect 563792 219908 563852 220086
rect 564617 220083 564683 220086
rect 569910 220086 572362 220146
rect 569910 220010 569970 220086
rect 573038 220010 573098 220222
rect 573449 220219 573515 220222
rect 573909 220284 573975 220285
rect 573909 220280 573956 220284
rect 574020 220282 574026 220284
rect 582741 220282 582807 220285
rect 591849 220282 591915 220285
rect 573909 220224 573914 220280
rect 573909 220220 573956 220224
rect 574020 220222 574066 220282
rect 582741 220280 591915 220282
rect 582741 220224 582746 220280
rect 582802 220224 591854 220280
rect 591910 220224 591915 220280
rect 582741 220222 591915 220224
rect 574020 220220 574026 220222
rect 573909 220219 573975 220220
rect 582741 220219 582807 220222
rect 591849 220219 591915 220222
rect 637665 220146 637731 220149
rect 671478 220146 671538 220494
rect 673821 220491 673887 220494
rect 673545 220282 673611 220285
rect 673545 220280 676292 220282
rect 673545 220224 673550 220280
rect 673606 220224 676292 220280
rect 673545 220222 676292 220224
rect 673545 220219 673611 220222
rect 637665 220144 671538 220146
rect 637665 220088 637670 220144
rect 637726 220088 671538 220144
rect 637665 220086 671538 220088
rect 637665 220083 637731 220086
rect 564758 219950 569970 220010
rect 572440 219950 573098 220010
rect 573265 220010 573331 220013
rect 582005 220010 582071 220013
rect 573265 220008 582071 220010
rect 573265 219952 573270 220008
rect 573326 219952 582010 220008
rect 582066 219952 582071 220008
rect 573265 219950 582071 219952
rect 563010 219848 563852 219908
rect 564065 219908 564131 219911
rect 564758 219908 564818 219950
rect 564065 219906 564818 219908
rect 564065 219850 564070 219906
rect 564126 219850 564818 219906
rect 564065 219848 564818 219850
rect 570873 219908 570939 219911
rect 572440 219908 572500 219950
rect 573265 219947 573331 219950
rect 582005 219947 582071 219950
rect 582557 220010 582623 220013
rect 592033 220010 592099 220013
rect 582557 220008 592099 220010
rect 582557 219952 582562 220008
rect 582618 219952 592038 220008
rect 592094 219952 592099 220008
rect 582557 219950 592099 219952
rect 582557 219947 582623 219950
rect 592033 219947 592099 219950
rect 570873 219906 572500 219908
rect 570873 219850 570878 219906
rect 570934 219850 572500 219906
rect 570873 219848 572500 219850
rect 671245 219874 671311 219877
rect 673913 219874 673979 219877
rect 683481 219874 683547 219877
rect 671245 219872 673979 219874
rect 564065 219845 564131 219848
rect 570873 219845 570939 219848
rect 671245 219816 671250 219872
rect 671306 219816 673918 219872
rect 673974 219816 673979 219872
rect 671245 219814 673979 219816
rect 683468 219872 683547 219874
rect 683468 219816 683486 219872
rect 683542 219816 683547 219872
rect 683468 219814 683547 219816
rect 671245 219811 671311 219814
rect 673913 219811 673979 219814
rect 683481 219811 683547 219814
rect 494881 219738 494947 219741
rect 630765 219738 630831 219741
rect 494881 219736 630831 219738
rect 494881 219680 494886 219736
rect 494942 219680 630770 219736
rect 630826 219680 630831 219736
rect 494881 219678 630831 219680
rect 494881 219675 494947 219678
rect 630765 219675 630831 219678
rect 484853 219602 484919 219605
rect 663425 219602 663491 219605
rect 671245 219602 671311 219605
rect 484853 219600 489930 219602
rect 484853 219544 484858 219600
rect 484914 219544 489930 219600
rect 484853 219542 489930 219544
rect 484853 219539 484919 219542
rect 489870 219466 489930 219542
rect 663425 219600 671311 219602
rect 663425 219544 663430 219600
rect 663486 219544 671250 219600
rect 671306 219544 671311 219600
rect 663425 219542 671311 219544
rect 663425 219539 663491 219542
rect 671245 219539 671311 219542
rect 631225 219466 631291 219469
rect 489870 219464 631291 219466
rect 489870 219408 631230 219464
rect 631286 219408 631291 219464
rect 489870 219406 631291 219408
rect 631225 219403 631291 219406
rect 671889 219466 671955 219469
rect 671889 219464 676292 219466
rect 671889 219408 671894 219464
rect 671950 219408 676292 219464
rect 671889 219406 676292 219408
rect 671889 219403 671955 219406
rect 487429 219332 487495 219333
rect 487429 219328 487476 219332
rect 487540 219330 487546 219332
rect 487429 219272 487434 219328
rect 487429 219268 487476 219272
rect 487540 219270 487586 219330
rect 487540 219268 487546 219270
rect 487429 219267 487495 219268
rect 503161 219194 503227 219197
rect 507209 219194 507275 219197
rect 503161 219192 507275 219194
rect 503161 219136 503166 219192
rect 503222 219136 507214 219192
rect 507270 219136 507275 219192
rect 503161 219134 507275 219136
rect 503161 219131 503227 219134
rect 507209 219131 507275 219134
rect 507393 219194 507459 219197
rect 509233 219194 509299 219197
rect 507393 219192 509299 219194
rect 507393 219136 507398 219192
rect 507454 219136 509238 219192
rect 509294 219136 509299 219192
rect 507393 219134 509299 219136
rect 507393 219131 507459 219134
rect 509233 219131 509299 219134
rect 509509 219194 509575 219197
rect 518985 219194 519051 219197
rect 509509 219192 519051 219194
rect 509509 219136 509514 219192
rect 509570 219136 518990 219192
rect 519046 219136 519051 219192
rect 509509 219134 519051 219136
rect 509509 219131 509575 219134
rect 518985 219131 519051 219134
rect 519169 219194 519235 219197
rect 617333 219194 617399 219197
rect 519169 219192 617399 219194
rect 519169 219136 519174 219192
rect 519230 219136 617338 219192
rect 617394 219136 617399 219192
rect 519169 219134 617399 219136
rect 519169 219131 519235 219134
rect 617333 219131 617399 219134
rect 655237 219194 655303 219197
rect 672073 219194 672139 219197
rect 655237 219192 672139 219194
rect 655237 219136 655242 219192
rect 655298 219136 672078 219192
rect 672134 219136 672139 219192
rect 655237 219134 672139 219136
rect 655237 219131 655303 219134
rect 672073 219131 672139 219134
rect 675017 219058 675083 219061
rect 675017 219056 676292 219058
rect 675017 219000 675022 219056
rect 675078 219000 676292 219056
rect 675017 218998 676292 219000
rect 675017 218995 675083 218998
rect 505185 218922 505251 218925
rect 509233 218922 509299 218925
rect 505185 218920 509299 218922
rect 505185 218864 505190 218920
rect 505246 218864 509238 218920
rect 509294 218864 509299 218920
rect 505185 218862 509299 218864
rect 505185 218859 505251 218862
rect 509233 218859 509299 218862
rect 518847 218922 518913 218925
rect 606201 218922 606267 218925
rect 612733 218922 612799 218925
rect 518847 218920 606267 218922
rect 518847 218864 518852 218920
rect 518908 218864 606206 218920
rect 606262 218864 606267 218920
rect 518847 218862 606267 218864
rect 518847 218859 518913 218862
rect 606201 218859 606267 218862
rect 606526 218920 612799 218922
rect 606526 218864 612738 218920
rect 612794 218864 612799 218920
rect 606526 218862 612799 218864
rect 149329 218786 149395 218789
rect 153929 218786 153995 218789
rect 518709 218786 518775 218789
rect 149329 218784 153995 218786
rect 149329 218728 149334 218784
rect 149390 218728 153934 218784
rect 153990 218728 153995 218784
rect 149329 218726 153995 218728
rect 149329 218723 149395 218726
rect 153929 218723 153995 218726
rect 509558 218784 518775 218786
rect 509558 218728 518714 218784
rect 518770 218728 518775 218784
rect 509558 218726 518775 218728
rect 140221 218650 140287 218653
rect 143625 218650 143691 218653
rect 140221 218648 143691 218650
rect 140221 218592 140226 218648
rect 140282 218592 143630 218648
rect 143686 218592 143691 218648
rect 140221 218590 143691 218592
rect 140221 218587 140287 218590
rect 143625 218587 143691 218590
rect 489913 218650 489979 218653
rect 491201 218652 491267 218653
rect 491150 218650 491156 218652
rect 489913 218648 491156 218650
rect 491220 218650 491267 218652
rect 497457 218650 497523 218653
rect 509558 218650 509618 218726
rect 518709 218723 518775 218726
rect 491220 218648 491312 218650
rect 489913 218592 489918 218648
rect 489974 218592 491156 218648
rect 491262 218592 491312 218648
rect 489913 218590 491156 218592
rect 489913 218587 489979 218590
rect 491150 218588 491156 218590
rect 491220 218590 491312 218592
rect 497457 218648 509618 218650
rect 497457 218592 497462 218648
rect 497518 218592 509618 218648
rect 497457 218590 509618 218592
rect 518847 218650 518913 218653
rect 528553 218650 528619 218653
rect 518847 218648 528619 218650
rect 518847 218592 518852 218648
rect 518908 218592 528558 218648
rect 528614 218592 528619 218648
rect 518847 218590 528619 218592
rect 491220 218588 491267 218590
rect 491201 218587 491267 218588
rect 497457 218587 497523 218590
rect 518847 218587 518913 218590
rect 528553 218587 528619 218590
rect 528737 218650 528803 218653
rect 534073 218650 534139 218653
rect 528737 218648 534139 218650
rect 528737 218592 528742 218648
rect 528798 218592 534078 218648
rect 534134 218592 534139 218648
rect 528737 218590 534139 218592
rect 528737 218587 528803 218590
rect 534073 218587 534139 218590
rect 534257 218650 534323 218653
rect 606526 218650 606586 218862
rect 612733 218859 612799 218862
rect 640425 218922 640491 218925
rect 670601 218922 670667 218925
rect 640425 218920 670667 218922
rect 640425 218864 640430 218920
rect 640486 218864 670606 218920
rect 670662 218864 670667 218920
rect 640425 218862 670667 218864
rect 640425 218859 640491 218862
rect 670601 218859 670667 218862
rect 671245 218922 671311 218925
rect 674782 218922 674788 218924
rect 671245 218920 674788 218922
rect 671245 218864 671250 218920
rect 671306 218864 674788 218920
rect 671245 218862 674788 218864
rect 671245 218859 671311 218862
rect 674782 218860 674788 218862
rect 674852 218860 674858 218924
rect 534257 218648 606586 218650
rect 534257 218592 534262 218648
rect 534318 218592 606586 218648
rect 534257 218590 606586 218592
rect 606753 218650 606819 218653
rect 627729 218650 627795 218653
rect 606753 218648 627795 218650
rect 606753 218592 606758 218648
rect 606814 218592 627734 218648
rect 627790 218592 627795 218648
rect 606753 218590 627795 218592
rect 534257 218587 534323 218590
rect 606753 218587 606819 218590
rect 627729 218587 627795 218590
rect 645485 218650 645551 218653
rect 673126 218650 673132 218652
rect 645485 218648 673132 218650
rect 645485 218592 645490 218648
rect 645546 218592 673132 218648
rect 645485 218590 673132 218592
rect 645485 218587 645551 218590
rect 673126 218588 673132 218590
rect 673196 218588 673202 218652
rect 675518 218588 675524 218652
rect 675588 218650 675594 218652
rect 675588 218590 676292 218650
rect 675588 218588 675594 218590
rect 161565 218378 161631 218381
rect 162301 218378 162367 218381
rect 161565 218376 162367 218378
rect 161565 218320 161570 218376
rect 161626 218320 162306 218376
rect 162362 218320 162367 218376
rect 161565 218318 162367 218320
rect 161565 218315 161631 218318
rect 162301 218315 162367 218318
rect 500401 218378 500467 218381
rect 554037 218378 554103 218381
rect 500401 218376 554103 218378
rect 500401 218320 500406 218376
rect 500462 218320 554042 218376
rect 554098 218320 554103 218376
rect 500401 218318 554103 218320
rect 500401 218315 500467 218318
rect 554037 218315 554103 218318
rect 554221 218378 554287 218381
rect 572110 218378 572116 218380
rect 554221 218376 572116 218378
rect 554221 218320 554226 218376
rect 554282 218320 572116 218376
rect 554221 218318 572116 218320
rect 554221 218315 554287 218318
rect 572110 218316 572116 218318
rect 572180 218316 572186 218380
rect 572345 218378 572411 218381
rect 601417 218378 601483 218381
rect 572345 218376 601483 218378
rect 572345 218320 572350 218376
rect 572406 218320 601422 218376
rect 601478 218320 601483 218376
rect 572345 218318 601483 218320
rect 572345 218315 572411 218318
rect 601417 218315 601483 218318
rect 601601 218378 601667 218381
rect 623957 218378 624023 218381
rect 601601 218376 624023 218378
rect 601601 218320 601606 218376
rect 601662 218320 623962 218376
rect 624018 218320 624023 218376
rect 601601 218318 624023 218320
rect 601601 218315 601667 218318
rect 623957 218315 624023 218318
rect 670601 218378 670667 218381
rect 675845 218378 675911 218381
rect 670601 218376 675911 218378
rect 670601 218320 670606 218376
rect 670662 218320 675850 218376
rect 675906 218320 675911 218376
rect 670601 218318 675911 218320
rect 670601 218315 670667 218318
rect 675845 218315 675911 218318
rect 676024 218180 676030 218244
rect 676094 218242 676100 218244
rect 676094 218182 676292 218242
rect 676094 218180 676100 218182
rect 490649 218106 490715 218109
rect 572529 218106 572595 218109
rect 582097 218106 582163 218109
rect 490649 218104 572224 218106
rect 490649 218048 490654 218104
rect 490710 218048 572224 218104
rect 490649 218046 572224 218048
rect 490649 218043 490715 218046
rect 35525 217970 35591 217973
rect 53097 217970 53163 217973
rect 35525 217968 53163 217970
rect 35525 217912 35530 217968
rect 35586 217912 53102 217968
rect 53158 217912 53163 217968
rect 35525 217910 53163 217912
rect 35525 217907 35591 217910
rect 53097 217907 53163 217910
rect 572164 217837 572224 218046
rect 572529 218104 582163 218106
rect 572529 218048 572534 218104
rect 572590 218048 582102 218104
rect 582158 218048 582163 218104
rect 572529 218046 582163 218048
rect 572529 218043 572595 218046
rect 582097 218043 582163 218046
rect 582557 218106 582623 218109
rect 601417 218106 601483 218109
rect 606753 218106 606819 218109
rect 582557 218104 601483 218106
rect 582557 218048 582562 218104
rect 582618 218048 601422 218104
rect 601478 218048 601483 218104
rect 582557 218046 601483 218048
rect 582557 218043 582623 218046
rect 601417 218043 601483 218046
rect 601650 218104 606819 218106
rect 601650 218048 606758 218104
rect 606814 218048 606819 218104
rect 601650 218046 606819 218048
rect 502977 217834 503043 217837
rect 503621 217834 503687 217837
rect 508037 217834 508103 217837
rect 502977 217832 508103 217834
rect 502977 217776 502982 217832
rect 503038 217776 503626 217832
rect 503682 217776 508042 217832
rect 508098 217776 508103 217832
rect 502977 217774 508103 217776
rect 502977 217771 503043 217774
rect 503621 217771 503687 217774
rect 508037 217771 508103 217774
rect 508221 217834 508287 217837
rect 509325 217834 509391 217837
rect 508221 217832 509391 217834
rect 508221 217776 508226 217832
rect 508282 217776 509330 217832
rect 509386 217776 509391 217832
rect 508221 217774 509391 217776
rect 508221 217771 508287 217774
rect 509325 217771 509391 217774
rect 509509 217834 509575 217837
rect 528645 217834 528711 217837
rect 509509 217832 528711 217834
rect 509509 217776 509514 217832
rect 509570 217776 528650 217832
rect 528706 217776 528711 217832
rect 509509 217774 528711 217776
rect 509509 217771 509575 217774
rect 528645 217771 528711 217774
rect 529105 217834 529171 217837
rect 571885 217834 571951 217837
rect 529105 217832 571951 217834
rect 529105 217776 529110 217832
rect 529166 217776 571890 217832
rect 571946 217776 571951 217832
rect 529105 217774 571951 217776
rect 529105 217771 529171 217774
rect 571885 217771 571951 217774
rect 572161 217832 572227 217837
rect 572161 217776 572166 217832
rect 572222 217776 572227 217832
rect 572161 217771 572227 217776
rect 572897 217834 572963 217837
rect 582557 217834 582623 217837
rect 572897 217832 582623 217834
rect 572897 217776 572902 217832
rect 572958 217776 582562 217832
rect 582618 217776 582623 217832
rect 572897 217774 582623 217776
rect 572897 217771 572963 217774
rect 582557 217771 582623 217774
rect 582741 217834 582807 217837
rect 601650 217834 601710 218046
rect 606753 218043 606819 218046
rect 582741 217832 601710 217834
rect 582741 217776 582746 217832
rect 582802 217776 601710 217832
rect 582741 217774 601710 217776
rect 649901 217834 649967 217837
rect 672022 217834 672028 217836
rect 649901 217832 672028 217834
rect 649901 217776 649906 217832
rect 649962 217776 672028 217832
rect 649901 217774 672028 217776
rect 582741 217771 582807 217774
rect 649901 217771 649967 217774
rect 672022 217772 672028 217774
rect 672092 217772 672098 217836
rect 674833 217834 674899 217837
rect 674833 217832 676292 217834
rect 674833 217776 674838 217832
rect 674894 217776 676292 217832
rect 674833 217774 676292 217776
rect 674833 217771 674899 217774
rect 494697 217698 494763 217701
rect 495157 217698 495223 217701
rect 494697 217696 495223 217698
rect 494697 217640 494702 217696
rect 494758 217640 495162 217696
rect 495218 217640 495223 217696
rect 494697 217638 495223 217640
rect 494697 217635 494763 217638
rect 495157 217635 495223 217638
rect 501321 217562 501387 217565
rect 501689 217562 501755 217565
rect 501321 217560 501755 217562
rect 501321 217504 501326 217560
rect 501382 217504 501694 217560
rect 501750 217504 501755 217560
rect 501321 217502 501755 217504
rect 501321 217499 501387 217502
rect 501689 217499 501755 217502
rect 505093 217562 505159 217565
rect 591941 217562 592007 217565
rect 505093 217560 592007 217562
rect 505093 217504 505098 217560
rect 505154 217504 591946 217560
rect 592002 217504 592007 217560
rect 505093 217502 592007 217504
rect 505093 217499 505159 217502
rect 591941 217499 592007 217502
rect 592350 217500 592356 217564
rect 592420 217562 592426 217564
rect 596357 217562 596423 217565
rect 592420 217560 596423 217562
rect 592420 217504 596362 217560
rect 596418 217504 596423 217560
rect 592420 217502 596423 217504
rect 592420 217500 592426 217502
rect 596357 217499 596423 217502
rect 601647 217562 601713 217565
rect 603257 217562 603323 217565
rect 601647 217560 603323 217562
rect 601647 217504 601652 217560
rect 601708 217504 603262 217560
rect 603318 217504 603323 217560
rect 601647 217502 603323 217504
rect 601647 217499 601713 217502
rect 603257 217499 603323 217502
rect 646865 217562 646931 217565
rect 675661 217562 675727 217565
rect 646865 217560 675727 217562
rect 646865 217504 646870 217560
rect 646926 217504 675666 217560
rect 675722 217504 675727 217560
rect 646865 217502 675727 217504
rect 646865 217499 646931 217502
rect 675661 217499 675727 217502
rect 675894 217366 676292 217426
rect 488901 217292 488967 217293
rect 488901 217290 488948 217292
rect 488856 217288 488948 217290
rect 488856 217232 488906 217288
rect 488856 217230 488948 217232
rect 488901 217228 488948 217230
rect 489012 217228 489018 217292
rect 498837 217290 498903 217293
rect 518985 217290 519051 217293
rect 498837 217288 519051 217290
rect 498837 217232 498842 217288
rect 498898 217232 518990 217288
rect 519046 217232 519051 217288
rect 498837 217230 519051 217232
rect 488901 217227 488967 217228
rect 498837 217227 498903 217230
rect 518985 217227 519051 217230
rect 519169 217290 519235 217293
rect 528277 217290 528343 217293
rect 519169 217288 528343 217290
rect 519169 217232 519174 217288
rect 519230 217232 528282 217288
rect 528338 217232 528343 217288
rect 519169 217230 528343 217232
rect 519169 217227 519235 217230
rect 528277 217227 528343 217230
rect 528461 217290 528527 217293
rect 534073 217290 534139 217293
rect 528461 217288 534139 217290
rect 528461 217232 528466 217288
rect 528522 217232 534078 217288
rect 534134 217232 534139 217288
rect 528461 217230 534139 217232
rect 528461 217227 528527 217230
rect 534073 217227 534139 217230
rect 534257 217290 534323 217293
rect 543457 217290 543523 217293
rect 534257 217288 543523 217290
rect 534257 217232 534262 217288
rect 534318 217232 543462 217288
rect 543518 217232 543523 217288
rect 534257 217230 543523 217232
rect 534257 217227 534323 217230
rect 543457 217227 543523 217230
rect 543641 217290 543707 217293
rect 591982 217290 591988 217292
rect 543641 217288 591988 217290
rect 543641 217232 543646 217288
rect 543702 217232 591988 217288
rect 543641 217230 591988 217232
rect 543641 217227 543707 217230
rect 591982 217228 591988 217230
rect 592052 217228 592058 217292
rect 596817 217290 596883 217293
rect 592174 217288 596883 217290
rect 592174 217232 596822 217288
rect 596878 217232 596883 217288
rect 592174 217230 596883 217232
rect 501321 217018 501387 217021
rect 592174 217018 592234 217230
rect 596817 217227 596883 217230
rect 666829 217290 666895 217293
rect 675894 217290 675954 217366
rect 666829 217288 675954 217290
rect 666829 217232 666834 217288
rect 666890 217232 675954 217288
rect 666829 217230 675954 217232
rect 666829 217227 666895 217230
rect 601509 217154 601575 217157
rect 601785 217154 601851 217157
rect 601509 217152 601851 217154
rect 601509 217096 601514 217152
rect 601570 217096 601790 217152
rect 601846 217096 601851 217152
rect 601509 217094 601851 217096
rect 601509 217091 601575 217094
rect 601785 217091 601851 217094
rect 501321 217016 592234 217018
rect 501321 216960 501326 217016
rect 501382 216960 592234 217016
rect 501321 216958 592234 216960
rect 597461 217018 597527 217021
rect 600957 217018 601023 217021
rect 597461 217016 601023 217018
rect 597461 216960 597466 217016
rect 597522 216960 600962 217016
rect 601018 216960 601023 217016
rect 597461 216958 601023 216960
rect 501321 216955 501387 216958
rect 597461 216955 597527 216958
rect 600957 216955 601023 216958
rect 675886 216956 675892 217020
rect 675956 217018 675962 217020
rect 675956 216958 676292 217018
rect 675956 216956 675962 216958
rect 601325 216882 601391 216885
rect 601785 216882 601851 216885
rect 675385 216882 675451 216885
rect 601325 216880 601851 216882
rect 601325 216824 601330 216880
rect 601386 216824 601790 216880
rect 601846 216824 601851 216880
rect 601325 216822 601851 216824
rect 601325 216819 601391 216822
rect 601785 216819 601851 216822
rect 675158 216880 675451 216882
rect 675158 216824 675390 216880
rect 675446 216824 675451 216880
rect 675158 216822 675451 216824
rect 495157 216746 495223 216749
rect 590101 216746 590167 216749
rect 495157 216744 590167 216746
rect 495157 216688 495162 216744
rect 495218 216688 590106 216744
rect 590162 216688 590167 216744
rect 495157 216686 590167 216688
rect 495157 216683 495223 216686
rect 590101 216683 590167 216686
rect 540145 216474 540211 216477
rect 557073 216474 557139 216477
rect 540145 216472 557139 216474
rect 540145 216416 540150 216472
rect 540206 216416 557078 216472
rect 557134 216416 557139 216472
rect 540145 216414 557139 216416
rect 540145 216411 540211 216414
rect 557073 216411 557139 216414
rect 557717 216474 557783 216477
rect 558545 216474 558611 216477
rect 602521 216474 602587 216477
rect 557717 216472 557826 216474
rect 557717 216416 557722 216472
rect 557778 216416 557826 216472
rect 557717 216411 557826 216416
rect 558545 216472 602587 216474
rect 558545 216416 558550 216472
rect 558606 216416 602526 216472
rect 602582 216416 602587 216472
rect 558545 216414 602587 216416
rect 558545 216411 558611 216414
rect 602521 216411 602587 216414
rect 646589 216474 646655 216477
rect 675158 216474 675218 216822
rect 675385 216819 675451 216822
rect 675385 216610 675451 216613
rect 675385 216608 676292 216610
rect 675385 216552 675390 216608
rect 675446 216552 676292 216608
rect 675385 216550 676292 216552
rect 675385 216547 675451 216550
rect 646589 216472 675218 216474
rect 646589 216416 646594 216472
rect 646650 216416 675218 216472
rect 646589 216414 675218 216416
rect 646589 216411 646655 216414
rect 557766 216202 557826 216411
rect 626625 216202 626691 216205
rect 557766 216200 626691 216202
rect 557766 216144 626630 216200
rect 626686 216144 626691 216200
rect 557766 216142 626691 216144
rect 626625 216139 626691 216142
rect 651097 216202 651163 216205
rect 672165 216202 672231 216205
rect 651097 216200 672231 216202
rect 651097 216144 651102 216200
rect 651158 216144 672170 216200
rect 672226 216144 672231 216200
rect 651097 216142 672231 216144
rect 651097 216139 651163 216142
rect 672165 216139 672231 216142
rect 674557 216202 674623 216205
rect 674557 216200 676292 216202
rect 674557 216144 674562 216200
rect 674618 216144 676292 216200
rect 674557 216142 676292 216144
rect 674557 216139 674623 216142
rect 643001 215930 643067 215933
rect 643001 215928 659670 215930
rect 643001 215872 643006 215928
rect 643062 215872 659670 215928
rect 643001 215870 659670 215872
rect 643001 215867 643067 215870
rect 659610 215522 659670 215870
rect 670601 215794 670667 215797
rect 670601 215792 676292 215794
rect 670601 215736 670606 215792
rect 670662 215736 676292 215792
rect 670601 215734 676292 215736
rect 670601 215731 670667 215734
rect 675150 215522 675156 215524
rect 659610 215462 675156 215522
rect 675150 215460 675156 215462
rect 675220 215460 675226 215524
rect 675702 215324 675708 215388
rect 675772 215386 675778 215388
rect 675772 215326 676292 215386
rect 675772 215324 675778 215326
rect 664897 215114 664963 215117
rect 676029 215114 676095 215117
rect 664897 215112 676095 215114
rect 664897 215056 664902 215112
rect 664958 215056 676034 215112
rect 676090 215056 676095 215112
rect 676254 215086 676260 215150
rect 676324 215086 676330 215150
rect 664897 215054 676095 215056
rect 664897 215051 664963 215054
rect 676029 215051 676095 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 676262 214948 676322 215086
rect 41492 214918 44883 214920
rect 44817 214915 44883 214918
rect 648521 214570 648587 214573
rect 675201 214570 675267 214573
rect 648521 214568 675267 214570
rect 35758 214301 35818 214540
rect 648521 214512 648526 214568
rect 648582 214512 675206 214568
rect 675262 214512 675267 214568
rect 648521 214510 675267 214512
rect 648521 214507 648587 214510
rect 675201 214507 675267 214510
rect 675661 214570 675727 214573
rect 675661 214568 676292 214570
rect 675661 214512 675666 214568
rect 675722 214512 676292 214568
rect 675661 214510 676292 214512
rect 675661 214507 675727 214510
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 35574 214132 35634 214235
rect 575982 214026 576042 214404
rect 672073 214162 672139 214165
rect 672073 214160 676292 214162
rect 672073 214104 672078 214160
rect 672134 214104 676292 214160
rect 672073 214102 676292 214104
rect 672073 214099 672139 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 42793 213754 42859 213757
rect 41492 213752 42859 213754
rect 41492 213696 42798 213752
rect 42854 213696 42859 213752
rect 41492 213694 42859 213696
rect 42793 213691 42859 213694
rect 664713 213754 664779 213757
rect 673085 213754 673151 213757
rect 664713 213752 672826 213754
rect 664713 213696 664718 213752
rect 664774 213696 672826 213752
rect 664713 213694 672826 213696
rect 664713 213691 664779 213694
rect 661493 213482 661559 213485
rect 672766 213482 672826 213694
rect 673085 213752 676292 213754
rect 673085 213696 673090 213752
rect 673146 213696 676292 213752
rect 673085 213694 676292 213696
rect 673085 213691 673151 213694
rect 676029 213482 676095 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 672766 213480 676095 213482
rect 672766 213424 676034 213480
rect 676090 213424 676095 213480
rect 672766 213422 676095 213424
rect 661493 213419 661559 213422
rect 43437 213346 43503 213349
rect 41492 213344 43503 213346
rect 41492 213288 43442 213344
rect 43498 213288 43503 213344
rect 41492 213286 43503 213288
rect 43437 213283 43503 213286
rect 575606 213148 575612 213212
rect 575676 213210 575682 213212
rect 594793 213210 594859 213213
rect 575676 213208 594859 213210
rect 575676 213152 594798 213208
rect 594854 213152 594859 213208
rect 575676 213150 594859 213152
rect 575676 213148 575682 213150
rect 594793 213147 594859 213150
rect 647141 213210 647207 213213
rect 669270 213210 669330 213422
rect 676029 213419 676095 213422
rect 683297 213346 683363 213349
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 683297 213283 683363 213286
rect 676029 213210 676095 213213
rect 647141 213208 663810 213210
rect 647141 213152 647146 213208
rect 647202 213152 663810 213208
rect 647141 213150 663810 213152
rect 669270 213208 676095 213210
rect 669270 213152 676034 213208
rect 676090 213152 676095 213208
rect 669270 213150 676095 213152
rect 647141 213147 647207 213150
rect 43621 212938 43687 212941
rect 41492 212936 43687 212938
rect 41492 212880 43626 212936
rect 43682 212880 43687 212936
rect 41492 212878 43687 212880
rect 663750 212938 663810 213150
rect 676029 213147 676095 213150
rect 674097 212938 674163 212941
rect 663750 212936 674163 212938
rect 663750 212880 674102 212936
rect 674158 212880 674163 212936
rect 663750 212878 674163 212880
rect 43621 212875 43687 212878
rect 674097 212875 674163 212878
rect 683070 212533 683130 212908
rect 47945 212530 48011 212533
rect 41492 212528 48011 212530
rect 41492 212472 47950 212528
rect 48006 212472 48011 212528
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 41492 212470 48011 212472
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 47945 212467 48011 212470
rect 683113 212467 683179 212470
rect 667974 212332 667980 212396
rect 668044 212394 668050 212396
rect 669221 212394 669287 212397
rect 668044 212392 669287 212394
rect 668044 212336 669226 212392
rect 669282 212336 669287 212392
rect 668044 212334 669287 212336
rect 668044 212332 668050 212334
rect 669221 212331 669287 212334
rect 42977 212122 43043 212125
rect 41492 212120 43043 212122
rect 41492 212064 42982 212120
rect 43038 212064 43043 212120
rect 41492 212062 43043 212064
rect 42977 212059 43043 212062
rect 575982 211714 576042 212228
rect 674097 212122 674163 212125
rect 674097 212120 676292 212122
rect 674097 212064 674102 212120
rect 674158 212064 676292 212120
rect 674097 212062 676292 212064
rect 674097 212059 674163 212062
rect 669221 211986 669287 211989
rect 672717 211986 672783 211989
rect 669221 211984 672783 211986
rect 669221 211928 669226 211984
rect 669282 211928 672722 211984
rect 672778 211928 672783 211984
rect 669221 211926 672783 211928
rect 669221 211923 669287 211926
rect 672717 211923 672783 211926
rect 669037 211850 669103 211853
rect 669037 211848 669146 211850
rect 669037 211792 669042 211848
rect 669098 211792 669146 211848
rect 669037 211787 669146 211792
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 35758 211445 35818 211684
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 669086 211578 669146 211787
rect 668902 211518 669146 211578
rect 35758 211440 35867 211445
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211382 35867 211384
rect 35801 211379 35867 211382
rect 668902 211309 668962 211518
rect 675661 211442 675727 211445
rect 676438 211442 676444 211444
rect 675661 211440 676444 211442
rect 675661 211384 675666 211440
rect 675722 211384 676444 211440
rect 675661 211382 676444 211384
rect 675661 211379 675727 211382
rect 676438 211380 676444 211382
rect 676508 211380 676514 211444
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 668902 211304 669011 211309
rect 668902 211248 668950 211304
rect 669006 211248 669011 211304
rect 668902 211246 669011 211248
rect 44173 211243 44239 211246
rect 668945 211243 669011 211246
rect 672717 211170 672783 211173
rect 683113 211170 683179 211173
rect 672717 211168 683179 211170
rect 672717 211112 672722 211168
rect 672778 211112 683118 211168
rect 683174 211112 683179 211168
rect 672717 211110 683179 211112
rect 672717 211107 672783 211110
rect 683113 211107 683179 211110
rect 45001 210898 45067 210901
rect 41492 210896 45067 210898
rect 41492 210840 45006 210896
rect 45062 210840 45067 210896
rect 41492 210838 45067 210840
rect 45001 210835 45067 210838
rect 44173 210490 44239 210493
rect 41492 210488 44239 210490
rect 41492 210432 44178 210488
rect 44234 210432 44239 210488
rect 41492 210430 44239 210432
rect 44173 210427 44239 210430
rect 672441 210490 672507 210493
rect 673126 210490 673132 210492
rect 672441 210488 673132 210490
rect 672441 210432 672446 210488
rect 672502 210432 673132 210488
rect 672441 210430 673132 210432
rect 672441 210427 672507 210430
rect 673126 210428 673132 210430
rect 673196 210428 673202 210492
rect 675518 210428 675524 210492
rect 675588 210490 675594 210492
rect 675886 210490 675892 210492
rect 675588 210430 675892 210490
rect 675588 210428 675594 210430
rect 675886 210428 675892 210430
rect 675956 210428 675962 210492
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 672717 210218 672783 210221
rect 678930 210218 678990 210294
rect 683297 210291 683363 210294
rect 672717 210216 678990 210218
rect 672717 210160 672722 210216
rect 672778 210160 678990 210216
rect 672717 210158 678990 210160
rect 672717 210155 672783 210158
rect 42006 210082 42012 210084
rect 41492 210022 42012 210082
rect 42006 210020 42012 210022
rect 42076 210020 42082 210084
rect 575982 209810 576042 210052
rect 579245 209810 579311 209813
rect 575982 209808 579311 209810
rect 575982 209752 579250 209808
rect 579306 209752 579311 209808
rect 575982 209750 579311 209752
rect 579245 209747 579311 209750
rect 42793 209674 42859 209677
rect 41492 209672 42859 209674
rect 41492 209616 42798 209672
rect 42854 209616 42859 209672
rect 41492 209614 42859 209616
rect 42793 209611 42859 209614
rect 673913 209674 673979 209677
rect 676673 209674 676739 209677
rect 673913 209672 676739 209674
rect 673913 209616 673918 209672
rect 673974 209616 676678 209672
rect 676734 209616 676739 209672
rect 673913 209614 676739 209616
rect 673913 209611 673979 209614
rect 676673 209611 676739 209614
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 41689 208994 41755 208997
rect 49509 208994 49575 208997
rect 41689 208992 49575 208994
rect 41689 208936 41694 208992
rect 41750 208936 49514 208992
rect 49570 208936 49575 208992
rect 41689 208934 49575 208936
rect 41689 208931 41755 208934
rect 49509 208931 49575 208934
rect 41462 208586 41522 208828
rect 44357 208586 44423 208589
rect 41462 208584 44423 208586
rect 41462 208528 44362 208584
rect 44418 208528 44423 208584
rect 41462 208526 44423 208528
rect 44357 208523 44423 208526
rect 40726 208180 40786 208420
rect 40718 208116 40724 208180
rect 40788 208116 40794 208180
rect 43253 208042 43319 208045
rect 41492 208040 43319 208042
rect 41492 207984 43258 208040
rect 43314 207984 43319 208040
rect 41492 207982 43319 207984
rect 43253 207979 43319 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40033 207770 40099 207773
rect 41638 207770 41644 207772
rect 40033 207768 41644 207770
rect 40033 207712 40038 207768
rect 40094 207712 41644 207768
rect 40033 207710 41644 207712
rect 40033 207707 40099 207710
rect 41638 207708 41644 207710
rect 41708 207708 41714 207772
rect 40910 207364 40970 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40902 207300 40908 207364
rect 40972 207300 40978 207364
rect 675845 207226 675911 207229
rect 669270 207224 675911 207226
rect 40542 206956 40602 207196
rect 666326 207090 666386 207196
rect 669270 207168 675850 207224
rect 675906 207168 675911 207224
rect 669270 207166 675911 207168
rect 669270 207090 669330 207166
rect 675845 207163 675911 207166
rect 666326 207030 669330 207090
rect 40534 206892 40540 206956
rect 40604 206892 40610 206956
rect 673729 206954 673795 206957
rect 677777 206954 677843 206957
rect 673729 206952 677843 206954
rect 673729 206896 673734 206952
rect 673790 206896 677782 206952
rect 677838 206896 677843 206952
rect 673729 206894 677843 206896
rect 673729 206891 673795 206894
rect 677777 206891 677843 206894
rect 43621 206818 43687 206821
rect 41492 206816 43687 206818
rect 41492 206760 43626 206816
rect 43682 206760 43687 206816
rect 41492 206758 43687 206760
rect 43621 206755 43687 206758
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 43437 206274 43503 206277
rect 49325 206274 49391 206277
rect 43437 206272 49391 206274
rect 43437 206216 43442 206272
rect 43498 206216 49330 206272
rect 49386 206216 49391 206272
rect 43437 206214 49391 206216
rect 43437 206211 43503 206214
rect 49325 206211 49391 206214
rect 44541 206002 44607 206005
rect 41492 206000 44607 206002
rect 41492 205944 44546 206000
rect 44602 205944 44607 206000
rect 41492 205942 44607 205944
rect 44541 205939 44607 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 43805 205594 43871 205597
rect 41492 205592 43871 205594
rect 41492 205536 43810 205592
rect 43866 205536 43871 205592
rect 41492 205534 43871 205536
rect 43805 205531 43871 205534
rect 675753 205594 675819 205597
rect 676622 205594 676628 205596
rect 675753 205592 676628 205594
rect 675753 205536 675758 205592
rect 675814 205536 676628 205592
rect 675753 205534 676628 205536
rect 675753 205531 675819 205534
rect 676622 205532 676628 205534
rect 676692 205532 676698 205596
rect 43989 205186 44055 205189
rect 41492 205184 44055 205186
rect 41492 205128 43994 205184
rect 44050 205128 44055 205184
rect 41492 205126 44055 205128
rect 43989 205123 44055 205126
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 35574 204101 35634 204340
rect 35574 204096 35683 204101
rect 35574 204040 35622 204096
rect 35678 204040 35683 204096
rect 35574 204038 35683 204040
rect 35617 204035 35683 204038
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 41462 203282 41522 203524
rect 50705 203282 50771 203285
rect 41462 203280 50771 203282
rect 41462 203224 50710 203280
rect 50766 203224 50771 203280
rect 41462 203222 50771 203224
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 666326 203282 666386 203932
rect 673913 203282 673979 203285
rect 666326 203280 673979 203282
rect 666326 203224 673918 203280
rect 673974 203224 673979 203280
rect 666326 203222 673979 203224
rect 50705 203219 50771 203222
rect 578325 203219 578391 203222
rect 673913 203219 673979 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 672257 203010 672323 203013
rect 673310 203010 673316 203012
rect 672257 203008 673316 203010
rect 672257 202952 672262 203008
rect 672318 202952 673316 203008
rect 672257 202950 673316 202952
rect 672257 202947 672323 202950
rect 673310 202948 673316 202950
rect 673380 202948 673386 203012
rect 35617 202194 35683 202197
rect 43437 202194 43503 202197
rect 35617 202192 43503 202194
rect 35617 202136 35622 202192
rect 35678 202136 43442 202192
rect 43498 202136 43503 202192
rect 35617 202134 43503 202136
rect 35617 202131 35683 202134
rect 43437 202131 43503 202134
rect 666326 201650 666386 202300
rect 674465 201922 674531 201925
rect 675385 201922 675451 201925
rect 674465 201920 675451 201922
rect 674465 201864 674470 201920
rect 674526 201864 675390 201920
rect 675446 201864 675451 201920
rect 674465 201862 675451 201864
rect 674465 201859 674531 201862
rect 675385 201859 675451 201862
rect 673729 201650 673795 201653
rect 666326 201648 673795 201650
rect 666326 201592 673734 201648
rect 673790 201592 673795 201648
rect 666326 201590 673795 201592
rect 673729 201587 673795 201590
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 670601 201378 670667 201381
rect 675385 201378 675451 201381
rect 670601 201376 675451 201378
rect 575982 200834 576042 201348
rect 670601 201320 670606 201376
rect 670662 201320 675390 201376
rect 675446 201320 675451 201376
rect 670601 201318 675451 201320
rect 670601 201315 670667 201318
rect 675385 201315 675451 201318
rect 672073 201106 672139 201109
rect 674833 201106 674899 201109
rect 672073 201104 674899 201106
rect 672073 201048 672078 201104
rect 672134 201048 674838 201104
rect 674894 201048 674899 201104
rect 672073 201046 674899 201048
rect 672073 201043 672139 201046
rect 674833 201043 674899 201046
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 675753 200834 675819 200837
rect 676438 200834 676444 200836
rect 675753 200832 676444 200834
rect 675753 200776 675758 200832
rect 675814 200776 676444 200832
rect 675753 200774 676444 200776
rect 675753 200771 675819 200774
rect 676438 200772 676444 200774
rect 676508 200772 676514 200836
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 575982 198930 576042 199172
rect 670785 199066 670851 199069
rect 666356 199064 670851 199066
rect 666356 199008 670790 199064
rect 670846 199008 670851 199064
rect 666356 199006 670851 199008
rect 670785 199003 670851 199006
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 666829 198386 666895 198389
rect 675385 198386 675451 198389
rect 666829 198384 675451 198386
rect 666829 198328 666834 198384
rect 666890 198328 675390 198384
rect 675446 198328 675451 198384
rect 666829 198326 675451 198328
rect 666829 198323 666895 198326
rect 675385 198323 675451 198326
rect 590377 198250 590443 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 590377 198187 590443 198190
rect 37917 197842 37983 197845
rect 41822 197842 41828 197844
rect 37917 197840 41828 197842
rect 37917 197784 37922 197840
rect 37978 197784 41828 197840
rect 37917 197782 41828 197784
rect 37917 197779 37983 197782
rect 41822 197780 41828 197782
rect 41892 197780 41898 197844
rect 674833 197570 674899 197573
rect 675477 197570 675543 197573
rect 674833 197568 675543 197570
rect 674833 197512 674838 197568
rect 674894 197512 675482 197568
rect 675538 197512 675543 197568
rect 674833 197510 675543 197512
rect 674833 197507 674899 197510
rect 675477 197507 675543 197510
rect 668025 197434 668091 197437
rect 666356 197432 668091 197434
rect 666356 197376 668030 197432
rect 668086 197376 668091 197432
rect 666356 197374 668091 197376
rect 668025 197371 668091 197374
rect 40718 197100 40724 197164
rect 40788 197162 40794 197164
rect 41781 197162 41847 197165
rect 40788 197160 41847 197162
rect 40788 197104 41786 197160
rect 41842 197104 41847 197160
rect 40788 197102 41847 197104
rect 40788 197100 40794 197102
rect 41781 197099 41847 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49509 196482 49575 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49509 196480 52164 196482
rect 49509 196424 49514 196480
rect 49570 196424 52164 196480
rect 49509 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49509 196419 49575 196422
rect 578509 196419 578575 196422
rect 673085 196482 673151 196485
rect 675385 196482 675451 196485
rect 673085 196480 675451 196482
rect 673085 196424 673090 196480
rect 673146 196424 675390 196480
rect 675446 196424 675451 196480
rect 673085 196422 675451 196424
rect 673085 196419 673151 196422
rect 675385 196419 675451 196422
rect 41873 195804 41939 195805
rect 41822 195802 41828 195804
rect 41782 195742 41828 195802
rect 41892 195800 41939 195804
rect 41934 195744 41939 195800
rect 41822 195740 41828 195742
rect 41892 195740 41939 195744
rect 41873 195739 41939 195740
rect 40902 195468 40908 195532
rect 40972 195530 40978 195532
rect 42609 195530 42675 195533
rect 40972 195528 42675 195530
rect 40972 195472 42614 195528
rect 42670 195472 42675 195528
rect 40972 195470 42675 195472
rect 40972 195468 40978 195470
rect 42609 195467 42675 195470
rect 41965 195260 42031 195261
rect 675661 195260 675727 195261
rect 41965 195256 42012 195260
rect 42076 195258 42082 195260
rect 41965 195200 41970 195256
rect 41965 195196 42012 195200
rect 42076 195198 42122 195258
rect 675661 195256 675708 195260
rect 675772 195258 675778 195260
rect 675661 195200 675666 195256
rect 42076 195196 42082 195198
rect 675661 195196 675708 195200
rect 675772 195198 675818 195258
rect 675772 195196 675778 195198
rect 41965 195195 42031 195196
rect 675661 195195 675727 195196
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 40534 194516 40540 194580
rect 40604 194578 40610 194580
rect 41454 194578 41460 194580
rect 40604 194518 41460 194578
rect 40604 194516 40610 194518
rect 41454 194516 41460 194518
rect 41524 194516 41530 194580
rect 48589 194442 48655 194445
rect 48589 194440 52164 194442
rect 48589 194384 48594 194440
rect 48650 194384 52164 194440
rect 48589 194382 52164 194384
rect 48589 194379 48655 194382
rect 668117 194170 668183 194173
rect 666356 194168 668183 194170
rect 666356 194112 668122 194168
rect 668178 194112 668183 194168
rect 666356 194110 668183 194112
rect 668117 194107 668183 194110
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42425 193218 42491 193221
rect 43621 193218 43687 193221
rect 42425 193216 43687 193218
rect 42425 193160 42430 193216
rect 42486 193160 43626 193216
rect 43682 193160 43687 193216
rect 42425 193158 43687 193160
rect 42425 193155 42491 193158
rect 43621 193155 43687 193158
rect 675661 193218 675727 193221
rect 675886 193218 675892 193220
rect 675661 193216 675892 193218
rect 675661 193160 675666 193216
rect 675722 193160 675892 193216
rect 675661 193158 675892 193160
rect 675661 193155 675727 193158
rect 675886 193156 675892 193158
rect 675956 193156 675962 193220
rect 42374 192884 42380 192948
rect 42444 192946 42450 192948
rect 42609 192946 42675 192949
rect 42444 192944 42675 192946
rect 42444 192888 42614 192944
rect 42670 192888 42675 192944
rect 42444 192886 42675 192888
rect 42444 192884 42450 192886
rect 42609 192883 42675 192886
rect 47945 192402 48011 192405
rect 47945 192400 52164 192402
rect 47945 192344 47950 192400
rect 48006 192344 52164 192400
rect 47945 192342 52164 192344
rect 47945 192339 48011 192342
rect 575982 192266 576042 192644
rect 668025 192538 668091 192541
rect 666356 192536 668091 192538
rect 666356 192480 668030 192536
rect 668086 192480 668091 192536
rect 666356 192478 668091 192480
rect 668025 192475 668091 192478
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 668117 192266 668183 192269
rect 673269 192266 673335 192269
rect 668117 192264 673335 192266
rect 668117 192208 668122 192264
rect 668178 192208 673274 192264
rect 673330 192208 673335 192264
rect 668117 192206 673335 192208
rect 668117 192203 668183 192206
rect 673269 192203 673335 192206
rect 42333 191722 42399 191725
rect 43989 191722 44055 191725
rect 42333 191720 44055 191722
rect 42333 191664 42338 191720
rect 42394 191664 43994 191720
rect 44050 191664 44055 191720
rect 42333 191662 44055 191664
rect 42333 191659 42399 191662
rect 43989 191659 44055 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43805 190498 43871 190501
rect 42425 190496 43871 190498
rect 42425 190440 42430 190496
rect 42486 190440 43810 190496
rect 43866 190440 43871 190496
rect 42425 190438 43871 190440
rect 42425 190435 42491 190438
rect 43805 190435 43871 190438
rect 49325 190498 49391 190501
rect 49325 190496 52164 190498
rect 49325 190440 49330 190496
rect 49386 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 49325 190438 52164 190440
rect 49325 190435 49391 190438
rect 669221 190362 669287 190365
rect 675293 190362 675359 190365
rect 669221 190360 675359 190362
rect 669221 190304 669226 190360
rect 669282 190304 675298 190360
rect 675354 190304 675359 190360
rect 669221 190302 675359 190304
rect 669221 190299 669287 190302
rect 675293 190299 675359 190302
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 44357 189954 44423 189957
rect 42425 189952 44423 189954
rect 42425 189896 42430 189952
rect 42486 189896 44362 189952
rect 44418 189896 44423 189952
rect 42425 189894 44423 189896
rect 42425 189891 42491 189894
rect 44357 189891 44423 189894
rect 669129 189274 669195 189277
rect 666356 189272 669195 189274
rect 666356 189216 669134 189272
rect 669190 189216 669195 189272
rect 666356 189214 669195 189216
rect 669129 189211 669195 189214
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 44541 187642 44607 187645
rect 668117 187642 668183 187645
rect 42425 187640 44607 187642
rect 42425 187584 42430 187640
rect 42486 187584 44546 187640
rect 44602 187584 44607 187640
rect 42425 187582 44607 187584
rect 666356 187640 668183 187642
rect 666356 187584 668122 187640
rect 668178 187584 668183 187640
rect 666356 187582 668183 187584
rect 42425 187579 42491 187582
rect 44541 187579 44607 187582
rect 668117 187579 668183 187582
rect 41454 187172 41460 187236
rect 41524 187234 41530 187236
rect 41781 187234 41847 187237
rect 41524 187232 41847 187234
rect 41524 187176 41786 187232
rect 41842 187176 41847 187232
rect 41524 187174 41847 187176
rect 41524 187172 41530 187174
rect 41781 187171 41847 187174
rect 666461 186962 666527 186965
rect 683113 186962 683179 186965
rect 666461 186960 683179 186962
rect 666461 186904 666466 186960
rect 666522 186904 683118 186960
rect 683174 186904 683179 186960
rect 666461 186902 683179 186904
rect 666461 186899 666527 186902
rect 683113 186899 683179 186902
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 42333 186284 42399 186285
rect 42333 186282 42380 186284
rect 42288 186280 42380 186282
rect 42288 186224 42338 186280
rect 42288 186222 42380 186224
rect 42333 186220 42380 186222
rect 42444 186220 42450 186284
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 42333 186219 42399 186220
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41781 185876 41847 185877
rect 41781 185872 41828 185876
rect 41892 185874 41898 185876
rect 41781 185816 41786 185872
rect 41781 185812 41828 185816
rect 41892 185814 41938 185874
rect 41892 185812 41898 185814
rect 41781 185811 41847 185812
rect 669129 185602 669195 185605
rect 672533 185602 672599 185605
rect 669129 185600 672599 185602
rect 669129 185544 669134 185600
rect 669190 185544 672538 185600
rect 672594 185544 672599 185600
rect 669129 185542 672599 185544
rect 669129 185539 669195 185542
rect 672533 185539 672599 185542
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 42425 184922 42491 184925
rect 44173 184922 44239 184925
rect 42425 184920 44239 184922
rect 42425 184864 42430 184920
rect 42486 184864 44178 184920
rect 44234 184864 44239 184920
rect 42425 184862 44239 184864
rect 42425 184859 42491 184862
rect 44173 184859 44239 184862
rect 579521 184378 579587 184381
rect 668025 184378 668091 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 666356 184376 668091 184378
rect 666356 184320 668030 184376
rect 668086 184320 668091 184376
rect 666356 184318 668091 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 668025 184315 668091 184318
rect 589457 183562 589523 183565
rect 672257 183562 672323 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672257 183560 672948 183562
rect 672257 183504 672262 183560
rect 672318 183504 672948 183560
rect 672257 183502 672948 183504
rect 589457 183499 589523 183502
rect 672257 183499 672323 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 43253 183154 43319 183157
rect 42425 183152 43319 183154
rect 42425 183096 42430 183152
rect 42486 183096 43258 183152
rect 43314 183096 43319 183152
rect 42425 183094 43319 183096
rect 42425 183091 42491 183094
rect 43253 183091 43319 183094
rect 668301 182746 668367 182749
rect 666356 182744 668367 182746
rect 666356 182688 668306 182744
rect 668362 182688 668367 182744
rect 666356 182686 668367 182688
rect 668301 182683 668367 182686
rect 672073 182066 672139 182069
rect 673126 182066 673132 182068
rect 672073 182064 673132 182066
rect 672073 182008 672078 182064
rect 672134 182008 673132 182064
rect 672073 182006 673132 182008
rect 672073 182003 672139 182006
rect 673126 182004 673132 182006
rect 673196 182004 673202 182068
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667381 181386 667447 181389
rect 676489 181386 676555 181389
rect 667381 181384 676555 181386
rect 667381 181328 667386 181384
rect 667442 181328 676494 181384
rect 676550 181328 676555 181384
rect 667381 181326 676555 181328
rect 667381 181323 667447 181326
rect 676489 181323 676555 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 674281 179482 674347 179485
rect 666356 179480 674347 179482
rect 666356 179424 674286 179480
rect 674342 179424 674347 179480
rect 666356 179422 674347 179424
rect 674281 179419 674347 179422
rect 666645 178802 666711 178805
rect 683113 178802 683179 178805
rect 666645 178800 675770 178802
rect 666645 178744 666650 178800
rect 666706 178744 675770 178800
rect 666645 178742 675770 178744
rect 666645 178739 666711 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 675710 177986 675770 178742
rect 683070 178800 683179 178802
rect 683070 178744 683118 178800
rect 683174 178744 683179 178800
rect 683070 178739 683179 178744
rect 683070 178500 683130 178739
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 675710 177926 675954 177986
rect 672901 177850 672967 177853
rect 666356 177848 672967 177850
rect 666356 177792 672906 177848
rect 672962 177792 672967 177848
rect 666356 177790 672967 177792
rect 672901 177787 672967 177790
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 675894 177714 675954 177926
rect 675894 177654 676292 177714
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 674649 177306 674715 177309
rect 674649 177304 676292 177306
rect 674649 177248 674654 177304
rect 674710 177248 676292 177304
rect 674649 177246 676292 177248
rect 674649 177243 674715 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673361 176898 673427 176901
rect 673361 176896 676292 176898
rect 673361 176840 673366 176896
rect 673422 176840 676292 176896
rect 673361 176838 676292 176840
rect 673361 176835 673427 176838
rect 667841 176490 667907 176493
rect 667841 176488 676292 176490
rect 667841 176432 667846 176488
rect 667902 176432 676292 176488
rect 667841 176430 676292 176432
rect 667841 176427 667907 176430
rect 673177 176082 673243 176085
rect 673177 176080 676292 176082
rect 673177 176024 673182 176080
rect 673238 176024 676292 176080
rect 673177 176022 676292 176024
rect 673177 176019 673243 176022
rect 673545 175674 673611 175677
rect 673545 175672 676292 175674
rect 673545 175616 673550 175672
rect 673606 175616 676292 175672
rect 673545 175614 676292 175616
rect 673545 175611 673611 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674649 175266 674715 175269
rect 674649 175264 676292 175266
rect 575982 175130 576042 175236
rect 674649 175208 674654 175264
rect 674710 175208 676292 175264
rect 674649 175206 676292 175208
rect 674649 175203 674715 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 671889 174858 671955 174861
rect 671889 174856 676292 174858
rect 671889 174800 671894 174856
rect 671950 174800 676292 174856
rect 671889 174798 676292 174800
rect 671889 174795 671955 174798
rect 667933 174586 667999 174589
rect 666356 174584 667999 174586
rect 666356 174528 667938 174584
rect 667994 174528 667999 174584
rect 666356 174526 667999 174528
rect 667933 174523 667999 174526
rect 674373 174450 674439 174453
rect 674373 174448 676292 174450
rect 674373 174392 674378 174448
rect 674434 174392 676292 174448
rect 674373 174390 676292 174392
rect 674373 174387 674439 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 680997 173226 681063 173229
rect 680997 173224 681076 173226
rect 680997 173168 681002 173224
rect 681058 173168 681076 173224
rect 680997 173166 681076 173168
rect 680997 173163 681063 173166
rect 671705 172954 671771 172957
rect 666356 172952 671771 172954
rect 666356 172896 671710 172952
rect 671766 172896 671771 172952
rect 666356 172894 671771 172896
rect 671705 172891 671771 172894
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 670601 172002 670667 172005
rect 670601 172000 676292 172002
rect 670601 171944 670606 172000
rect 670662 171944 676292 172000
rect 670601 171942 676292 171944
rect 670601 171939 670667 171942
rect 678237 171594 678303 171597
rect 678237 171592 678316 171594
rect 678237 171536 678242 171592
rect 678298 171536 678316 171592
rect 678237 171534 678316 171536
rect 678237 171531 678303 171534
rect 679617 171186 679683 171189
rect 679604 171184 679683 171186
rect 679604 171128 679622 171184
rect 679678 171128 679683 171184
rect 679604 171126 679683 171128
rect 679617 171123 679683 171126
rect 579521 171050 579587 171053
rect 575798 171048 579587 171050
rect 575798 170992 579526 171048
rect 579582 170992 579587 171048
rect 575798 170990 579587 170992
rect 575798 170884 575858 170990
rect 579521 170987 579587 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589457 170506 589523 170509
rect 589457 170504 592572 170506
rect 589457 170448 589462 170504
rect 589518 170448 592572 170504
rect 589457 170446 592572 170448
rect 589457 170443 589523 170446
rect 675702 170308 675708 170372
rect 675772 170370 675778 170372
rect 675772 170310 676292 170370
rect 675772 170308 675778 170310
rect 671889 169962 671955 169965
rect 671889 169960 676292 169962
rect 671889 169904 671894 169960
rect 671950 169904 676292 169960
rect 671889 169902 676292 169904
rect 671889 169899 671955 169902
rect 669129 169690 669195 169693
rect 666356 169688 669195 169690
rect 666356 169632 669134 169688
rect 669190 169632 669195 169688
rect 666356 169630 669195 169632
rect 669129 169627 669195 169630
rect 669773 169554 669839 169557
rect 669773 169552 676292 169554
rect 669773 169496 669778 169552
rect 669834 169496 676292 169552
rect 669773 169494 676292 169496
rect 669773 169491 669839 169494
rect 578325 169282 578391 169285
rect 575798 169280 578391 169282
rect 575798 169224 578330 169280
rect 578386 169224 578391 169280
rect 575798 169222 578391 169224
rect 575798 168708 575858 169222
rect 578325 169219 578391 169222
rect 672993 169146 673059 169149
rect 672993 169144 676292 169146
rect 672993 169088 672998 169144
rect 673054 169088 676292 169144
rect 672993 169086 676292 169088
rect 672993 169083 673059 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673913 168738 673979 168741
rect 673913 168736 676292 168738
rect 673913 168680 673918 168736
rect 673974 168680 676292 168736
rect 673913 168678 676292 168680
rect 673913 168675 673979 168678
rect 669589 168330 669655 168333
rect 669589 168328 676292 168330
rect 669589 168272 669594 168328
rect 669650 168272 676292 168328
rect 669589 168270 676292 168272
rect 669589 168267 669655 168270
rect 669037 168058 669103 168061
rect 666356 168056 669103 168058
rect 666356 168000 669042 168056
rect 669098 168000 669103 168056
rect 666356 167998 669103 168000
rect 669037 167995 669103 167998
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675886 167452 675892 167516
rect 675956 167514 675962 167516
rect 675956 167454 676292 167514
rect 675956 167452 675962 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578969 166970 579035 166973
rect 575798 166968 579035 166970
rect 575798 166912 578974 166968
rect 579030 166912 579035 166968
rect 575798 166910 579035 166912
rect 575798 166532 575858 166910
rect 578969 166907 579035 166910
rect 671705 166970 671771 166973
rect 676170 166970 676230 167046
rect 671705 166968 676230 166970
rect 671705 166912 671710 166968
rect 671766 166912 676230 166968
rect 671705 166910 676230 166912
rect 671705 166907 671771 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 670141 165610 670207 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 670141 165608 676095 165610
rect 670141 165552 670146 165608
rect 670202 165552 676034 165608
rect 676090 165552 676095 165608
rect 670141 165550 676095 165552
rect 589457 165547 589523 165550
rect 670141 165547 670207 165550
rect 676029 165547 676095 165550
rect 668025 164794 668091 164797
rect 666356 164792 668091 164794
rect 666356 164736 668030 164792
rect 668086 164736 668091 164792
rect 666356 164734 668091 164736
rect 668025 164731 668091 164734
rect 578877 164522 578943 164525
rect 575798 164520 578943 164522
rect 575798 164464 578882 164520
rect 578938 164464 578943 164520
rect 575798 164462 578943 164464
rect 575798 164356 575858 164462
rect 578877 164459 578943 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668945 163162 669011 163165
rect 666356 163160 669011 163162
rect 666356 163104 668950 163160
rect 669006 163104 669011 163160
rect 666356 163102 669011 163104
rect 668945 163099 669011 163102
rect 579429 162482 579495 162485
rect 575798 162480 579495 162482
rect 575798 162424 579434 162480
rect 579490 162424 579495 162480
rect 575798 162422 579495 162424
rect 575798 162180 575858 162422
rect 579429 162419 579495 162422
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675201 161938 675267 161941
rect 675845 161938 675911 161941
rect 675201 161936 675911 161938
rect 675201 161880 675206 161936
rect 675262 161880 675850 161936
rect 675906 161880 675911 161936
rect 675201 161878 675911 161880
rect 675201 161875 675267 161878
rect 675845 161875 675911 161878
rect 675518 161332 675524 161396
rect 675588 161394 675594 161396
rect 676029 161394 676095 161397
rect 675588 161392 676095 161394
rect 675588 161336 676034 161392
rect 676090 161336 676095 161392
rect 675588 161334 676095 161336
rect 675588 161332 675594 161334
rect 676029 161331 676095 161334
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 666185 160170 666251 160173
rect 666142 160168 666251 160170
rect 666142 160112 666190 160168
rect 666246 160112 666251 160168
rect 666142 160107 666251 160112
rect 575982 159898 576042 160004
rect 579245 159898 579311 159901
rect 575982 159896 579311 159898
rect 575982 159840 579250 159896
rect 579306 159840 579311 159896
rect 666142 159868 666202 160107
rect 575982 159838 579311 159840
rect 579245 159835 579311 159838
rect 675753 159490 675819 159493
rect 676438 159490 676444 159492
rect 675753 159488 676444 159490
rect 675753 159432 675758 159488
rect 675814 159432 676444 159488
rect 675753 159430 676444 159432
rect 675753 159427 675819 159430
rect 676438 159428 676444 159430
rect 676508 159428 676514 159492
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 579153 158266 579219 158269
rect 671521 158266 671587 158269
rect 575798 158264 579219 158266
rect 575798 158208 579158 158264
rect 579214 158208 579219 158264
rect 575798 158206 579219 158208
rect 666356 158264 671587 158266
rect 666356 158208 671526 158264
rect 671582 158208 671587 158264
rect 666356 158206 671587 158208
rect 575798 157828 575858 158206
rect 579153 158203 579219 158206
rect 671521 158203 671587 158206
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589457 157450 589523 157453
rect 589457 157448 592572 157450
rect 589457 157392 589462 157448
rect 589518 157392 592572 157448
rect 589457 157390 592572 157392
rect 589457 157387 589523 157390
rect 675569 157044 675635 157045
rect 675518 156980 675524 157044
rect 675588 157042 675635 157044
rect 675588 157040 675680 157042
rect 675630 156984 675680 157040
rect 675588 156982 675680 156984
rect 675588 156980 675635 156982
rect 675569 156979 675635 156980
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 579521 155954 579587 155957
rect 575798 155952 579587 155954
rect 575798 155896 579526 155952
rect 579582 155896 579587 155952
rect 575798 155894 579587 155896
rect 575798 155652 575858 155894
rect 579521 155891 579587 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 666326 154594 666386 154972
rect 674046 154594 674052 154596
rect 666326 154534 674052 154594
rect 674046 154532 674052 154534
rect 674116 154532 674122 154596
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578233 154050 578299 154053
rect 575798 154048 578299 154050
rect 575798 153992 578238 154048
rect 578294 153992 578299 154048
rect 575798 153990 578299 153992
rect 575798 153476 575858 153990
rect 578233 153987 578299 153990
rect 668761 153370 668827 153373
rect 666356 153368 668827 153370
rect 666356 153312 668766 153368
rect 668822 153312 668827 153368
rect 666356 153310 668827 153312
rect 668761 153307 668827 153310
rect 672993 153098 673059 153101
rect 675109 153098 675175 153101
rect 672993 153096 675175 153098
rect 672993 153040 672998 153096
rect 673054 153040 675114 153096
rect 675170 153040 675175 153096
rect 672993 153038 675175 153040
rect 672993 153035 673059 153038
rect 675109 153035 675175 153038
rect 675753 153098 675819 153101
rect 676254 153098 676260 153100
rect 675753 153096 676260 153098
rect 675753 153040 675758 153096
rect 675814 153040 676260 153096
rect 675753 153038 676260 153040
rect 675753 153035 675819 153038
rect 676254 153036 676260 153038
rect 676324 153036 676330 153100
rect 669773 152690 669839 152693
rect 675293 152690 675359 152693
rect 669773 152688 675359 152690
rect 669773 152632 669778 152688
rect 669834 152632 675298 152688
rect 675354 152632 675359 152688
rect 669773 152630 675359 152632
rect 669773 152627 669839 152630
rect 675293 152627 675359 152630
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 671889 151738 671955 151741
rect 675109 151738 675175 151741
rect 671889 151736 675175 151738
rect 671889 151680 671894 151736
rect 671950 151680 675114 151736
rect 675170 151680 675175 151736
rect 671889 151678 675175 151680
rect 671889 151675 671955 151678
rect 675109 151675 675175 151678
rect 673913 151058 673979 151061
rect 675109 151058 675175 151061
rect 673913 151056 675175 151058
rect 673913 151000 673918 151056
rect 673974 151000 675114 151056
rect 675170 151000 675175 151056
rect 673913 150998 675175 151000
rect 673913 150995 673979 150998
rect 675109 150995 675175 150998
rect 589457 150922 589523 150925
rect 589457 150920 592572 150922
rect 589457 150864 589462 150920
rect 589518 150864 592572 150920
rect 589457 150862 592572 150864
rect 589457 150859 589523 150862
rect 675753 150380 675819 150381
rect 675702 150378 675708 150380
rect 675662 150318 675708 150378
rect 675772 150376 675819 150380
rect 675814 150320 675819 150376
rect 675702 150316 675708 150318
rect 675772 150316 675819 150320
rect 675753 150315 675819 150316
rect 668669 150106 668735 150109
rect 666356 150104 668735 150106
rect 666356 150048 668674 150104
rect 668730 150048 668735 150104
rect 666356 150046 668735 150048
rect 668669 150043 668735 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589181 149290 589247 149293
rect 589181 149288 592572 149290
rect 589181 149232 589186 149288
rect 589242 149232 592572 149288
rect 589181 149230 592572 149232
rect 589181 149227 589247 149230
rect 670601 149018 670667 149021
rect 675293 149018 675359 149021
rect 670601 149016 675359 149018
rect 670601 148960 670606 149016
rect 670662 148960 675298 149016
rect 675354 148960 675359 149016
rect 670601 148958 675359 148960
rect 670601 148955 670667 148958
rect 675293 148955 675359 148958
rect 668485 148474 668551 148477
rect 666356 148472 668551 148474
rect 666356 148416 668490 148472
rect 668546 148416 668551 148472
rect 666356 148414 668551 148416
rect 668485 148411 668551 148414
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 668761 147794 668827 147797
rect 673310 147794 673316 147796
rect 668761 147792 673316 147794
rect 668761 147736 668766 147792
rect 668822 147736 673316 147792
rect 668761 147734 673316 147736
rect 668761 147731 668827 147734
rect 673310 147732 673316 147734
rect 673380 147732 673386 147796
rect 589365 147658 589431 147661
rect 675661 147658 675727 147661
rect 675886 147658 675892 147660
rect 589365 147656 592572 147658
rect 589365 147600 589370 147656
rect 589426 147600 592572 147656
rect 589365 147598 592572 147600
rect 675661 147656 675892 147658
rect 675661 147600 675666 147656
rect 675722 147600 675892 147656
rect 675661 147598 675892 147600
rect 589365 147595 589431 147598
rect 675661 147595 675727 147598
rect 675886 147596 675892 147598
rect 675956 147596 675962 147660
rect 579521 147250 579587 147253
rect 575798 147248 579587 147250
rect 575798 147192 579526 147248
rect 579582 147192 579587 147248
rect 575798 147190 579587 147192
rect 575798 146948 575858 147190
rect 579521 147187 579587 147190
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 671286 145210 671292 145212
rect 666356 145150 671292 145210
rect 671286 145148 671292 145150
rect 671356 145148 671362 145212
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589917 144394 589983 144397
rect 589917 144392 592572 144394
rect 589917 144336 589922 144392
rect 589978 144336 592572 144392
rect 589917 144334 592572 144336
rect 589917 144331 589983 144334
rect 673678 143578 673684 143580
rect 666356 143518 673684 143578
rect 673678 143516 673684 143518
rect 673748 143516 673754 143580
rect 578509 143034 578575 143037
rect 575798 143032 578575 143034
rect 575798 142976 578514 143032
rect 578570 142976 578575 143032
rect 575798 142974 578575 142976
rect 575798 142596 575858 142974
rect 578509 142971 578575 142974
rect 589457 142762 589523 142765
rect 589457 142760 592572 142762
rect 589457 142704 589462 142760
rect 589518 142704 592572 142760
rect 589457 142702 592572 142704
rect 589457 142699 589523 142702
rect 589089 141130 589155 141133
rect 589089 141128 592572 141130
rect 589089 141072 589094 141128
rect 589150 141072 592572 141128
rect 589089 141070 592572 141072
rect 589089 141067 589155 141070
rect 579521 140586 579587 140589
rect 575798 140584 579587 140586
rect 575798 140528 579526 140584
rect 579582 140528 579587 140584
rect 575798 140526 579587 140528
rect 575798 140420 575858 140526
rect 579521 140523 579587 140526
rect 672257 140314 672323 140317
rect 666356 140312 672323 140314
rect 666356 140256 672262 140312
rect 672318 140256 672323 140312
rect 666356 140254 672323 140256
rect 672257 140251 672323 140254
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578693 138818 578759 138821
rect 575798 138816 578759 138818
rect 575798 138760 578698 138816
rect 578754 138760 578759 138816
rect 575798 138758 578759 138760
rect 575798 138244 575858 138758
rect 578693 138755 578759 138758
rect 669129 138682 669195 138685
rect 666356 138680 669195 138682
rect 666356 138624 669134 138680
rect 669190 138624 669195 138680
rect 666356 138622 669195 138624
rect 669129 138619 669195 138622
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589273 136234 589339 136237
rect 589273 136232 592572 136234
rect 589273 136176 589278 136232
rect 589334 136176 592572 136232
rect 589273 136174 592572 136176
rect 589273 136171 589339 136174
rect 667565 135962 667631 135965
rect 683113 135962 683179 135965
rect 667565 135960 683179 135962
rect 667565 135904 667570 135960
rect 667626 135904 683118 135960
rect 683174 135904 683179 135960
rect 667565 135902 683179 135904
rect 667565 135899 667631 135902
rect 683113 135899 683179 135902
rect 667933 135418 667999 135421
rect 666356 135416 667999 135418
rect 666356 135360 667938 135416
rect 667994 135360 667999 135416
rect 666356 135358 667999 135360
rect 667933 135355 667999 135358
rect 589457 134602 589523 134605
rect 667197 134602 667263 134605
rect 675845 134602 675911 134605
rect 589457 134600 592572 134602
rect 589457 134544 589462 134600
rect 589518 134544 592572 134600
rect 589457 134542 592572 134544
rect 667197 134600 675911 134602
rect 667197 134544 667202 134600
rect 667258 134544 675850 134600
rect 675906 134544 675911 134600
rect 667197 134542 675911 134544
rect 589457 134539 589523 134542
rect 667197 134539 667263 134542
rect 675845 134539 675911 134542
rect 578325 134466 578391 134469
rect 575798 134464 578391 134466
rect 575798 134408 578330 134464
rect 578386 134408 578391 134464
rect 575798 134406 578391 134408
rect 575798 133892 575858 134406
rect 578325 134403 578391 134406
rect 672073 133786 672139 133789
rect 666356 133784 672139 133786
rect 666356 133728 672078 133784
rect 672134 133728 672139 133784
rect 666356 133726 672139 133728
rect 672073 133723 672139 133726
rect 667013 133106 667079 133109
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 667013 133104 676322 133106
rect 667013 133048 667018 133104
rect 667074 133048 676322 133104
rect 667013 133046 676322 133048
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 667013 133043 667079 133046
rect 676446 133043 676555 133048
rect 588537 132970 588603 132973
rect 588537 132968 592572 132970
rect 588537 132912 588542 132968
rect 588598 132912 592572 132968
rect 676446 132940 676506 133043
rect 588537 132910 592572 132912
rect 588537 132907 588603 132910
rect 683113 132698 683179 132701
rect 682886 132696 683179 132698
rect 682886 132640 683118 132696
rect 683174 132640 683179 132696
rect 682886 132638 683179 132640
rect 682886 132532 682946 132638
rect 683113 132635 683179 132638
rect 578233 132290 578299 132293
rect 575798 132288 578299 132290
rect 575798 132232 578238 132288
rect 578294 132232 578299 132288
rect 575798 132230 578299 132232
rect 575798 131716 575858 132230
rect 578233 132227 578299 132230
rect 673361 132154 673427 132157
rect 673361 132152 676292 132154
rect 673361 132096 673366 132152
rect 673422 132096 676292 132152
rect 673361 132094 676292 132096
rect 673361 132091 673427 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 590101 131338 590167 131341
rect 673177 131338 673243 131341
rect 590101 131336 592572 131338
rect 590101 131280 590106 131336
rect 590162 131280 592572 131336
rect 590101 131278 592572 131280
rect 673177 131336 676292 131338
rect 673177 131280 673182 131336
rect 673238 131280 676292 131336
rect 673177 131278 676292 131280
rect 590101 131275 590167 131278
rect 673177 131275 673243 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130522 667980 130524
rect 666356 130462 667980 130522
rect 667974 130460 667980 130462
rect 668044 130460 668050 130524
rect 674649 130522 674715 130525
rect 674649 130520 676292 130522
rect 674649 130464 674654 130520
rect 674710 130464 676292 130520
rect 674649 130462 676292 130464
rect 674649 130459 674715 130462
rect 675937 130114 676003 130117
rect 675937 130112 676292 130114
rect 675937 130056 675942 130112
rect 675998 130056 676292 130112
rect 675937 130054 676292 130056
rect 675937 130051 676003 130054
rect 579521 129706 579587 129709
rect 575798 129704 579587 129706
rect 575798 129648 579526 129704
rect 579582 129648 579587 129704
rect 575798 129646 579587 129648
rect 575798 129540 575858 129646
rect 579521 129643 579587 129646
rect 589457 129706 589523 129709
rect 674373 129706 674439 129709
rect 589457 129704 592572 129706
rect 589457 129648 589462 129704
rect 589518 129648 592572 129704
rect 589457 129646 592572 129648
rect 674373 129704 676292 129706
rect 674373 129648 674378 129704
rect 674434 129648 676292 129704
rect 674373 129646 676292 129648
rect 589457 129643 589523 129646
rect 674373 129643 674439 129646
rect 674465 129298 674531 129301
rect 674465 129296 676292 129298
rect 674465 129240 674470 129296
rect 674526 129240 676292 129296
rect 674465 129238 676292 129240
rect 674465 129235 674531 129238
rect 666326 128482 666386 128860
rect 676630 128620 676690 128860
rect 676622 128556 676628 128620
rect 676692 128556 676698 128620
rect 673494 128482 673500 128484
rect 666326 128422 673500 128482
rect 673494 128420 673500 128422
rect 673564 128420 673570 128484
rect 674281 128346 674347 128349
rect 675937 128346 676003 128349
rect 674281 128344 676003 128346
rect 674281 128288 674286 128344
rect 674342 128288 675942 128344
rect 675998 128288 676003 128344
rect 674281 128286 676003 128288
rect 674281 128283 674347 128286
rect 675937 128283 676003 128286
rect 668577 128210 668643 128213
rect 674097 128210 674163 128213
rect 668577 128208 674163 128210
rect 668577 128152 668582 128208
rect 668638 128152 674102 128208
rect 674158 128152 674163 128208
rect 668577 128150 674163 128152
rect 668577 128147 668643 128150
rect 674097 128147 674163 128150
rect 676070 128148 676076 128212
rect 676140 128210 676146 128212
rect 676262 128210 676322 128452
rect 676140 128150 676322 128210
rect 676140 128148 676146 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 682334 127805 682394 128044
rect 578325 127802 578391 127805
rect 575798 127800 578391 127802
rect 575798 127744 578330 127800
rect 578386 127744 578391 127800
rect 575798 127742 578391 127744
rect 682334 127800 682443 127805
rect 682334 127744 682382 127800
rect 682438 127744 682443 127800
rect 682334 127742 682443 127744
rect 575798 127364 575858 127742
rect 578325 127739 578391 127742
rect 682377 127739 682443 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 676254 126924 676260 126988
rect 676324 126924 676330 126988
rect 676262 126820 676322 126924
rect 589917 126442 589983 126445
rect 675017 126442 675083 126445
rect 589917 126440 592572 126442
rect 589917 126384 589922 126440
rect 589978 126384 592572 126440
rect 589917 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 589917 126379 589983 126382
rect 675017 126379 675083 126382
rect 672993 126034 673059 126037
rect 672993 126032 676292 126034
rect 672993 125976 672998 126032
rect 673054 125976 676292 126032
rect 672993 125974 676292 125976
rect 672993 125971 673059 125974
rect 668761 125626 668827 125629
rect 666356 125624 668827 125626
rect 666356 125568 668766 125624
rect 668822 125568 668827 125624
rect 666356 125566 668827 125568
rect 668761 125563 668827 125566
rect 674649 125626 674715 125629
rect 674649 125624 676292 125626
rect 674649 125568 674654 125624
rect 674710 125568 676292 125624
rect 674649 125566 676292 125568
rect 674649 125563 674715 125566
rect 579245 125354 579311 125357
rect 575798 125352 579311 125354
rect 575798 125296 579250 125352
rect 579306 125296 579311 125352
rect 575798 125294 579311 125296
rect 575798 125188 575858 125294
rect 579245 125291 579311 125294
rect 674097 125218 674163 125221
rect 674097 125216 676292 125218
rect 674097 125160 674102 125216
rect 674158 125160 676292 125216
rect 674097 125158 676292 125160
rect 674097 125155 674163 125158
rect 589457 124810 589523 124813
rect 589457 124808 592572 124810
rect 589457 124752 589462 124808
rect 589518 124752 592572 124808
rect 589457 124750 592572 124752
rect 589457 124747 589523 124750
rect 676446 124540 676506 124780
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 673177 124402 673243 124405
rect 673177 124400 676292 124402
rect 673177 124344 673182 124400
rect 673238 124344 676292 124400
rect 673177 124342 676292 124344
rect 673177 124339 673243 124342
rect 672717 123994 672783 123997
rect 666356 123992 672783 123994
rect 666356 123936 672722 123992
rect 672778 123936 672783 123992
rect 666356 123934 672783 123936
rect 672717 123931 672783 123934
rect 672950 123934 676292 123994
rect 672533 123722 672599 123725
rect 672950 123722 673010 123934
rect 672533 123720 673010 123722
rect 672533 123664 672538 123720
rect 672594 123664 673010 123720
rect 672533 123662 673010 123664
rect 672533 123659 672599 123662
rect 579245 123586 579311 123589
rect 575798 123584 579311 123586
rect 575798 123528 579250 123584
rect 579306 123528 579311 123584
rect 575798 123526 579311 123528
rect 575798 123012 575858 123526
rect 579245 123523 579311 123526
rect 673361 123586 673427 123589
rect 673361 123584 676292 123586
rect 673361 123528 673366 123584
rect 673422 123528 676292 123584
rect 673361 123526 676292 123528
rect 673361 123523 673427 123526
rect 589457 123178 589523 123181
rect 672349 123178 672415 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672349 123176 676292 123178
rect 672349 123120 672354 123176
rect 672410 123120 676292 123176
rect 672349 123118 676292 123120
rect 589457 123115 589523 123118
rect 672349 123115 672415 123118
rect 669957 122770 670023 122773
rect 669957 122768 676292 122770
rect 669957 122712 669962 122768
rect 670018 122712 676292 122768
rect 669957 122710 676292 122712
rect 669957 122707 670023 122710
rect 675702 122300 675708 122364
rect 675772 122362 675778 122364
rect 675772 122302 676292 122362
rect 675772 122300 675778 122302
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589457 121546 589523 121549
rect 589457 121544 592572 121546
rect 589457 121488 589462 121544
rect 589518 121488 592572 121544
rect 589457 121486 592572 121488
rect 589457 121483 589523 121486
rect 672717 121410 672783 121413
rect 675894 121410 675954 121622
rect 672717 121408 675954 121410
rect 672717 121352 672722 121408
rect 672778 121352 675954 121408
rect 672717 121350 675954 121352
rect 672717 121347 672783 121350
rect 579061 121138 579127 121141
rect 575798 121136 579127 121138
rect 575798 121080 579066 121136
rect 579122 121080 579127 121136
rect 575798 121078 579127 121080
rect 575798 120836 575858 121078
rect 579061 121075 579127 121078
rect 668577 120730 668643 120733
rect 666356 120728 668643 120730
rect 666356 120672 668582 120728
rect 668638 120672 668643 120728
rect 666356 120670 668643 120672
rect 668577 120667 668643 120670
rect 668669 120186 668735 120189
rect 672349 120186 672415 120189
rect 668669 120184 672415 120186
rect 668669 120128 668674 120184
rect 668730 120128 672354 120184
rect 672410 120128 672415 120184
rect 668669 120126 672415 120128
rect 668669 120123 668735 120126
rect 672349 120123 672415 120126
rect 590101 119914 590167 119917
rect 590101 119912 592572 119914
rect 590101 119856 590106 119912
rect 590162 119856 592572 119912
rect 590101 119854 592572 119856
rect 590101 119851 590167 119854
rect 669221 119098 669287 119101
rect 666356 119096 669287 119098
rect 666356 119040 669226 119096
rect 669282 119040 669287 119096
rect 666356 119038 669287 119040
rect 669221 119035 669287 119038
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 668025 117466 668091 117469
rect 666356 117464 668091 117466
rect 666356 117408 668030 117464
rect 668086 117408 668091 117464
rect 666356 117406 668091 117408
rect 668025 117403 668091 117406
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 671705 115834 671771 115837
rect 666356 115832 671771 115834
rect 666356 115776 671710 115832
rect 671766 115776 671771 115832
rect 666356 115774 671771 115776
rect 671705 115771 671771 115774
rect 589825 115018 589891 115021
rect 589825 115016 592572 115018
rect 589825 114960 589830 115016
rect 589886 114960 592572 115016
rect 589825 114958 592572 114960
rect 589825 114955 589891 114958
rect 579521 114474 579587 114477
rect 575798 114472 579587 114474
rect 575798 114416 579526 114472
rect 579582 114416 579587 114472
rect 575798 114414 579587 114416
rect 575798 114308 575858 114414
rect 579521 114411 579587 114414
rect 668669 114202 668735 114205
rect 666356 114200 668735 114202
rect 666356 114144 668674 114200
rect 668730 114144 668735 114200
rect 666356 114142 668735 114144
rect 668669 114139 668735 114142
rect 590561 113386 590627 113389
rect 590561 113384 592572 113386
rect 590561 113328 590566 113384
rect 590622 113328 592572 113384
rect 590561 113326 592572 113328
rect 590561 113323 590627 113326
rect 675293 113114 675359 113117
rect 676622 113114 676628 113116
rect 675293 113112 676628 113114
rect 675293 113056 675298 113112
rect 675354 113056 676628 113112
rect 675293 113054 676628 113056
rect 675293 113051 675359 113054
rect 676622 113052 676628 113054
rect 676692 113052 676698 113116
rect 579521 112706 579587 112709
rect 575798 112704 579587 112706
rect 575798 112648 579526 112704
rect 579582 112648 579587 112704
rect 575798 112646 579587 112648
rect 575798 112132 575858 112646
rect 579521 112643 579587 112646
rect 668117 112570 668183 112573
rect 666356 112568 668183 112570
rect 666356 112512 668122 112568
rect 668178 112512 668183 112568
rect 666356 112510 668183 112512
rect 668117 112507 668183 112510
rect 668301 111890 668367 111893
rect 674465 111890 674531 111893
rect 668301 111888 674531 111890
rect 668301 111832 668306 111888
rect 668362 111832 674470 111888
rect 674526 111832 674531 111888
rect 668301 111830 674531 111832
rect 668301 111827 668367 111830
rect 674465 111827 674531 111830
rect 589365 111754 589431 111757
rect 589365 111752 592572 111754
rect 589365 111696 589370 111752
rect 589426 111696 592572 111752
rect 589365 111694 592572 111696
rect 589365 111691 589431 111694
rect 672993 111482 673059 111485
rect 675109 111482 675175 111485
rect 672993 111480 675175 111482
rect 672993 111424 672998 111480
rect 673054 111424 675114 111480
rect 675170 111424 675175 111480
rect 672993 111422 675175 111424
rect 672993 111419 673059 111422
rect 675109 111419 675175 111422
rect 672717 110938 672783 110941
rect 666356 110936 672783 110938
rect 666356 110880 672722 110936
rect 672778 110880 672783 110936
rect 666356 110878 672783 110880
rect 672717 110875 672783 110878
rect 673177 110394 673243 110397
rect 675109 110394 675175 110397
rect 673177 110392 675175 110394
rect 673177 110336 673182 110392
rect 673238 110336 675114 110392
rect 675170 110336 675175 110392
rect 673177 110334 675175 110336
rect 673177 110331 673243 110334
rect 675109 110331 675175 110334
rect 579429 110258 579495 110261
rect 575798 110256 579495 110258
rect 575798 110200 579434 110256
rect 579490 110200 579495 110256
rect 575798 110198 579495 110200
rect 575798 109956 575858 110198
rect 579429 110195 579495 110198
rect 589641 110122 589707 110125
rect 589641 110120 592572 110122
rect 589641 110064 589646 110120
rect 589702 110064 592572 110120
rect 589641 110062 592572 110064
rect 589641 110059 589707 110062
rect 668025 109306 668091 109309
rect 666356 109304 668091 109306
rect 666356 109248 668030 109304
rect 668086 109248 668091 109304
rect 666356 109246 668091 109248
rect 668025 109243 668091 109246
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 671521 107674 671587 107677
rect 666356 107672 671587 107674
rect 666356 107616 671526 107672
rect 671582 107616 671587 107672
rect 666356 107614 671587 107616
rect 671521 107611 671587 107614
rect 589917 106858 589983 106861
rect 589917 106856 592572 106858
rect 589917 106800 589922 106856
rect 589978 106800 592572 106856
rect 589917 106798 592572 106800
rect 589917 106795 589983 106798
rect 672533 106314 672599 106317
rect 675109 106314 675175 106317
rect 672533 106312 675175 106314
rect 672533 106256 672538 106312
rect 672594 106256 675114 106312
rect 675170 106256 675175 106312
rect 672533 106254 675175 106256
rect 672533 106251 672599 106254
rect 675109 106251 675175 106254
rect 675753 106178 675819 106181
rect 676438 106178 676444 106180
rect 675753 106176 676444 106178
rect 675753 106120 675758 106176
rect 675814 106120 676444 106176
rect 675753 106118 676444 106120
rect 675753 106115 675819 106118
rect 676438 106116 676444 106118
rect 676508 106116 676514 106180
rect 666645 106042 666711 106045
rect 667197 106042 667263 106045
rect 666356 106040 667263 106042
rect 666356 105984 666650 106040
rect 666706 105984 667202 106040
rect 667258 105984 667263 106040
rect 666356 105982 667263 105984
rect 666645 105979 666711 105982
rect 667197 105979 667263 105982
rect 578325 105906 578391 105909
rect 575798 105904 578391 105906
rect 575798 105848 578330 105904
rect 578386 105848 578391 105904
rect 575798 105846 578391 105848
rect 575798 105604 575858 105846
rect 578325 105843 578391 105846
rect 673361 105634 673427 105637
rect 675109 105634 675175 105637
rect 673361 105632 675175 105634
rect 673361 105576 673366 105632
rect 673422 105576 675114 105632
rect 675170 105576 675175 105632
rect 673361 105574 675175 105576
rect 673361 105571 673427 105574
rect 675109 105571 675175 105574
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 674097 104682 674163 104685
rect 675109 104682 675175 104685
rect 674097 104680 675175 104682
rect 674097 104624 674102 104680
rect 674158 104624 675114 104680
rect 675170 104624 675175 104680
rect 674097 104622 675175 104624
rect 674097 104619 674163 104622
rect 675109 104619 675175 104622
rect 668301 104410 668367 104413
rect 666356 104408 668367 104410
rect 666356 104352 668306 104408
rect 668362 104352 668367 104408
rect 666356 104350 668367 104352
rect 668301 104347 668367 104350
rect 590101 103594 590167 103597
rect 590101 103592 592572 103594
rect 590101 103536 590106 103592
rect 590162 103536 592572 103592
rect 590101 103534 592572 103536
rect 590101 103531 590167 103534
rect 575982 103322 576042 103428
rect 579521 103322 579587 103325
rect 575982 103320 579587 103322
rect 575982 103264 579526 103320
rect 579582 103264 579587 103320
rect 575982 103262 579587 103264
rect 579521 103259 579587 103262
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 666326 102234 666386 102748
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 668485 102234 668551 102237
rect 674281 102234 674347 102237
rect 666326 102232 674347 102234
rect 666326 102176 668490 102232
rect 668546 102176 674286 102232
rect 674342 102176 674347 102232
rect 666326 102174 674347 102176
rect 668485 102171 668551 102174
rect 674281 102171 674347 102174
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579245 101826 579311 101829
rect 575798 101824 579311 101826
rect 575798 101768 579250 101824
rect 579306 101768 579311 101824
rect 575798 101766 579311 101768
rect 575798 101252 575858 101766
rect 579245 101763 579311 101766
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 579521 97474 579587 97477
rect 575798 97472 579587 97474
rect 575798 97416 579526 97472
rect 579582 97416 579587 97472
rect 575798 97414 579587 97416
rect 575798 96900 575858 97414
rect 579521 97411 579587 97414
rect 634854 96868 634860 96932
rect 634924 96930 634930 96932
rect 635733 96930 635799 96933
rect 634924 96928 635799 96930
rect 634924 96872 635738 96928
rect 635794 96872 635799 96928
rect 634924 96870 635799 96872
rect 634924 96868 634930 96870
rect 635733 96867 635799 96870
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 626441 95434 626507 95437
rect 626441 95432 628268 95434
rect 626441 95376 626446 95432
rect 626502 95376 628268 95432
rect 626441 95374 628268 95376
rect 626441 95371 626507 95374
rect 643185 95162 643251 95165
rect 642958 95160 643251 95162
rect 642958 95104 643190 95160
rect 643246 95104 643251 95160
rect 642958 95102 643251 95104
rect 578693 95026 578759 95029
rect 575798 95024 578759 95026
rect 575798 94968 578698 95024
rect 578754 94968 578759 95024
rect 575798 94966 578759 94968
rect 575798 94724 575858 94966
rect 578693 94963 578759 94966
rect 642958 94588 643018 95102
rect 643185 95099 643251 95102
rect 626257 94482 626323 94485
rect 626257 94480 628268 94482
rect 626257 94424 626262 94480
rect 626318 94424 628268 94480
rect 626257 94422 628268 94424
rect 626257 94419 626323 94422
rect 655237 94210 655303 94213
rect 655237 94208 656788 94210
rect 655237 94152 655242 94208
rect 655298 94152 656788 94208
rect 655237 94150 656788 94152
rect 655237 94147 655303 94150
rect 626441 93530 626507 93533
rect 626441 93528 628268 93530
rect 626441 93472 626446 93528
rect 626502 93472 628268 93528
rect 626441 93470 628268 93472
rect 626441 93467 626507 93470
rect 655053 93394 655119 93397
rect 665541 93394 665607 93397
rect 655053 93392 656788 93394
rect 655053 93336 655058 93392
rect 655114 93336 656788 93392
rect 655053 93334 656788 93336
rect 663596 93392 665607 93394
rect 663596 93336 665546 93392
rect 665602 93336 665607 93392
rect 663596 93334 665607 93336
rect 655053 93331 655119 93334
rect 665541 93331 665607 93334
rect 579521 93122 579587 93125
rect 575798 93120 579587 93122
rect 575798 93064 579526 93120
rect 579582 93064 579587 93120
rect 575798 93062 579587 93064
rect 575798 92548 575858 93062
rect 579521 93059 579587 93062
rect 625429 93122 625495 93125
rect 625429 93120 628298 93122
rect 625429 93064 625434 93120
rect 625490 93064 628298 93120
rect 625429 93062 628298 93064
rect 625429 93059 625495 93062
rect 628238 92548 628298 93062
rect 654869 92578 654935 92581
rect 665173 92578 665239 92581
rect 654869 92576 656788 92578
rect 654869 92520 654874 92576
rect 654930 92520 656788 92576
rect 654869 92518 656788 92520
rect 663596 92576 665239 92578
rect 663596 92520 665178 92576
rect 665234 92520 665239 92576
rect 663596 92518 665239 92520
rect 654869 92515 654935 92518
rect 665173 92515 665239 92518
rect 644933 92170 644999 92173
rect 642988 92168 644999 92170
rect 642988 92112 644938 92168
rect 644994 92112 644999 92168
rect 642988 92110 644999 92112
rect 644933 92107 644999 92110
rect 663701 92034 663767 92037
rect 663382 92032 663767 92034
rect 663382 91976 663706 92032
rect 663762 91976 663767 92032
rect 663382 91974 663767 91976
rect 663382 91732 663442 91974
rect 663701 91971 663767 91974
rect 625429 91626 625495 91629
rect 625429 91624 628268 91626
rect 625429 91568 625434 91624
rect 625490 91568 628268 91624
rect 625429 91566 628268 91568
rect 625429 91563 625495 91566
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 579061 90946 579127 90949
rect 575798 90944 579127 90946
rect 575798 90888 579066 90944
rect 579122 90888 579127 90944
rect 575798 90886 579127 90888
rect 575798 90372 575858 90886
rect 579061 90883 579127 90886
rect 626441 90674 626507 90677
rect 654133 90674 654199 90677
rect 665357 90674 665423 90677
rect 626441 90672 628268 90674
rect 626441 90616 626446 90672
rect 626502 90616 628268 90672
rect 626441 90614 628268 90616
rect 654133 90672 656788 90674
rect 654133 90616 654138 90672
rect 654194 90616 656788 90672
rect 654133 90614 656788 90616
rect 663596 90672 665423 90674
rect 663596 90616 665362 90672
rect 665418 90616 665423 90672
rect 663596 90614 665423 90616
rect 626441 90611 626507 90614
rect 654133 90611 654199 90614
rect 665357 90611 665423 90614
rect 655789 89858 655855 89861
rect 664621 89858 664687 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664687 89858
rect 663596 89800 664626 89856
rect 664682 89800 664687 89856
rect 663596 89798 664687 89800
rect 655789 89795 655855 89798
rect 664621 89795 664687 89798
rect 625797 89722 625863 89725
rect 644013 89722 644079 89725
rect 625797 89720 628268 89722
rect 625797 89664 625802 89720
rect 625858 89664 628268 89720
rect 625797 89662 628268 89664
rect 642988 89720 644079 89722
rect 642988 89664 644018 89720
rect 644074 89664 644079 89720
rect 642988 89662 644079 89664
rect 625797 89659 625863 89662
rect 644013 89659 644079 89662
rect 664161 89042 664227 89045
rect 663596 89040 664227 89042
rect 663596 88984 664166 89040
rect 664222 88984 664227 89040
rect 663596 88982 664227 88984
rect 664161 88979 664227 88982
rect 626441 88906 626507 88909
rect 626441 88904 628268 88906
rect 626441 88848 626446 88904
rect 626502 88848 628268 88904
rect 626441 88846 628268 88848
rect 626441 88843 626507 88846
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 643461 87138 643527 87141
rect 642988 87136 643527 87138
rect 642988 87080 643466 87136
rect 643522 87080 643527 87136
rect 642988 87078 643527 87080
rect 643461 87075 643527 87078
rect 625613 87002 625679 87005
rect 625613 87000 628268 87002
rect 625613 86944 625618 87000
rect 625674 86944 628268 87000
rect 625613 86942 628268 86944
rect 625613 86939 625679 86942
rect 578601 86458 578667 86461
rect 575798 86456 578667 86458
rect 575798 86400 578606 86456
rect 578662 86400 578667 86456
rect 575798 86398 578667 86400
rect 575798 86020 575858 86398
rect 578601 86395 578667 86398
rect 626441 86050 626507 86053
rect 626441 86048 628268 86050
rect 626441 85992 626446 86048
rect 626502 85992 628268 86048
rect 626441 85990 628268 85992
rect 626441 85987 626507 85990
rect 626441 85098 626507 85101
rect 626441 85096 628268 85098
rect 626441 85040 626446 85096
rect 626502 85040 628268 85096
rect 626441 85038 628268 85040
rect 626441 85035 626507 85038
rect 644749 84690 644815 84693
rect 642988 84688 644815 84690
rect 642988 84632 644754 84688
rect 644810 84632 644815 84688
rect 642988 84630 644815 84632
rect 644749 84627 644815 84630
rect 625613 84146 625679 84149
rect 625613 84144 628268 84146
rect 625613 84088 625618 84144
rect 625674 84088 628268 84144
rect 625613 84086 628268 84088
rect 625613 84083 625679 84086
rect 579245 84010 579311 84013
rect 575798 84008 579311 84010
rect 575798 83952 579250 84008
rect 579306 83952 579311 84008
rect 575798 83950 579311 83952
rect 575798 83844 575858 83950
rect 579245 83947 579311 83950
rect 624417 82922 624483 82925
rect 628238 82922 628298 83164
rect 624417 82920 628298 82922
rect 624417 82864 624422 82920
rect 624478 82864 628298 82920
rect 624417 82862 628298 82864
rect 624417 82859 624483 82862
rect 643737 82786 643803 82789
rect 642958 82784 643803 82786
rect 642958 82728 643742 82784
rect 643798 82728 643803 82784
rect 642958 82726 643803 82728
rect 579245 82242 579311 82245
rect 575798 82240 579311 82242
rect 575798 82184 579250 82240
rect 579306 82184 579311 82240
rect 642958 82212 643018 82726
rect 643737 82723 643803 82726
rect 575798 82182 579311 82184
rect 575798 81668 575858 82182
rect 579245 82179 579311 82182
rect 628606 81701 628666 82212
rect 628606 81696 628715 81701
rect 628606 81640 628654 81696
rect 628710 81640 628715 81696
rect 628606 81638 628715 81640
rect 628649 81635 628715 81638
rect 628790 80882 628850 81396
rect 629201 80882 629267 80885
rect 628790 80880 629267 80882
rect 628790 80824 629206 80880
rect 629262 80824 629267 80880
rect 628790 80822 629267 80824
rect 629201 80819 629267 80822
rect 633893 80474 633959 80477
rect 634854 80474 634860 80476
rect 633893 80472 634860 80474
rect 633893 80416 633898 80472
rect 633954 80416 634860 80472
rect 633893 80414 634860 80416
rect 633893 80411 633959 80414
rect 634854 80412 634860 80414
rect 634924 80412 634930 80476
rect 578785 80066 578851 80069
rect 575798 80064 578851 80066
rect 575798 80008 578790 80064
rect 578846 80008 578851 80064
rect 575798 80006 578851 80008
rect 575798 79492 575858 80006
rect 578785 80003 578851 80006
rect 578969 77890 579035 77893
rect 575798 77888 579035 77890
rect 575798 77832 578974 77888
rect 579030 77832 579035 77888
rect 575798 77830 579035 77832
rect 575798 77316 575858 77830
rect 578969 77827 579035 77830
rect 585777 77890 585843 77893
rect 637062 77890 637068 77892
rect 585777 77888 637068 77890
rect 585777 77832 585782 77888
rect 585838 77832 637068 77888
rect 585777 77830 637068 77832
rect 585777 77827 585843 77830
rect 637062 77828 637068 77830
rect 637132 77890 637138 77892
rect 639597 77890 639663 77893
rect 637132 77888 639663 77890
rect 637132 77832 639602 77888
rect 639658 77832 639663 77888
rect 637132 77830 639663 77832
rect 637132 77828 637138 77830
rect 639597 77827 639663 77830
rect 578693 75442 578759 75445
rect 575798 75440 578759 75442
rect 575798 75384 578698 75440
rect 578754 75384 578759 75440
rect 575798 75382 578759 75384
rect 575798 75140 575858 75382
rect 578693 75379 578759 75382
rect 647049 74490 647115 74493
rect 646668 74488 647115 74490
rect 646668 74432 647054 74488
rect 647110 74432 647115 74488
rect 646668 74430 647115 74432
rect 647049 74427 647115 74430
rect 578509 73130 578575 73133
rect 575798 73128 578575 73130
rect 575798 73072 578514 73128
rect 578570 73072 578575 73128
rect 575798 73070 578575 73072
rect 575798 72964 575858 73070
rect 578509 73067 578575 73070
rect 646865 72994 646931 72997
rect 646668 72992 646931 72994
rect 646668 72936 646870 72992
rect 646926 72936 646931 72992
rect 646668 72934 646931 72936
rect 646865 72931 646931 72934
rect 648981 71498 649047 71501
rect 646668 71496 649047 71498
rect 646668 71440 648986 71496
rect 649042 71440 649047 71496
rect 646668 71438 649047 71440
rect 648981 71435 649047 71438
rect 579153 71362 579219 71365
rect 575798 71360 579219 71362
rect 575798 71304 579158 71360
rect 579214 71304 579219 71360
rect 575798 71302 579219 71304
rect 575798 70788 575858 71302
rect 579153 71299 579219 71302
rect 647325 70002 647391 70005
rect 646668 70000 647391 70002
rect 646668 69944 647330 70000
rect 647386 69944 647391 70000
rect 646668 69942 647391 69944
rect 647325 69939 647391 69942
rect 646221 68914 646287 68917
rect 646221 68912 646330 68914
rect 646221 68856 646226 68912
rect 646282 68856 646330 68912
rect 646221 68851 646330 68856
rect 575982 68098 576042 68612
rect 646270 68476 646330 68851
rect 579521 68098 579587 68101
rect 575982 68096 579587 68098
rect 575982 68040 579526 68096
rect 579582 68040 579587 68096
rect 575982 68038 579587 68040
rect 579521 68035 579587 68038
rect 649165 67010 649231 67013
rect 646668 67008 649231 67010
rect 646668 66952 649170 67008
rect 649226 66952 649231 67008
rect 646668 66950 649231 66952
rect 649165 66947 649231 66950
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 647509 65514 647575 65517
rect 646668 65512 647575 65514
rect 646668 65456 647514 65512
rect 647570 65456 647575 65512
rect 646668 65454 647575 65456
rect 647509 65451 647575 65454
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 646086 63988 646146 64363
rect 575982 61842 576042 62084
rect 578509 61842 578575 61845
rect 575982 61840 578575 61842
rect 575982 61784 578514 61840
rect 578570 61784 578575 61840
rect 575982 61782 578575 61784
rect 578509 61779 578575 61782
rect 579521 60346 579587 60349
rect 575798 60344 579587 60346
rect 575798 60288 579526 60344
rect 579582 60288 579587 60344
rect 575798 60286 579587 60288
rect 575798 59908 575858 60286
rect 579521 60283 579587 60286
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 579521 56130 579587 56133
rect 575798 56128 579587 56130
rect 575798 56072 579526 56128
rect 579582 56072 579587 56128
rect 575798 56070 579587 56072
rect 575798 55556 575858 56070
rect 579521 56067 579587 56070
rect 461710 54980 461716 55044
rect 461780 55042 461786 55044
rect 581637 55042 581703 55045
rect 461780 55040 581703 55042
rect 461780 54984 581642 55040
rect 581698 54984 581703 55040
rect 461780 54982 581703 54984
rect 461780 54980 461786 54982
rect 581637 54979 581703 54982
rect 580257 54770 580323 54773
rect 460798 54768 580323 54770
rect 460798 54712 580262 54768
rect 580318 54712 580323 54768
rect 460798 54710 580323 54712
rect 460798 53685 460858 54710
rect 580257 54707 580323 54710
rect 594057 54498 594123 54501
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 460982 54496 594123 54498
rect 460982 54440 594062 54496
rect 594118 54440 594123 54496
rect 460982 54438 594123 54440
rect 460749 53619 460815 53622
rect 459921 53410 459987 53413
rect 460982 53410 461042 54438
rect 594057 54435 594123 54438
rect 577681 54226 577747 54229
rect 466410 54224 577747 54226
rect 466410 54168 577686 54224
rect 577742 54168 577747 54224
rect 466410 54166 577747 54168
rect 461710 53892 461716 53956
rect 461780 53892 461786 53956
rect 466410 53954 466470 54166
rect 577681 54163 577747 54166
rect 462638 53894 466470 53954
rect 461718 53685 461778 53892
rect 462638 53685 462698 53894
rect 461669 53680 461778 53685
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462589 53680 462698 53685
rect 462589 53624 462594 53680
rect 462650 53624 462698 53680
rect 462589 53622 462698 53624
rect 463693 53682 463759 53685
rect 472249 53682 472315 53685
rect 463693 53680 472315 53682
rect 463693 53624 463698 53680
rect 463754 53624 472254 53680
rect 472310 53624 472315 53680
rect 463693 53622 472315 53624
rect 461669 53619 461735 53622
rect 462589 53619 462655 53622
rect 463693 53619 463759 53622
rect 472249 53619 472315 53622
rect 459921 53408 461042 53410
rect 459921 53352 459926 53408
rect 459982 53352 461042 53408
rect 459921 53350 461042 53352
rect 459921 53347 459987 53350
rect 462957 53274 463023 53277
rect 471881 53274 471947 53277
rect 462957 53272 471947 53274
rect 462957 53216 462962 53272
rect 463018 53216 471886 53272
rect 471942 53216 471947 53272
rect 462957 53214 471947 53216
rect 462957 53211 463023 53214
rect 471881 53211 471947 53214
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 308990 49676 308996 49740
rect 309060 49738 309066 49740
rect 309685 49738 309751 49741
rect 309060 49736 309751 49738
rect 309060 49680 309690 49736
rect 309746 49680 309751 49736
rect 309060 49678 309751 49680
rect 309060 49676 309066 49678
rect 309685 49675 309751 49678
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 663977 48514 664043 48517
rect 662094 48512 664043 48514
rect 661480 48456 663982 48512
rect 664038 48456 664043 48512
rect 661480 48454 664043 48456
rect 661480 48452 662154 48454
rect 663977 48451 664043 48454
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 663793 47834 663859 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661910 47832 663859 47834
rect 661910 47791 663798 47832
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47776 663798 47791
rect 663854 47776 663859 47832
rect 661388 47774 663859 47776
rect 661388 47731 661970 47774
rect 663793 47771 663859 47774
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 461342 44372 461348 44436
rect 461412 44434 461418 44436
rect 461945 44434 462011 44437
rect 461412 44432 462011 44434
rect 461412 44376 461950 44432
rect 462006 44376 462011 44432
rect 461412 44374 462011 44376
rect 461412 44372 461418 44374
rect 461945 44371 462011 44374
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462497 44434 462563 44437
rect 462332 44432 462563 44434
rect 462332 44376 462502 44432
rect 462558 44376 462563 44432
rect 462332 44374 462563 44376
rect 462332 44372 462338 44374
rect 462497 44371 462563 44374
rect 310421 44162 310487 44165
rect 364885 44162 364951 44165
rect 463693 44162 463759 44165
rect 310421 44160 354690 44162
rect 310421 44104 310426 44160
rect 310482 44104 354690 44160
rect 310421 44102 354690 44104
rect 310421 44099 310487 44102
rect 354630 43890 354690 44102
rect 364885 44160 463759 44162
rect 364885 44104 364890 44160
rect 364946 44104 463698 44160
rect 463754 44104 463759 44160
rect 364885 44102 463759 44104
rect 364885 44099 364951 44102
rect 463693 44099 463759 44102
rect 440182 43890 440188 43892
rect 354630 43830 440188 43890
rect 440182 43828 440188 43830
rect 440252 43828 440258 43892
rect 440918 43828 440924 43892
rect 440988 43890 440994 43892
rect 462957 43890 463023 43893
rect 440988 43888 463023 43890
rect 440988 43832 462962 43888
rect 463018 43832 463023 43888
rect 440988 43830 463023 43832
rect 440988 43828 440994 43830
rect 462957 43827 463023 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463693 42938 463759 42941
rect 461761 42936 463759 42938
rect 461761 42880 461766 42936
rect 461822 42880 463698 42936
rect 463754 42880 463759 42936
rect 461761 42878 463759 42880
rect 461761 42875 461827 42878
rect 463693 42875 463759 42878
rect 308949 42804 309015 42805
rect 518801 42804 518867 42805
rect 308949 42800 308996 42804
rect 309060 42802 309066 42804
rect 518750 42802 518756 42804
rect 308949 42744 308954 42800
rect 308949 42740 308996 42744
rect 309060 42742 309106 42802
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 309060 42740 309066 42742
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 308949 42739 309015 42740
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 443545 42258 443611 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 443545 42256 461183 42258
rect 443545 42200 443550 42256
rect 443606 42200 461122 42256
rect 461178 42200 461183 42256
rect 443545 42198 461183 42200
rect 443545 42195 443611 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 443545 41578 443611 41581
rect 427770 41576 443611 41578
rect 427770 41520 443550 41576
rect 443606 41520 443611 41576
rect 427770 41518 443611 41520
rect 443545 41515 443611 41518
rect 141693 40490 141759 40493
rect 142613 40490 142679 40493
rect 141693 40488 142679 40490
rect 141693 40432 141698 40488
rect 141754 40432 142618 40488
rect 142674 40432 142679 40488
rect 141693 40430 142679 40432
rect 141693 40427 141759 40430
rect 142613 40427 142679 40430
<< via3 >>
rect 192524 997188 192588 997252
rect 388116 997188 388180 997252
rect 504588 997732 504652 997796
rect 476436 997188 476500 997252
rect 529060 997188 529124 997252
rect 89852 996916 89916 996980
rect 140268 996508 140332 996572
rect 183692 996372 183756 996436
rect 89852 995420 89916 995484
rect 140268 995420 140332 995484
rect 187924 995828 187988 995892
rect 238524 996372 238588 996436
rect 191788 995752 191852 995756
rect 191788 995696 191802 995752
rect 191802 995696 191852 995752
rect 191788 995692 191852 995696
rect 192524 995752 192588 995756
rect 192524 995696 192538 995752
rect 192538 995696 192588 995752
rect 192524 995692 192588 995696
rect 183692 995344 183756 995348
rect 183692 995288 183706 995344
rect 183706 995288 183756 995344
rect 183692 995284 183756 995288
rect 188476 995284 188540 995348
rect 238524 995344 238588 995348
rect 238524 995288 238574 995344
rect 238574 995288 238588 995344
rect 238524 995284 238588 995288
rect 630812 996916 630876 996980
rect 291332 996644 291396 996708
rect 384988 996644 385052 996708
rect 476804 996644 476868 996708
rect 629708 996644 629772 996708
rect 481220 996372 481284 996436
rect 291332 995344 291396 995348
rect 291332 995288 291382 995344
rect 291382 995288 291396 995344
rect 291332 995284 291396 995288
rect 384988 995752 385052 995756
rect 384988 995696 385038 995752
rect 385038 995696 385052 995752
rect 384988 995692 385052 995696
rect 388116 995480 388180 995484
rect 388116 995424 388166 995480
rect 388166 995424 388180 995480
rect 388116 995420 388180 995424
rect 485636 995752 485700 995756
rect 485636 995696 485650 995752
rect 485650 995696 485700 995752
rect 485636 995692 485700 995696
rect 481220 995616 481284 995620
rect 503668 995828 503732 995892
rect 481220 995560 481270 995616
rect 481270 995560 481284 995616
rect 481220 995556 481284 995560
rect 476436 995344 476500 995348
rect 476436 995288 476486 995344
rect 476486 995288 476500 995344
rect 476436 995284 476500 995288
rect 476804 995284 476868 995348
rect 529060 995752 529124 995756
rect 529060 995696 529110 995752
rect 529110 995696 529124 995752
rect 529060 995692 529124 995696
rect 533476 995752 533540 995756
rect 533476 995696 533526 995752
rect 533526 995696 533540 995752
rect 533476 995692 533540 995696
rect 629708 995752 629772 995756
rect 629708 995696 629758 995752
rect 629758 995696 629772 995752
rect 629708 995692 629772 995696
rect 630812 995752 630876 995756
rect 630812 995696 630862 995752
rect 630862 995696 630876 995752
rect 630812 995692 630876 995696
rect 243308 994528 243372 994532
rect 243308 994472 243322 994528
rect 243322 994472 243372 994528
rect 243308 994468 243372 994472
rect 226380 994196 226444 994260
rect 278636 994196 278700 994260
rect 41460 967132 41524 967196
rect 675708 966512 675772 966516
rect 675708 966456 675722 966512
rect 675722 966456 675772 966512
rect 675708 966452 675772 966456
rect 676076 965092 676140 965156
rect 676812 964684 676876 964748
rect 675524 963384 675588 963388
rect 675524 963328 675538 963384
rect 675538 963328 675588 963384
rect 675524 963324 675588 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 41276 959788 41340 959852
rect 40540 959108 40604 959172
rect 675524 959108 675588 959172
rect 41828 957808 41892 957812
rect 41828 957752 41842 957808
rect 41842 957752 41892 957808
rect 41828 957748 41892 957752
rect 676628 957748 676692 957812
rect 676996 956388 677060 956452
rect 40724 955436 40788 955500
rect 675708 954620 675772 954684
rect 41828 952852 41892 952916
rect 41460 952444 41524 952508
rect 41644 952172 41708 952236
rect 41276 951628 41340 951692
rect 676812 950676 676876 950740
rect 676076 949452 676140 949516
rect 39804 943800 39868 943804
rect 39804 943744 39818 943800
rect 39818 943744 39868 943800
rect 39804 943740 39868 943744
rect 40724 943740 40788 943804
rect 42012 943740 42076 943804
rect 41782 939388 41846 939452
rect 674604 938028 674668 938092
rect 674972 937620 675036 937684
rect 41828 936532 41892 936596
rect 676996 931908 677060 931972
rect 676628 931500 676692 931564
rect 42012 911916 42076 911980
rect 42196 911644 42260 911708
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 676076 875876 676140 875940
rect 675892 873972 675956 874036
rect 676812 871932 676876 871996
rect 673868 869484 673932 869548
rect 674420 854312 674484 854316
rect 674420 854256 674470 854312
rect 674470 854256 674484 854312
rect 674420 854252 674484 854256
rect 39988 814234 40052 814298
rect 41828 813180 41892 813244
rect 40908 805428 40972 805492
rect 40540 805352 40604 805356
rect 40540 805296 40590 805352
rect 40590 805296 40604 805352
rect 40540 805292 40604 805296
rect 40724 805080 40788 805084
rect 40724 805024 40774 805080
rect 40774 805024 40788 805080
rect 40724 805020 40788 805024
rect 42012 804748 42076 804812
rect 41644 804476 41708 804540
rect 40724 794956 40788 795020
rect 40908 794140 40972 794204
rect 40540 792508 40604 792572
rect 41644 788972 41708 789036
rect 41828 788624 41892 788628
rect 41828 788568 41842 788624
rect 41842 788568 41892 788624
rect 41828 788564 41892 788568
rect 41460 788156 41524 788220
rect 674788 787264 674852 787268
rect 674788 787208 674838 787264
rect 674838 787208 674852 787264
rect 674788 787204 674852 787208
rect 674972 786660 675036 786724
rect 674972 783320 675036 783324
rect 674972 783264 674986 783320
rect 674986 783264 675036 783320
rect 674972 783260 675036 783264
rect 674788 782716 674852 782780
rect 676996 780540 677060 780604
rect 675892 772652 675956 772716
rect 41460 769796 41524 769860
rect 676076 768708 676140 768772
rect 675892 766532 675956 766596
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 676076 765036 676140 765100
rect 40724 764900 40788 764964
rect 41644 764492 41708 764556
rect 676996 761832 677060 761836
rect 676628 761788 676692 761792
rect 676628 761732 676642 761788
rect 676642 761732 676692 761788
rect 676628 761728 676692 761732
rect 676996 761776 677010 761832
rect 677010 761776 677060 761832
rect 676996 761772 677060 761776
rect 41828 757692 41892 757756
rect 40356 757284 40420 757348
rect 42012 756332 42076 756396
rect 673868 754700 673932 754764
rect 40356 754428 40420 754492
rect 42012 754080 42076 754084
rect 42012 754024 42026 754080
rect 42026 754024 42076 754080
rect 42012 754020 42076 754024
rect 674420 753748 674484 753812
rect 40724 752116 40788 752180
rect 40908 751028 40972 751092
rect 40540 749396 40604 749460
rect 41644 745044 41708 745108
rect 41828 744772 41892 744836
rect 41460 743684 41524 743748
rect 674420 741508 674484 741572
rect 674604 738108 674668 738172
rect 670740 734088 670804 734092
rect 670740 734032 670754 734088
rect 670754 734032 670804 734088
rect 670740 734028 670804 734032
rect 674236 732804 674300 732868
rect 675892 728724 675956 728788
rect 676812 728724 676876 728788
rect 670740 728512 670804 728516
rect 670740 728456 670754 728512
rect 670754 728456 670804 728512
rect 670740 728452 670804 728456
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 40356 721708 40420 721772
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 718524 40604 718588
rect 40356 716756 40420 716820
rect 40908 716756 40972 716820
rect 41828 714716 41892 714780
rect 42012 714640 42076 714644
rect 42012 714584 42026 714640
rect 42026 714584 42076 714640
rect 42012 714580 42076 714584
rect 675892 711996 675956 712060
rect 42012 709880 42076 709884
rect 42012 709824 42026 709880
rect 42026 709824 42076 709880
rect 42012 709820 42076 709824
rect 40908 708460 40972 708524
rect 40724 706692 40788 706756
rect 673316 705060 673380 705124
rect 40540 704244 40604 704308
rect 41828 701796 41892 701860
rect 41644 701524 41708 701588
rect 41460 700436 41524 700500
rect 676996 694044 677060 694108
rect 674788 689692 674852 689756
rect 674788 688800 674852 688804
rect 674788 688744 674802 688800
rect 674802 688744 674852 688800
rect 674788 688740 674852 688744
rect 42196 683572 42260 683636
rect 42012 682756 42076 682820
rect 674420 682348 674484 682412
rect 674236 680988 674300 681052
rect 40540 678928 40604 678992
rect 40908 678928 40972 678992
rect 41828 678268 41892 678332
rect 41828 677588 41892 677652
rect 42196 677588 42260 677652
rect 40356 671196 40420 671260
rect 41828 670924 41892 670988
rect 42196 669292 42260 669356
rect 42196 667856 42260 667860
rect 42196 667800 42246 667856
rect 42246 667800 42260 667856
rect 42196 667796 42260 667800
rect 40356 667524 40420 667588
rect 40908 666980 40972 667044
rect 42012 666980 42076 667044
rect 674420 666300 674484 666364
rect 673500 665756 673564 665820
rect 673684 665620 673748 665684
rect 40724 665348 40788 665412
rect 673684 665076 673748 665140
rect 674420 665076 674484 665140
rect 673684 664260 673748 664324
rect 42012 664048 42076 664052
rect 42012 663992 42026 664048
rect 42026 663992 42076 664048
rect 42012 663988 42076 663992
rect 40540 662628 40604 662692
rect 674604 662220 674668 662284
rect 41644 658548 41708 658612
rect 41828 658276 41892 658340
rect 41460 657188 41524 657252
rect 675340 652896 675404 652900
rect 675340 652840 675390 652896
rect 675390 652840 675404 652896
rect 675340 652836 675404 652840
rect 675524 651536 675588 651540
rect 675524 651480 675538 651536
rect 675538 651480 675588 651536
rect 675524 651476 675588 651480
rect 674236 648892 674300 648956
rect 674604 645084 674668 645148
rect 676812 644676 676876 644740
rect 41460 640596 41524 640660
rect 675156 640460 675220 640524
rect 41828 639168 41892 639232
rect 41644 638556 41708 638620
rect 675340 638012 675404 638076
rect 675524 637800 675588 637804
rect 675524 637744 675574 637800
rect 675574 637744 675588 637800
rect 675524 637740 675588 637744
rect 675156 637664 675220 637668
rect 675156 637608 675206 637664
rect 675206 637608 675220 637664
rect 675156 637604 675220 637608
rect 40540 634884 40604 634948
rect 675156 632980 675220 633044
rect 676076 631348 676140 631412
rect 675524 629716 675588 629780
rect 42012 626588 42076 626652
rect 42196 625016 42260 625020
rect 42196 624960 42246 625016
rect 42246 624960 42260 625016
rect 42196 624956 42260 624960
rect 42012 624472 42076 624476
rect 42012 624416 42062 624472
rect 42062 624416 42076 624472
rect 42012 624412 42076 624416
rect 40540 622100 40604 622164
rect 42196 620196 42260 620260
rect 676996 619108 677060 619172
rect 41460 615980 41524 616044
rect 41828 615768 41892 615772
rect 41828 615712 41842 615768
rect 41842 615712 41892 615768
rect 41828 615708 41892 615712
rect 41828 612776 41892 612780
rect 41828 612720 41842 612776
rect 41842 612720 41892 612776
rect 41828 612716 41892 612720
rect 674420 602924 674484 602988
rect 42012 597212 42076 597276
rect 675708 596668 675772 596732
rect 41828 596396 41892 596460
rect 676996 594084 677060 594148
rect 675524 593812 675588 593876
rect 675156 592860 675220 592924
rect 674236 592588 674300 592652
rect 41828 592316 41892 592380
rect 675708 592316 675772 592380
rect 43852 591500 43916 591564
rect 676076 590548 676140 590612
rect 40540 589656 40604 589660
rect 40540 589600 40554 589656
rect 40554 589600 40604 589656
rect 40540 589596 40604 589600
rect 41276 589596 41340 589660
rect 41828 589596 41892 589660
rect 40908 589324 40972 589388
rect 40356 585924 40420 585988
rect 41828 585652 41892 585716
rect 42380 585244 42444 585308
rect 41092 584564 41156 584628
rect 42012 584564 42076 584628
rect 40356 582524 40420 582588
rect 40908 580620 40972 580684
rect 41092 580212 41156 580276
rect 40724 579940 40788 580004
rect 40540 576812 40604 576876
rect 42196 576540 42260 576604
rect 676996 576404 677060 576468
rect 42012 573200 42076 573204
rect 42012 573144 42026 573200
rect 42026 573144 42076 573200
rect 42012 573140 42076 573144
rect 676812 572732 676876 572796
rect 41460 571644 41524 571708
rect 41828 571372 41892 571436
rect 41644 570964 41708 571028
rect 675524 562728 675588 562732
rect 675524 562672 675538 562728
rect 675538 562672 675588 562728
rect 675524 562668 675588 562672
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676260 557636 676324 557700
rect 676812 553964 676876 554028
rect 41828 553208 41892 553212
rect 41828 553152 41842 553208
rect 41842 553152 41892 553208
rect 41828 553148 41892 553152
rect 41828 552740 41892 552804
rect 675892 550428 675956 550492
rect 676996 550156 677060 550220
rect 675892 547632 675956 547636
rect 675892 547576 675942 547632
rect 675942 547576 675956 547632
rect 675892 547572 675956 547576
rect 676260 547572 676324 547636
rect 41644 546348 41708 546412
rect 40724 545668 40788 545732
rect 40540 545396 40604 545460
rect 675340 544912 675404 544916
rect 675340 544856 675354 544912
rect 675354 544856 675404 544912
rect 675340 544852 675404 544856
rect 675524 544444 675588 544508
rect 40724 538188 40788 538252
rect 40540 534924 40604 534988
rect 674420 533836 674484 533900
rect 41460 530572 41524 530636
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 41644 529076 41708 529140
rect 676996 503644 677060 503708
rect 676812 503372 676876 503436
rect 675892 488820 675956 488884
rect 674604 475356 674668 475420
rect 673316 474872 673380 474876
rect 673316 474816 673330 474872
rect 673330 474816 673380 474872
rect 673316 474812 673380 474816
rect 675340 453732 675404 453796
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 41644 418780 41708 418844
rect 40540 418704 40604 418708
rect 40540 418648 40554 418704
rect 40554 418648 40604 418704
rect 40540 418644 40604 418648
rect 40724 418508 40788 418572
rect 675340 410484 675404 410548
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 41460 401780 41524 401844
rect 676812 401236 676876 401300
rect 41828 398848 41892 398852
rect 41828 398792 41842 398848
rect 41842 398792 41892 398848
rect 41828 398788 41892 398792
rect 675892 398788 675956 398852
rect 676628 396748 676692 396812
rect 676260 395116 676324 395180
rect 676444 394708 676508 394772
rect 676076 393076 676140 393140
rect 675708 387636 675772 387700
rect 676628 384916 676692 384980
rect 41460 381788 41524 381852
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 41828 378524 41892 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 40908 377708 40972 377772
rect 676260 377300 676324 377364
rect 41644 376484 41708 376548
rect 40356 375668 40420 375732
rect 675892 374988 675956 375052
rect 676076 372948 676140 373012
rect 674788 372540 674852 372604
rect 40356 368596 40420 368660
rect 40908 364244 40972 364308
rect 40724 363564 40788 363628
rect 41828 362944 41892 362948
rect 41828 362888 41842 362944
rect 41842 362888 41892 362944
rect 41828 362884 41892 362888
rect 40540 360028 40604 360092
rect 41460 358668 41524 358732
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43852 354240 43916 354244
rect 43852 354184 43902 354240
rect 43902 354184 43916 354240
rect 43852 354180 43916 354184
rect 675340 354180 675404 354244
rect 44220 353772 44284 353836
rect 675524 352956 675588 353020
rect 675892 351868 675956 351932
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675892 349208 675956 349212
rect 675892 349152 675942 349208
rect 675942 349152 675956 349208
rect 675892 349148 675956 349152
rect 44404 342892 44468 342956
rect 44220 342620 44284 342684
rect 44404 342076 44468 342140
rect 43668 340444 43732 340508
rect 676628 340172 676692 340236
rect 675340 339008 675404 339012
rect 675340 338952 675390 339008
rect 675390 338952 675404 339008
rect 675340 338948 675404 338952
rect 41460 337724 41524 337788
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 42932 337452 42996 337516
rect 43116 337180 43180 337244
rect 676444 336636 676508 336700
rect 40540 336500 40604 336564
rect 43300 336364 43364 336428
rect 41828 336092 41892 336156
rect 42748 335684 42812 335748
rect 40724 335276 40788 335340
rect 42748 334596 42812 334660
rect 43300 334596 43364 334660
rect 40908 333644 40972 333708
rect 676260 332284 676324 332348
rect 41644 328340 41708 328404
rect 676076 328340 676140 328404
rect 41460 326708 41524 326772
rect 40908 325348 40972 325412
rect 41460 324804 41524 324868
rect 40724 317460 40788 317524
rect 40540 316644 40604 316708
rect 43116 315964 43180 316028
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 42932 312700 42996 312764
rect 44588 311476 44652 311540
rect 44404 311264 44468 311268
rect 44404 311208 44418 311264
rect 44418 311208 44468 311264
rect 44404 311204 44468 311208
rect 675708 308756 675772 308820
rect 675892 306716 675956 306780
rect 675892 302636 675956 302700
rect 676444 301608 676508 301612
rect 676444 301552 676494 301608
rect 676494 301552 676508 301608
rect 676444 301548 676508 301552
rect 676628 301472 676692 301476
rect 676628 301416 676678 301472
rect 676678 301416 676692 301472
rect 676628 301412 676692 301416
rect 675708 298012 675772 298076
rect 43668 297604 43732 297668
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676260 295156 676324 295220
rect 40540 292528 40604 292592
rect 40908 292528 40972 292592
rect 41828 292496 41892 292500
rect 41828 292440 41842 292496
rect 41842 292440 41892 292496
rect 41828 292436 41892 292440
rect 676444 291484 676508 291548
rect 41828 290456 41892 290460
rect 41828 290400 41842 290456
rect 41842 290400 41892 290456
rect 41828 290396 41892 290400
rect 676628 286996 676692 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 40724 278428 40788 278492
rect 40908 277884 40972 277948
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 674972 263604 675036 263668
rect 676076 262380 676140 262444
rect 676996 261564 677060 261628
rect 676812 259932 676876 259996
rect 40724 251364 40788 251428
rect 676996 250276 677060 250340
rect 676076 249868 676140 249932
rect 40540 249732 40604 249796
rect 674788 249596 674852 249660
rect 674788 245516 674852 245580
rect 675892 245516 675956 245580
rect 676812 245516 676876 245580
rect 675340 245244 675404 245308
rect 675892 242252 675956 242316
rect 675340 240272 675404 240276
rect 675340 240216 675390 240272
rect 675390 240216 675404 240272
rect 675340 240212 675404 240216
rect 40724 240076 40788 240140
rect 673316 239940 673380 240004
rect 42012 237356 42076 237420
rect 674788 237220 674852 237284
rect 674052 237084 674116 237148
rect 40540 235860 40604 235924
rect 673316 235180 673380 235244
rect 671292 233140 671356 233204
rect 669268 231372 669332 231436
rect 673316 228924 673380 228988
rect 669452 228788 669516 228852
rect 672948 228576 673012 228580
rect 672948 228520 672962 228576
rect 672962 228520 673012 228576
rect 672948 228516 673012 228520
rect 674788 228516 674852 228580
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 671108 227156 671172 227220
rect 671660 226748 671724 226812
rect 673132 226748 673196 226812
rect 671844 226672 671908 226676
rect 671844 226616 671894 226672
rect 671894 226616 671908 226672
rect 671844 226612 671908 226616
rect 672028 226536 672092 226540
rect 672028 226480 672032 226536
rect 672032 226480 672088 226536
rect 672088 226480 672092 226536
rect 672028 226476 672092 226480
rect 675156 226476 675220 226540
rect 673684 226204 673748 226268
rect 671844 225116 671908 225180
rect 673316 224844 673380 224908
rect 671660 224164 671724 224228
rect 671108 223892 671172 223956
rect 673500 223620 673564 223684
rect 562364 222048 562428 222052
rect 562364 221992 562378 222048
rect 562378 221992 562428 222048
rect 562364 221988 562428 221992
rect 564572 221988 564636 222052
rect 572852 221988 572916 222052
rect 572852 220628 572916 220692
rect 572116 220356 572180 220420
rect 578188 220416 578252 220420
rect 578188 220360 578238 220416
rect 578238 220360 578252 220416
rect 578188 220356 578252 220360
rect 573956 220280 574020 220284
rect 573956 220224 573970 220280
rect 573970 220224 574020 220280
rect 573956 220220 574020 220224
rect 487476 219328 487540 219332
rect 487476 219272 487490 219328
rect 487490 219272 487540 219328
rect 487476 219268 487540 219272
rect 491156 218648 491220 218652
rect 491156 218592 491206 218648
rect 491206 218592 491220 218648
rect 491156 218588 491220 218592
rect 674788 218860 674852 218924
rect 673132 218588 673196 218652
rect 675524 218588 675588 218652
rect 572116 218316 572180 218380
rect 676030 218180 676094 218244
rect 672028 217772 672092 217836
rect 592356 217500 592420 217564
rect 488948 217288 489012 217292
rect 488948 217232 488962 217288
rect 488962 217232 489012 217288
rect 488948 217228 489012 217232
rect 591988 217228 592052 217292
rect 675892 216956 675956 217020
rect 675156 215460 675220 215524
rect 675708 215324 675772 215388
rect 676260 215086 676324 215150
rect 575612 213148 575676 213212
rect 667980 212332 668044 212396
rect 676444 211380 676508 211444
rect 673132 210428 673196 210492
rect 675524 210428 675588 210492
rect 675892 210428 675956 210492
rect 42012 210020 42076 210084
rect 40724 208116 40788 208180
rect 41644 207708 41708 207772
rect 40908 207300 40972 207364
rect 40540 206892 40604 206956
rect 676628 205532 676692 205596
rect 673316 202948 673380 203012
rect 676444 200772 676508 200836
rect 41828 197780 41892 197844
rect 40724 197100 40788 197164
rect 676260 197100 676324 197164
rect 41828 195800 41892 195804
rect 41828 195744 41878 195800
rect 41878 195744 41892 195800
rect 41828 195740 41892 195744
rect 40908 195468 40972 195532
rect 42012 195256 42076 195260
rect 42012 195200 42026 195256
rect 42026 195200 42076 195256
rect 42012 195196 42076 195200
rect 675708 195256 675772 195260
rect 675708 195200 675722 195256
rect 675722 195200 675772 195256
rect 675708 195196 675772 195200
rect 40540 194516 40604 194580
rect 41460 194516 41524 194580
rect 675892 193156 675956 193220
rect 42380 192884 42444 192948
rect 676076 191524 676140 191588
rect 41460 187172 41524 187236
rect 42380 186280 42444 186284
rect 42380 186224 42394 186280
rect 42394 186224 42444 186280
rect 42380 186220 42444 186224
rect 41828 185872 41892 185876
rect 41828 185816 41842 185872
rect 41842 185816 41892 185872
rect 41828 185812 41892 185816
rect 672948 183500 673012 183564
rect 673132 182004 673196 182068
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675708 170308 675772 170372
rect 675892 167452 675956 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 675524 161332 675588 161396
rect 676444 159428 676508 159492
rect 675524 157040 675588 157044
rect 675524 156984 675574 157040
rect 675574 156984 675588 157040
rect 675524 156980 675588 156984
rect 676628 156300 676692 156364
rect 674052 154532 674116 154596
rect 676260 153036 676324 153100
rect 675708 150376 675772 150380
rect 675708 150320 675758 150376
rect 675758 150320 675772 150376
rect 675708 150316 675772 150320
rect 676076 148412 676140 148476
rect 673316 147732 673380 147796
rect 675892 147596 675956 147660
rect 671292 145148 671356 145212
rect 673684 143516 673748 143580
rect 667980 130460 668044 130524
rect 676628 128556 676692 128620
rect 673500 128420 673564 128484
rect 676076 128148 676140 128212
rect 675892 127196 675956 127260
rect 676260 126924 676324 126988
rect 676444 124476 676508 124540
rect 675708 122300 675772 122364
rect 676628 113052 676692 113116
rect 675892 108020 675956 108084
rect 676444 106116 676508 106180
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676260 101356 676324 101420
rect 634860 96868 634924 96932
rect 637252 96868 637316 96932
rect 634860 80412 634924 80476
rect 637068 77828 637132 77892
rect 461716 54980 461780 55044
rect 461716 53892 461780 53956
rect 194364 50220 194428 50284
rect 308996 49676 309060 49740
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 461348 44372 461412 44436
rect 462268 44372 462332 44436
rect 440188 43828 440252 43892
rect 440924 43828 440988 43892
rect 308996 42800 309060 42804
rect 308996 42744 309010 42800
rect 309010 42744 309060 42800
rect 308996 42740 309060 42744
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
<< metal4 >>
rect 504587 997796 504653 997797
rect 504587 997732 504588 997796
rect 504652 997732 504653 997796
rect 504587 997731 504653 997732
rect 192523 997252 192589 997253
rect 192523 997188 192524 997252
rect 192588 997188 192589 997252
rect 192523 997187 192589 997188
rect 89851 996980 89917 996981
rect 89851 996916 89852 996980
rect 89916 996916 89917 996980
rect 89851 996915 89917 996916
rect 89854 995485 89914 996915
rect 140267 996572 140333 996573
rect 140267 996508 140268 996572
rect 140332 996508 140333 996572
rect 140267 996507 140333 996508
rect 140270 995485 140330 996507
rect 183691 996436 183757 996437
rect 183691 996372 183692 996436
rect 183756 996372 183757 996436
rect 183691 996371 183757 996372
rect 89851 995484 89917 995485
rect 89851 995420 89852 995484
rect 89916 995420 89917 995484
rect 89851 995419 89917 995420
rect 140267 995484 140333 995485
rect 140267 995420 140268 995484
rect 140332 995420 140333 995484
rect 140267 995419 140333 995420
rect 183694 995349 183754 996371
rect 187923 995892 187989 995893
rect 187923 995828 187924 995892
rect 187988 995890 187989 995892
rect 187988 995830 188538 995890
rect 187988 995828 187989 995830
rect 187923 995827 187989 995828
rect 188478 995349 188538 995830
rect 191790 995757 191850 997102
rect 192526 995757 192586 997187
rect 388115 997252 388181 997253
rect 388115 997188 388116 997252
rect 388180 997188 388181 997252
rect 388115 997187 388181 997188
rect 476435 997252 476501 997253
rect 476435 997188 476436 997252
rect 476500 997188 476501 997252
rect 476435 997187 476501 997188
rect 191787 995756 191853 995757
rect 191787 995692 191788 995756
rect 191852 995692 191853 995756
rect 191787 995691 191853 995692
rect 192523 995756 192589 995757
rect 192523 995692 192524 995756
rect 192588 995692 192589 995756
rect 192523 995691 192589 995692
rect 183691 995348 183757 995349
rect 183691 995284 183692 995348
rect 183756 995284 183757 995348
rect 183691 995283 183757 995284
rect 188475 995348 188541 995349
rect 188475 995284 188476 995348
rect 188540 995284 188541 995348
rect 188475 995283 188541 995284
rect 226382 994261 226442 997102
rect 238523 996436 238589 996437
rect 238523 996372 238524 996436
rect 238588 996372 238589 996436
rect 238523 996371 238589 996372
rect 238526 995349 238586 996371
rect 238523 995348 238589 995349
rect 238523 995284 238524 995348
rect 238588 995284 238589 995348
rect 238523 995283 238589 995284
rect 243310 994533 243370 997102
rect 243307 994532 243373 994533
rect 243307 994468 243308 994532
rect 243372 994468 243373 994532
rect 243307 994467 243373 994468
rect 278638 994261 278698 997102
rect 291331 996708 291397 996709
rect 291331 996644 291332 996708
rect 291396 996644 291397 996708
rect 291331 996643 291397 996644
rect 384987 996708 385053 996709
rect 384987 996644 384988 996708
rect 385052 996644 385053 996708
rect 384987 996643 385053 996644
rect 291334 995349 291394 996643
rect 384990 995757 385050 996643
rect 384987 995756 385053 995757
rect 384987 995692 384988 995756
rect 385052 995692 385053 995756
rect 384987 995691 385053 995692
rect 388118 995485 388178 997187
rect 388115 995484 388181 995485
rect 388115 995420 388116 995484
rect 388180 995420 388181 995484
rect 388115 995419 388181 995420
rect 476438 995349 476498 997187
rect 504590 997250 504650 997731
rect 504590 997190 505238 997250
rect 529059 997252 529125 997253
rect 529059 997188 529060 997252
rect 529124 997188 529125 997252
rect 529059 997187 529125 997188
rect 476803 996708 476869 996709
rect 476803 996644 476804 996708
rect 476868 996644 476869 996708
rect 476803 996643 476869 996644
rect 476806 995349 476866 996643
rect 481219 996436 481285 996437
rect 481219 996372 481220 996436
rect 481284 996372 481285 996436
rect 481219 996371 481285 996372
rect 481222 995621 481282 996371
rect 485638 995757 485698 997102
rect 503670 995893 503730 997102
rect 503667 995892 503733 995893
rect 503667 995828 503668 995892
rect 503732 995828 503733 995892
rect 503667 995827 503733 995828
rect 529062 995757 529122 997187
rect 533478 995757 533538 997102
rect 630811 996980 630877 996981
rect 630811 996916 630812 996980
rect 630876 996916 630877 996980
rect 630811 996915 630877 996916
rect 629707 996708 629773 996709
rect 629707 996644 629708 996708
rect 629772 996644 629773 996708
rect 629707 996643 629773 996644
rect 629710 995757 629770 996643
rect 630814 995757 630874 996915
rect 485635 995756 485701 995757
rect 485635 995692 485636 995756
rect 485700 995692 485701 995756
rect 485635 995691 485701 995692
rect 529059 995756 529125 995757
rect 529059 995692 529060 995756
rect 529124 995692 529125 995756
rect 529059 995691 529125 995692
rect 533475 995756 533541 995757
rect 533475 995692 533476 995756
rect 533540 995692 533541 995756
rect 533475 995691 533541 995692
rect 629707 995756 629773 995757
rect 629707 995692 629708 995756
rect 629772 995692 629773 995756
rect 629707 995691 629773 995692
rect 630811 995756 630877 995757
rect 630811 995692 630812 995756
rect 630876 995692 630877 995756
rect 630811 995691 630877 995692
rect 481219 995620 481285 995621
rect 481219 995556 481220 995620
rect 481284 995556 481285 995620
rect 481219 995555 481285 995556
rect 291331 995348 291397 995349
rect 291331 995284 291332 995348
rect 291396 995284 291397 995348
rect 291331 995283 291397 995284
rect 476435 995348 476501 995349
rect 476435 995284 476436 995348
rect 476500 995284 476501 995348
rect 476435 995283 476501 995284
rect 476803 995348 476869 995349
rect 476803 995284 476804 995348
rect 476868 995284 476869 995348
rect 476803 995283 476869 995284
rect 226379 994260 226445 994261
rect 226379 994196 226380 994260
rect 226444 994196 226445 994260
rect 226379 994195 226445 994196
rect 278635 994260 278701 994261
rect 278635 994196 278636 994260
rect 278700 994196 278701 994260
rect 278635 994195 278701 994196
rect 41459 967196 41525 967197
rect 41459 967132 41460 967196
rect 41524 967132 41525 967196
rect 41459 967131 41525 967132
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 945330 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 39806 945270 40602 945330
rect 39806 943805 39866 945270
rect 40726 943805 40786 955435
rect 41278 951693 41338 959787
rect 41462 952509 41522 967131
rect 675707 966516 675773 966517
rect 675707 966452 675708 966516
rect 675772 966452 675773 966516
rect 675707 966451 675773 966452
rect 675523 963388 675589 963389
rect 675523 963324 675524 963388
rect 675588 963324 675589 963388
rect 675523 963323 675589 963324
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 959130 41890 962099
rect 675526 959173 675586 963323
rect 41646 959070 41890 959130
rect 675523 959172 675589 959173
rect 675523 959108 675524 959172
rect 675588 959108 675589 959172
rect 675523 959107 675589 959108
rect 41459 952508 41525 952509
rect 41459 952444 41460 952508
rect 41524 952444 41525 952508
rect 41459 952443 41525 952444
rect 41646 952237 41706 959070
rect 41827 957812 41893 957813
rect 41827 957748 41828 957812
rect 41892 957748 41893 957812
rect 41827 957747 41893 957748
rect 41830 952917 41890 957747
rect 675710 954685 675770 966451
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675707 954684 675773 954685
rect 675707 954620 675708 954684
rect 675772 954620 675773 954684
rect 675707 954619 675773 954620
rect 41827 952916 41893 952917
rect 41827 952852 41828 952916
rect 41892 952852 41893 952916
rect 41827 952851 41893 952852
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 41275 951692 41341 951693
rect 41275 951628 41276 951692
rect 41340 951628 41341 951692
rect 41275 951627 41341 951628
rect 676078 949517 676138 965091
rect 676811 964748 676877 964749
rect 676811 964684 676812 964748
rect 676876 964684 676877 964748
rect 676811 964683 676877 964684
rect 676627 957812 676693 957813
rect 676627 957748 676628 957812
rect 676692 957748 676693 957812
rect 676627 957747 676693 957748
rect 676075 949516 676141 949517
rect 676075 949452 676076 949516
rect 676140 949452 676141 949516
rect 676075 949451 676141 949452
rect 39803 943804 39869 943805
rect 39803 943740 39804 943804
rect 39868 943740 39869 943804
rect 39803 943739 39869 943740
rect 40723 943804 40789 943805
rect 40723 943740 40724 943804
rect 40788 943740 40789 943804
rect 40723 943739 40789 943740
rect 42011 943804 42077 943805
rect 42011 943740 42012 943804
rect 42076 943740 42077 943804
rect 42011 943739 42077 943740
rect 41781 939452 41847 939453
rect 41781 939450 41782 939452
rect 39990 939390 41782 939450
rect 39990 814299 40050 939390
rect 41781 939388 41782 939390
rect 41846 939388 41847 939452
rect 41781 939387 41847 939388
rect 42014 937050 42074 943739
rect 674603 938092 674669 938093
rect 674603 938028 674604 938092
rect 674668 938090 674669 938092
rect 674668 938030 675034 938090
rect 674668 938028 674669 938030
rect 674603 938027 674669 938028
rect 674974 937685 675034 938030
rect 674971 937684 675037 937685
rect 674971 937620 674972 937684
rect 675036 937620 675037 937684
rect 674971 937619 675037 937620
rect 41830 936990 42074 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 676630 931565 676690 957747
rect 676814 950741 676874 964683
rect 676995 956452 677061 956453
rect 676995 956388 676996 956452
rect 677060 956388 677061 956452
rect 676995 956387 677061 956388
rect 676811 950740 676877 950741
rect 676811 950676 676812 950740
rect 676876 950676 676877 950740
rect 676811 950675 676877 950676
rect 676998 931973 677058 956387
rect 676995 931972 677061 931973
rect 676995 931908 676996 931972
rect 677060 931908 677061 931972
rect 676995 931907 677061 931908
rect 676627 931564 676693 931565
rect 676627 931500 676628 931564
rect 676692 931500 676693 931564
rect 676627 931499 676693 931500
rect 42011 911980 42077 911981
rect 42011 911916 42012 911980
rect 42076 911916 42077 911980
rect 42011 911915 42077 911916
rect 42014 885461 42074 911915
rect 42195 911708 42261 911709
rect 42195 911644 42196 911708
rect 42260 911644 42261 911708
rect 42195 911643 42261 911644
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911643
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675891 874036 675957 874037
rect 675891 873972 675892 874036
rect 675956 873972 675957 874036
rect 675891 873971 675957 873972
rect 673867 869548 673933 869549
rect 673867 869484 673868 869548
rect 673932 869484 673933 869548
rect 673867 869483 673933 869484
rect 39987 814298 40053 814299
rect 39987 814234 39988 814298
rect 40052 814234 40053 814298
rect 39987 814233 40053 814234
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40907 805492 40973 805493
rect 40907 805428 40908 805492
rect 40972 805428 40973 805492
rect 40907 805427 40973 805428
rect 40539 805356 40605 805357
rect 40539 805292 40540 805356
rect 40604 805292 40605 805356
rect 40539 805291 40605 805292
rect 40542 792573 40602 805291
rect 40723 805084 40789 805085
rect 40723 805020 40724 805084
rect 40788 805020 40789 805084
rect 40723 805019 40789 805020
rect 40726 795021 40786 805019
rect 40723 795020 40789 795021
rect 40723 794956 40724 795020
rect 40788 794956 40789 795020
rect 40723 794955 40789 794956
rect 40910 794205 40970 805427
rect 40907 794204 40973 794205
rect 40907 794140 40908 794204
rect 40972 794140 40973 794204
rect 40907 794139 40973 794140
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 788221 41522 812910
rect 42011 804812 42077 804813
rect 42011 804748 42012 804812
rect 42076 804748 42077 804812
rect 42011 804747 42077 804748
rect 41643 804540 41709 804541
rect 41643 804476 41644 804540
rect 41708 804476 41709 804540
rect 41643 804475 41709 804476
rect 41646 789037 41706 804475
rect 42014 794910 42074 804747
rect 41830 794850 42074 794910
rect 41643 789036 41709 789037
rect 41643 788972 41644 789036
rect 41708 788972 41709 789036
rect 41643 788971 41709 788972
rect 41830 788629 41890 794850
rect 41827 788628 41893 788629
rect 41827 788564 41828 788628
rect 41892 788564 41893 788628
rect 41827 788563 41893 788564
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757348 40421 757349
rect 40355 757284 40356 757348
rect 40420 757284 40421 757348
rect 40355 757283 40421 757284
rect 40358 754493 40418 757283
rect 40355 754492 40421 754493
rect 40355 754428 40356 754492
rect 40420 754428 40421 754492
rect 40355 754427 40421 754428
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 752181 40786 764899
rect 40723 752180 40789 752181
rect 40723 752116 40724 752180
rect 40788 752116 40789 752180
rect 40723 752115 40789 752116
rect 40910 751093 40970 765715
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 743749 41522 769795
rect 41643 764556 41709 764557
rect 41643 764492 41644 764556
rect 41708 764492 41709 764556
rect 41643 764491 41709 764492
rect 41646 745109 41706 764491
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41643 745108 41709 745109
rect 41643 745044 41644 745108
rect 41708 745044 41709 745108
rect 41643 745043 41709 745044
rect 41830 744837 41890 757691
rect 42011 756396 42077 756397
rect 42011 756332 42012 756396
rect 42076 756332 42077 756396
rect 42011 756331 42077 756332
rect 42014 754085 42074 756331
rect 673870 754765 673930 869483
rect 674419 854316 674485 854317
rect 674419 854252 674420 854316
rect 674484 854252 674485 854316
rect 674419 854251 674485 854252
rect 673867 754764 673933 754765
rect 673867 754700 673868 754764
rect 673932 754700 673933 754764
rect 673867 754699 673933 754700
rect 42011 754084 42077 754085
rect 42011 754020 42012 754084
rect 42076 754020 42077 754084
rect 42011 754019 42077 754020
rect 674422 753813 674482 854251
rect 674787 787268 674853 787269
rect 674787 787204 674788 787268
rect 674852 787204 674853 787268
rect 674787 787203 674853 787204
rect 674790 782781 674850 787203
rect 674971 786724 675037 786725
rect 674971 786660 674972 786724
rect 675036 786660 675037 786724
rect 674971 786659 675037 786660
rect 674974 783325 675034 786659
rect 674971 783324 675037 783325
rect 674971 783260 674972 783324
rect 675036 783260 675037 783324
rect 674971 783259 675037 783260
rect 674787 782780 674853 782781
rect 674787 782716 674788 782780
rect 674852 782716 674853 782780
rect 674787 782715 674853 782716
rect 675894 772717 675954 873971
rect 675891 772716 675957 772717
rect 675891 772652 675892 772716
rect 675956 772652 675957 772716
rect 675891 772651 675957 772652
rect 676078 768773 676138 875875
rect 676811 871996 676877 871997
rect 676811 871932 676812 871996
rect 676876 871932 676877 871996
rect 676811 871931 676877 871932
rect 676075 768772 676141 768773
rect 676075 768708 676076 768772
rect 676140 768708 676141 768772
rect 676075 768707 676141 768708
rect 675891 766596 675957 766597
rect 675891 766532 675892 766596
rect 675956 766532 675957 766596
rect 675891 766531 675957 766532
rect 674419 753812 674485 753813
rect 674419 753748 674420 753812
rect 674484 753748 674485 753812
rect 674419 753747 674485 753748
rect 41827 744836 41893 744837
rect 41827 744772 41828 744836
rect 41892 744772 41893 744836
rect 41827 744771 41893 744772
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674419 741572 674485 741573
rect 674419 741508 674420 741572
rect 674484 741508 674485 741572
rect 674419 741507 674485 741508
rect 670739 734092 670805 734093
rect 670739 734028 670740 734092
rect 670804 734028 670805 734092
rect 670739 734027 670805 734028
rect 670742 728517 670802 734027
rect 674235 732868 674301 732869
rect 674235 732804 674236 732868
rect 674300 732804 674301 732868
rect 674235 732803 674301 732804
rect 670739 728516 670805 728517
rect 670739 728452 670740 728516
rect 670804 728452 670805 728516
rect 670739 728451 670805 728452
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40355 721772 40421 721773
rect 40355 721708 40356 721772
rect 40420 721708 40421 721772
rect 40355 721707 40421 721708
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40358 716821 40418 721707
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40355 716820 40421 716821
rect 40355 716756 40356 716820
rect 40420 716756 40421 716820
rect 40355 716755 40421 716756
rect 40542 704309 40602 718523
rect 40726 706757 40786 721707
rect 40907 716820 40973 716821
rect 40907 716756 40908 716820
rect 40972 716756 40973 716820
rect 40907 716755 40973 716756
rect 40910 708525 40970 716755
rect 40907 708524 40973 708525
rect 40907 708460 40908 708524
rect 40972 708460 40973 708524
rect 40907 708459 40973 708460
rect 40723 706756 40789 706757
rect 40723 706692 40724 706756
rect 40788 706692 40789 706756
rect 40723 706691 40789 706692
rect 40539 704308 40605 704309
rect 40539 704244 40540 704308
rect 40604 704244 40605 704308
rect 40539 704243 40605 704244
rect 41462 700501 41522 726550
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41646 701589 41706 721707
rect 41827 714780 41893 714781
rect 41827 714716 41828 714780
rect 41892 714716 41893 714780
rect 41827 714715 41893 714716
rect 41830 701861 41890 714715
rect 42011 714644 42077 714645
rect 42011 714580 42012 714644
rect 42076 714580 42077 714644
rect 42011 714579 42077 714580
rect 42014 709885 42074 714579
rect 42011 709884 42077 709885
rect 42011 709820 42012 709884
rect 42076 709820 42077 709884
rect 42011 709819 42077 709820
rect 673315 705124 673381 705125
rect 673315 705060 673316 705124
rect 673380 705060 673381 705124
rect 673315 705059 673381 705060
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41643 701588 41709 701589
rect 41643 701524 41644 701588
rect 41708 701524 41709 701588
rect 41643 701523 41709 701524
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 42195 683636 42261 683637
rect 42195 683572 42196 683636
rect 42260 683572 42261 683636
rect 42195 683571 42261 683572
rect 42011 682820 42077 682821
rect 42011 682756 42012 682820
rect 42076 682756 42077 682820
rect 42011 682755 42077 682756
rect 40726 679222 41154 679282
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40355 671260 40421 671261
rect 40355 671196 40356 671260
rect 40420 671196 40421 671260
rect 40355 671195 40421 671196
rect 40358 667589 40418 671195
rect 40355 667588 40421 667589
rect 40355 667524 40356 667588
rect 40420 667524 40421 667588
rect 40355 667523 40421 667524
rect 40542 662693 40602 678927
rect 40726 665413 40786 679222
rect 40907 678992 40973 678993
rect 40907 678928 40908 678992
rect 40972 678928 40973 678992
rect 40907 678927 40973 678928
rect 40910 667045 40970 678927
rect 41094 678330 41154 679222
rect 41827 678332 41893 678333
rect 41827 678330 41828 678332
rect 41094 678270 41828 678330
rect 41827 678268 41828 678270
rect 41892 678268 41893 678332
rect 41827 678267 41893 678268
rect 41827 677652 41893 677653
rect 41827 677650 41828 677652
rect 41462 677590 41828 677650
rect 40907 667044 40973 667045
rect 40907 666980 40908 667044
rect 40972 666980 40973 667044
rect 40907 666979 40973 666980
rect 40723 665412 40789 665413
rect 40723 665348 40724 665412
rect 40788 665348 40789 665412
rect 40723 665347 40789 665348
rect 40539 662692 40605 662693
rect 40539 662628 40540 662692
rect 40604 662628 40605 662692
rect 40539 662627 40605 662628
rect 41462 657253 41522 677590
rect 41827 677588 41828 677590
rect 41892 677588 41893 677652
rect 41827 677587 41893 677588
rect 42014 676230 42074 682755
rect 42198 677653 42258 683571
rect 42195 677652 42261 677653
rect 42195 677588 42196 677652
rect 42260 677588 42261 677652
rect 42195 677587 42261 677588
rect 41646 676170 42074 676230
rect 41646 658613 41706 676170
rect 41827 670988 41893 670989
rect 41827 670924 41828 670988
rect 41892 670924 41893 670988
rect 41827 670923 41893 670924
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 670923
rect 42195 669356 42261 669357
rect 42195 669292 42196 669356
rect 42260 669292 42261 669356
rect 42195 669291 42261 669292
rect 42198 667861 42258 669291
rect 42195 667860 42261 667861
rect 42195 667796 42196 667860
rect 42260 667796 42261 667860
rect 42195 667795 42261 667796
rect 42011 667044 42077 667045
rect 42011 666980 42012 667044
rect 42076 666980 42077 667044
rect 42011 666979 42077 666980
rect 42014 664053 42074 666979
rect 42011 664052 42077 664053
rect 42011 663988 42012 664052
rect 42076 663988 42077 664052
rect 42011 663987 42077 663988
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 634948 40605 634949
rect 40539 634884 40540 634948
rect 40604 634884 40605 634948
rect 40539 634883 40605 634884
rect 40542 622165 40602 634883
rect 40539 622164 40605 622165
rect 40539 622100 40540 622164
rect 40604 622100 40605 622164
rect 40539 622099 40605 622100
rect 41462 616045 41522 640595
rect 41827 639232 41893 639233
rect 41827 639168 41828 639232
rect 41892 639168 41893 639232
rect 41827 639167 41893 639168
rect 41643 638620 41709 638621
rect 41643 638556 41644 638620
rect 41708 638556 41709 638620
rect 41643 638555 41709 638556
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41646 615510 41706 638555
rect 41830 615773 41890 639167
rect 42011 626652 42077 626653
rect 42011 626588 42012 626652
rect 42076 626588 42077 626652
rect 42011 626587 42077 626588
rect 42014 624477 42074 626587
rect 42195 625020 42261 625021
rect 42195 624956 42196 625020
rect 42260 624956 42261 625020
rect 42195 624955 42261 624956
rect 42011 624476 42077 624477
rect 42011 624412 42012 624476
rect 42076 624412 42077 624476
rect 42011 624411 42077 624412
rect 42198 620261 42258 624955
rect 42195 620260 42261 620261
rect 42195 620196 42196 620260
rect 42260 620196 42261 620260
rect 42195 620195 42261 620196
rect 41827 615772 41893 615773
rect 41827 615708 41828 615772
rect 41892 615708 41893 615772
rect 41827 615707 41893 615708
rect 41646 615450 41890 615510
rect 41830 612781 41890 615450
rect 41827 612780 41893 612781
rect 41827 612716 41828 612780
rect 41892 612716 41893 612780
rect 41827 612715 41893 612716
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 596460 41893 596461
rect 41827 596396 41828 596460
rect 41892 596396 41893 596460
rect 41827 596395 41893 596396
rect 41830 596050 41890 596395
rect 41646 595990 41890 596050
rect 40726 589870 41338 589930
rect 40539 589660 40605 589661
rect 40539 589596 40540 589660
rect 40604 589596 40605 589660
rect 40539 589595 40605 589596
rect 40355 585988 40421 585989
rect 40355 585924 40356 585988
rect 40420 585924 40421 585988
rect 40355 585923 40421 585924
rect 40358 582589 40418 585923
rect 40355 582588 40421 582589
rect 40355 582524 40356 582588
rect 40420 582524 40421 582588
rect 40355 582523 40421 582524
rect 40542 576877 40602 589595
rect 40726 580005 40786 589870
rect 41278 589661 41338 589870
rect 41275 589660 41341 589661
rect 41275 589596 41276 589660
rect 41340 589596 41341 589660
rect 41275 589595 41341 589596
rect 40907 589388 40973 589389
rect 40907 589324 40908 589388
rect 40972 589324 40973 589388
rect 40907 589323 40973 589324
rect 40910 580685 40970 589323
rect 41646 589290 41706 595990
rect 41827 592380 41893 592381
rect 41827 592316 41828 592380
rect 41892 592316 41893 592380
rect 41827 592315 41893 592316
rect 41830 589661 41890 592315
rect 41827 589660 41893 589661
rect 41827 589596 41828 589660
rect 41892 589596 41893 589660
rect 41827 589595 41893 589596
rect 42014 589290 42074 597211
rect 43851 591564 43917 591565
rect 43851 591500 43852 591564
rect 43916 591500 43917 591564
rect 43851 591499 43917 591500
rect 41462 589230 41706 589290
rect 41830 589230 42074 589290
rect 41091 584628 41157 584629
rect 41091 584564 41092 584628
rect 41156 584564 41157 584628
rect 41091 584563 41157 584564
rect 40907 580684 40973 580685
rect 40907 580620 40908 580684
rect 40972 580620 40973 580684
rect 40907 580619 40973 580620
rect 41094 580277 41154 584563
rect 41091 580276 41157 580277
rect 41091 580212 41092 580276
rect 41156 580212 41157 580276
rect 41091 580211 41157 580212
rect 40723 580004 40789 580005
rect 40723 579940 40724 580004
rect 40788 579940 40789 580004
rect 40723 579939 40789 579940
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 571709 41522 589230
rect 41830 587210 41890 589230
rect 41646 587150 41890 587210
rect 41459 571708 41525 571709
rect 41459 571644 41460 571708
rect 41524 571644 41525 571708
rect 41459 571643 41525 571644
rect 41646 571029 41706 587150
rect 41827 585716 41893 585717
rect 41827 585652 41828 585716
rect 41892 585652 41893 585716
rect 41827 585651 41893 585652
rect 41830 571437 41890 585651
rect 42379 585308 42445 585309
rect 42379 585244 42380 585308
rect 42444 585244 42445 585308
rect 42379 585243 42445 585244
rect 42011 584628 42077 584629
rect 42011 584564 42012 584628
rect 42076 584564 42077 584628
rect 42011 584563 42077 584564
rect 42014 573205 42074 584563
rect 42382 578250 42442 585243
rect 42198 578190 42442 578250
rect 42198 576605 42258 578190
rect 42195 576604 42261 576605
rect 42195 576540 42196 576604
rect 42260 576540 42261 576604
rect 42195 576539 42261 576540
rect 42011 573204 42077 573205
rect 42011 573140 42012 573204
rect 42076 573140 42077 573204
rect 42011 573139 42077 573140
rect 41827 571436 41893 571437
rect 41827 571372 41828 571436
rect 41892 571372 41893 571436
rect 41827 571371 41893 571372
rect 41643 571028 41709 571029
rect 41643 570964 41644 571028
rect 41708 570964 41709 571028
rect 41643 570963 41709 570964
rect 41827 553212 41893 553213
rect 41827 553210 41828 553212
rect 41462 553150 41828 553210
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 534989 40602 545395
rect 40726 538253 40786 545667
rect 40723 538252 40789 538253
rect 40723 538188 40724 538252
rect 40788 538188 40789 538252
rect 40723 538187 40789 538188
rect 40539 534988 40605 534989
rect 40539 534924 40540 534988
rect 40604 534924 40605 534988
rect 40539 534923 40605 534924
rect 41462 530637 41522 553150
rect 41827 553148 41828 553150
rect 41892 553148 41893 553212
rect 41827 553147 41893 553148
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 530636 41525 530637
rect 41459 530572 41460 530636
rect 41524 530572 41525 530636
rect 41459 530571 41525 530572
rect 41646 529141 41706 546347
rect 41830 529413 41890 552739
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 41643 529140 41709 529141
rect 41643 529076 41644 529140
rect 41708 529076 41709 529140
rect 41643 529075 41709 529076
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41462 424630 41890 424690
rect 40539 418708 40605 418709
rect 40539 418644 40540 418708
rect 40604 418644 40605 418708
rect 40539 418643 40605 418644
rect 40542 403885 40602 418643
rect 40723 418572 40789 418573
rect 40723 418508 40724 418572
rect 40788 418508 40789 418572
rect 40723 418507 40789 418508
rect 40726 409461 40786 418507
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 401845 41522 424630
rect 41643 418844 41709 418845
rect 41643 418780 41644 418844
rect 41708 418780 41709 418844
rect 41643 418779 41709 418780
rect 41646 402990 41706 418779
rect 42014 408510 42074 424763
rect 41830 408450 42074 408510
rect 41830 406333 41890 408450
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41459 401844 41525 401845
rect 41459 401780 41460 401844
rect 41524 401780 41525 401844
rect 41459 401779 41525 401780
rect 41830 398853 41890 402930
rect 41827 398852 41893 398853
rect 41827 398788 41828 398852
rect 41892 398788 41893 398852
rect 41827 398787 41893 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40355 375732 40421 375733
rect 40355 375668 40356 375732
rect 40420 375668 40421 375732
rect 40355 375667 40421 375668
rect 40358 368661 40418 375667
rect 40355 368660 40421 368661
rect 40355 368596 40356 368660
rect 40420 368596 40421 368660
rect 40355 368595 40421 368596
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363629 40786 378115
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364309 40970 377707
rect 40907 364308 40973 364309
rect 40907 364244 40908 364308
rect 40972 364244 40973 364308
rect 40907 364243 40973 364244
rect 40723 363628 40789 363629
rect 40723 363564 40724 363628
rect 40788 363564 40789 363628
rect 40723 363563 40789 363564
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 358733 41522 381787
rect 41827 378588 41893 378589
rect 41827 378524 41828 378588
rect 41892 378524 41893 378588
rect 41827 378523 41893 378524
rect 41643 376548 41709 376549
rect 41643 376484 41644 376548
rect 41708 376484 41709 376548
rect 41643 376483 41709 376484
rect 41646 360210 41706 376483
rect 41830 362949 41890 378523
rect 41827 362948 41893 362949
rect 41827 362884 41828 362948
rect 41892 362884 41893 362948
rect 41827 362883 41893 362884
rect 41646 360150 41890 360210
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 41830 355741 41890 360150
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43854 354245 43914 591499
rect 673318 474877 673378 705059
rect 674238 681053 674298 732803
rect 674422 682413 674482 741507
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674419 682412 674485 682413
rect 674419 682348 674420 682412
rect 674484 682348 674485 682412
rect 674419 682347 674485 682348
rect 674235 681052 674301 681053
rect 674235 680988 674236 681052
rect 674300 680988 674301 681052
rect 674235 680987 674301 680988
rect 674419 666364 674485 666365
rect 674419 666300 674420 666364
rect 674484 666300 674485 666364
rect 674419 666299 674485 666300
rect 673499 665820 673565 665821
rect 673499 665756 673500 665820
rect 673564 665756 673565 665820
rect 673499 665755 673565 665756
rect 673502 664730 673562 665755
rect 673683 665684 673749 665685
rect 673683 665620 673684 665684
rect 673748 665620 673749 665684
rect 673683 665619 673749 665620
rect 673686 665141 673746 665619
rect 674422 665141 674482 666299
rect 673683 665140 673749 665141
rect 673683 665076 673684 665140
rect 673748 665076 673749 665140
rect 673683 665075 673749 665076
rect 674419 665140 674485 665141
rect 674419 665076 674420 665140
rect 674484 665076 674485 665140
rect 674419 665075 674485 665076
rect 673502 664670 673746 664730
rect 673686 664325 673746 664670
rect 673683 664324 673749 664325
rect 673683 664260 673684 664324
rect 673748 664260 673749 664324
rect 673683 664259 673749 664260
rect 674606 662285 674666 738107
rect 675894 728789 675954 766531
rect 676075 765100 676141 765101
rect 676075 765036 676076 765100
rect 676140 765036 676141 765100
rect 676075 765035 676141 765036
rect 675891 728788 675957 728789
rect 675891 728724 675892 728788
rect 675956 728724 675957 728788
rect 675891 728723 675957 728724
rect 676078 725797 676138 765035
rect 676627 761792 676693 761793
rect 676627 761728 676628 761792
rect 676692 761790 676693 761792
rect 676814 761790 676874 871931
rect 676995 780604 677061 780605
rect 676995 780540 676996 780604
rect 677060 780540 677061 780604
rect 676995 780539 677061 780540
rect 676998 761837 677058 780539
rect 676692 761730 676874 761790
rect 676995 761836 677061 761837
rect 676995 761772 676996 761836
rect 677060 761772 677061 761836
rect 676995 761771 677061 761772
rect 676692 761728 676693 761730
rect 676627 761727 676693 761728
rect 676811 728788 676877 728789
rect 676811 728724 676812 728788
rect 676876 728724 676877 728788
rect 676811 728723 676877 728724
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712110 676874 728723
rect 675894 712061 676874 712110
rect 675891 712060 676874 712061
rect 675891 711996 675892 712060
rect 675956 712050 676874 712060
rect 675956 711996 675957 712050
rect 675891 711995 675957 711996
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 674787 689756 674853 689757
rect 674787 689692 674788 689756
rect 674852 689692 674853 689756
rect 674787 689691 674853 689692
rect 674790 688805 674850 689691
rect 674787 688804 674853 688805
rect 674787 688740 674788 688804
rect 674852 688740 674853 688804
rect 674787 688739 674853 688740
rect 674603 662284 674669 662285
rect 674603 662220 674604 662284
rect 674668 662220 674669 662284
rect 674603 662219 674669 662220
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674235 648956 674301 648957
rect 674235 648892 674236 648956
rect 674300 648892 674301 648956
rect 674235 648891 674301 648892
rect 674238 592653 674298 648891
rect 674603 645148 674669 645149
rect 674603 645084 674604 645148
rect 674668 645084 674669 645148
rect 674603 645083 674669 645084
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674235 592652 674301 592653
rect 674235 592588 674236 592652
rect 674300 592588 674301 592652
rect 674235 592587 674301 592588
rect 674422 533901 674482 602923
rect 674419 533900 674485 533901
rect 674419 533836 674420 533900
rect 674484 533836 674485 533900
rect 674419 533835 674485 533836
rect 674606 475421 674666 645083
rect 675155 640524 675221 640525
rect 675155 640460 675156 640524
rect 675220 640460 675221 640524
rect 675155 640459 675221 640460
rect 675158 637669 675218 640459
rect 675342 638077 675402 652835
rect 675523 651540 675589 651541
rect 675523 651476 675524 651540
rect 675588 651476 675589 651540
rect 675523 651475 675589 651476
rect 675339 638076 675405 638077
rect 675339 638012 675340 638076
rect 675404 638012 675405 638076
rect 675339 638011 675405 638012
rect 675526 637805 675586 651475
rect 676811 644740 676877 644741
rect 676811 644676 676812 644740
rect 676876 644676 676877 644740
rect 676811 644675 676877 644676
rect 675523 637804 675589 637805
rect 675523 637740 675524 637804
rect 675588 637740 675589 637804
rect 675523 637739 675589 637740
rect 675155 637668 675221 637669
rect 675155 637604 675156 637668
rect 675220 637604 675221 637668
rect 675155 637603 675221 637604
rect 675155 633044 675221 633045
rect 675155 632980 675156 633044
rect 675220 632980 675221 633044
rect 675155 632979 675221 632980
rect 675158 592925 675218 632979
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 675523 629780 675589 629781
rect 675523 629716 675524 629780
rect 675588 629716 675589 629780
rect 675523 629715 675589 629716
rect 675526 593877 675586 629715
rect 675707 596732 675773 596733
rect 675707 596668 675708 596732
rect 675772 596668 675773 596732
rect 675707 596667 675773 596668
rect 675523 593876 675589 593877
rect 675523 593812 675524 593876
rect 675588 593812 675589 593876
rect 675523 593811 675589 593812
rect 675155 592924 675221 592925
rect 675155 592860 675156 592924
rect 675220 592860 675221 592924
rect 675155 592859 675221 592860
rect 675710 592381 675770 596667
rect 675707 592380 675773 592381
rect 675707 592316 675708 592380
rect 675772 592316 675773 592380
rect 675707 592315 675773 592316
rect 676078 590613 676138 631347
rect 676075 590612 676141 590613
rect 676075 590548 676076 590612
rect 676140 590548 676141 590612
rect 676075 590547 676141 590548
rect 676814 572797 676874 644675
rect 676998 619173 677058 694043
rect 676995 619172 677061 619173
rect 676995 619108 676996 619172
rect 677060 619108 677061 619172
rect 676995 619107 677061 619108
rect 676995 594148 677061 594149
rect 676995 594084 676996 594148
rect 677060 594084 677061 594148
rect 676995 594083 677061 594084
rect 676998 576469 677058 594083
rect 676995 576468 677061 576469
rect 676995 576404 676996 576468
rect 677060 576404 677061 576468
rect 676995 576403 677061 576404
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 675523 562732 675589 562733
rect 675523 562730 675524 562732
rect 675342 562670 675524 562730
rect 675342 544917 675402 562670
rect 675523 562668 675524 562670
rect 675588 562668 675589 562732
rect 675523 562667 675589 562668
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 675339 544916 675405 544917
rect 675339 544852 675340 544916
rect 675404 544852 675405 544916
rect 675339 544851 675405 544852
rect 675526 544509 675586 561171
rect 676259 557700 676325 557701
rect 676259 557636 676260 557700
rect 676324 557636 676325 557700
rect 676259 557635 676325 557636
rect 675891 550492 675957 550493
rect 675891 550428 675892 550492
rect 675956 550428 675957 550492
rect 675891 550427 675957 550428
rect 675894 547637 675954 550427
rect 676262 547637 676322 557635
rect 676811 554028 676877 554029
rect 676811 553964 676812 554028
rect 676876 553964 676877 554028
rect 676811 553963 676877 553964
rect 675891 547636 675957 547637
rect 675891 547572 675892 547636
rect 675956 547572 675957 547636
rect 675891 547571 675957 547572
rect 676259 547636 676325 547637
rect 676259 547572 676260 547636
rect 676324 547572 676325 547636
rect 676259 547571 676325 547572
rect 675523 544508 675589 544509
rect 675523 544444 675524 544508
rect 675588 544444 675589 544508
rect 675523 544443 675589 544444
rect 676814 503437 676874 553963
rect 676995 550220 677061 550221
rect 676995 550156 676996 550220
rect 677060 550156 677061 550220
rect 676995 550155 677061 550156
rect 676998 503709 677058 550155
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 503436 676877 503437
rect 676811 503372 676812 503436
rect 676876 503372 676877 503436
rect 676811 503371 676877 503372
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 675894 488610 675954 488819
rect 675894 488550 676874 488610
rect 674603 475420 674669 475421
rect 674603 475356 674604 475420
rect 674668 475356 674669 475420
rect 674603 475355 674669 475356
rect 673315 474876 673381 474877
rect 673315 474812 673316 474876
rect 673380 474812 673381 474876
rect 673315 474811 673381 474812
rect 675339 453796 675405 453797
rect 675339 453732 675340 453796
rect 675404 453732 675405 453796
rect 675339 453731 675405 453732
rect 675342 410549 675402 453731
rect 675339 410548 675405 410549
rect 675339 410484 675340 410548
rect 675404 410484 675405 410548
rect 675339 410483 675405 410484
rect 676814 401301 676874 488550
rect 676811 401300 676877 401301
rect 676811 401236 676812 401300
rect 676876 401236 676877 401300
rect 676811 401235 676877 401236
rect 675891 398852 675957 398853
rect 675891 398788 675892 398852
rect 675956 398788 675957 398852
rect 675891 398787 675957 398788
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 674790 372605 674850 377979
rect 675894 375053 675954 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676075 393140 676141 393141
rect 676075 393076 676076 393140
rect 676140 393076 676141 393140
rect 676075 393075 676141 393076
rect 675891 375052 675957 375053
rect 675891 374988 675892 375052
rect 675956 374988 675957 375052
rect 675891 374987 675957 374988
rect 676078 373013 676138 393075
rect 676262 377365 676322 395115
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676446 380629 676506 394707
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 676075 373012 676141 373013
rect 676075 372948 676076 373012
rect 676140 372948 676141 373012
rect 676075 372947 676141 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 43851 354244 43917 354245
rect 43851 354180 43852 354244
rect 43916 354180 43917 354244
rect 43851 354179 43917 354180
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 44219 353836 44285 353837
rect 44219 353772 44220 353836
rect 44284 353772 44285 353836
rect 44219 353771 44285 353772
rect 44222 342685 44282 353771
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 342684 44285 342685
rect 44219 342620 44220 342684
rect 44284 342620 44285 342684
rect 44219 342619 44285 342620
rect 44406 342410 44466 342891
rect 44222 342350 44466 342410
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 41459 337788 41525 337789
rect 41459 337724 41460 337788
rect 41524 337724 41525 337788
rect 41459 337723 41525 337724
rect 40539 336564 40605 336565
rect 40539 336500 40540 336564
rect 40604 336500 40605 336564
rect 40539 336499 40605 336500
rect 40542 316709 40602 336499
rect 40723 335340 40789 335341
rect 40723 335276 40724 335340
rect 40788 335276 40789 335340
rect 40723 335275 40789 335276
rect 40726 317525 40786 335275
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40910 325413 40970 333643
rect 41462 326773 41522 337723
rect 42931 337516 42997 337517
rect 42931 337452 42932 337516
rect 42996 337452 42997 337516
rect 42931 337451 42997 337452
rect 41827 336156 41893 336157
rect 41827 336092 41828 336156
rect 41892 336092 41893 336156
rect 41827 336091 41893 336092
rect 41643 328404 41709 328405
rect 41643 328340 41644 328404
rect 41708 328340 41709 328404
rect 41643 328339 41709 328340
rect 41459 326772 41525 326773
rect 41459 326708 41460 326772
rect 41524 326708 41525 326772
rect 41459 326707 41525 326708
rect 41646 325710 41706 328339
rect 41462 325650 41706 325710
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41462 324869 41522 325650
rect 41459 324868 41525 324869
rect 41459 324804 41460 324868
rect 41524 324804 41525 324868
rect 41459 324803 41525 324804
rect 40723 317524 40789 317525
rect 40723 317460 40724 317524
rect 40788 317460 40789 317524
rect 40723 317459 40789 317460
rect 40539 316708 40605 316709
rect 40539 316644 40540 316708
rect 40604 316644 40605 316708
rect 40539 316643 40605 316644
rect 41830 315621 41890 336091
rect 42747 335748 42813 335749
rect 42747 335684 42748 335748
rect 42812 335684 42813 335748
rect 42747 335683 42813 335684
rect 42750 334661 42810 335683
rect 42747 334660 42813 334661
rect 42747 334596 42748 334660
rect 42812 334596 42813 334660
rect 42747 334595 42813 334596
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 42934 312765 42994 337451
rect 43115 337244 43181 337245
rect 43115 337180 43116 337244
rect 43180 337180 43181 337244
rect 43115 337179 43181 337180
rect 43118 316029 43178 337179
rect 43299 336428 43365 336429
rect 43299 336364 43300 336428
rect 43364 336364 43365 336428
rect 43299 336363 43365 336364
rect 43302 334661 43362 336363
rect 43299 334660 43365 334661
rect 43299 334596 43300 334660
rect 43364 334596 43365 334660
rect 43299 334595 43365 334596
rect 43115 316028 43181 316029
rect 43115 315964 43116 316028
rect 43180 315964 43181 316028
rect 43115 315963 43181 315964
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 43670 297669 43730 340443
rect 44222 316050 44282 342350
rect 44403 342140 44469 342141
rect 44403 342076 44404 342140
rect 44468 342076 44469 342140
rect 44403 342075 44469 342076
rect 44406 325710 44466 342075
rect 675342 339013 675402 354179
rect 675523 353020 675589 353021
rect 675523 352956 675524 353020
rect 675588 352956 675589 353020
rect 675523 352955 675589 352956
rect 675339 339012 675405 339013
rect 675339 338948 675340 339012
rect 675404 338948 675405 339012
rect 675339 338947 675405 338948
rect 675526 337789 675586 352955
rect 675891 351932 675957 351933
rect 675891 351868 675892 351932
rect 675956 351930 675957 351932
rect 675956 351870 676322 351930
rect 675956 351868 675957 351870
rect 675891 351867 675957 351868
rect 676262 351250 676322 351870
rect 676262 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675891 349212 675957 349213
rect 675891 349148 675892 349212
rect 675956 349210 675957 349212
rect 675956 349150 676138 349210
rect 675956 349148 675957 349150
rect 675891 349147 675957 349148
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 676078 328405 676138 349150
rect 676262 332349 676322 349830
rect 676446 336701 676506 350510
rect 676630 340237 676690 351190
rect 676627 340236 676693 340237
rect 676627 340172 676628 340236
rect 676692 340172 676693 340236
rect 676627 340171 676693 340172
rect 676443 336700 676509 336701
rect 676443 336636 676444 336700
rect 676508 336636 676509 336700
rect 676443 336635 676509 336636
rect 676259 332348 676325 332349
rect 676259 332284 676260 332348
rect 676324 332284 676325 332348
rect 676259 332283 676325 332284
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 44406 325650 44650 325710
rect 44222 315990 44466 316050
rect 44406 311269 44466 315990
rect 44590 311541 44650 325650
rect 44587 311540 44653 311541
rect 44587 311476 44588 311540
rect 44652 311476 44653 311540
rect 44587 311475 44653 311476
rect 44403 311268 44469 311269
rect 44403 311204 44404 311268
rect 44468 311204 44469 311268
rect 44403 311203 44469 311204
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 303650 675770 308755
rect 675891 306780 675957 306781
rect 675891 306716 675892 306780
rect 675956 306716 675957 306780
rect 675891 306715 675957 306716
rect 675894 305010 675954 306715
rect 675894 304950 676322 305010
rect 675710 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 675707 298076 675773 298077
rect 675707 298012 675708 298076
rect 675772 298012 675773 298076
rect 675707 298011 675773 298012
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 292770 41890 295563
rect 40726 292710 41890 292770
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 40726 278493 40786 292710
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 40907 292527 40973 292528
rect 40723 278492 40789 278493
rect 40723 278428 40724 278492
rect 40788 278428 40789 278492
rect 40723 278427 40789 278428
rect 40910 277949 40970 292527
rect 41827 292500 41893 292501
rect 41827 292436 41828 292500
rect 41892 292436 41893 292500
rect 41827 292435 41893 292436
rect 41830 292090 41890 292435
rect 41646 292030 41890 292090
rect 41646 289830 41706 292030
rect 41827 290460 41893 290461
rect 41827 290396 41828 290460
rect 41892 290396 41893 290460
rect 41827 290395 41893 290396
rect 41462 289770 41706 289830
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 289770
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 290395
rect 42014 281485 42074 296379
rect 675710 281621 675770 298011
rect 675894 282845 675954 302635
rect 676078 283661 676138 303590
rect 676262 295221 676322 304950
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676259 295220 676325 295221
rect 676259 295156 676260 295220
rect 676324 295156 676325 295220
rect 676259 295155 676325 295156
rect 676446 291549 676506 301547
rect 676627 301476 676693 301477
rect 676627 301412 676628 301476
rect 676692 301412 676693 301476
rect 676627 301411 676693 301412
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676630 287061 676690 301411
rect 676627 287060 676693 287061
rect 676627 286996 676628 287060
rect 676692 286996 676693 287060
rect 676627 286995 676693 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 674971 263668 675037 263669
rect 674971 263604 674972 263668
rect 675036 263604 675037 263668
rect 674971 263603 675037 263604
rect 674974 253950 675034 263603
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 674790 253890 675034 253950
rect 40723 251428 40789 251429
rect 40723 251364 40724 251428
rect 40788 251364 40789 251428
rect 40723 251363 40789 251364
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 235925 40602 249731
rect 40726 240141 40786 251363
rect 674790 249661 674850 253890
rect 676078 249933 676138 262379
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 676075 249932 676141 249933
rect 676075 249868 676076 249932
rect 676140 249868 676141 249932
rect 676075 249867 676141 249868
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676814 245581 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 674787 245580 674853 245581
rect 674787 245516 674788 245580
rect 674852 245516 674853 245580
rect 674787 245515 674853 245516
rect 675891 245580 675957 245581
rect 675891 245516 675892 245580
rect 675956 245516 675957 245580
rect 675891 245515 675957 245516
rect 676811 245580 676877 245581
rect 676811 245516 676812 245580
rect 676876 245516 676877 245580
rect 676811 245515 676877 245516
rect 40723 240140 40789 240141
rect 40723 240076 40724 240140
rect 40788 240076 40789 240140
rect 40723 240075 40789 240076
rect 673315 240004 673381 240005
rect 673315 239940 673316 240004
rect 673380 239940 673381 240004
rect 673315 239939 673381 239940
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 40539 235924 40605 235925
rect 40539 235860 40540 235924
rect 40604 235860 40605 235924
rect 40539 235859 40605 235860
rect 42014 227357 42074 237355
rect 673318 235245 673378 239939
rect 674790 237285 674850 245515
rect 675339 245308 675405 245309
rect 675339 245244 675340 245308
rect 675404 245244 675405 245308
rect 675339 245243 675405 245244
rect 675342 240277 675402 245243
rect 675894 242317 675954 245515
rect 675891 242316 675957 242317
rect 675891 242252 675892 242316
rect 675956 242252 675957 242316
rect 675891 242251 675957 242252
rect 675339 240276 675405 240277
rect 675339 240212 675340 240276
rect 675404 240212 675405 240276
rect 675339 240211 675405 240212
rect 674787 237284 674853 237285
rect 674787 237220 674788 237284
rect 674852 237220 674853 237284
rect 674787 237219 674853 237220
rect 674051 237148 674117 237149
rect 674051 237084 674052 237148
rect 674116 237084 674117 237148
rect 674051 237083 674117 237084
rect 673315 235244 673381 235245
rect 673315 235180 673316 235244
rect 673380 235180 673381 235244
rect 673315 235179 673381 235180
rect 671291 233204 671357 233205
rect 671291 233140 671292 233204
rect 671356 233140 671357 233204
rect 671291 233139 671357 233140
rect 669267 231436 669333 231437
rect 669267 231372 669268 231436
rect 669332 231372 669333 231436
rect 669267 231371 669333 231372
rect 669270 230890 669330 231371
rect 669270 230830 669514 230890
rect 669454 228853 669514 230830
rect 669451 228852 669517 228853
rect 669451 228788 669452 228852
rect 669516 228788 669517 228852
rect 669451 228787 669517 228788
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 671107 227220 671173 227221
rect 671107 227156 671108 227220
rect 671172 227156 671173 227220
rect 671107 227155 671173 227156
rect 671110 223957 671170 227155
rect 671107 223956 671173 223957
rect 671107 223892 671108 223956
rect 671172 223892 671173 223956
rect 671107 223891 671173 223892
rect 562363 222052 562429 222053
rect 562363 221988 562364 222052
rect 562428 222050 562429 222052
rect 564571 222052 564637 222053
rect 564571 222050 564572 222052
rect 562428 221990 564572 222050
rect 562428 221988 562429 221990
rect 562363 221987 562429 221988
rect 564571 221988 564572 221990
rect 564636 221988 564637 222052
rect 564571 221987 564637 221988
rect 572851 222052 572917 222053
rect 572851 221988 572852 222052
rect 572916 221988 572917 222052
rect 572851 221987 572917 221988
rect 572854 221370 572914 221987
rect 572118 221310 572914 221370
rect 572118 220421 572178 221310
rect 572851 220692 572917 220693
rect 572851 220628 572852 220692
rect 572916 220628 572917 220692
rect 572851 220627 572917 220628
rect 572115 220420 572181 220421
rect 572115 220356 572116 220420
rect 572180 220356 572181 220420
rect 572115 220355 572181 220356
rect 572854 218650 572914 220627
rect 578187 220420 578253 220421
rect 578187 220356 578188 220420
rect 578252 220356 578253 220420
rect 578187 220355 578253 220356
rect 573955 220284 574021 220285
rect 573955 220220 573956 220284
rect 574020 220220 574021 220284
rect 573955 220219 574021 220220
rect 573958 219418 574018 220219
rect 578190 218738 578250 220355
rect 572118 218590 572914 218650
rect 572118 218381 572178 218590
rect 572115 218380 572181 218381
rect 572115 218316 572116 218380
rect 572180 218316 572181 218380
rect 572115 218315 572181 218316
rect 592355 217564 592421 217565
rect 592355 217500 592356 217564
rect 592420 217500 592421 217564
rect 592355 217499 592421 217500
rect 591987 217292 592053 217293
rect 591987 217228 591988 217292
rect 592052 217290 592053 217292
rect 592358 217290 592418 217499
rect 592052 217230 592418 217290
rect 592052 217228 592053 217230
rect 591987 217227 592053 217228
rect 575614 213213 575674 217142
rect 575611 213212 575677 213213
rect 575611 213148 575612 213212
rect 575676 213148 575677 213212
rect 575611 213147 575677 213148
rect 667979 212396 668045 212397
rect 667979 212332 667980 212396
rect 668044 212332 668045 212396
rect 667979 212331 668045 212332
rect 42011 210084 42077 210085
rect 42011 210020 42012 210084
rect 42076 210020 42077 210084
rect 42011 210019 42077 210020
rect 40723 208180 40789 208181
rect 40723 208116 40724 208180
rect 40788 208116 40789 208180
rect 40723 208115 40789 208116
rect 40539 206956 40605 206957
rect 40539 206892 40540 206956
rect 40604 206892 40605 206956
rect 40539 206891 40605 206892
rect 40542 194581 40602 206891
rect 40726 197165 40786 208115
rect 41643 207772 41709 207773
rect 41643 207708 41644 207772
rect 41708 207708 41709 207772
rect 41643 207707 41709 207708
rect 40907 207364 40973 207365
rect 40907 207300 40908 207364
rect 40972 207300 40973 207364
rect 40907 207299 40973 207300
rect 40723 197164 40789 197165
rect 40723 197100 40724 197164
rect 40788 197100 40789 197164
rect 40723 197099 40789 197100
rect 40910 195533 40970 207299
rect 40907 195532 40973 195533
rect 40907 195468 40908 195532
rect 40972 195468 40973 195532
rect 40907 195467 40973 195468
rect 40539 194580 40605 194581
rect 40539 194516 40540 194580
rect 40604 194516 40605 194580
rect 40539 194515 40605 194516
rect 41459 194580 41525 194581
rect 41459 194516 41460 194580
rect 41524 194516 41525 194580
rect 41459 194515 41525 194516
rect 41462 187237 41522 194515
rect 41646 190470 41706 207707
rect 41827 197844 41893 197845
rect 41827 197780 41828 197844
rect 41892 197780 41893 197844
rect 41827 197779 41893 197780
rect 41830 195805 41890 197779
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 42014 195261 42074 210019
rect 42011 195260 42077 195261
rect 42011 195196 42012 195260
rect 42076 195196 42077 195260
rect 42011 195195 42077 195196
rect 42379 192948 42445 192949
rect 42379 192884 42380 192948
rect 42444 192884 42445 192948
rect 42379 192883 42445 192884
rect 41646 190410 41890 190470
rect 41459 187236 41525 187237
rect 41459 187172 41460 187236
rect 41524 187172 41525 187236
rect 41459 187171 41525 187172
rect 41830 185877 41890 190410
rect 42382 186285 42442 192883
rect 42379 186284 42445 186285
rect 42379 186220 42380 186284
rect 42444 186220 42445 186284
rect 42379 186219 42445 186220
rect 41827 185876 41893 185877
rect 41827 185812 41828 185876
rect 41892 185812 41893 185876
rect 41827 185811 41893 185812
rect 667982 130525 668042 212331
rect 671294 145213 671354 233139
rect 673315 228988 673381 228989
rect 673315 228924 673316 228988
rect 673380 228924 673381 228988
rect 673315 228923 673381 228924
rect 672947 228580 673013 228581
rect 672947 228516 672948 228580
rect 673012 228516 673013 228580
rect 672947 228515 673013 228516
rect 671659 226812 671725 226813
rect 671659 226748 671660 226812
rect 671724 226748 671725 226812
rect 671659 226747 671725 226748
rect 671662 224229 671722 226747
rect 671843 226676 671909 226677
rect 671843 226612 671844 226676
rect 671908 226612 671909 226676
rect 671843 226611 671909 226612
rect 671846 225181 671906 226611
rect 672027 226540 672093 226541
rect 672027 226476 672028 226540
rect 672092 226476 672093 226540
rect 672027 226475 672093 226476
rect 671843 225180 671909 225181
rect 671843 225116 671844 225180
rect 671908 225116 671909 225180
rect 671843 225115 671909 225116
rect 671659 224228 671725 224229
rect 671659 224164 671660 224228
rect 671724 224164 671725 224228
rect 671659 224163 671725 224164
rect 672030 217837 672090 226475
rect 672027 217836 672093 217837
rect 672027 217772 672028 217836
rect 672092 217772 672093 217836
rect 672027 217771 672093 217772
rect 672950 183565 673010 228515
rect 673131 226812 673197 226813
rect 673131 226748 673132 226812
rect 673196 226748 673197 226812
rect 673131 226747 673197 226748
rect 673134 218653 673194 226747
rect 673318 224909 673378 228923
rect 673683 226268 673749 226269
rect 673683 226204 673684 226268
rect 673748 226204 673749 226268
rect 673683 226203 673749 226204
rect 673315 224908 673381 224909
rect 673315 224844 673316 224908
rect 673380 224844 673381 224908
rect 673315 224843 673381 224844
rect 673499 223684 673565 223685
rect 673499 223620 673500 223684
rect 673564 223620 673565 223684
rect 673499 223619 673565 223620
rect 673131 218652 673197 218653
rect 673131 218588 673132 218652
rect 673196 218588 673197 218652
rect 673131 218587 673197 218588
rect 673131 210492 673197 210493
rect 673131 210428 673132 210492
rect 673196 210428 673197 210492
rect 673131 210427 673197 210428
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 673134 182069 673194 210427
rect 673315 203012 673381 203013
rect 673315 202948 673316 203012
rect 673380 202948 673381 203012
rect 673315 202947 673381 202948
rect 673131 182068 673197 182069
rect 673131 182004 673132 182068
rect 673196 182004 673197 182068
rect 673131 182003 673197 182004
rect 673318 147797 673378 202947
rect 673315 147796 673381 147797
rect 673315 147732 673316 147796
rect 673380 147732 673381 147796
rect 673315 147731 673381 147732
rect 671291 145212 671357 145213
rect 671291 145148 671292 145212
rect 671356 145148 671357 145212
rect 671291 145147 671357 145148
rect 667979 130524 668045 130525
rect 667979 130460 667980 130524
rect 668044 130460 668045 130524
rect 667979 130459 668045 130460
rect 673502 128485 673562 223619
rect 673686 143581 673746 226203
rect 674054 154597 674114 237083
rect 674787 228580 674853 228581
rect 674787 228516 674788 228580
rect 674852 228516 674853 228580
rect 674787 228515 674853 228516
rect 674790 218925 674850 228515
rect 675155 226540 675221 226541
rect 675155 226476 675156 226540
rect 675220 226476 675221 226540
rect 675155 226475 675221 226476
rect 674787 218924 674853 218925
rect 674787 218860 674788 218924
rect 674852 218860 674853 218924
rect 674787 218859 674853 218860
rect 675158 215525 675218 226475
rect 675523 218652 675589 218653
rect 675523 218588 675524 218652
rect 675588 218588 675589 218652
rect 675523 218587 675589 218588
rect 675155 215524 675221 215525
rect 675155 215460 675156 215524
rect 675220 215460 675221 215524
rect 675155 215459 675221 215460
rect 675526 210493 675586 218587
rect 676029 218244 676095 218245
rect 676029 218180 676030 218244
rect 676094 218180 676095 218244
rect 676029 218179 676095 218180
rect 676032 217970 676092 218179
rect 676032 217910 676322 217970
rect 676262 217290 676322 217910
rect 676262 217230 677058 217290
rect 675891 217020 675957 217021
rect 675891 216956 675892 217020
rect 675956 216956 675957 217020
rect 675891 216955 675957 216956
rect 675707 215388 675773 215389
rect 675707 215324 675708 215388
rect 675772 215324 675773 215388
rect 675707 215323 675773 215324
rect 675523 210492 675589 210493
rect 675523 210428 675524 210492
rect 675588 210428 675589 210492
rect 675523 210427 675589 210428
rect 675710 195261 675770 215323
rect 675894 211170 675954 216955
rect 676259 215150 676325 215151
rect 676259 215086 676260 215150
rect 676324 215086 676325 215150
rect 676259 215085 676325 215086
rect 675894 211110 676138 211170
rect 675891 210492 675957 210493
rect 675891 210428 675892 210492
rect 675956 210428 675957 210492
rect 675891 210427 675957 210428
rect 675707 195260 675773 195261
rect 675707 195196 675708 195260
rect 675772 195196 675773 195260
rect 675707 195195 675773 195196
rect 675894 193221 675954 210427
rect 675891 193220 675957 193221
rect 675891 193156 675892 193220
rect 675956 193156 675957 193220
rect 675891 193155 675957 193156
rect 676078 191589 676138 211110
rect 676262 197165 676322 215085
rect 676998 212550 677058 217230
rect 676630 212490 677058 212550
rect 676443 211444 676509 211445
rect 676443 211380 676444 211444
rect 676508 211380 676509 211444
rect 676443 211379 676509 211380
rect 676446 200837 676506 211379
rect 676630 205597 676690 212490
rect 676627 205596 676693 205597
rect 676627 205532 676628 205596
rect 676692 205532 676693 205596
rect 676627 205531 676693 205532
rect 676443 200836 676509 200837
rect 676443 200772 676444 200836
rect 676508 200772 676509 200836
rect 676443 200771 676509 200772
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675710 171050 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675710 170990 676138 171050
rect 675707 170372 675773 170373
rect 675707 170308 675708 170372
rect 675772 170308 675773 170372
rect 675707 170307 675773 170308
rect 675523 161396 675589 161397
rect 675523 161332 675524 161396
rect 675588 161332 675589 161396
rect 675523 161331 675589 161332
rect 675526 157045 675586 161331
rect 675523 157044 675589 157045
rect 675523 156980 675524 157044
rect 675588 156980 675589 157044
rect 675523 156979 675589 156980
rect 674051 154596 674117 154597
rect 674051 154532 674052 154596
rect 674116 154532 674117 154596
rect 674051 154531 674117 154532
rect 675710 150381 675770 170307
rect 675891 167516 675957 167517
rect 675891 167452 675892 167516
rect 675956 167452 675957 167516
rect 675891 167451 675957 167452
rect 675707 150380 675773 150381
rect 675707 150316 675708 150380
rect 675772 150316 675773 150380
rect 675707 150315 675773 150316
rect 675894 147661 675954 167451
rect 676078 148477 676138 170990
rect 676262 153101 676322 172350
rect 676446 159493 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159492 676509 159493
rect 676443 159428 676444 159492
rect 676508 159428 676509 159492
rect 676443 159427 676509 159428
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 153100 676325 153101
rect 676259 153036 676260 153100
rect 676324 153036 676325 153100
rect 676259 153035 676325 153036
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675891 147660 675957 147661
rect 675891 147596 675892 147660
rect 675956 147596 675957 147660
rect 675891 147595 675957 147596
rect 673683 143580 673749 143581
rect 673683 143516 673684 143580
rect 673748 143516 673749 143580
rect 673683 143515 673749 143516
rect 676627 128620 676693 128621
rect 676627 128556 676628 128620
rect 676692 128556 676693 128620
rect 676627 128555 676693 128556
rect 673499 128484 673565 128485
rect 673499 128420 673500 128484
rect 673564 128420 673565 128484
rect 673499 128419 673565 128420
rect 676075 128212 676141 128213
rect 676075 128148 676076 128212
rect 676140 128148 676141 128212
rect 676075 128147 676141 128148
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 122364 675773 122365
rect 675707 122300 675708 122364
rect 675772 122300 675773 122364
rect 675707 122299 675773 122300
rect 675710 102645 675770 122299
rect 675894 108085 675954 127195
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 128147
rect 676259 126988 676325 126989
rect 676259 126924 676260 126988
rect 676324 126924 676325 126988
rect 676259 126923 676325 126924
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676262 101421 676322 126923
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 106181 676506 124475
rect 676630 113117 676690 128555
rect 676627 113116 676693 113117
rect 676627 113052 676628 113116
rect 676692 113052 676693 113116
rect 676627 113051 676693 113052
rect 676443 106180 676509 106181
rect 676443 106116 676444 106180
rect 676508 106116 676509 106180
rect 676443 106115 676509 106116
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 634859 96932 634925 96933
rect 634859 96868 634860 96932
rect 634924 96868 634925 96932
rect 634859 96867 634925 96868
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 634862 80477 634922 96867
rect 637254 84210 637314 96867
rect 637070 84150 637314 84210
rect 634859 80476 634925 80477
rect 634859 80412 634860 80476
rect 634924 80412 634925 80476
rect 634859 80411 634925 80412
rect 637070 77893 637130 84150
rect 637067 77892 637133 77893
rect 637067 77828 637068 77892
rect 637132 77828 637133 77892
rect 637067 77827 637133 77828
rect 461715 55044 461781 55045
rect 461715 54980 461716 55044
rect 461780 54980 461781 55044
rect 461715 54979 461781 54980
rect 461718 53957 461778 54979
rect 461715 53956 461781 53957
rect 461715 53892 461716 53956
rect 461780 53892 461781 53956
rect 461715 53891 461781 53892
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 194366 42125 194426 50219
rect 308995 49740 309061 49741
rect 308995 49676 308996 49740
rect 309060 49676 309061 49740
rect 308995 49675 309061 49676
rect 308998 42805 309058 49675
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 461347 44436 461413 44437
rect 461347 44372 461348 44436
rect 461412 44372 461413 44436
rect 461347 44371 461413 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 440187 43892 440253 43893
rect 440187 43828 440188 43892
rect 440252 43890 440253 43892
rect 440923 43892 440989 43893
rect 440923 43890 440924 43892
rect 440252 43830 440924 43890
rect 440252 43828 440253 43830
rect 440187 43827 440253 43828
rect 440923 43828 440924 43830
rect 440988 43828 440989 43892
rect 440923 43827 440989 43828
rect 308995 42804 309061 42805
rect 308995 42740 308996 42804
rect 309060 42740 309061 42804
rect 308995 42739 309061 42740
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 421974 41850 422034 42059
rect 461350 41938 461410 44371
rect 462270 41938 462330 44371
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 421974 41790 422162 41850
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
<< via4 >>
rect 191702 997102 191938 997338
rect 226294 997102 226530 997338
rect 243222 997102 243458 997338
rect 278550 997102 278786 997338
rect 485550 997102 485786 997338
rect 503582 997102 503818 997338
rect 505238 997102 505474 997338
rect 533390 997102 533626 997338
rect 487390 219332 487626 219418
rect 487390 219268 487476 219332
rect 487476 219268 487540 219332
rect 487540 219268 487626 219332
rect 487390 219182 487626 219268
rect 491070 218652 491306 218738
rect 491070 218588 491156 218652
rect 491156 218588 491220 218652
rect 491220 218588 491306 218652
rect 573870 219182 574106 219418
rect 491070 218502 491306 218588
rect 578102 218502 578338 218738
rect 488862 217292 489098 217378
rect 488862 217228 488948 217292
rect 488948 217228 489012 217292
rect 489012 217228 489098 217292
rect 488862 217142 489098 217228
rect 575526 217142 575762 217378
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 191660 997338 226572 997380
rect 191660 997102 191702 997338
rect 191938 997102 226294 997338
rect 226530 997102 226572 997338
rect 191660 997060 226572 997102
rect 243180 997338 278828 997380
rect 243180 997102 243222 997338
rect 243458 997102 278550 997338
rect 278786 997102 278828 997338
rect 243180 997060 278828 997102
rect 485508 997338 503860 997380
rect 485508 997102 485550 997338
rect 485786 997102 503582 997338
rect 503818 997102 503860 997338
rect 485508 997060 503860 997102
rect 505196 997338 533668 997380
rect 505196 997102 505238 997338
rect 505474 997102 533390 997338
rect 533626 997102 533668 997338
rect 505196 997060 533668 997102
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 487348 219418 574148 219460
rect 487348 219182 487390 219418
rect 487626 219182 573870 219418
rect 574106 219182 574148 219418
rect 487348 219140 574148 219182
rect 491028 218738 578380 218780
rect 491028 218502 491070 218738
rect 491306 218502 578102 218738
rect 578338 218502 578380 218738
rect 491028 218460 578380 218502
rect 488820 217378 575804 217420
rect 488820 217142 488862 217378
rect 489098 217142 575526 217378
rect 575762 217142 575804 217378
rect 488820 217100 575804 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo
timestamp 0
transform 1 0 269370 0 1 5100
box 0 0 1 1
use caravel_motto  caravel_motto
timestamp 0
transform 1 0 -54372 0 1 -4446
box 0 0 1 1
use copyright_block  copyright_block
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206098 0 1 2054
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1665958328
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1665958328
transform 1 0 626764 0 1 63284
box 136 70 20000 12000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1665958328
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1665958328
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1665958328
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1665958328
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1665958328
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use simple_por  por
timestamp 1665958328
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1665958328
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1665958328
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1665958328
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1665958328
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1665958328
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1665958328
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1665958328
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1665958328
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1665958328
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1665958328
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1665958328
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1665958328
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1665958328
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1665958328
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1665958328
transform 1 0 588632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1665958328
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1665958328
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1665958328
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1665958328
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1665958328
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1665958328
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1665958328
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1665958328
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1665958328
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1665958328
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1665958328
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1665958328
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1665958328
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1665958328
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1665958328
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1665958328
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1665958328
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1665958328
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1665958328
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1665958328
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1665958328
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1665958328
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1665958328
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1665958328
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1665958328
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1665958328
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1665958328
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1665958328
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1665958328
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1665958328
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1665958328
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1665958328
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1665958328
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1665958328
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1665958328
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1665958328
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1665958328
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1665958328
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1665958328
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1665958328
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1665958328
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1665958328
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1665958328
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1665958328
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1665958328
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1665958328
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1665958328
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1665958328
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1665958328
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1665958328
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1665958328
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1665958328
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1665958328
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1665958328
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1665958328
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1665958328
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1665958328
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1665958328
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1665958328
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1665958328
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1665958328
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1665958328
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1665958328
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1665958328
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1665958328
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1665958328
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1665958328
transform 1 0 0 0 1 0
box 6022 33900 711814 1031696
use user_project_wrapper  mprj
timestamp 1665958328
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1665958328
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering  sigbuf
timestamp 1665958328
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal3 s 418245 997803 418551 997897 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal3 s 417057 997799 417363 997893 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
