magic
tech sky130A
magscale 1 2
timestamp 1666432150
<< metal1 >>
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 652018 896996 652024 897048
rect 652076 897036 652082 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 652076 897008 663794 897036
rect 652076 896996 652082 897008
rect 654778 895772 654784 895824
rect 654836 895812 654842 895824
rect 675846 895812 675852 895824
rect 654836 895784 675852 895812
rect 654836 895772 654842 895784
rect 675846 895772 675852 895784
rect 675904 895772 675910 895824
rect 672718 895636 672724 895688
rect 672776 895676 672782 895688
rect 676030 895676 676036 895688
rect 672776 895648 676036 895676
rect 672776 895636 672782 895648
rect 676030 895636 676036 895648
rect 676088 895636 676094 895688
rect 671982 894412 671988 894464
rect 672040 894452 672046 894464
rect 676030 894452 676036 894464
rect 672040 894424 676036 894452
rect 672040 894412 672046 894424
rect 676030 894412 676036 894424
rect 676088 894412 676094 894464
rect 671430 894276 671436 894328
rect 671488 894316 671494 894328
rect 675846 894316 675852 894328
rect 671488 894288 675852 894316
rect 671488 894276 671494 894288
rect 675846 894276 675852 894288
rect 675904 894276 675910 894328
rect 672350 892984 672356 893036
rect 672408 893024 672414 893036
rect 675846 893024 675852 893036
rect 672408 892996 675852 893024
rect 672408 892984 672414 892996
rect 675846 892984 675852 892996
rect 675904 892984 675910 893036
rect 673362 892848 673368 892900
rect 673420 892888 673426 892900
rect 676030 892888 676036 892900
rect 673420 892860 676036 892888
rect 673420 892848 673426 892860
rect 676030 892848 676036 892860
rect 676088 892848 676094 892900
rect 676214 891488 676220 891540
rect 676272 891528 676278 891540
rect 676858 891528 676864 891540
rect 676272 891500 676864 891528
rect 676272 891488 676278 891500
rect 676858 891488 676864 891500
rect 676916 891488 676922 891540
rect 676030 889992 676036 890044
rect 676088 890032 676094 890044
rect 677042 890032 677048 890044
rect 676088 890004 677048 890032
rect 676088 889992 676094 890004
rect 677042 889992 677048 890004
rect 677100 889992 677106 890044
rect 674374 888904 674380 888956
rect 674432 888944 674438 888956
rect 676030 888944 676036 888956
rect 674432 888916 676036 888944
rect 674432 888904 674438 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 674834 888700 674840 888752
rect 674892 888740 674898 888752
rect 675662 888740 675668 888752
rect 674892 888712 675668 888740
rect 674892 888700 674898 888712
rect 675662 888700 675668 888712
rect 675720 888700 675726 888752
rect 674650 888496 674656 888548
rect 674708 888536 674714 888548
rect 676030 888536 676036 888548
rect 674708 888508 676036 888536
rect 674708 888496 674714 888508
rect 676030 888496 676036 888508
rect 676088 888496 676094 888548
rect 674190 888088 674196 888140
rect 674248 888128 674254 888140
rect 676030 888128 676036 888140
rect 674248 888100 676036 888128
rect 674248 888088 674254 888100
rect 676030 888088 676036 888100
rect 676088 888088 676094 888140
rect 671798 886864 671804 886916
rect 671856 886904 671862 886916
rect 675478 886904 675484 886916
rect 671856 886876 675484 886904
rect 671856 886864 671862 886876
rect 675478 886864 675484 886876
rect 675536 886864 675542 886916
rect 673178 885640 673184 885692
rect 673236 885680 673242 885692
rect 676030 885680 676036 885692
rect 673236 885652 676036 885680
rect 673236 885640 673242 885652
rect 676030 885640 676036 885652
rect 676088 885640 676094 885692
rect 675202 881084 675208 881136
rect 675260 881124 675266 881136
rect 683298 881124 683304 881136
rect 675260 881096 683304 881124
rect 675260 881084 675266 881096
rect 683298 881084 683304 881096
rect 683356 881084 683362 881136
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 675570 880512 675576 880524
rect 653456 880484 675576 880512
rect 653456 880472 653462 880484
rect 675570 880472 675576 880484
rect 675628 880472 675634 880524
rect 675938 880132 675944 880184
rect 675996 880172 676002 880184
rect 679618 880172 679624 880184
rect 675996 880144 679624 880172
rect 675996 880132 676002 880144
rect 679618 880132 679624 880144
rect 679676 880132 679682 880184
rect 675754 879316 675760 879368
rect 675812 879356 675818 879368
rect 677042 879356 677048 879368
rect 675812 879328 677048 879356
rect 675812 879316 675818 879328
rect 677042 879316 677048 879328
rect 677100 879316 677106 879368
rect 674926 879112 674932 879164
rect 674984 879152 674990 879164
rect 678238 879152 678244 879164
rect 674984 879124 678244 879152
rect 674984 879112 674990 879124
rect 678238 879112 678244 879124
rect 678296 879112 678302 879164
rect 675386 878976 675392 879028
rect 675444 879016 675450 879028
rect 676858 879016 676864 879028
rect 675444 878988 676864 879016
rect 675444 878976 675450 878988
rect 676858 878976 676864 878988
rect 676916 878976 676922 879028
rect 675754 878364 675760 878416
rect 675812 878364 675818 878416
rect 675772 878200 675800 878364
rect 675588 878172 675800 878200
rect 675588 877384 675616 878172
rect 675496 877356 675616 877384
rect 675496 877260 675524 877356
rect 675478 877208 675484 877260
rect 675536 877208 675542 877260
rect 674190 873604 674196 873656
rect 674248 873644 674254 873656
rect 675110 873644 675116 873656
rect 674248 873616 675116 873644
rect 674248 873604 674254 873616
rect 675110 873604 675116 873616
rect 675168 873604 675174 873656
rect 674834 872380 674840 872432
rect 674892 872420 674898 872432
rect 675294 872420 675300 872432
rect 674892 872392 675300 872420
rect 674892 872380 674898 872392
rect 675294 872380 675300 872392
rect 675352 872380 675358 872432
rect 674650 869796 674656 869848
rect 674708 869836 674714 869848
rect 675202 869836 675208 869848
rect 674708 869808 675208 869836
rect 674708 869796 674714 869808
rect 675202 869796 675208 869808
rect 675260 869796 675266 869848
rect 674374 869592 674380 869644
rect 674432 869632 674438 869644
rect 674834 869632 674840 869644
rect 674432 869604 674840 869632
rect 674432 869592 674438 869604
rect 674834 869592 674840 869604
rect 674892 869592 674898 869644
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 675018 869428 675024 869440
rect 657596 869400 675024 869428
rect 657596 869388 657602 869400
rect 675018 869388 675024 869400
rect 675076 869388 675082 869440
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 674742 868068 674748 868080
rect 654192 868040 674748 868068
rect 654192 868028 654198 868040
rect 674742 868028 674748 868040
rect 674800 868028 674806 868080
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 46198 817136 46204 817148
rect 35860 817108 46204 817136
rect 35860 817096 35866 817108
rect 46198 817096 46204 817108
rect 46256 817096 46262 817148
rect 35618 816960 35624 817012
rect 35676 817000 35682 817012
rect 61378 817000 61384 817012
rect 35676 816972 61384 817000
rect 35676 816960 35682 816972
rect 61378 816960 61384 816972
rect 61436 816960 61442 817012
rect 35802 815736 35808 815788
rect 35860 815776 35866 815788
rect 44266 815776 44272 815788
rect 35860 815748 44272 815776
rect 35860 815736 35866 815748
rect 44266 815736 44272 815748
rect 44324 815736 44330 815788
rect 35434 815600 35440 815652
rect 35492 815640 35498 815652
rect 44818 815640 44824 815652
rect 35492 815612 44824 815640
rect 35492 815600 35498 815612
rect 44818 815600 44824 815612
rect 44876 815600 44882 815652
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 44542 814416 44548 814428
rect 35676 814388 44548 814416
rect 35676 814376 35682 814388
rect 44542 814376 44548 814388
rect 44600 814376 44606 814428
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 45094 814280 45100 814292
rect 35860 814252 45100 814280
rect 35860 814240 35866 814252
rect 45094 814240 45100 814252
rect 45152 814240 45158 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 43346 812852 43352 812864
rect 41380 812824 43352 812852
rect 41380 812812 41386 812824
rect 43346 812812 43352 812824
rect 43404 812812 43410 812864
rect 40954 810704 40960 810756
rect 41012 810744 41018 810756
rect 42518 810744 42524 810756
rect 41012 810716 42524 810744
rect 41012 810704 41018 810716
rect 42518 810704 42524 810716
rect 42576 810704 42582 810756
rect 41138 807440 41144 807492
rect 41196 807480 41202 807492
rect 43162 807480 43168 807492
rect 41196 807452 43168 807480
rect 41196 807440 41202 807452
rect 43162 807440 43168 807452
rect 43220 807440 43226 807492
rect 40954 807304 40960 807356
rect 41012 807344 41018 807356
rect 45278 807344 45284 807356
rect 41012 807316 45284 807344
rect 41012 807304 41018 807316
rect 45278 807304 45284 807316
rect 45336 807304 45342 807356
rect 31754 806624 31760 806676
rect 31812 806664 31818 806676
rect 35618 806664 35624 806676
rect 31812 806636 35624 806664
rect 31812 806624 31818 806636
rect 35618 806624 35624 806636
rect 35676 806624 35682 806676
rect 44818 806556 44824 806608
rect 44876 806596 44882 806608
rect 62758 806596 62764 806608
rect 44876 806568 62764 806596
rect 44876 806556 44882 806568
rect 62758 806556 62764 806568
rect 62816 806556 62822 806608
rect 44910 806420 44916 806472
rect 44968 806460 44974 806472
rect 45278 806460 45284 806472
rect 44968 806432 45284 806460
rect 44968 806420 44974 806432
rect 45278 806420 45284 806432
rect 45336 806420 45342 806472
rect 41322 805944 41328 805996
rect 41380 805984 41386 805996
rect 43806 805984 43812 805996
rect 41380 805956 43812 805984
rect 41380 805944 41386 805956
rect 43806 805944 43812 805956
rect 43864 805944 43870 805996
rect 35618 802612 35624 802664
rect 35676 802652 35682 802664
rect 42334 802652 42340 802664
rect 35676 802624 42340 802652
rect 35676 802612 35682 802624
rect 42334 802612 42340 802624
rect 42392 802612 42398 802664
rect 33042 802408 33048 802460
rect 33100 802448 33106 802460
rect 42150 802448 42156 802460
rect 33100 802420 42156 802448
rect 33100 802408 33106 802420
rect 42150 802408 42156 802420
rect 42208 802408 42214 802460
rect 33778 801252 33784 801304
rect 33836 801292 33842 801304
rect 39850 801292 39856 801304
rect 33836 801264 39856 801292
rect 33836 801252 33842 801264
rect 39850 801252 39856 801264
rect 39908 801252 39914 801304
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 40678 801088 40684 801100
rect 31076 801060 40684 801088
rect 31076 801048 31082 801060
rect 40678 801048 40684 801060
rect 40736 801048 40742 801100
rect 43530 799076 43536 799128
rect 43588 799116 43594 799128
rect 53098 799116 53104 799128
rect 43588 799088 53104 799116
rect 43588 799076 43594 799088
rect 53098 799076 53104 799088
rect 53156 799076 53162 799128
rect 42886 797648 42892 797700
rect 42944 797688 42950 797700
rect 57238 797688 57244 797700
rect 42944 797660 57244 797688
rect 42944 797648 42950 797660
rect 57238 797648 57244 797660
rect 57296 797648 57302 797700
rect 42242 796288 42248 796340
rect 42300 796328 42306 796340
rect 42886 796328 42892 796340
rect 42300 796300 42892 796328
rect 42300 796288 42306 796300
rect 42886 796288 42892 796300
rect 42944 796288 42950 796340
rect 43530 794996 43536 795048
rect 43588 795036 43594 795048
rect 44910 795036 44916 795048
rect 43588 795008 44916 795036
rect 43588 794996 43594 795008
rect 44910 794996 44916 795008
rect 44968 794996 44974 795048
rect 42242 794792 42248 794844
rect 42300 794832 42306 794844
rect 43070 794832 43076 794844
rect 42300 794804 43076 794832
rect 42300 794792 42306 794804
rect 43070 794792 43076 794804
rect 43128 794792 43134 794844
rect 42334 793772 42340 793824
rect 42392 793812 42398 793824
rect 43438 793812 43444 793824
rect 42392 793784 43444 793812
rect 42392 793772 42398 793784
rect 43438 793772 43444 793784
rect 43496 793772 43502 793824
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 671614 789352 671620 789404
rect 671672 789392 671678 789404
rect 675110 789392 675116 789404
rect 671672 789364 675116 789392
rect 671672 789352 671678 789364
rect 675110 789352 675116 789364
rect 675168 789352 675174 789404
rect 57238 789148 57244 789200
rect 57296 789188 57302 789200
rect 62114 789188 62120 789200
rect 57296 789160 62120 789188
rect 57296 789148 57302 789160
rect 62114 789148 62120 789160
rect 62172 789148 62178 789200
rect 42702 786632 42708 786684
rect 42760 786672 42766 786684
rect 62114 786672 62120 786684
rect 42760 786644 62120 786672
rect 42760 786632 42766 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 46198 785136 46204 785188
rect 46256 785176 46262 785188
rect 62114 785176 62120 785188
rect 46256 785148 62120 785176
rect 46256 785136 46262 785148
rect 62114 785136 62120 785148
rect 62172 785136 62178 785188
rect 672994 783844 673000 783896
rect 673052 783884 673058 783896
rect 675110 783884 675116 783896
rect 673052 783856 675116 783884
rect 673052 783844 673058 783856
rect 675110 783844 675116 783856
rect 675168 783844 675174 783896
rect 673730 782620 673736 782672
rect 673788 782660 673794 782672
rect 675110 782660 675116 782672
rect 673788 782632 675116 782660
rect 673788 782620 673794 782632
rect 675110 782620 675116 782632
rect 675168 782620 675174 782672
rect 669222 782484 669228 782536
rect 669280 782524 669286 782536
rect 675294 782524 675300 782536
rect 669280 782496 675300 782524
rect 669280 782484 669286 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 655514 781192 655520 781244
rect 655572 781232 655578 781244
rect 675018 781232 675024 781244
rect 655572 781204 675024 781232
rect 655572 781192 655578 781204
rect 675018 781192 675024 781204
rect 675076 781192 675082 781244
rect 673914 779968 673920 780020
rect 673972 780008 673978 780020
rect 675110 780008 675116 780020
rect 673972 779980 675116 780008
rect 673972 779968 673978 779980
rect 675110 779968 675116 779980
rect 675168 779968 675174 780020
rect 673546 778540 673552 778592
rect 673604 778580 673610 778592
rect 675294 778580 675300 778592
rect 673604 778552 675300 778580
rect 673604 778540 673610 778552
rect 675294 778540 675300 778552
rect 675352 778540 675358 778592
rect 655054 778336 655060 778388
rect 655112 778376 655118 778388
rect 675110 778376 675116 778388
rect 655112 778348 675116 778376
rect 655112 778336 655118 778348
rect 675110 778336 675116 778348
rect 675168 778336 675174 778388
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 674282 776976 674288 777028
rect 674340 777016 674346 777028
rect 675294 777016 675300 777028
rect 674340 776988 675300 777016
rect 674340 776976 674346 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 674650 775684 674656 775736
rect 674708 775724 674714 775736
rect 675110 775724 675116 775736
rect 674708 775696 675116 775724
rect 674708 775684 674714 775696
rect 675110 775684 675116 775696
rect 675168 775684 675174 775736
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 669958 775588 669964 775600
rect 651524 775560 669964 775588
rect 651524 775548 651530 775560
rect 669958 775548 669964 775560
rect 670016 775548 670022 775600
rect 672166 775548 672172 775600
rect 672224 775588 672230 775600
rect 675018 775588 675024 775600
rect 672224 775560 675024 775588
rect 672224 775548 672230 775560
rect 675018 775548 675024 775560
rect 675076 775548 675082 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 669774 774256 669780 774308
rect 669832 774296 669838 774308
rect 675110 774296 675116 774308
rect 669832 774268 675116 774296
rect 669832 774256 669838 774268
rect 675110 774256 675116 774268
rect 675168 774256 675174 774308
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 59998 774228 60004 774240
rect 42116 774200 60004 774228
rect 42116 774188 42122 774200
rect 59998 774188 60004 774200
rect 60056 774188 60062 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655054 773820 655060 773832
rect 651524 773792 655060 773820
rect 651524 773780 651530 773792
rect 655054 773780 655060 773792
rect 655112 773780 655118 773832
rect 35802 773304 35808 773356
rect 35860 773344 35866 773356
rect 41690 773344 41696 773356
rect 35860 773316 41696 773344
rect 35860 773304 35866 773316
rect 41690 773304 41696 773316
rect 41748 773304 41754 773356
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 41046 773140 41052 773152
rect 35860 773112 41052 773140
rect 35860 773100 35866 773112
rect 41046 773100 41052 773112
rect 41104 773100 41110 773152
rect 35618 772964 35624 773016
rect 35676 773004 35682 773016
rect 41506 773004 41512 773016
rect 35676 772976 41512 773004
rect 35676 772964 35682 772976
rect 41506 772964 41512 772976
rect 41564 772964 41570 773016
rect 35434 772828 35440 772880
rect 35492 772868 35498 772880
rect 41322 772868 41328 772880
rect 35492 772840 41328 772868
rect 35492 772828 35498 772840
rect 41322 772828 41328 772840
rect 41380 772828 41386 772880
rect 42058 772828 42064 772880
rect 42116 772868 42122 772880
rect 61378 772868 61384 772880
rect 42116 772840 61384 772868
rect 42116 772828 42122 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 35526 771808 35532 771860
rect 35584 771848 35590 771860
rect 39758 771848 39764 771860
rect 35584 771820 39764 771848
rect 35584 771808 35590 771820
rect 39758 771808 39764 771820
rect 39816 771808 39822 771860
rect 42058 771604 42064 771656
rect 42116 771644 42122 771656
rect 45094 771644 45100 771656
rect 42116 771616 45100 771644
rect 42116 771604 42122 771616
rect 45094 771604 45100 771616
rect 45152 771604 45158 771656
rect 35802 771536 35808 771588
rect 35860 771576 35866 771588
rect 41690 771576 41696 771588
rect 35860 771548 41696 771576
rect 35860 771536 35866 771548
rect 41690 771536 41696 771548
rect 41748 771536 41754 771588
rect 35342 771400 35348 771452
rect 35400 771440 35406 771452
rect 41690 771440 41696 771452
rect 35400 771412 41696 771440
rect 35400 771400 35406 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 42058 771400 42064 771452
rect 42116 771440 42122 771452
rect 44542 771440 44548 771452
rect 42116 771412 44548 771440
rect 42116 771400 42122 771412
rect 44542 771400 44548 771412
rect 44600 771400 44606 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 40310 770488 40316 770500
rect 35860 770460 40316 770488
rect 35860 770448 35866 770460
rect 40310 770448 40316 770460
rect 40368 770448 40374 770500
rect 41690 770284 41696 770296
rect 41386 770256 41696 770284
rect 35618 770176 35624 770228
rect 35676 770216 35682 770228
rect 41386 770216 41414 770256
rect 41690 770244 41696 770256
rect 41748 770244 41754 770296
rect 42058 770244 42064 770296
rect 42116 770284 42122 770296
rect 43254 770284 43260 770296
rect 42116 770256 43260 770284
rect 42116 770244 42122 770256
rect 43254 770244 43260 770256
rect 43312 770244 43318 770296
rect 35676 770188 41414 770216
rect 35676 770176 35682 770188
rect 35802 770040 35808 770092
rect 35860 770080 35866 770092
rect 41690 770080 41696 770092
rect 35860 770052 41696 770080
rect 35860 770040 35866 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44266 770080 44272 770092
rect 42116 770052 44272 770080
rect 42116 770040 42122 770052
rect 44266 770040 44272 770052
rect 44324 770040 44330 770092
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 39574 768992 39580 769004
rect 35860 768964 39580 768992
rect 35860 768952 35866 768964
rect 39574 768952 39580 768964
rect 39632 768952 39638 769004
rect 35526 768816 35532 768868
rect 35584 768856 35590 768868
rect 40678 768856 40684 768868
rect 35584 768828 40684 768856
rect 35584 768816 35590 768828
rect 40678 768816 40684 768828
rect 40736 768816 40742 768868
rect 35342 768680 35348 768732
rect 35400 768720 35406 768732
rect 41690 768720 41696 768732
rect 35400 768692 41696 768720
rect 35400 768680 35406 768692
rect 41690 768680 41696 768692
rect 41748 768680 41754 768732
rect 35802 767524 35808 767576
rect 35860 767564 35866 767576
rect 35860 767524 35894 767564
rect 35866 767496 35894 767524
rect 35866 767468 40080 767496
rect 35802 767320 35808 767372
rect 35860 767360 35866 767372
rect 36538 767360 36544 767372
rect 35860 767332 36544 767360
rect 35860 767320 35866 767332
rect 36538 767320 36544 767332
rect 36596 767320 36602 767372
rect 40052 767292 40080 767468
rect 41690 767292 41696 767304
rect 40052 767264 41696 767292
rect 41690 767252 41696 767264
rect 41748 767252 41754 767304
rect 35802 766096 35808 766148
rect 35860 766136 35866 766148
rect 41230 766136 41236 766148
rect 35860 766108 41236 766136
rect 35860 766096 35866 766108
rect 41230 766096 41236 766108
rect 41288 766096 41294 766148
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 40862 764844 40868 764856
rect 35860 764816 40868 764844
rect 35860 764804 35866 764816
rect 40862 764804 40868 764816
rect 40920 764804 40926 764856
rect 35802 764532 35808 764584
rect 35860 764572 35866 764584
rect 41506 764572 41512 764584
rect 35860 764544 41512 764572
rect 35860 764532 35866 764544
rect 41506 764532 41512 764544
rect 41564 764532 41570 764584
rect 35802 763308 35808 763360
rect 35860 763348 35866 763360
rect 39298 763348 39304 763360
rect 35860 763320 39304 763348
rect 35860 763308 35866 763320
rect 39298 763308 39304 763320
rect 39356 763308 39362 763360
rect 41506 763280 41512 763292
rect 39500 763252 41512 763280
rect 35618 763172 35624 763224
rect 35676 763212 35682 763224
rect 39500 763212 39528 763252
rect 41506 763240 41512 763252
rect 41564 763240 41570 763292
rect 35676 763184 39528 763212
rect 35676 763172 35682 763184
rect 35802 761880 35808 761932
rect 35860 761920 35866 761932
rect 38930 761920 38936 761932
rect 35860 761892 38936 761920
rect 35860 761880 35866 761892
rect 38930 761880 38936 761892
rect 38988 761880 38994 761932
rect 33042 760996 33048 761048
rect 33100 761036 33106 761048
rect 41506 761036 41512 761048
rect 33100 761008 41512 761036
rect 33100 760996 33106 761008
rect 41506 760996 41512 761008
rect 41564 760996 41570 761048
rect 35158 759636 35164 759688
rect 35216 759676 35222 759688
rect 40034 759676 40040 759688
rect 35216 759648 40040 759676
rect 35216 759636 35222 759648
rect 40034 759636 40040 759648
rect 40092 759636 40098 759688
rect 39298 757732 39304 757784
rect 39356 757772 39362 757784
rect 41598 757772 41604 757784
rect 39356 757744 41604 757772
rect 39356 757732 39362 757744
rect 41598 757732 41604 757744
rect 41656 757732 41662 757784
rect 44726 755488 44732 755540
rect 44784 755528 44790 755540
rect 62758 755528 62764 755540
rect 44784 755500 62764 755528
rect 44784 755488 44790 755500
rect 62758 755488 62764 755500
rect 62816 755488 62822 755540
rect 43438 754876 43444 754928
rect 43496 754916 43502 754928
rect 45278 754916 45284 754928
rect 43496 754888 45284 754916
rect 43496 754876 43502 754888
rect 45278 754876 45284 754888
rect 45336 754876 45342 754928
rect 42242 754264 42248 754316
rect 42300 754304 42306 754316
rect 44726 754304 44732 754316
rect 42300 754276 44732 754304
rect 42300 754264 42306 754276
rect 44726 754264 44732 754276
rect 44784 754264 44790 754316
rect 42242 753856 42248 753908
rect 42300 753896 42306 753908
rect 42978 753896 42984 753908
rect 42300 753868 42984 753896
rect 42300 753856 42306 753868
rect 42978 753856 42984 753868
rect 43036 753856 43042 753908
rect 43622 753652 43628 753704
rect 43680 753692 43686 753704
rect 45094 753692 45100 753704
rect 43680 753664 45100 753692
rect 43680 753652 43686 753664
rect 45094 753652 45100 753664
rect 45152 753652 45158 753704
rect 61378 746988 61384 747040
rect 61436 747028 61442 747040
rect 62390 747028 62396 747040
rect 61436 747000 62396 747028
rect 61436 746988 61442 747000
rect 62390 746988 62396 747000
rect 62448 746988 62454 747040
rect 45094 746512 45100 746564
rect 45152 746552 45158 746564
rect 62114 746552 62120 746564
rect 45152 746524 62120 746552
rect 45152 746512 45158 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 670786 745220 670792 745272
rect 670844 745260 670850 745272
rect 675018 745260 675024 745272
rect 670844 745232 675024 745260
rect 670844 745220 670850 745232
rect 675018 745220 675024 745232
rect 675076 745220 675082 745272
rect 42702 743996 42708 744048
rect 42760 744036 42766 744048
rect 42760 744008 45554 744036
rect 42760 743996 42766 744008
rect 45526 743900 45554 744008
rect 62114 743900 62120 743912
rect 45526 743872 62120 743900
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 671246 743792 671252 743844
rect 671304 743832 671310 743844
rect 675110 743832 675116 743844
rect 671304 743804 675116 743832
rect 671304 743792 671310 743804
rect 675110 743792 675116 743804
rect 675168 743792 675174 743844
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 59998 742364 60004 742416
rect 60056 742404 60062 742416
rect 62114 742404 62120 742416
rect 60056 742376 62120 742404
rect 60056 742364 60062 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 670142 739100 670148 739152
rect 670200 739140 670206 739152
rect 675386 739140 675392 739152
rect 670200 739112 675392 739140
rect 670200 739100 670206 739112
rect 675386 739100 675392 739112
rect 675444 739100 675450 739152
rect 674190 738624 674196 738676
rect 674248 738664 674254 738676
rect 675386 738664 675392 738676
rect 674248 738636 675392 738664
rect 674248 738624 674254 738636
rect 675386 738624 675392 738636
rect 675444 738624 675450 738676
rect 668394 736924 668400 736976
rect 668452 736964 668458 736976
rect 675294 736964 675300 736976
rect 668452 736936 675300 736964
rect 668452 736924 668458 736936
rect 675294 736924 675300 736936
rect 675352 736924 675358 736976
rect 652018 736176 652024 736228
rect 652076 736216 652082 736228
rect 653398 736216 653404 736228
rect 652076 736188 653404 736216
rect 652076 736176 652082 736188
rect 653398 736176 653404 736188
rect 653456 736176 653462 736228
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 667474 735604 667480 735616
rect 657596 735576 667480 735604
rect 657596 735564 657602 735576
rect 667474 735564 667480 735576
rect 667532 735564 667538 735616
rect 667474 734816 667480 734868
rect 667532 734856 667538 734868
rect 675202 734856 675208 734868
rect 667532 734828 675208 734856
rect 667532 734816 667538 734828
rect 675202 734816 675208 734828
rect 675260 734816 675266 734868
rect 673638 734272 673644 734324
rect 673696 734312 673702 734324
rect 675294 734312 675300 734324
rect 673696 734284 675300 734312
rect 673696 734272 673702 734284
rect 675294 734272 675300 734284
rect 675352 734272 675358 734324
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 670970 734176 670976 734188
rect 654836 734148 670976 734176
rect 654836 734136 654842 734148
rect 670970 734136 670976 734148
rect 671028 734136 671034 734188
rect 675294 733592 675300 733644
rect 675352 733592 675358 733644
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668578 733428 668584 733440
rect 651524 733400 668584 733428
rect 651524 733388 651530 733400
rect 668578 733388 668584 733400
rect 668636 733388 668642 733440
rect 675312 733304 675340 733592
rect 675294 733252 675300 733304
rect 675352 733252 675358 733304
rect 651466 732776 651472 732828
rect 651524 732816 651530 732828
rect 661678 732816 661684 732828
rect 651524 732788 661684 732816
rect 651524 732776 651530 732788
rect 661678 732776 661684 732788
rect 661736 732776 661742 732828
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 651466 731280 651472 731332
rect 651524 731320 651530 731332
rect 671246 731320 671252 731332
rect 651524 731292 671252 731320
rect 651524 731280 651530 731292
rect 671246 731280 671252 731292
rect 671304 731280 671310 731332
rect 672534 730464 672540 730516
rect 672592 730504 672598 730516
rect 675202 730504 675208 730516
rect 672592 730476 675208 730504
rect 672592 730464 672598 730476
rect 675202 730464 675208 730476
rect 675260 730464 675266 730516
rect 43438 730328 43444 730380
rect 43496 730368 43502 730380
rect 61378 730368 61384 730380
rect 43496 730340 61384 730368
rect 43496 730328 43502 730340
rect 61378 730328 61384 730340
rect 61436 730328 61442 730380
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 667842 729920 667848 729972
rect 667900 729960 667906 729972
rect 675202 729960 675208 729972
rect 667900 729932 675208 729960
rect 667900 729920 667906 729932
rect 675202 729920 675208 729932
rect 675260 729920 675266 729972
rect 42242 729308 42248 729360
rect 42300 729348 42306 729360
rect 62758 729348 62764 729360
rect 42300 729320 62764 729348
rect 42300 729308 42306 729320
rect 62758 729308 62764 729320
rect 62816 729308 62822 729360
rect 41322 729036 41328 729088
rect 41380 729076 41386 729088
rect 41690 729076 41696 729088
rect 41380 729048 41696 729076
rect 41380 729036 41386 729048
rect 41690 729036 41696 729048
rect 41748 729036 41754 729088
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 43070 728668 43076 728680
rect 42116 728640 43076 728668
rect 42116 728628 42122 728640
rect 43070 728628 43076 728640
rect 43128 728628 43134 728680
rect 670326 728628 670332 728680
rect 670384 728668 670390 728680
rect 675294 728668 675300 728680
rect 670384 728640 675300 728668
rect 670384 728628 670390 728640
rect 675294 728628 675300 728640
rect 675352 728628 675358 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 673178 728288 673184 728340
rect 673236 728328 673242 728340
rect 673236 728300 674176 728328
rect 673236 728288 673242 728300
rect 671798 728084 671804 728136
rect 671856 728124 671862 728136
rect 671856 728096 674058 728124
rect 671856 728084 671862 728096
rect 674650 727880 674656 727932
rect 674708 727920 674714 727932
rect 683298 727920 683304 727932
rect 674708 727892 683304 727920
rect 674708 727880 674714 727892
rect 683298 727880 683304 727892
rect 683356 727880 683362 727932
rect 672810 727812 672816 727864
rect 672868 727852 672874 727864
rect 673454 727852 673460 727864
rect 672868 727824 673460 727852
rect 672868 727812 672874 727824
rect 673454 727812 673460 727824
rect 673512 727812 673518 727864
rect 675110 727744 675116 727796
rect 675168 727784 675174 727796
rect 677318 727784 677324 727796
rect 675168 727756 677324 727784
rect 675168 727744 675174 727756
rect 677318 727744 677324 727756
rect 677376 727744 677382 727796
rect 675018 727608 675024 727660
rect 675076 727608 675082 727660
rect 40862 727404 40868 727456
rect 40920 727444 40926 727456
rect 41690 727444 41696 727456
rect 40920 727416 41696 727444
rect 40920 727404 40926 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 44542 727444 44548 727456
rect 42116 727416 44548 727444
rect 42116 727404 42122 727416
rect 44542 727404 44548 727416
rect 44600 727404 44606 727456
rect 674834 727404 674840 727456
rect 674892 727444 674898 727456
rect 675036 727444 675064 727608
rect 674892 727416 675064 727444
rect 674892 727404 674898 727416
rect 41322 727268 41328 727320
rect 41380 727308 41386 727320
rect 41690 727308 41696 727320
rect 41380 727280 41696 727308
rect 41380 727268 41386 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 45002 727308 45008 727320
rect 42116 727280 45008 727308
rect 42116 727268 42122 727280
rect 45002 727268 45008 727280
rect 45060 727268 45066 727320
rect 674650 727268 674656 727320
rect 674708 727308 674714 727320
rect 675018 727308 675024 727320
rect 674708 727280 675024 727308
rect 674708 727268 674714 727280
rect 675018 727268 675024 727280
rect 675076 727268 675082 727320
rect 674374 726588 674380 726640
rect 674432 726628 674438 726640
rect 683482 726628 683488 726640
rect 674432 726600 683488 726628
rect 674432 726588 674438 726600
rect 683482 726588 683488 726600
rect 683540 726588 683546 726640
rect 41322 726180 41328 726232
rect 41380 726220 41386 726232
rect 41690 726220 41696 726232
rect 41380 726192 41696 726220
rect 41380 726180 41386 726192
rect 41690 726180 41696 726192
rect 41748 726180 41754 726232
rect 41138 725908 41144 725960
rect 41196 725948 41202 725960
rect 41598 725948 41604 725960
rect 41196 725920 41604 725948
rect 41196 725908 41202 725920
rect 41598 725908 41604 725920
rect 41656 725908 41662 725960
rect 672810 723120 672816 723172
rect 672868 723160 672874 723172
rect 673546 723160 673552 723172
rect 672868 723132 673552 723160
rect 672868 723120 672874 723132
rect 673546 723120 673552 723132
rect 673604 723120 673610 723172
rect 673730 722168 673736 722220
rect 673788 722168 673794 722220
rect 673748 722084 673776 722168
rect 673730 722032 673736 722084
rect 673788 722032 673794 722084
rect 673914 721964 673920 722016
rect 673972 721964 673978 722016
rect 673932 721812 673960 721964
rect 673914 721760 673920 721812
rect 673972 721760 673978 721812
rect 675754 721692 675760 721744
rect 675812 721692 675818 721744
rect 675938 721692 675944 721744
rect 675996 721692 676002 721744
rect 675772 721268 675800 721692
rect 675956 721268 675984 721692
rect 675754 721216 675760 721268
rect 675812 721216 675818 721268
rect 675938 721216 675944 721268
rect 675996 721216 676002 721268
rect 675754 720808 675760 720860
rect 675812 720808 675818 720860
rect 675938 720808 675944 720860
rect 675996 720808 676002 720860
rect 673914 720536 673920 720588
rect 673972 720536 673978 720588
rect 673932 720452 673960 720536
rect 675772 720520 675800 720808
rect 675956 720520 675984 720808
rect 675754 720468 675760 720520
rect 675812 720468 675818 720520
rect 675938 720468 675944 720520
rect 675996 720468 676002 720520
rect 673914 720400 673920 720452
rect 673972 720400 673978 720452
rect 43070 719720 43076 719772
rect 43128 719720 43134 719772
rect 42886 719516 42892 719568
rect 42944 719556 42950 719568
rect 43088 719556 43116 719720
rect 42944 719528 43116 719556
rect 42944 719516 42950 719528
rect 42702 719380 42708 719432
rect 42760 719420 42766 719432
rect 43070 719420 43076 719432
rect 42760 719392 43076 719420
rect 42760 719380 42766 719392
rect 43070 719380 43076 719392
rect 43128 719380 43134 719432
rect 674282 716456 674288 716508
rect 674340 716496 674346 716508
rect 676030 716496 676036 716508
rect 674340 716468 676036 716496
rect 674340 716456 674346 716468
rect 676030 716456 676036 716468
rect 676088 716456 676094 716508
rect 653398 716252 653404 716304
rect 653456 716292 653462 716304
rect 674006 716292 674012 716304
rect 653456 716264 674012 716292
rect 653456 716252 653462 716264
rect 674006 716252 674012 716264
rect 674064 716252 674070 716304
rect 35158 715776 35164 715828
rect 35216 715816 35222 715828
rect 41690 715816 41696 715828
rect 35216 715788 41696 715816
rect 35216 715776 35222 715788
rect 41690 715776 41696 715788
rect 41748 715776 41754 715828
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 674006 715748 674012 715760
rect 670016 715720 674012 715748
rect 670016 715708 670022 715720
rect 674006 715708 674012 715720
rect 674064 715708 674070 715760
rect 33778 715640 33784 715692
rect 33836 715680 33842 715692
rect 40402 715680 40408 715692
rect 33836 715652 40408 715680
rect 33836 715640 33842 715652
rect 40402 715640 40408 715652
rect 40460 715640 40466 715692
rect 32950 715504 32956 715556
rect 33008 715544 33014 715556
rect 40586 715544 40592 715556
rect 33008 715516 40592 715544
rect 33008 715504 33014 715516
rect 40586 715504 40592 715516
rect 40644 715504 40650 715556
rect 671430 715300 671436 715352
rect 671488 715340 671494 715352
rect 674006 715340 674012 715352
rect 671488 715312 674012 715340
rect 671488 715300 671494 715312
rect 674006 715300 674012 715312
rect 674064 715300 674070 715352
rect 671062 714960 671068 715012
rect 671120 715000 671126 715012
rect 674006 715000 674012 715012
rect 671120 714972 674012 715000
rect 671120 714960 671126 714972
rect 674006 714960 674012 714972
rect 674064 714960 674070 715012
rect 674282 714892 674288 714944
rect 674340 714932 674346 714944
rect 676030 714932 676036 714944
rect 674340 714904 676036 714932
rect 674340 714892 674346 714904
rect 676030 714892 676036 714904
rect 676088 714892 676094 714944
rect 660298 714824 660304 714876
rect 660356 714864 660362 714876
rect 674006 714864 674012 714876
rect 660356 714836 674012 714864
rect 660356 714824 660362 714836
rect 674006 714824 674012 714836
rect 674064 714824 674070 714876
rect 671982 714484 671988 714536
rect 672040 714524 672046 714536
rect 674006 714524 674012 714536
rect 672040 714496 674012 714524
rect 672040 714484 672046 714496
rect 674006 714484 674012 714496
rect 674064 714484 674070 714536
rect 672350 713668 672356 713720
rect 672408 713708 672414 713720
rect 674006 713708 674012 713720
rect 672408 713680 674012 713708
rect 672408 713668 672414 713680
rect 674006 713668 674012 713680
rect 674064 713668 674070 713720
rect 671338 713192 671344 713244
rect 671396 713232 671402 713244
rect 674006 713232 674012 713244
rect 671396 713204 674012 713232
rect 671396 713192 671402 713204
rect 674006 713192 674012 713204
rect 674064 713192 674070 713244
rect 671154 712376 671160 712428
rect 671212 712416 671218 712428
rect 674006 712416 674012 712428
rect 671212 712388 674012 712416
rect 671212 712376 671218 712388
rect 674006 712376 674012 712388
rect 674064 712376 674070 712428
rect 42886 712104 42892 712156
rect 42944 712144 42950 712156
rect 50338 712144 50344 712156
rect 42944 712116 50344 712144
rect 42944 712104 42950 712116
rect 50338 712104 50344 712116
rect 50396 712104 50402 712156
rect 676214 712036 676220 712088
rect 676272 712076 676278 712088
rect 677318 712076 677324 712088
rect 676272 712048 677324 712076
rect 676272 712036 676278 712048
rect 677318 712036 677324 712048
rect 677376 712036 677382 712088
rect 672166 709996 672172 710048
rect 672224 710036 672230 710048
rect 674006 710036 674012 710048
rect 672224 710008 674012 710036
rect 672224 709996 672230 710008
rect 674006 709996 674012 710008
rect 674064 709996 674070 710048
rect 42242 709724 42248 709776
rect 42300 709764 42306 709776
rect 44634 709764 44640 709776
rect 42300 709736 44640 709764
rect 42300 709724 42306 709736
rect 44634 709724 44640 709736
rect 44692 709724 44698 709776
rect 671614 709588 671620 709640
rect 671672 709628 671678 709640
rect 674006 709628 674012 709640
rect 671672 709600 674012 709628
rect 671672 709588 671678 709600
rect 674006 709588 674012 709600
rect 674064 709588 674070 709640
rect 674282 709520 674288 709572
rect 674340 709560 674346 709572
rect 676030 709560 676036 709572
rect 674340 709532 676036 709560
rect 674340 709520 674346 709532
rect 676030 709520 676036 709532
rect 676088 709520 676094 709572
rect 669222 709316 669228 709368
rect 669280 709356 669286 709368
rect 674006 709356 674012 709368
rect 669280 709328 674012 709356
rect 669280 709316 669286 709328
rect 674006 709316 674012 709328
rect 674064 709316 674070 709368
rect 42242 707956 42248 708008
rect 42300 707996 42306 708008
rect 44634 707996 44640 708008
rect 42300 707968 44640 707996
rect 42300 707956 42306 707968
rect 44634 707956 44640 707968
rect 44692 707956 44698 708008
rect 674282 707956 674288 708008
rect 674340 707996 674346 708008
rect 675846 707996 675852 708008
rect 674340 707968 675852 707996
rect 674340 707956 674346 707968
rect 675846 707956 675852 707968
rect 675904 707956 675910 708008
rect 674466 707548 674472 707600
rect 674524 707588 674530 707600
rect 676030 707588 676036 707600
rect 674524 707560 676036 707588
rect 674524 707548 674530 707560
rect 676030 707548 676036 707560
rect 676088 707548 676094 707600
rect 674650 707140 674656 707192
rect 674708 707180 674714 707192
rect 676030 707180 676036 707192
rect 674708 707152 676036 707180
rect 674708 707140 674714 707152
rect 676030 707140 676036 707152
rect 676088 707140 676094 707192
rect 42242 705508 42248 705560
rect 42300 705548 42306 705560
rect 43622 705548 43628 705560
rect 42300 705520 43628 705548
rect 42300 705508 42306 705520
rect 43622 705508 43628 705520
rect 43680 705508 43686 705560
rect 669774 705372 669780 705424
rect 669832 705412 669838 705424
rect 674006 705412 674012 705424
rect 669832 705384 674012 705412
rect 669832 705372 669838 705384
rect 674006 705372 674012 705384
rect 674064 705372 674070 705424
rect 674282 705304 674288 705356
rect 674340 705344 674346 705356
rect 683114 705344 683120 705356
rect 674340 705316 683120 705344
rect 674340 705304 674346 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 50338 705100 50344 705152
rect 50396 705140 50402 705152
rect 62114 705140 62120 705152
rect 50396 705112 62120 705140
rect 50396 705100 50402 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 669222 703808 669228 703860
rect 669280 703848 669286 703860
rect 674006 703848 674012 703860
rect 669280 703820 674012 703848
rect 669280 703808 669286 703820
rect 674006 703808 674012 703820
rect 674064 703808 674070 703860
rect 674282 703808 674288 703860
rect 674340 703848 674346 703860
rect 676030 703848 676036 703860
rect 674340 703820 676036 703848
rect 674340 703808 674346 703820
rect 676030 703808 676036 703820
rect 676088 703808 676094 703860
rect 44450 703740 44456 703792
rect 44508 703780 44514 703792
rect 62114 703780 62120 703792
rect 44508 703752 62120 703780
rect 44508 703740 44514 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 673454 701428 673460 701480
rect 673512 701468 673518 701480
rect 673914 701468 673920 701480
rect 673512 701440 673920 701468
rect 673512 701428 673518 701440
rect 673914 701428 673920 701440
rect 673972 701428 673978 701480
rect 666462 701224 666468 701276
rect 666520 701264 666526 701276
rect 674006 701264 674012 701276
rect 666520 701236 674012 701264
rect 666520 701224 666526 701236
rect 674006 701224 674012 701236
rect 674064 701224 674070 701276
rect 674282 701224 674288 701276
rect 674340 701264 674346 701276
rect 675110 701264 675116 701276
rect 674340 701236 675116 701264
rect 674340 701224 674346 701236
rect 675110 701224 675116 701236
rect 675168 701224 675174 701276
rect 42702 701020 42708 701072
rect 42760 701060 42766 701072
rect 62206 701060 62212 701072
rect 42760 701032 62212 701060
rect 42760 701020 42766 701032
rect 62206 701020 62212 701032
rect 62264 701020 62270 701072
rect 654778 701020 654784 701072
rect 654836 701060 654842 701072
rect 674006 701060 674012 701072
rect 654836 701032 674012 701060
rect 654836 701020 654842 701032
rect 674006 701020 674012 701032
rect 674064 701020 674070 701072
rect 674282 701020 674288 701072
rect 674340 701060 674346 701072
rect 675386 701060 675392 701072
rect 674340 701032 675392 701060
rect 674340 701020 674346 701032
rect 675386 701020 675392 701032
rect 675444 701020 675450 701072
rect 42886 700408 42892 700460
rect 42944 700408 42950 700460
rect 42904 700244 42932 700408
rect 43070 700340 43076 700392
rect 43128 700380 43134 700392
rect 43128 700352 43300 700380
rect 43128 700340 43134 700352
rect 43070 700244 43076 700256
rect 42904 700216 43076 700244
rect 43070 700204 43076 700216
rect 43128 700204 43134 700256
rect 42886 700068 42892 700120
rect 42944 700108 42950 700120
rect 43272 700108 43300 700352
rect 42944 700080 43300 700108
rect 42944 700068 42950 700080
rect 46198 698164 46204 698216
rect 46256 698204 46262 698216
rect 62114 698204 62120 698216
rect 46256 698176 62120 698204
rect 46256 698164 46262 698176
rect 62114 698164 62120 698176
rect 62172 698164 62178 698216
rect 666278 696940 666284 696992
rect 666336 696980 666342 696992
rect 673730 696980 673736 696992
rect 666336 696952 673736 696980
rect 666336 696940 666342 696952
rect 673730 696940 673736 696952
rect 673788 696940 673794 696992
rect 674466 693472 674472 693524
rect 674524 693512 674530 693524
rect 675386 693512 675392 693524
rect 674524 693484 675392 693512
rect 674524 693472 674530 693484
rect 675386 693472 675392 693484
rect 675444 693472 675450 693524
rect 674282 692996 674288 693048
rect 674340 693036 674346 693048
rect 675110 693036 675116 693048
rect 674340 693008 675116 693036
rect 674340 692996 674346 693008
rect 675110 692996 675116 693008
rect 675168 692996 675174 693048
rect 656434 690072 656440 690124
rect 656492 690112 656498 690124
rect 673730 690112 673736 690124
rect 656492 690084 673736 690112
rect 656492 690072 656498 690084
rect 673730 690072 673736 690084
rect 673788 690072 673794 690124
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 673730 688820 673736 688832
rect 652812 688792 673736 688820
rect 652812 688780 652818 688792
rect 673730 688780 673736 688792
rect 673788 688780 673794 688832
rect 651466 688644 651472 688696
rect 651524 688684 651530 688696
rect 657538 688684 657544 688696
rect 651524 688656 657544 688684
rect 651524 688644 651530 688656
rect 657538 688644 657544 688656
rect 657596 688644 657602 688696
rect 42702 687284 42708 687336
rect 42760 687324 42766 687336
rect 42760 687296 51074 687324
rect 42760 687284 42766 687296
rect 51046 687256 51074 687296
rect 61378 687256 61384 687268
rect 51046 687228 61384 687256
rect 61378 687216 61384 687228
rect 61436 687216 61442 687268
rect 651466 687216 651472 687268
rect 651524 687256 651530 687268
rect 669958 687256 669964 687268
rect 651524 687228 669964 687256
rect 651524 687216 651530 687228
rect 669958 687216 669964 687228
rect 670016 687216 670022 687268
rect 651466 687012 651472 687064
rect 651524 687052 651530 687064
rect 654778 687052 654784 687064
rect 651524 687024 654784 687052
rect 651524 687012 651530 687024
rect 654778 687012 654784 687024
rect 654836 687012 654842 687064
rect 43438 686468 43444 686520
rect 43496 686508 43502 686520
rect 62758 686508 62764 686520
rect 43496 686480 62764 686508
rect 43496 686468 43502 686480
rect 62758 686468 62764 686480
rect 62816 686468 62822 686520
rect 651650 686468 651656 686520
rect 651708 686508 651714 686520
rect 667198 686508 667204 686520
rect 651708 686480 667204 686508
rect 651708 686468 651714 686480
rect 667198 686468 667204 686480
rect 667256 686468 667262 686520
rect 41322 686264 41328 686316
rect 41380 686304 41386 686316
rect 41690 686304 41696 686316
rect 41380 686276 41696 686304
rect 41380 686264 41386 686276
rect 41690 686264 41696 686276
rect 41748 686264 41754 686316
rect 42058 686264 42064 686316
rect 42116 686304 42122 686316
rect 43070 686304 43076 686316
rect 42116 686276 43076 686304
rect 42116 686264 42122 686276
rect 43070 686264 43076 686276
rect 43128 686264 43134 686316
rect 41138 686060 41144 686112
rect 41196 686100 41202 686112
rect 41690 686100 41696 686112
rect 41196 686072 41696 686100
rect 41196 686060 41202 686072
rect 41690 686060 41696 686072
rect 41748 686060 41754 686112
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 45186 686100 45192 686112
rect 42116 686072 45192 686100
rect 42116 686060 42122 686072
rect 45186 686060 45192 686072
rect 45244 686060 45250 686112
rect 40862 685856 40868 685908
rect 40920 685896 40926 685908
rect 41690 685896 41696 685908
rect 40920 685868 41696 685896
rect 40920 685856 40926 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45186 685896 45192 685908
rect 42116 685868 45192 685896
rect 42116 685856 42122 685868
rect 45186 685856 45192 685868
rect 45244 685856 45250 685908
rect 668762 685856 668768 685908
rect 668820 685896 668826 685908
rect 672166 685896 672172 685908
rect 668820 685868 672172 685896
rect 668820 685856 668826 685868
rect 672166 685856 672172 685868
rect 672224 685856 672230 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656434 685556 656440 685568
rect 651524 685528 656440 685556
rect 651524 685516 651530 685528
rect 656434 685516 656440 685528
rect 656492 685516 656498 685568
rect 41046 684700 41052 684752
rect 41104 684740 41110 684752
rect 41690 684740 41696 684752
rect 41104 684712 41696 684740
rect 41104 684700 41110 684712
rect 41690 684700 41696 684712
rect 41748 684700 41754 684752
rect 41322 683408 41328 683460
rect 41380 683448 41386 683460
rect 41690 683448 41696 683460
rect 41380 683420 41696 683448
rect 41380 683408 41386 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 42058 683408 42064 683460
rect 42116 683448 42122 683460
rect 42702 683448 42708 683460
rect 42116 683420 42708 683448
rect 42116 683408 42122 683420
rect 42702 683408 42708 683420
rect 42760 683408 42766 683460
rect 41138 683272 41144 683324
rect 41196 683312 41202 683324
rect 41690 683312 41696 683324
rect 41196 683284 41696 683312
rect 41196 683272 41202 683284
rect 41690 683272 41696 683284
rect 41748 683272 41754 683324
rect 42058 683272 42064 683324
rect 42116 683312 42122 683324
rect 44266 683312 44272 683324
rect 42116 683284 44272 683312
rect 42116 683272 42122 683284
rect 44266 683272 44272 683284
rect 44324 683272 44330 683324
rect 40770 683136 40776 683188
rect 40828 683176 40834 683188
rect 41690 683176 41696 683188
rect 40828 683148 41696 683176
rect 40828 683136 40834 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 42058 683136 42064 683188
rect 42116 683176 42122 683188
rect 45002 683176 45008 683188
rect 42116 683148 45008 683176
rect 42116 683136 42122 683148
rect 45002 683136 45008 683148
rect 45060 683136 45066 683188
rect 674558 682388 674564 682440
rect 674616 682428 674622 682440
rect 683206 682428 683212 682440
rect 674616 682400 683212 682428
rect 674616 682388 674622 682400
rect 683206 682388 683212 682400
rect 683264 682388 683270 682440
rect 41322 681980 41328 682032
rect 41380 682020 41386 682032
rect 41690 682020 41696 682032
rect 41380 681992 41696 682020
rect 41380 681980 41386 681992
rect 41690 681980 41696 681992
rect 41748 681980 41754 682032
rect 42058 681980 42064 682032
rect 42116 682020 42122 682032
rect 42518 682020 42524 682032
rect 42116 681992 42524 682020
rect 42116 681980 42122 681992
rect 42518 681980 42524 681992
rect 42576 681980 42582 682032
rect 40954 679124 40960 679176
rect 41012 679164 41018 679176
rect 41322 679164 41328 679176
rect 41012 679136 41328 679164
rect 41012 679124 41018 679136
rect 41322 679124 41328 679136
rect 41380 679124 41386 679176
rect 41138 678988 41144 679040
rect 41196 679028 41202 679040
rect 41690 679028 41696 679040
rect 41196 679000 41696 679028
rect 41196 678988 41202 679000
rect 41690 678988 41696 679000
rect 41748 678988 41754 679040
rect 42058 678988 42064 679040
rect 42116 679028 42122 679040
rect 45002 679028 45008 679040
rect 42116 679000 45008 679028
rect 42116 678988 42122 679000
rect 45002 678988 45008 679000
rect 45060 678988 45066 679040
rect 40954 677696 40960 677748
rect 41012 677736 41018 677748
rect 41598 677736 41604 677748
rect 41012 677708 41604 677736
rect 41012 677696 41018 677708
rect 41598 677696 41604 677708
rect 41656 677696 41662 677748
rect 35158 672868 35164 672920
rect 35216 672908 35222 672920
rect 38838 672908 38844 672920
rect 35216 672880 38844 672908
rect 35216 672868 35222 672880
rect 38838 672868 38844 672880
rect 38896 672868 38902 672920
rect 33778 672732 33784 672784
rect 33836 672772 33842 672784
rect 37918 672772 37924 672784
rect 33836 672744 37924 672772
rect 33836 672732 33842 672744
rect 37918 672732 37924 672744
rect 37976 672732 37982 672784
rect 42426 671508 42432 671560
rect 42484 671508 42490 671560
rect 42444 671412 42472 671508
rect 42444 671384 42564 671412
rect 42536 671140 42564 671384
rect 42702 671140 42708 671152
rect 42536 671112 42708 671140
rect 42702 671100 42708 671112
rect 42760 671100 42766 671152
rect 668578 671100 668584 671152
rect 668636 671140 668642 671152
rect 673914 671140 673920 671152
rect 668636 671112 673920 671140
rect 668636 671100 668642 671112
rect 673914 671100 673920 671112
rect 673972 671100 673978 671152
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673546 670732 673552 670744
rect 661736 670704 673552 670732
rect 661736 670692 661742 670704
rect 673546 670692 673552 670704
rect 673604 670692 673610 670744
rect 670970 670080 670976 670132
rect 671028 670120 671034 670132
rect 673914 670120 673920 670132
rect 671028 670092 673920 670120
rect 671028 670080 671034 670092
rect 673914 670080 673920 670092
rect 673972 670080 673978 670132
rect 658918 669468 658924 669520
rect 658976 669508 658982 669520
rect 673546 669508 673552 669520
rect 658976 669480 673552 669508
rect 658976 669468 658982 669480
rect 673546 669468 673552 669480
rect 673604 669468 673610 669520
rect 45370 669332 45376 669384
rect 45428 669372 45434 669384
rect 53098 669372 53104 669384
rect 45428 669344 53104 669372
rect 45428 669332 45434 669344
rect 53098 669332 53104 669344
rect 53156 669332 53162 669384
rect 669590 669332 669596 669384
rect 669648 669372 669654 669384
rect 673914 669372 673920 669384
rect 669648 669344 673920 669372
rect 669648 669332 669654 669344
rect 673914 669332 673920 669344
rect 673972 669332 673978 669384
rect 671338 668516 671344 668568
rect 671396 668556 671402 668568
rect 673914 668556 673920 668568
rect 671396 668528 673920 668556
rect 671396 668516 671402 668528
rect 673914 668516 673920 668528
rect 673972 668516 673978 668568
rect 671522 668176 671528 668228
rect 671580 668216 671586 668228
rect 673546 668216 673552 668228
rect 671580 668188 673552 668216
rect 671580 668176 671586 668188
rect 673546 668176 673552 668188
rect 673604 668176 673610 668228
rect 45738 667904 45744 667956
rect 45796 667944 45802 667956
rect 57238 667944 57244 667956
rect 45796 667916 57244 667944
rect 45796 667904 45802 667916
rect 57238 667904 57244 667916
rect 57296 667904 57302 667956
rect 671338 667904 671344 667956
rect 671396 667944 671402 667956
rect 673914 667944 673920 667956
rect 671396 667916 673920 667944
rect 671396 667904 671402 667916
rect 673914 667904 673920 667916
rect 673972 667904 673978 667956
rect 42242 667428 42248 667480
rect 42300 667468 42306 667480
rect 45370 667468 45376 667480
rect 42300 667440 45376 667468
rect 42300 667428 42306 667440
rect 45370 667428 45376 667440
rect 45428 667428 45434 667480
rect 671154 666884 671160 666936
rect 671212 666924 671218 666936
rect 673914 666924 673920 666936
rect 671212 666896 673920 666924
rect 671212 666884 671218 666896
rect 673914 666884 673920 666896
rect 673972 666884 673978 666936
rect 669406 666544 669412 666596
rect 669464 666584 669470 666596
rect 673546 666584 673552 666596
rect 669464 666556 673552 666584
rect 669464 666544 669470 666556
rect 673546 666544 673552 666556
rect 673604 666544 673610 666596
rect 670878 666000 670884 666052
rect 670936 666040 670942 666052
rect 673914 666040 673920 666052
rect 670936 666012 673920 666040
rect 670936 666000 670942 666012
rect 673914 666000 673920 666012
rect 673972 666000 673978 666052
rect 42334 665796 42340 665848
rect 42392 665836 42398 665848
rect 45738 665836 45744 665848
rect 42392 665808 45744 665836
rect 42392 665796 42398 665808
rect 45738 665796 45744 665808
rect 45796 665796 45802 665848
rect 42242 665388 42248 665440
rect 42300 665428 42306 665440
rect 43990 665428 43996 665440
rect 42300 665400 43996 665428
rect 42300 665388 42306 665400
rect 43990 665388 43996 665400
rect 44048 665388 44054 665440
rect 672534 665388 672540 665440
rect 672592 665428 672598 665440
rect 673546 665428 673552 665440
rect 672592 665400 673552 665428
rect 672592 665388 672598 665400
rect 673546 665388 673552 665400
rect 673604 665388 673610 665440
rect 668946 665184 668952 665236
rect 669004 665224 669010 665236
rect 673914 665224 673920 665236
rect 669004 665196 673920 665224
rect 669004 665184 669010 665196
rect 673914 665184 673920 665196
rect 673972 665184 673978 665236
rect 670326 664436 670332 664488
rect 670384 664476 670390 664488
rect 673914 664476 673920 664488
rect 670384 664448 673920 664476
rect 670384 664436 670390 664448
rect 673914 664436 673920 664448
rect 673972 664436 673978 664488
rect 670142 663960 670148 664012
rect 670200 664000 670206 664012
rect 673914 664000 673920 664012
rect 670200 663972 673920 664000
rect 670200 663960 670206 663972
rect 673914 663960 673920 663972
rect 673972 663960 673978 664012
rect 674926 663960 674932 664012
rect 674984 664000 674990 664012
rect 676214 664000 676220 664012
rect 674984 663972 676220 664000
rect 674984 663960 674990 663972
rect 676214 663960 676220 663972
rect 676272 663960 676278 664012
rect 42426 663552 42432 663604
rect 42484 663552 42490 663604
rect 42444 663128 42472 663552
rect 42426 663076 42432 663128
rect 42484 663076 42490 663128
rect 668394 661920 668400 661972
rect 668452 661960 668458 661972
rect 673914 661960 673920 661972
rect 668452 661932 673920 661960
rect 668452 661920 668458 661932
rect 673914 661920 673920 661932
rect 673972 661920 673978 661972
rect 670510 661580 670516 661632
rect 670568 661620 670574 661632
rect 673914 661620 673920 661632
rect 670568 661592 673920 661620
rect 670568 661580 670574 661592
rect 673914 661580 673920 661592
rect 673972 661580 673978 661632
rect 667382 661104 667388 661156
rect 667440 661144 667446 661156
rect 673914 661144 673920 661156
rect 667440 661116 673920 661144
rect 667440 661104 667446 661116
rect 673914 661104 673920 661116
rect 673972 661104 673978 661156
rect 53098 660900 53104 660952
rect 53156 660940 53162 660952
rect 62114 660940 62120 660952
rect 53156 660912 62120 660940
rect 53156 660900 53162 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43622 660532 43628 660544
rect 42208 660504 43628 660532
rect 42208 660492 42214 660504
rect 43622 660492 43628 660504
rect 43680 660492 43686 660544
rect 667842 660152 667848 660204
rect 667900 660192 667906 660204
rect 673914 660192 673920 660204
rect 667900 660164 673920 660192
rect 667900 660152 667906 660164
rect 673914 660152 673920 660164
rect 673972 660152 673978 660204
rect 674558 659812 674564 659864
rect 674616 659852 674622 659864
rect 683114 659852 683120 659864
rect 674616 659824 683120 659852
rect 674616 659812 674622 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 672166 659676 672172 659728
rect 672224 659716 672230 659728
rect 673914 659716 673920 659728
rect 672224 659688 673920 659716
rect 672224 659676 672230 659688
rect 673914 659676 673920 659688
rect 673972 659676 673978 659728
rect 57238 659540 57244 659592
rect 57296 659580 57302 659592
rect 62114 659580 62120 659592
rect 57296 659552 62120 659580
rect 57296 659540 57302 659552
rect 62114 659540 62120 659552
rect 62172 659540 62178 659592
rect 62114 657540 62120 657552
rect 45526 657512 62120 657540
rect 42518 657228 42524 657280
rect 42576 657268 42582 657280
rect 45526 657268 45554 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 42576 657240 45554 657268
rect 42576 657228 42582 657240
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 673914 655568 673920 655580
rect 653456 655540 673920 655568
rect 653456 655528 653462 655540
rect 673914 655528 673920 655540
rect 673972 655528 673978 655580
rect 44818 655460 44824 655512
rect 44876 655500 44882 655512
rect 62114 655500 62120 655512
rect 44876 655472 62120 655500
rect 44876 655460 44882 655472
rect 62114 655460 62120 655472
rect 62172 655460 62178 655512
rect 667566 647232 667572 647284
rect 667624 647272 667630 647284
rect 674006 647272 674012 647284
rect 667624 647244 674012 647272
rect 667624 647232 667630 647244
rect 674006 647232 674012 647244
rect 674064 647232 674070 647284
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 670970 645912 670976 645924
rect 655572 645884 670976 645912
rect 655572 645872 655578 645884
rect 670970 645872 670976 645884
rect 671028 645872 671034 645924
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 41690 644484 41696 644496
rect 35860 644456 41696 644484
rect 35860 644444 35866 644456
rect 41690 644444 41696 644456
rect 41748 644444 41754 644496
rect 42058 644444 42064 644496
rect 42116 644484 42122 644496
rect 59998 644484 60004 644496
rect 42116 644456 60004 644484
rect 42116 644444 42122 644456
rect 59998 644444 60004 644456
rect 60056 644444 60062 644496
rect 674926 643560 674932 643612
rect 674984 643560 674990 643612
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 40494 643532 40500 643544
rect 35860 643504 40500 643532
rect 35860 643492 35866 643504
rect 40494 643492 40500 643504
rect 40552 643492 40558 643544
rect 674944 643476 674972 643560
rect 675110 643492 675116 643544
rect 675168 643492 675174 643544
rect 674926 643424 674932 643476
rect 674984 643424 674990 643476
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 45186 643328 45192 643340
rect 42116 643300 45192 643328
rect 42116 643288 42122 643300
rect 45186 643288 45192 643300
rect 45244 643288 45250 643340
rect 674742 643288 674748 643340
rect 674800 643328 674806 643340
rect 675128 643328 675156 643492
rect 674800 643300 675156 643328
rect 674800 643288 674806 643300
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 61378 643124 61384 643136
rect 42116 643096 61384 643124
rect 42116 643084 42122 643096
rect 61378 643084 61384 643096
rect 61436 643084 61442 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 674006 643124 674012 643136
rect 655388 643096 674012 643124
rect 655388 643084 655394 643096
rect 674006 643084 674012 643096
rect 674064 643084 674070 643136
rect 674558 642744 674564 642796
rect 674616 642784 674622 642796
rect 675294 642784 675300 642796
rect 674616 642756 675300 642784
rect 674616 642744 674622 642756
rect 675294 642744 675300 642756
rect 675352 642744 675358 642796
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62758 642376 62764 642388
rect 42116 642348 62764 642376
rect 42116 642336 42122 642348
rect 62758 642336 62764 642348
rect 62816 642336 62822 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 658918 642376 658924 642388
rect 651524 642348 658924 642376
rect 651524 642336 651530 642348
rect 658918 642336 658924 642348
rect 658976 642336 658982 642388
rect 35618 641996 35624 642048
rect 35676 642036 35682 642048
rect 39574 642036 39580 642048
rect 35676 642008 39580 642036
rect 35676 641996 35682 642008
rect 39574 641996 39580 642008
rect 39632 641996 39638 642048
rect 35802 641724 35808 641776
rect 35860 641764 35866 641776
rect 41690 641764 41696 641776
rect 35860 641736 41696 641764
rect 35860 641724 35866 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 44634 641764 44640 641776
rect 42116 641736 44640 641764
rect 42116 641724 42122 641736
rect 44634 641724 44640 641736
rect 44692 641724 44698 641776
rect 35802 640704 35808 640756
rect 35860 640744 35866 640756
rect 39942 640744 39948 640756
rect 35860 640716 39948 640744
rect 35860 640704 35866 640716
rect 39942 640704 39948 640716
rect 40000 640704 40006 640756
rect 41690 640540 41696 640552
rect 41386 640512 41696 640540
rect 35342 640432 35348 640484
rect 35400 640472 35406 640484
rect 41386 640472 41414 640512
rect 41690 640500 41696 640512
rect 41748 640500 41754 640552
rect 42058 640500 42064 640552
rect 42116 640540 42122 640552
rect 44634 640540 44640 640552
rect 42116 640512 44640 640540
rect 42116 640500 42122 640512
rect 44634 640500 44640 640512
rect 44692 640500 44698 640552
rect 35400 640444 41414 640472
rect 35400 640432 35406 640444
rect 35526 640296 35532 640348
rect 35584 640336 35590 640348
rect 41690 640336 41696 640348
rect 35584 640308 41696 640336
rect 35584 640296 35590 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 44266 640336 44272 640348
rect 42116 640308 44272 640336
rect 42116 640296 42122 640308
rect 44266 640296 44272 640308
rect 44324 640296 44330 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 668578 640336 668584 640348
rect 651524 640308 668584 640336
rect 651524 640296 651530 640308
rect 668578 640296 668584 640308
rect 668636 640296 668642 640348
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 37918 639112 37924 639124
rect 35866 639084 37924 639112
rect 37918 639072 37924 639084
rect 37976 639072 37982 639124
rect 39224 639016 40080 639044
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 39224 638976 39252 639016
rect 35860 638948 39252 638976
rect 35860 638936 35866 638948
rect 40052 638908 40080 639016
rect 41690 638908 41696 638920
rect 40052 638880 41696 638908
rect 41690 638868 41696 638880
rect 41748 638868 41754 638920
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 36538 637616 36544 637628
rect 35860 637588 36544 637616
rect 35860 637576 35866 637588
rect 36538 637576 36544 637588
rect 36596 637576 36602 637628
rect 35618 636828 35624 636880
rect 35676 636868 35682 636880
rect 39114 636868 39120 636880
rect 35676 636840 39120 636868
rect 35676 636828 35682 636840
rect 39114 636828 39120 636840
rect 39172 636828 39178 636880
rect 674282 636828 674288 636880
rect 674340 636868 674346 636880
rect 683298 636868 683304 636880
rect 674340 636840 683304 636868
rect 674340 636828 674346 636840
rect 683298 636828 683304 636840
rect 683356 636828 683362 636880
rect 35526 636488 35532 636540
rect 35584 636528 35590 636540
rect 39758 636528 39764 636540
rect 35584 636500 39764 636528
rect 35584 636488 35590 636500
rect 39758 636488 39764 636500
rect 39816 636488 39822 636540
rect 35802 636216 35808 636268
rect 35860 636256 35866 636268
rect 39942 636256 39948 636268
rect 35860 636228 39948 636256
rect 35860 636216 35866 636228
rect 39942 636216 39948 636228
rect 40000 636216 40006 636268
rect 669590 635604 669596 635656
rect 669648 635644 669654 635656
rect 670234 635644 670240 635656
rect 669648 635616 670240 635644
rect 669648 635604 669654 635616
rect 670234 635604 670240 635616
rect 670292 635604 670298 635656
rect 35802 634924 35808 634976
rect 35860 634964 35866 634976
rect 41414 634964 41420 634976
rect 35860 634936 41420 634964
rect 35860 634924 35866 634936
rect 41414 634924 41420 634936
rect 41472 634924 41478 634976
rect 35802 633700 35808 633752
rect 35860 633740 35866 633752
rect 39114 633740 39120 633752
rect 35860 633712 39120 633740
rect 35860 633700 35866 633712
rect 39114 633700 39120 633712
rect 39172 633700 39178 633752
rect 35802 633428 35808 633480
rect 35860 633468 35866 633480
rect 40402 633468 40408 633480
rect 35860 633440 40408 633468
rect 35860 633428 35866 633440
rect 40402 633428 40408 633440
rect 40460 633428 40466 633480
rect 669406 633088 669412 633140
rect 669464 633128 669470 633140
rect 671154 633128 671160 633140
rect 669464 633100 671160 633128
rect 669464 633088 669470 633100
rect 671154 633088 671160 633100
rect 671212 633088 671218 633140
rect 669498 631320 669504 631372
rect 669556 631360 669562 631372
rect 669866 631360 669872 631372
rect 669556 631332 669872 631360
rect 669556 631320 669562 631332
rect 669866 631320 669872 631332
rect 669924 631320 669930 631372
rect 36538 630708 36544 630760
rect 36596 630748 36602 630760
rect 41506 630748 41512 630760
rect 36596 630720 41512 630748
rect 36596 630708 36602 630720
rect 41506 630708 41512 630720
rect 41564 630708 41570 630760
rect 32030 629892 32036 629944
rect 32088 629932 32094 629944
rect 37734 629932 37740 629944
rect 32088 629904 37740 629932
rect 32088 629892 32094 629904
rect 37734 629892 37740 629904
rect 37792 629892 37798 629944
rect 42058 629484 42064 629536
rect 42116 629524 42122 629536
rect 42702 629524 42708 629536
rect 42116 629496 42708 629524
rect 42116 629484 42122 629496
rect 42702 629484 42708 629496
rect 42760 629484 42766 629536
rect 674282 627852 674288 627904
rect 674340 627892 674346 627904
rect 675386 627892 675392 627904
rect 674340 627864 675392 627892
rect 674340 627852 674346 627864
rect 675386 627852 675392 627864
rect 675444 627852 675450 627904
rect 670050 625948 670056 626000
rect 670108 625988 670114 626000
rect 673546 625988 673552 626000
rect 670108 625960 673552 625988
rect 670108 625948 670114 625960
rect 673546 625948 673552 625960
rect 673604 625948 673610 626000
rect 45738 625812 45744 625864
rect 45796 625852 45802 625864
rect 62942 625852 62948 625864
rect 45796 625824 62948 625852
rect 45796 625812 45802 625824
rect 62942 625812 62948 625824
rect 63000 625812 63006 625864
rect 667198 625676 667204 625728
rect 667256 625716 667262 625728
rect 674006 625716 674012 625728
rect 667256 625688 674012 625716
rect 667256 625676 667262 625688
rect 674006 625676 674012 625688
rect 674064 625676 674070 625728
rect 674926 625676 674932 625728
rect 674984 625716 674990 625728
rect 676490 625716 676496 625728
rect 674984 625688 676496 625716
rect 674984 625676 674990 625688
rect 676490 625676 676496 625688
rect 676548 625676 676554 625728
rect 657538 625132 657544 625184
rect 657596 625172 657602 625184
rect 674006 625172 674012 625184
rect 657596 625144 674012 625172
rect 657596 625132 657602 625144
rect 674006 625132 674012 625144
rect 674064 625132 674070 625184
rect 670142 624656 670148 624708
rect 670200 624696 670206 624708
rect 674006 624696 674012 624708
rect 670200 624668 674012 624696
rect 670200 624656 670206 624668
rect 674006 624656 674012 624668
rect 674064 624656 674070 624708
rect 42334 624452 42340 624504
rect 42392 624492 42398 624504
rect 44358 624492 44364 624504
rect 42392 624464 44364 624492
rect 42392 624452 42398 624464
rect 44358 624452 44364 624464
rect 44416 624452 44422 624504
rect 671522 624316 671528 624368
rect 671580 624356 671586 624368
rect 674006 624356 674012 624368
rect 671580 624328 674012 624356
rect 671580 624316 671586 624328
rect 674006 624316 674012 624328
rect 674064 624316 674070 624368
rect 671614 623840 671620 623892
rect 671672 623880 671678 623892
rect 674006 623880 674012 623892
rect 671672 623852 674012 623880
rect 671672 623840 671678 623852
rect 674006 623840 674012 623852
rect 674064 623840 674070 623892
rect 671338 623500 671344 623552
rect 671396 623540 671402 623552
rect 674006 623540 674012 623552
rect 671396 623512 674012 623540
rect 671396 623500 671402 623512
rect 674006 623500 674012 623512
rect 674064 623500 674070 623552
rect 669958 623024 669964 623076
rect 670016 623064 670022 623076
rect 674006 623064 674012 623076
rect 670016 623036 674012 623064
rect 670016 623024 670022 623036
rect 674006 623024 674012 623036
rect 674064 623024 674070 623076
rect 669498 622888 669504 622940
rect 669556 622888 669562 622940
rect 669516 622804 669544 622888
rect 669498 622752 669504 622804
rect 669556 622752 669562 622804
rect 670326 622208 670332 622260
rect 670384 622248 670390 622260
rect 674006 622248 674012 622260
rect 670384 622220 674012 622248
rect 670384 622208 670390 622220
rect 674006 622208 674012 622220
rect 674064 622208 674070 622260
rect 668210 621732 668216 621784
rect 668268 621772 668274 621784
rect 674006 621772 674012 621784
rect 668268 621744 674012 621772
rect 668268 621732 668274 621744
rect 674006 621732 674012 621744
rect 674064 621732 674070 621784
rect 666462 621052 666468 621104
rect 666520 621092 666526 621104
rect 674006 621092 674012 621104
rect 666520 621064 674012 621092
rect 666520 621052 666526 621064
rect 674006 621052 674012 621064
rect 674064 621052 674070 621104
rect 674374 620848 674380 620900
rect 674432 620888 674438 620900
rect 675386 620888 675392 620900
rect 674432 620860 675392 620888
rect 674432 620848 674438 620860
rect 675386 620848 675392 620860
rect 675444 620848 675450 620900
rect 668762 620236 668768 620288
rect 668820 620276 668826 620288
rect 674006 620276 674012 620288
rect 668820 620248 674012 620276
rect 668820 620236 668826 620248
rect 674006 620236 674012 620248
rect 674064 620236 674070 620288
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 44174 619664 44180 619676
rect 42300 619636 44180 619664
rect 42300 619624 42306 619636
rect 44174 619624 44180 619636
rect 44232 619624 44238 619676
rect 666278 619624 666284 619676
rect 666336 619664 666342 619676
rect 673638 619664 673644 619676
rect 666336 619636 673644 619664
rect 666336 619624 666342 619636
rect 673638 619624 673644 619636
rect 673696 619624 673702 619676
rect 672350 619012 672356 619064
rect 672408 619052 672414 619064
rect 674006 619052 674012 619064
rect 672408 619024 674012 619052
rect 672408 619012 672414 619024
rect 674006 619012 674012 619024
rect 674064 619012 674070 619064
rect 42150 617244 42156 617296
rect 42208 617284 42214 617296
rect 42702 617284 42708 617296
rect 42208 617256 42708 617284
rect 42208 617244 42214 617256
rect 42702 617244 42708 617256
rect 42760 617244 42766 617296
rect 668026 616904 668032 616956
rect 668084 616944 668090 616956
rect 674006 616944 674012 616956
rect 668084 616916 674012 616944
rect 668084 616904 668090 616916
rect 674006 616904 674012 616916
rect 674064 616904 674070 616956
rect 44358 616768 44364 616820
rect 44416 616808 44422 616820
rect 62114 616808 62120 616820
rect 44416 616780 62120 616808
rect 44416 616768 44422 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 670694 616564 670700 616616
rect 670752 616604 670758 616616
rect 674006 616604 674012 616616
rect 670752 616576 674012 616604
rect 670752 616564 670758 616576
rect 674006 616564 674012 616576
rect 674064 616564 674070 616616
rect 669774 615476 669780 615528
rect 669832 615516 669838 615528
rect 674006 615516 674012 615528
rect 669832 615488 674012 615516
rect 669832 615476 669838 615488
rect 674006 615476 674012 615488
rect 674064 615476 674070 615528
rect 675110 615476 675116 615528
rect 675168 615516 675174 615528
rect 683114 615516 683120 615528
rect 675168 615488 683120 615516
rect 675168 615476 675174 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 670694 614864 670700 614916
rect 670752 614904 670758 614916
rect 674006 614904 674012 614916
rect 670752 614876 674012 614904
rect 670752 614864 670758 614876
rect 674006 614864 674012 614876
rect 674064 614864 674070 614916
rect 43070 614252 43076 614304
rect 43128 614292 43134 614304
rect 44450 614292 44456 614304
rect 43128 614264 44456 614292
rect 43128 614252 43134 614264
rect 44450 614252 44456 614264
rect 44508 614252 44514 614304
rect 42610 614116 42616 614168
rect 42668 614156 42674 614168
rect 62114 614156 62120 614168
rect 42668 614128 62120 614156
rect 42668 614116 42674 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 43898 612688 43904 612740
rect 43956 612688 43962 612740
rect 43916 612592 43944 612688
rect 59998 612620 60004 612672
rect 60056 612660 60062 612672
rect 62114 612660 62120 612672
rect 60056 612632 62120 612660
rect 60056 612620 60062 612632
rect 62114 612620 62120 612632
rect 62172 612620 62178 612672
rect 43548 612564 43944 612592
rect 43548 612510 43576 612564
rect 44082 612388 44088 612400
rect 43663 612360 44088 612388
rect 43663 612306 43691 612360
rect 44082 612348 44088 612360
rect 44140 612348 44146 612400
rect 43766 612196 43818 612202
rect 43766 612138 43818 612144
rect 44082 612048 44088 612060
rect 43887 612020 44088 612048
rect 43887 611966 43915 612020
rect 44082 612008 44088 612020
rect 44140 612008 44146 612060
rect 43996 611788 44048 611794
rect 43996 611730 44048 611736
rect 44266 611600 44272 611652
rect 44324 611640 44330 611652
rect 44324 611612 45048 611640
rect 44324 611600 44330 611612
rect 44088 611584 44140 611590
rect 44088 611526 44140 611532
rect 44205 611328 44211 611380
rect 44263 611328 44269 611380
rect 44818 611232 44824 611244
rect 44447 611204 44824 611232
rect 44312 611124 44318 611176
rect 44370 611124 44376 611176
rect 44447 610946 44475 611204
rect 44818 611192 44824 611204
rect 44876 611192 44882 611244
rect 45020 611028 45048 611612
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 674006 611368 674012 611380
rect 653456 611340 674012 611368
rect 653456 611328 653462 611340
rect 674006 611328 674012 611340
rect 674064 611328 674070 611380
rect 44560 611000 45048 611028
rect 44560 610742 44588 611000
rect 674834 604528 674840 604580
rect 674892 604568 674898 604580
rect 675294 604568 675300 604580
rect 674892 604540 675300 604568
rect 674892 604528 674898 604540
rect 675294 604528 675300 604540
rect 675352 604528 675358 604580
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 36538 601712 36544 601724
rect 35860 601684 36544 601712
rect 35860 601672 35866 601684
rect 36538 601672 36544 601684
rect 36596 601672 36602 601724
rect 657538 600312 657544 600364
rect 657596 600352 657602 600364
rect 673822 600352 673828 600364
rect 657596 600324 673828 600352
rect 657596 600312 657602 600324
rect 673822 600312 673828 600324
rect 673880 600312 673886 600364
rect 673822 599468 673828 599480
rect 663766 599440 673828 599468
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 663766 598992 663794 599440
rect 673822 599428 673828 599440
rect 673880 599428 673886 599480
rect 654836 598964 663794 598992
rect 654836 598952 654842 598964
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 667198 597564 667204 597576
rect 651524 597536 667204 597564
rect 651524 597524 651530 597536
rect 667198 597524 667204 597536
rect 667256 597524 667262 597576
rect 42886 597388 42892 597440
rect 42944 597388 42950 597440
rect 42904 597032 42932 597388
rect 42886 596980 42892 597032
rect 42944 596980 42950 597032
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 660298 596204 660304 596216
rect 651524 596176 660304 596204
rect 651524 596164 651530 596176
rect 660298 596164 660304 596176
rect 660356 596164 660362 596216
rect 39942 595756 39948 595808
rect 40000 595796 40006 595808
rect 41690 595796 41696 595808
rect 40000 595768 41696 595796
rect 40000 595756 40006 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595416 651656 595468
rect 651708 595456 651714 595468
rect 653398 595456 653404 595468
rect 651708 595428 653404 595456
rect 651708 595416 651714 595428
rect 653398 595416 653404 595428
rect 653456 595416 653462 595468
rect 675018 595212 675024 595264
rect 675076 595252 675082 595264
rect 675076 595224 675248 595252
rect 675076 595212 675082 595224
rect 675220 595060 675248 595224
rect 675202 595008 675208 595060
rect 675260 595008 675266 595060
rect 651466 594872 651472 594924
rect 651524 594912 651530 594924
rect 656158 594912 656164 594924
rect 651524 594884 656164 594912
rect 651524 594872 651530 594884
rect 656158 594872 656164 594884
rect 656216 594872 656222 594924
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 38562 594260 38568 594312
rect 38620 594300 38626 594312
rect 41598 594300 41604 594312
rect 38620 594272 41604 594300
rect 38620 594260 38626 594272
rect 41598 594260 41604 594272
rect 41656 594260 41662 594312
rect 36538 593036 36544 593088
rect 36596 593076 36602 593088
rect 41690 593076 41696 593088
rect 36596 593048 41696 593076
rect 36596 593036 36602 593048
rect 41690 593036 41696 593048
rect 41748 593036 41754 593088
rect 651466 593036 651472 593088
rect 651524 593076 651530 593088
rect 654778 593076 654784 593088
rect 651524 593048 654784 593076
rect 651524 593036 651530 593048
rect 654778 593036 654784 593048
rect 654836 593036 654842 593088
rect 675478 591404 675484 591456
rect 675536 591444 675542 591456
rect 683206 591444 683212 591456
rect 675536 591416 683212 591444
rect 675536 591404 675542 591416
rect 683206 591404 683212 591416
rect 683264 591404 683270 591456
rect 674374 591268 674380 591320
rect 674432 591308 674438 591320
rect 683390 591308 683396 591320
rect 674432 591280 683396 591308
rect 674432 591268 674438 591280
rect 683390 591268 683396 591280
rect 683448 591268 683454 591320
rect 35618 587256 35624 587308
rect 35676 587296 35682 587308
rect 39574 587296 39580 587308
rect 35676 587268 39580 587296
rect 35676 587256 35682 587268
rect 39574 587256 39580 587268
rect 39632 587256 39638 587308
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 41414 587160 41420 587172
rect 33100 587132 41420 587160
rect 33100 587120 33106 587132
rect 41414 587120 41420 587132
rect 41472 587120 41478 587172
rect 33778 585896 33784 585948
rect 33836 585936 33842 585948
rect 40218 585936 40224 585948
rect 33836 585908 40224 585936
rect 33836 585896 33842 585908
rect 40218 585896 40224 585908
rect 40276 585896 40282 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 39942 585800 39948 585812
rect 31076 585772 39948 585800
rect 31076 585760 31082 585772
rect 39942 585760 39948 585772
rect 40000 585760 40006 585812
rect 42150 585760 42156 585812
rect 42208 585800 42214 585812
rect 42702 585800 42708 585812
rect 42208 585772 42708 585800
rect 42208 585760 42214 585772
rect 42702 585760 42708 585772
rect 42760 585760 42766 585812
rect 652018 581000 652024 581052
rect 652076 581040 652082 581052
rect 674006 581040 674012 581052
rect 652076 581012 674012 581040
rect 652076 581000 652082 581012
rect 674006 581000 674012 581012
rect 674064 581000 674070 581052
rect 670142 580388 670148 580440
rect 670200 580428 670206 580440
rect 674006 580428 674012 580440
rect 670200 580400 674012 580428
rect 670200 580388 670206 580400
rect 674006 580388 674012 580400
rect 674064 580388 674070 580440
rect 668578 580252 668584 580304
rect 668636 580292 668642 580304
rect 674006 580292 674012 580304
rect 668636 580264 674012 580292
rect 668636 580252 668642 580264
rect 674006 580252 674012 580264
rect 674064 580252 674070 580304
rect 674282 580252 674288 580304
rect 674340 580292 674346 580304
rect 676398 580292 676404 580304
rect 674340 580264 676404 580292
rect 674340 580252 674346 580264
rect 676398 580252 676404 580264
rect 676456 580252 676462 580304
rect 674282 580116 674288 580168
rect 674340 580156 674346 580168
rect 676214 580156 676220 580168
rect 674340 580128 676220 580156
rect 674340 580116 674346 580128
rect 676214 580116 676220 580128
rect 676272 580116 676278 580168
rect 658918 579640 658924 579692
rect 658976 579680 658982 579692
rect 674006 579680 674012 579692
rect 658976 579652 674012 579680
rect 658976 579640 658982 579652
rect 674006 579640 674012 579652
rect 674064 579640 674070 579692
rect 669774 579232 669780 579284
rect 669832 579272 669838 579284
rect 674006 579272 674012 579284
rect 669832 579244 674012 579272
rect 669832 579232 669838 579244
rect 674006 579232 674012 579244
rect 674064 579232 674070 579284
rect 674282 579232 674288 579284
rect 674340 579272 674346 579284
rect 676214 579272 676220 579284
rect 674340 579244 676220 579272
rect 674340 579232 674346 579244
rect 676214 579232 676220 579244
rect 676272 579232 676278 579284
rect 671614 579028 671620 579080
rect 671672 579068 671678 579080
rect 674006 579068 674012 579080
rect 671672 579040 674012 579068
rect 671672 579028 671678 579040
rect 674006 579028 674012 579040
rect 674064 579028 674070 579080
rect 674282 578416 674288 578468
rect 674340 578456 674346 578468
rect 676214 578456 676220 578468
rect 674340 578428 676220 578456
rect 674340 578416 674346 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 671522 578280 671528 578332
rect 671580 578320 671586 578332
rect 674006 578320 674012 578332
rect 671580 578292 674012 578320
rect 671580 578280 671586 578292
rect 674006 578280 674012 578292
rect 674064 578280 674070 578332
rect 42242 578212 42248 578264
rect 42300 578252 42306 578264
rect 42702 578252 42708 578264
rect 42300 578224 42708 578252
rect 42300 578212 42306 578224
rect 42702 578212 42708 578224
rect 42760 578212 42766 578264
rect 669958 578076 669964 578128
rect 670016 578116 670022 578128
rect 674006 578116 674012 578128
rect 670016 578088 674012 578116
rect 670016 578076 670022 578088
rect 674006 578076 674012 578088
rect 674064 578076 674070 578128
rect 674282 578076 674288 578128
rect 674340 578116 674346 578128
rect 676214 578116 676220 578128
rect 674340 578088 676220 578116
rect 674340 578076 674346 578088
rect 676214 578076 676220 578088
rect 676272 578076 676278 578128
rect 674834 577872 674840 577924
rect 674892 577912 674898 577924
rect 675478 577912 675484 577924
rect 674892 577884 675484 577912
rect 674892 577872 674898 577884
rect 675478 577872 675484 577884
rect 675536 577872 675542 577924
rect 670326 577804 670332 577856
rect 670384 577844 670390 577856
rect 674006 577844 674012 577856
rect 670384 577816 674012 577844
rect 670384 577804 670390 577816
rect 674006 577804 674012 577816
rect 674064 577804 674070 577856
rect 674282 577736 674288 577788
rect 674340 577776 674346 577788
rect 675846 577776 675852 577788
rect 674340 577748 675852 577776
rect 674340 577736 674346 577748
rect 675846 577736 675852 577748
rect 675904 577736 675910 577788
rect 674282 577600 674288 577652
rect 674340 577640 674346 577652
rect 676214 577640 676220 577652
rect 674340 577612 676220 577640
rect 674340 577600 674346 577612
rect 676214 577600 676220 577612
rect 676272 577600 676278 577652
rect 670234 577464 670240 577516
rect 670292 577504 670298 577516
rect 674006 577504 674012 577516
rect 670292 577476 674012 577504
rect 670292 577464 670298 577476
rect 674006 577464 674012 577476
rect 674064 577464 674070 577516
rect 671154 576920 671160 576972
rect 671212 576960 671218 576972
rect 674006 576960 674012 576972
rect 671212 576932 674012 576960
rect 671212 576920 671218 576932
rect 674006 576920 674012 576932
rect 674064 576920 674070 576972
rect 674282 575968 674288 576020
rect 674340 576008 674346 576020
rect 676214 576008 676220 576020
rect 674340 575980 676220 576008
rect 674340 575968 674346 575980
rect 676214 575968 676220 575980
rect 676272 575968 676278 576020
rect 668394 575492 668400 575544
rect 668452 575532 668458 575544
rect 674006 575532 674012 575544
rect 668452 575504 674012 575532
rect 668452 575492 668458 575504
rect 674006 575492 674012 575504
rect 674064 575492 674070 575544
rect 44634 575424 44640 575476
rect 44692 575464 44698 575476
rect 62114 575464 62120 575476
rect 44692 575436 62120 575464
rect 44692 575424 44698 575436
rect 62114 575424 62120 575436
rect 62172 575424 62178 575476
rect 670970 574540 670976 574592
rect 671028 574580 671034 574592
rect 674006 574580 674012 574592
rect 671028 574552 674012 574580
rect 671028 574540 671034 574552
rect 674006 574540 674012 574552
rect 674064 574540 674070 574592
rect 671982 574268 671988 574320
rect 672040 574308 672046 574320
rect 674006 574308 674012 574320
rect 672040 574280 674012 574308
rect 672040 574268 672046 574280
rect 674006 574268 674012 574280
rect 674064 574268 674070 574320
rect 674282 574132 674288 574184
rect 674340 574172 674346 574184
rect 676214 574172 676220 574184
rect 674340 574144 676220 574172
rect 674340 574132 674346 574144
rect 676214 574132 676220 574144
rect 676272 574132 676278 574184
rect 667566 574064 667572 574116
rect 667624 574104 667630 574116
rect 674006 574104 674012 574116
rect 667624 574076 674012 574104
rect 667624 574064 667630 574076
rect 674006 574064 674012 574076
rect 674064 574064 674070 574116
rect 45554 573996 45560 574048
rect 45612 574036 45618 574048
rect 62114 574036 62120 574048
rect 45612 574008 62120 574036
rect 45612 573996 45618 574008
rect 62114 573996 62120 574008
rect 62172 573996 62178 574048
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 42610 573492 42616 573504
rect 42208 573464 42616 573492
rect 42208 573452 42214 573464
rect 42610 573452 42616 573464
rect 42668 573452 42674 573504
rect 669498 573044 669504 573096
rect 669556 573084 669562 573096
rect 674006 573084 674012 573096
rect 669556 573056 674012 573084
rect 669556 573044 669562 573056
rect 674006 573044 674012 573056
rect 674064 573044 674070 573096
rect 674282 572908 674288 572960
rect 674340 572948 674346 572960
rect 676214 572948 676220 572960
rect 674340 572920 676220 572948
rect 674340 572908 674346 572920
rect 676214 572908 676220 572920
rect 676272 572908 676278 572960
rect 667750 572704 667756 572756
rect 667808 572744 667814 572756
rect 674006 572744 674012 572756
rect 667808 572716 674012 572744
rect 667808 572704 667814 572716
rect 674006 572704 674012 572716
rect 674064 572704 674070 572756
rect 674282 571888 674288 571940
rect 674340 571928 674346 571940
rect 676214 571928 676220 571940
rect 674340 571900 676220 571928
rect 674340 571888 674346 571900
rect 676214 571888 676220 571900
rect 676272 571888 676278 571940
rect 670418 571412 670424 571464
rect 670476 571452 670482 571464
rect 674006 571452 674012 571464
rect 670476 571424 674012 571452
rect 670476 571412 670482 571424
rect 674006 571412 674012 571424
rect 674064 571412 674070 571464
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 674282 570052 674288 570104
rect 674340 570092 674346 570104
rect 676214 570092 676220 570104
rect 674340 570064 676220 570092
rect 674340 570052 674346 570064
rect 676214 570052 676220 570064
rect 676272 570052 676278 570104
rect 671982 569916 671988 569968
rect 672040 569956 672046 569968
rect 674006 569956 674012 569968
rect 672040 569928 674012 569956
rect 672040 569916 672046 569928
rect 674006 569916 674012 569928
rect 674064 569916 674070 569968
rect 674282 569236 674288 569288
rect 674340 569276 674346 569288
rect 676214 569276 676220 569288
rect 674340 569248 676220 569276
rect 674340 569236 674346 569248
rect 676214 569236 676220 569248
rect 676272 569236 676278 569288
rect 670050 568556 670056 568608
rect 670108 568596 670114 568608
rect 674006 568596 674012 568608
rect 670108 568568 674012 568596
rect 670108 568556 670114 568568
rect 674006 568556 674012 568568
rect 674064 568556 674070 568608
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 673822 565876 673828 565888
rect 653456 565848 673828 565876
rect 653456 565836 653462 565848
rect 673822 565836 673828 565848
rect 673880 565836 673886 565888
rect 674466 559308 674472 559360
rect 674524 559348 674530 559360
rect 675110 559348 675116 559360
rect 674524 559320 675116 559348
rect 674524 559308 674530 559320
rect 675110 559308 675116 559320
rect 675168 559308 675174 559360
rect 674282 558220 674288 558272
rect 674340 558260 674346 558272
rect 675386 558260 675392 558272
rect 674340 558232 675392 558260
rect 674340 558220 674346 558232
rect 675386 558220 675392 558232
rect 675444 558220 675450 558272
rect 674650 557540 674656 557592
rect 674708 557580 674714 557592
rect 675110 557580 675116 557592
rect 674708 557552 675116 557580
rect 674708 557540 674714 557552
rect 675110 557540 675116 557552
rect 675168 557540 675174 557592
rect 657814 554752 657820 554804
rect 657872 554792 657878 554804
rect 673822 554792 673828 554804
rect 657872 554764 673828 554792
rect 657872 554752 657878 554764
rect 673822 554752 673828 554764
rect 673880 554752 673886 554804
rect 674466 554684 674472 554736
rect 674524 554724 674530 554736
rect 675110 554724 675116 554736
rect 674524 554696 675116 554724
rect 674524 554684 674530 554696
rect 675110 554684 675116 554696
rect 675168 554684 675174 554736
rect 673822 553704 673828 553716
rect 663766 553676 673828 553704
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 663766 553432 663794 553676
rect 673822 553664 673828 553676
rect 673880 553664 673886 553716
rect 655204 553404 663794 553432
rect 655204 553392 655210 553404
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 651466 552032 651472 552084
rect 651524 552072 651530 552084
rect 658918 552072 658924 552084
rect 651524 552044 658924 552072
rect 651524 552032 651530 552044
rect 658918 552032 658924 552044
rect 658976 552032 658982 552084
rect 40034 550944 40040 550996
rect 40092 550984 40098 550996
rect 41690 550984 41696 550996
rect 40092 550956 41696 550984
rect 40092 550944 40098 550956
rect 41690 550944 41696 550956
rect 41748 550944 41754 550996
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 669590 550644 669596 550656
rect 651524 550616 669596 550644
rect 651524 550604 651530 550616
rect 669590 550604 669596 550616
rect 669648 550604 669654 550656
rect 651374 550332 651380 550384
rect 651432 550372 651438 550384
rect 653398 550372 653404 550384
rect 651432 550344 653404 550372
rect 651432 550332 651438 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 675018 549992 675024 550044
rect 675076 550032 675082 550044
rect 675076 550004 675340 550032
rect 675076 549992 675082 550004
rect 675312 549840 675340 550004
rect 675294 549788 675300 549840
rect 675352 549788 675358 549840
rect 651466 549040 651472 549092
rect 651524 549080 651530 549092
rect 657814 549080 657820 549092
rect 651524 549052 657820 549080
rect 651524 549040 651530 549052
rect 657814 549040 657820 549052
rect 657872 549040 657878 549092
rect 651466 548836 651472 548888
rect 651524 548876 651530 548888
rect 655146 548876 655152 548888
rect 651524 548848 655152 548876
rect 651524 548836 651530 548848
rect 655146 548836 655152 548848
rect 655204 548836 655210 548888
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 41598 547448 41604 547460
rect 31812 547420 41604 547448
rect 31812 547408 31818 547420
rect 41598 547408 41604 547420
rect 41656 547408 41662 547460
rect 675478 547136 675484 547188
rect 675536 547176 675542 547188
rect 684310 547176 684316 547188
rect 675536 547148 684316 547176
rect 675536 547136 675542 547148
rect 684310 547136 684316 547148
rect 684368 547136 684374 547188
rect 675110 546864 675116 546916
rect 675168 546864 675174 546916
rect 675128 546712 675156 546864
rect 675110 546660 675116 546712
rect 675168 546660 675174 546712
rect 676186 546536 678974 546564
rect 674834 546456 674840 546508
rect 674892 546496 674898 546508
rect 676186 546496 676214 546536
rect 674892 546468 676214 546496
rect 678946 546496 678974 546536
rect 680998 546496 681004 546508
rect 678946 546468 681004 546496
rect 674892 546456 674898 546468
rect 680998 546456 681004 546468
rect 681056 546456 681062 546508
rect 675662 545708 675668 545760
rect 675720 545748 675726 545760
rect 683298 545748 683304 545760
rect 675720 545720 683304 545748
rect 675720 545708 675726 545720
rect 683298 545708 683304 545720
rect 683356 545708 683362 545760
rect 34422 544348 34428 544400
rect 34480 544388 34486 544400
rect 37826 544388 37832 544400
rect 34480 544360 37832 544388
rect 34480 544348 34486 544360
rect 37826 544348 37832 544360
rect 37884 544348 37890 544400
rect 42978 538160 42984 538212
rect 43036 538160 43042 538212
rect 42794 537888 42800 537940
rect 42852 537928 42858 537940
rect 42996 537928 43024 538160
rect 42852 537900 43024 537928
rect 42852 537888 42858 537900
rect 667198 535644 667204 535696
rect 667256 535684 667262 535696
rect 674006 535684 674012 535696
rect 667256 535656 674012 535684
rect 667256 535644 667262 535656
rect 674006 535644 674012 535656
rect 674064 535644 674070 535696
rect 660298 535440 660304 535492
rect 660356 535480 660362 535492
rect 674006 535480 674012 535492
rect 660356 535452 674012 535480
rect 660356 535440 660362 535452
rect 674006 535440 674012 535452
rect 674064 535440 674070 535492
rect 669774 534964 669780 535016
rect 669832 535004 669838 535016
rect 672718 535004 672724 535016
rect 669832 534976 672724 535004
rect 669832 534964 669838 534976
rect 672718 534964 672724 534976
rect 672776 534964 672782 535016
rect 656158 534216 656164 534268
rect 656216 534256 656222 534268
rect 674006 534256 674012 534268
rect 656216 534228 674012 534256
rect 656216 534216 656222 534228
rect 674006 534216 674012 534228
rect 674064 534216 674070 534268
rect 670786 534080 670792 534132
rect 670844 534120 670850 534132
rect 674006 534120 674012 534132
rect 670844 534092 674012 534120
rect 670844 534080 670850 534092
rect 674006 534080 674012 534092
rect 674064 534080 674070 534132
rect 670234 532924 670240 532976
rect 670292 532964 670298 532976
rect 674006 532964 674012 532976
rect 670292 532936 674012 532964
rect 670292 532924 670298 532936
rect 674006 532924 674012 532936
rect 674064 532924 674070 532976
rect 42426 532720 42432 532772
rect 42484 532760 42490 532772
rect 43162 532760 43168 532772
rect 42484 532732 43168 532760
rect 42484 532720 42490 532732
rect 43162 532720 43168 532732
rect 43220 532720 43226 532772
rect 671614 532720 671620 532772
rect 671672 532760 671678 532772
rect 674006 532760 674012 532772
rect 671672 532732 674012 532760
rect 671672 532720 671678 532732
rect 674006 532720 674012 532732
rect 674064 532720 674070 532772
rect 671154 531700 671160 531752
rect 671212 531740 671218 531752
rect 674006 531740 674012 531752
rect 671212 531712 674012 531740
rect 671212 531700 671218 531712
rect 674006 531700 674012 531712
rect 674064 531700 674070 531752
rect 671154 531292 671160 531344
rect 671212 531332 671218 531344
rect 674006 531332 674012 531344
rect 671212 531304 674012 531332
rect 671212 531292 671218 531304
rect 674006 531292 674012 531304
rect 674064 531292 674070 531344
rect 44726 531224 44732 531276
rect 44784 531264 44790 531276
rect 62114 531264 62120 531276
rect 44784 531236 62120 531264
rect 44784 531224 44790 531236
rect 62114 531224 62120 531236
rect 62172 531224 62178 531276
rect 59998 531088 60004 531140
rect 60056 531128 60062 531140
rect 62298 531128 62304 531140
rect 60056 531100 62304 531128
rect 60056 531088 60062 531100
rect 62298 531088 62304 531100
rect 62356 531088 62362 531140
rect 667014 530476 667020 530528
rect 667072 530516 667078 530528
rect 674006 530516 674012 530528
rect 667072 530488 674012 530516
rect 667072 530476 667078 530488
rect 674006 530476 674012 530488
rect 674064 530476 674070 530528
rect 671798 530204 671804 530256
rect 671856 530244 671862 530256
rect 674006 530244 674012 530256
rect 671856 530216 674012 530244
rect 671856 530204 671862 530216
rect 674006 530204 674012 530216
rect 674064 530204 674070 530256
rect 42150 530068 42156 530120
rect 42208 530108 42214 530120
rect 42978 530108 42984 530120
rect 42208 530080 42984 530108
rect 42208 530068 42214 530080
rect 42978 530068 42984 530080
rect 43036 530068 43042 530120
rect 669038 530000 669044 530052
rect 669096 530040 669102 530052
rect 669096 530012 674052 530040
rect 669096 530000 669102 530012
rect 674024 529916 674052 530012
rect 674006 529864 674012 529916
rect 674064 529864 674070 529916
rect 671338 528708 671344 528760
rect 671396 528748 671402 528760
rect 674006 528748 674012 528760
rect 671396 528720 674012 528748
rect 671396 528708 671402 528720
rect 674006 528708 674012 528720
rect 674064 528708 674070 528760
rect 45094 528572 45100 528624
rect 45152 528612 45158 528624
rect 62114 528612 62120 528624
rect 45152 528584 62120 528612
rect 45152 528572 45158 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 668854 528572 668860 528624
rect 668912 528612 668918 528624
rect 674006 528612 674012 528624
rect 668912 528584 674012 528612
rect 668912 528572 668918 528584
rect 674006 528572 674012 528584
rect 674064 528572 674070 528624
rect 42058 527756 42064 527808
rect 42116 527796 42122 527808
rect 42610 527796 42616 527808
rect 42116 527768 42616 527796
rect 42116 527756 42122 527768
rect 42610 527756 42616 527768
rect 42668 527756 42674 527808
rect 672534 527348 672540 527400
rect 672592 527388 672598 527400
rect 674006 527388 674012 527400
rect 672592 527360 674012 527388
rect 672592 527348 672598 527360
rect 674006 527348 674012 527360
rect 674064 527348 674070 527400
rect 672350 527144 672356 527196
rect 672408 527184 672414 527196
rect 673638 527184 673644 527196
rect 672408 527156 673644 527184
rect 672408 527144 672414 527156
rect 673638 527144 673644 527156
rect 673696 527144 673702 527196
rect 680998 525716 681004 525768
rect 681056 525756 681062 525768
rect 683114 525756 683120 525768
rect 681056 525728 683120 525756
rect 681056 525716 681062 525728
rect 683114 525716 683120 525728
rect 683172 525716 683178 525768
rect 676858 518916 676864 518968
rect 676916 518956 676922 518968
rect 683298 518956 683304 518968
rect 676916 518928 683304 518956
rect 676916 518916 676922 518928
rect 683298 518916 683304 518928
rect 683356 518916 683362 518968
rect 677870 518820 677876 518832
rect 675496 518792 677876 518820
rect 675496 518696 675524 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 675478 518644 675484 518696
rect 675536 518644 675542 518696
rect 675662 503820 675668 503872
rect 675720 503860 675726 503872
rect 678238 503860 678244 503872
rect 675720 503832 678244 503860
rect 675720 503820 675726 503832
rect 678238 503820 678244 503832
rect 678296 503820 678302 503872
rect 674282 494708 674288 494760
rect 674340 494748 674346 494760
rect 683206 494748 683212 494760
rect 674340 494720 683212 494748
rect 674340 494708 674346 494720
rect 683206 494708 683212 494720
rect 683264 494708 683270 494760
rect 669590 491852 669596 491904
rect 669648 491892 669654 491904
rect 674006 491892 674012 491904
rect 669648 491864 674012 491892
rect 669648 491852 669654 491864
rect 674006 491852 674012 491864
rect 674064 491852 674070 491904
rect 674282 491784 674288 491836
rect 674340 491824 674346 491836
rect 675846 491824 675852 491836
rect 674340 491796 675852 491824
rect 674340 491784 674346 491796
rect 675846 491784 675852 491796
rect 675904 491784 675910 491836
rect 674282 491648 674288 491700
rect 674340 491688 674346 491700
rect 676030 491688 676036 491700
rect 674340 491660 676036 491688
rect 674340 491648 674346 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 665818 491444 665824 491496
rect 665876 491484 665882 491496
rect 674006 491484 674012 491496
rect 665876 491456 674012 491484
rect 665876 491444 665882 491456
rect 674006 491444 674012 491456
rect 674064 491444 674070 491496
rect 658918 491308 658924 491360
rect 658976 491348 658982 491360
rect 673822 491348 673828 491360
rect 658976 491320 673828 491348
rect 658976 491308 658982 491320
rect 673822 491308 673828 491320
rect 673880 491308 673886 491360
rect 670786 490900 670792 490952
rect 670844 490940 670850 490952
rect 674006 490940 674012 490952
rect 670844 490912 674012 490940
rect 670844 490900 670850 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 671614 489268 671620 489320
rect 671672 489308 671678 489320
rect 673914 489308 673920 489320
rect 671672 489280 673920 489308
rect 671672 489268 671678 489280
rect 673914 489268 673920 489280
rect 673972 489268 673978 489320
rect 671154 488452 671160 488504
rect 671212 488492 671218 488504
rect 673914 488492 673920 488504
rect 671212 488464 673920 488492
rect 671212 488452 671218 488464
rect 673914 488452 673920 488464
rect 673972 488452 673978 488504
rect 675202 488452 675208 488504
rect 675260 488492 675266 488504
rect 676030 488492 676036 488504
rect 675260 488464 676036 488492
rect 675260 488452 675266 488464
rect 676030 488452 676036 488464
rect 676088 488452 676094 488504
rect 668670 485800 668676 485852
rect 668728 485840 668734 485852
rect 673914 485840 673920 485852
rect 668728 485812 673920 485840
rect 668728 485800 668734 485812
rect 673914 485800 673920 485812
rect 673972 485800 673978 485852
rect 670970 485596 670976 485648
rect 671028 485636 671034 485648
rect 674006 485636 674012 485648
rect 671028 485608 674012 485636
rect 671028 485596 671034 485608
rect 674006 485596 674012 485608
rect 674064 485596 674070 485648
rect 667750 484372 667756 484424
rect 667808 484412 667814 484424
rect 674006 484412 674012 484424
rect 667808 484384 674012 484412
rect 667808 484372 667814 484384
rect 674006 484372 674012 484384
rect 674064 484372 674070 484424
rect 670418 483964 670424 484016
rect 670476 484004 670482 484016
rect 674006 484004 674012 484016
rect 670476 483976 674012 484004
rect 670476 483964 670482 483976
rect 674006 483964 674012 483976
rect 674064 483964 674070 484016
rect 674926 480428 674932 480480
rect 674984 480468 674990 480480
rect 683114 480468 683120 480480
rect 674984 480440 683120 480468
rect 674984 480428 674990 480440
rect 683114 480428 683120 480440
rect 683172 480428 683178 480480
rect 675294 475192 675300 475244
rect 675352 475232 675358 475244
rect 680354 475232 680360 475244
rect 675352 475204 680360 475232
rect 675352 475192 675358 475204
rect 680354 475192 680360 475204
rect 680412 475192 680418 475244
rect 669222 456560 669228 456612
rect 669280 456600 669286 456612
rect 669280 456572 673988 456600
rect 669280 456560 669286 456572
rect 673960 456246 673988 456572
rect 673362 455948 673368 456000
rect 673420 455988 673426 456000
rect 673420 455960 673854 455988
rect 673420 455948 673426 455960
rect 672166 455812 672172 455864
rect 672224 455852 672230 455864
rect 672224 455824 673762 455852
rect 672224 455812 672230 455824
rect 667382 455608 667388 455660
rect 667440 455648 667446 455660
rect 667440 455620 673624 455648
rect 667440 455608 667446 455620
rect 670602 455472 670608 455524
rect 670660 455512 670666 455524
rect 670660 455484 673454 455512
rect 670660 455472 670666 455484
rect 673270 455336 673276 455388
rect 673328 455336 673334 455388
rect 673426 455376 673454 455484
rect 673426 455348 673532 455376
rect 672074 455064 672080 455116
rect 672132 455104 672138 455116
rect 672132 455076 673224 455104
rect 672132 455064 672138 455076
rect 673196 454900 673224 455076
rect 673288 455022 673316 455336
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 674282 454996 674288 455048
rect 674340 455036 674346 455048
rect 675478 455036 675484 455048
rect 674340 455008 675484 455036
rect 674340 454996 674346 455008
rect 675478 454996 675484 455008
rect 675536 454996 675542 455048
rect 673176 454872 673224 454900
rect 673040 454792 673046 454844
rect 673098 454792 673104 454844
rect 673176 454818 673204 454872
rect 672902 454656 672908 454708
rect 672960 454696 672966 454708
rect 672960 454656 672994 454696
rect 672810 454384 672816 454436
rect 672868 454384 672874 454436
rect 672966 454410 672994 454656
rect 673058 454614 673086 454792
rect 674282 454724 674288 454776
rect 674340 454764 674346 454776
rect 676858 454764 676864 454776
rect 674340 454736 676864 454764
rect 674340 454724 674346 454736
rect 676858 454724 676864 454736
rect 676916 454724 676922 454776
rect 674282 454452 674288 454504
rect 674340 454492 674346 454504
rect 675662 454492 675668 454504
rect 674340 454464 675668 454492
rect 674340 454452 674346 454464
rect 675662 454452 675668 454464
rect 675720 454452 675726 454504
rect 672828 454206 672856 454384
rect 672442 453908 672448 453960
rect 672500 453948 672506 453960
rect 672500 453920 672750 453948
rect 672500 453908 672506 453920
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41690 429196 41696 429208
rect 35860 429168 41696 429196
rect 35860 429156 35866 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 41322 425076 41328 425128
rect 41380 425116 41386 425128
rect 41690 425116 41696 425128
rect 41380 425088 41696 425116
rect 41380 425076 41386 425088
rect 41690 425076 41696 425088
rect 41748 425076 41754 425128
rect 40954 424260 40960 424312
rect 41012 424300 41018 424312
rect 41506 424300 41512 424312
rect 41012 424272 41512 424300
rect 41012 424260 41018 424272
rect 41506 424260 41512 424272
rect 41564 424260 41570 424312
rect 32030 416168 32036 416220
rect 32088 416208 32094 416220
rect 41690 416208 41696 416220
rect 32088 416180 41696 416208
rect 32088 416168 32094 416180
rect 41690 416168 41696 416180
rect 41748 416168 41754 416220
rect 53834 404268 53840 404320
rect 53892 404308 53898 404320
rect 62114 404308 62120 404320
rect 53892 404280 62120 404308
rect 53892 404268 53898 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 674558 403248 674564 403300
rect 674616 403288 674622 403300
rect 676214 403288 676220 403300
rect 674616 403260 676220 403288
rect 674616 403248 674622 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 45278 402908 45284 402960
rect 45336 402948 45342 402960
rect 62114 402948 62120 402960
rect 45336 402920 62120 402948
rect 45336 402908 45342 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 59998 400052 60004 400104
rect 60056 400092 60062 400104
rect 62114 400092 62120 400104
rect 60056 400064 62120 400092
rect 60056 400052 60062 400064
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 674834 398828 674840 398880
rect 674892 398868 674898 398880
rect 676030 398868 676036 398880
rect 674892 398840 676036 398868
rect 674892 398828 674898 398840
rect 676030 398828 676036 398840
rect 676088 398828 676094 398880
rect 675018 396176 675024 396228
rect 675076 396216 675082 396228
rect 676214 396216 676220 396228
rect 675076 396188 676220 396216
rect 675076 396176 675082 396188
rect 676214 396176 676220 396188
rect 676272 396176 676278 396228
rect 674374 396040 674380 396092
rect 674432 396080 674438 396092
rect 676030 396080 676036 396092
rect 674432 396052 676036 396080
rect 674432 396040 674438 396052
rect 676030 396040 676036 396052
rect 676088 396040 676094 396092
rect 674650 395088 674656 395140
rect 674708 395128 674714 395140
rect 676214 395128 676220 395140
rect 674708 395100 676220 395128
rect 674708 395088 674714 395100
rect 676214 395088 676220 395100
rect 676272 395088 676278 395140
rect 675202 389104 675208 389156
rect 675260 389144 675266 389156
rect 679618 389144 679624 389156
rect 675260 389116 679624 389144
rect 675260 389104 675266 389116
rect 679618 389104 679624 389116
rect 679676 389104 679682 389156
rect 675202 386316 675208 386368
rect 675260 386356 675266 386368
rect 675260 386328 675524 386356
rect 675260 386316 675266 386328
rect 675496 386028 675524 386328
rect 675478 385976 675484 386028
rect 675536 385976 675542 386028
rect 674834 384752 674840 384804
rect 674892 384792 674898 384804
rect 675478 384792 675484 384804
rect 674892 384764 675484 384792
rect 674892 384752 674898 384764
rect 675478 384752 675484 384764
rect 675536 384752 675542 384804
rect 41322 382236 41328 382288
rect 41380 382276 41386 382288
rect 41690 382276 41696 382288
rect 41380 382248 41696 382276
rect 41380 382236 41386 382248
rect 41690 382236 41696 382248
rect 41748 382236 41754 382288
rect 674374 382168 674380 382220
rect 674432 382208 674438 382220
rect 675110 382208 675116 382220
rect 674432 382180 675116 382208
rect 674432 382168 674438 382180
rect 675110 382168 675116 382180
rect 675168 382168 675174 382220
rect 674374 378088 674380 378140
rect 674432 378128 674438 378140
rect 675110 378128 675116 378140
rect 674432 378100 675116 378128
rect 674432 378088 674438 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 40218 378020 40224 378072
rect 40276 378060 40282 378072
rect 41690 378060 41696 378072
rect 40276 378032 41696 378060
rect 40276 378020 40282 378032
rect 41690 378020 41696 378032
rect 41748 378020 41754 378072
rect 42058 377952 42064 378004
rect 42116 377992 42122 378004
rect 42702 377992 42708 378004
rect 42116 377964 42708 377992
rect 42116 377952 42122 377964
rect 42702 377952 42708 377964
rect 42760 377952 42766 378004
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 657538 373980 657544 373992
rect 651524 373952 657544 373980
rect 651524 373940 651530 373952
rect 657538 373940 657544 373952
rect 657596 373940 657602 373992
rect 35158 371832 35164 371884
rect 35216 371872 35222 371884
rect 41690 371872 41696 371884
rect 35216 371844 41696 371872
rect 35216 371832 35222 371844
rect 41690 371832 41696 371844
rect 41748 371832 41754 371884
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 42242 365236 42248 365288
rect 42300 365236 42306 365288
rect 42260 364948 42288 365236
rect 42242 364896 42248 364948
rect 42300 364896 42306 364948
rect 42242 364284 42248 364336
rect 42300 364284 42306 364336
rect 42260 364188 42288 364284
rect 42702 364188 42708 364200
rect 42260 364160 42708 364188
rect 42702 364148 42708 364160
rect 42760 364148 42766 364200
rect 46566 361496 46572 361548
rect 46624 361536 46630 361548
rect 62114 361536 62120 361548
rect 46624 361508 62120 361536
rect 46624 361496 46630 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 45370 360136 45376 360188
rect 45428 360176 45434 360188
rect 62114 360176 62120 360188
rect 45428 360148 62120 360176
rect 45428 360136 45434 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 44634 359592 44640 359644
rect 44692 359632 44698 359644
rect 45370 359632 45376 359644
rect 44692 359604 45376 359632
rect 44692 359592 44698 359604
rect 45370 359592 45376 359604
rect 45428 359592 45434 359644
rect 44818 359456 44824 359508
rect 44876 359496 44882 359508
rect 45462 359496 45468 359508
rect 44876 359468 45468 359496
rect 44876 359456 44882 359468
rect 45462 359456 45468 359468
rect 45520 359456 45526 359508
rect 51718 357416 51724 357468
rect 51776 357456 51782 357468
rect 62114 357456 62120 357468
rect 51776 357428 62120 357456
rect 51776 357416 51782 357428
rect 62114 357416 62120 357428
rect 62172 357416 62178 357468
rect 44640 354748 44692 354754
rect 44818 354696 44824 354748
rect 44876 354696 44882 354748
rect 44640 354690 44692 354696
rect 44836 354600 44864 354696
rect 44836 354572 45002 354600
rect 44732 354476 44784 354482
rect 44849 354424 44855 354476
rect 44907 354424 44913 354476
rect 44732 354418 44784 354424
rect 44867 354314 44895 354424
rect 44974 354110 45002 354572
rect 45830 353920 45836 353932
rect 45105 353892 45836 353920
rect 45830 353880 45836 353892
rect 45888 353880 45894 353932
rect 45830 353716 45836 353728
rect 45218 353688 45836 353716
rect 45830 353676 45836 353688
rect 45888 353676 45894 353728
rect 45303 353524 45355 353530
rect 45303 353466 45355 353472
rect 45422 353252 45474 353258
rect 45422 353194 45474 353200
rect 676030 347420 676036 347472
rect 676088 347460 676094 347472
rect 676490 347460 676496 347472
rect 676088 347432 676496 347460
rect 676088 347420 676094 347432
rect 676490 347420 676496 347432
rect 676548 347420 676554 347472
rect 35802 344564 35808 344616
rect 35860 344604 35866 344616
rect 39850 344604 39856 344616
rect 35860 344576 39856 344604
rect 35860 344564 35866 344576
rect 39850 344564 39856 344576
rect 39908 344564 39914 344616
rect 35618 343612 35624 343664
rect 35676 343652 35682 343664
rect 40034 343652 40040 343664
rect 35676 343624 40040 343652
rect 35676 343612 35682 343624
rect 40034 343612 40040 343624
rect 40092 343612 40098 343664
rect 35802 342184 35808 342236
rect 35860 342224 35866 342236
rect 40218 342224 40224 342236
rect 35860 342196 40224 342224
rect 35860 342184 35866 342196
rect 40218 342184 40224 342196
rect 40276 342184 40282 342236
rect 45462 342184 45468 342236
rect 45520 342224 45526 342236
rect 63126 342224 63132 342236
rect 45520 342196 63132 342224
rect 45520 342184 45526 342196
rect 63126 342184 63132 342196
rect 63184 342184 63190 342236
rect 35802 341504 35808 341556
rect 35860 341544 35866 341556
rect 40218 341544 40224 341556
rect 35860 341516 40224 341544
rect 35860 341504 35866 341516
rect 40218 341504 40224 341516
rect 40276 341504 40282 341556
rect 35802 341028 35808 341080
rect 35860 341068 35866 341080
rect 40126 341068 40132 341080
rect 35860 341040 40132 341068
rect 35860 341028 35866 341040
rect 40126 341028 40132 341040
rect 40184 341028 40190 341080
rect 35526 339600 35532 339652
rect 35584 339640 35590 339652
rect 37090 339640 37096 339652
rect 35584 339612 37096 339640
rect 35584 339600 35590 339612
rect 37090 339600 37096 339612
rect 37148 339600 37154 339652
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 38838 339504 38844 339516
rect 35860 339476 38844 339504
rect 35860 339464 35866 339476
rect 38838 339464 38844 339476
rect 38896 339464 38902 339516
rect 674834 339328 674840 339380
rect 674892 339368 674898 339380
rect 675478 339368 675484 339380
rect 674892 339340 675484 339368
rect 674892 339328 674898 339340
rect 675478 339328 675484 339340
rect 675536 339328 675542 339380
rect 674374 336540 674380 336592
rect 674432 336580 674438 336592
rect 675386 336580 675392 336592
rect 674432 336552 675392 336580
rect 674432 336540 674438 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 39850 335356 39856 335368
rect 35860 335328 39856 335356
rect 35860 335316 35866 335328
rect 39850 335316 39856 335328
rect 39908 335316 39914 335368
rect 35802 334092 35808 334144
rect 35860 334132 35866 334144
rect 40310 334132 40316 334144
rect 35860 334104 40316 334132
rect 35860 334092 35866 334104
rect 40310 334092 40316 334104
rect 40368 334092 40374 334144
rect 651374 328244 651380 328296
rect 651432 328284 651438 328296
rect 654778 328284 654784 328296
rect 651432 328256 654784 328284
rect 651432 328244 651438 328256
rect 654778 328244 654784 328256
rect 654836 328244 654842 328296
rect 651374 325592 651380 325644
rect 651432 325632 651438 325644
rect 653398 325632 653404 325644
rect 651432 325604 653404 325632
rect 651432 325592 651438 325604
rect 653398 325592 653404 325604
rect 653456 325592 653462 325644
rect 53834 317364 53840 317416
rect 53892 317404 53898 317416
rect 62114 317404 62120 317416
rect 53892 317376 62120 317404
rect 53892 317364 53898 317376
rect 62114 317364 62120 317376
rect 62172 317364 62178 317416
rect 53098 315936 53104 315988
rect 53156 315976 53162 315988
rect 62114 315976 62120 315988
rect 53156 315948 62120 315976
rect 53156 315936 53162 315948
rect 62114 315936 62120 315948
rect 62172 315936 62178 315988
rect 59906 314712 59912 314764
rect 59964 314752 59970 314764
rect 62114 314752 62120 314764
rect 59964 314724 62120 314752
rect 59964 314712 59970 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 676214 307776 676220 307828
rect 676272 307816 676278 307828
rect 676858 307816 676864 307828
rect 676272 307788 676864 307816
rect 676272 307776 676278 307788
rect 676858 307776 676864 307788
rect 676916 307776 676922 307828
rect 675846 304512 675852 304564
rect 675904 304552 675910 304564
rect 676214 304552 676220 304564
rect 675904 304524 676220 304552
rect 675904 304512 675910 304524
rect 676214 304512 676220 304524
rect 676272 304512 676278 304564
rect 651374 303492 651380 303544
rect 651432 303532 651438 303544
rect 653398 303532 653404 303544
rect 651432 303504 653404 303532
rect 651432 303492 651438 303504
rect 653398 303492 653404 303504
rect 653456 303492 653462 303544
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 664438 300812 664444 300824
rect 651524 300784 664444 300812
rect 651524 300772 651530 300784
rect 664438 300772 664444 300784
rect 664496 300772 664502 300824
rect 35618 298732 35624 298784
rect 35676 298772 35682 298784
rect 41598 298772 41604 298784
rect 35676 298744 41604 298772
rect 35676 298732 35682 298744
rect 41598 298732 41604 298744
rect 41656 298732 41662 298784
rect 35802 298256 35808 298308
rect 35860 298296 35866 298308
rect 41598 298296 41604 298308
rect 35860 298268 41604 298296
rect 35860 298256 35866 298268
rect 41598 298256 41604 298268
rect 41656 298256 41662 298308
rect 651466 298120 651472 298172
rect 651524 298160 651530 298172
rect 662414 298160 662420 298172
rect 651524 298132 662420 298160
rect 651524 298120 651530 298132
rect 662414 298120 662420 298132
rect 662472 298120 662478 298172
rect 676122 298052 676128 298104
rect 676180 298092 676186 298104
rect 676858 298092 676864 298104
rect 676180 298064 676864 298092
rect 676180 298052 676186 298064
rect 676858 298052 676864 298064
rect 676916 298052 676922 298104
rect 675938 297644 675944 297696
rect 675996 297684 676002 297696
rect 677594 297684 677600 297696
rect 675996 297656 677600 297684
rect 675996 297644 676002 297656
rect 677594 297644 677600 297656
rect 677652 297644 677658 297696
rect 675846 297168 675852 297220
rect 675904 297208 675910 297220
rect 679618 297208 679624 297220
rect 675904 297180 679624 297208
rect 675904 297168 675910 297180
rect 679618 297168 679624 297180
rect 679676 297168 679682 297220
rect 651466 297032 651472 297084
rect 651524 297072 651530 297084
rect 656158 297072 656164 297084
rect 651524 297044 656164 297072
rect 651524 297032 651530 297044
rect 656158 297032 656164 297044
rect 656216 297032 656222 297084
rect 652662 295944 652668 295996
rect 652720 295984 652726 295996
rect 665818 295984 665824 295996
rect 652720 295956 665824 295984
rect 652720 295944 652726 295956
rect 665818 295944 665824 295956
rect 665876 295944 665882 295996
rect 35802 295604 35808 295656
rect 35860 295644 35866 295656
rect 40678 295644 40684 295656
rect 35860 295616 40684 295644
rect 35860 295604 35866 295616
rect 40678 295604 40684 295616
rect 40736 295604 40742 295656
rect 35434 295468 35440 295520
rect 35492 295508 35498 295520
rect 40034 295508 40040 295520
rect 35492 295480 40040 295508
rect 35492 295468 35498 295480
rect 40034 295468 40040 295480
rect 40092 295468 40098 295520
rect 58618 295400 58624 295452
rect 58676 295440 58682 295452
rect 62114 295440 62120 295452
rect 58676 295412 62120 295440
rect 58676 295400 58682 295412
rect 62114 295400 62120 295412
rect 62172 295400 62178 295452
rect 35618 295332 35624 295384
rect 35676 295372 35682 295384
rect 41598 295372 41604 295384
rect 35676 295344 41604 295372
rect 35676 295332 35682 295344
rect 41598 295332 41604 295344
rect 41656 295332 41662 295384
rect 35802 294244 35808 294296
rect 35860 294284 35866 294296
rect 41690 294284 41696 294296
rect 35860 294256 41696 294284
rect 35860 294244 35866 294256
rect 41690 294244 41696 294256
rect 41748 294244 41754 294296
rect 57238 294040 57244 294092
rect 57296 294080 57302 294092
rect 62114 294080 62120 294092
rect 57296 294052 62120 294080
rect 57296 294040 57302 294052
rect 62114 294040 62120 294052
rect 62172 294040 62178 294092
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 35802 292884 35808 292936
rect 35860 292924 35866 292936
rect 35860 292884 35894 292924
rect 35866 292856 35894 292884
rect 41322 292856 41328 292868
rect 35866 292828 41328 292856
rect 41322 292816 41328 292828
rect 41380 292816 41386 292868
rect 35802 292544 35808 292596
rect 35860 292584 35866 292596
rect 39206 292584 39212 292596
rect 35860 292556 39212 292584
rect 35860 292544 35866 292556
rect 39206 292544 39212 292556
rect 39264 292544 39270 292596
rect 54478 292544 54484 292596
rect 54536 292584 54542 292596
rect 62298 292584 62304 292596
rect 54536 292556 62304 292584
rect 54536 292544 54542 292556
rect 62298 292544 62304 292556
rect 62356 292544 62362 292596
rect 651466 292544 651472 292596
rect 651524 292584 651530 292596
rect 663058 292584 663064 292596
rect 651524 292556 663064 292584
rect 651524 292544 651530 292556
rect 663058 292544 663064 292556
rect 663116 292544 663122 292596
rect 46198 292408 46204 292460
rect 46256 292448 46262 292460
rect 62114 292448 62120 292460
rect 46256 292420 62120 292448
rect 46256 292408 46262 292420
rect 62114 292408 62120 292420
rect 62172 292408 62178 292460
rect 40034 291320 40040 291372
rect 40092 291360 40098 291372
rect 41690 291360 41696 291372
rect 40092 291332 41696 291360
rect 40092 291320 40098 291332
rect 41690 291320 41696 291332
rect 41748 291320 41754 291372
rect 42058 291184 42064 291236
rect 42116 291224 42122 291236
rect 42610 291224 42616 291236
rect 42116 291196 42616 291224
rect 42116 291184 42122 291196
rect 42610 291184 42616 291196
rect 42668 291184 42674 291236
rect 53098 291116 53104 291168
rect 53156 291156 53162 291168
rect 62114 291156 62120 291168
rect 53156 291128 62120 291156
rect 53156 291116 53162 291128
rect 62114 291116 62120 291128
rect 62172 291116 62178 291168
rect 35802 289892 35808 289944
rect 35860 289932 35866 289944
rect 41690 289932 41696 289944
rect 35860 289904 41696 289932
rect 35860 289892 35866 289904
rect 41690 289892 41696 289904
rect 41748 289892 41754 289944
rect 42058 289824 42064 289876
rect 42116 289864 42122 289876
rect 43346 289864 43352 289876
rect 42116 289836 43352 289864
rect 42116 289824 42122 289836
rect 43346 289824 43352 289836
rect 43404 289824 43410 289876
rect 651466 289824 651472 289876
rect 651524 289864 651530 289876
rect 660298 289864 660304 289876
rect 651524 289836 660304 289864
rect 651524 289824 651530 289836
rect 660298 289824 660304 289836
rect 660356 289824 660362 289876
rect 35618 289076 35624 289128
rect 35676 289116 35682 289128
rect 41690 289116 41696 289128
rect 35676 289088 41696 289116
rect 35676 289076 35682 289088
rect 41690 289076 41696 289088
rect 41748 289076 41754 289128
rect 55858 288464 55864 288516
rect 55916 288504 55922 288516
rect 62114 288504 62120 288516
rect 55916 288476 62120 288504
rect 55916 288464 55922 288476
rect 62114 288464 62120 288476
rect 62172 288464 62178 288516
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 661678 288436 661684 288448
rect 651524 288408 661684 288436
rect 651524 288396 651530 288408
rect 661678 288396 661684 288408
rect 661736 288396 661742 288448
rect 651466 287036 651472 287088
rect 651524 287076 651530 287088
rect 672442 287076 672448 287088
rect 651524 287048 672448 287076
rect 651524 287036 651530 287048
rect 672442 287036 672448 287048
rect 672500 287036 672506 287088
rect 674374 286968 674380 287020
rect 674432 287008 674438 287020
rect 675110 287008 675116 287020
rect 674432 286980 675116 287008
rect 674432 286968 674438 286980
rect 675110 286968 675116 286980
rect 675168 286968 675174 287020
rect 33778 286288 33784 286340
rect 33836 286328 33842 286340
rect 41690 286328 41696 286340
rect 33836 286300 41696 286328
rect 33836 286288 33842 286300
rect 41690 286288 41696 286300
rect 41748 286288 41754 286340
rect 46198 285676 46204 285728
rect 46256 285716 46262 285728
rect 62114 285716 62120 285728
rect 46256 285688 62120 285716
rect 46256 285676 46262 285688
rect 62114 285676 62120 285688
rect 62172 285676 62178 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 672074 285716 672080 285728
rect 651524 285688 672080 285716
rect 651524 285676 651530 285688
rect 672074 285676 672080 285688
rect 672132 285676 672138 285728
rect 59998 284384 60004 284436
rect 60056 284424 60062 284436
rect 62114 284424 62120 284436
rect 60056 284396 62120 284424
rect 60056 284384 60062 284396
rect 62114 284384 62120 284396
rect 62172 284384 62178 284436
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672626 284356 672632 284368
rect 651524 284328 672632 284356
rect 651524 284316 651530 284328
rect 672626 284316 672632 284328
rect 672684 284316 672690 284368
rect 651466 282888 651472 282940
rect 651524 282928 651530 282940
rect 667198 282928 667204 282940
rect 651524 282900 667204 282928
rect 651524 282888 651530 282900
rect 667198 282888 667204 282900
rect 667256 282888 667262 282940
rect 42242 281732 42248 281784
rect 42300 281772 42306 281784
rect 42610 281772 42616 281784
rect 42300 281744 42616 281772
rect 42300 281732 42306 281744
rect 42610 281732 42616 281744
rect 42668 281732 42674 281784
rect 47762 280304 47768 280356
rect 47820 280344 47826 280356
rect 62114 280344 62120 280356
rect 47820 280316 62120 280344
rect 47820 280304 47826 280316
rect 62114 280304 62120 280316
rect 62172 280304 62178 280356
rect 651466 280168 651472 280220
rect 651524 280208 651530 280220
rect 667382 280208 667388 280220
rect 651524 280180 667388 280208
rect 651524 280168 651530 280180
rect 667382 280168 667388 280180
rect 667440 280168 667446 280220
rect 42242 280100 42248 280152
rect 42300 280140 42306 280152
rect 42978 280140 42984 280152
rect 42300 280112 42984 280140
rect 42300 280100 42306 280112
rect 42978 280100 42984 280112
rect 43036 280100 43042 280152
rect 482830 277312 482836 277364
rect 482888 277352 482894 277364
rect 557534 277352 557540 277364
rect 482888 277324 557540 277352
rect 482888 277312 482894 277324
rect 557534 277312 557540 277324
rect 557592 277312 557598 277364
rect 485682 277176 485688 277228
rect 485740 277216 485746 277228
rect 562318 277216 562324 277228
rect 485740 277188 562324 277216
rect 485740 277176 485746 277188
rect 562318 277176 562324 277188
rect 562376 277176 562382 277228
rect 495066 277040 495072 277092
rect 495124 277080 495130 277092
rect 576486 277080 576492 277092
rect 495124 277052 576492 277080
rect 495124 277040 495130 277052
rect 576486 277040 576492 277052
rect 576544 277040 576550 277092
rect 511626 276904 511632 276956
rect 511684 276944 511690 276956
rect 600130 276944 600136 276956
rect 511684 276916 600136 276944
rect 511684 276904 511690 276916
rect 600130 276904 600136 276916
rect 600188 276904 600194 276956
rect 42242 276768 42248 276820
rect 42300 276808 42306 276820
rect 42610 276808 42616 276820
rect 42300 276780 42616 276808
rect 42300 276768 42306 276780
rect 42610 276768 42616 276780
rect 42668 276768 42674 276820
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 518710 276632 518716 276684
rect 518768 276672 518774 276684
rect 609606 276672 609612 276684
rect 518768 276644 609612 276672
rect 518768 276632 518774 276644
rect 609606 276632 609612 276644
rect 609664 276632 609670 276684
rect 478506 276496 478512 276548
rect 478564 276536 478570 276548
rect 551646 276536 551652 276548
rect 478564 276508 551652 276536
rect 478564 276496 478570 276508
rect 551646 276496 551652 276508
rect 551704 276496 551710 276548
rect 477034 276360 477040 276412
rect 477092 276400 477098 276412
rect 550450 276400 550456 276412
rect 477092 276372 550456 276400
rect 477092 276360 477098 276372
rect 550450 276360 550456 276372
rect 550508 276360 550514 276412
rect 471606 276224 471612 276276
rect 471664 276264 471670 276276
rect 543366 276264 543372 276276
rect 471664 276236 543372 276264
rect 471664 276224 471670 276236
rect 543366 276224 543372 276236
rect 543424 276224 543430 276276
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 162118 275992 162124 276004
rect 107252 275964 162124 275992
rect 107252 275952 107258 275964
rect 162118 275952 162124 275964
rect 162176 275952 162182 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 454402 275952 454408 276004
rect 454460 275992 454466 276004
rect 454460 275964 454724 275992
rect 454460 275952 454466 275964
rect 100110 275816 100116 275868
rect 100168 275856 100174 275868
rect 161382 275856 161388 275868
rect 100168 275828 161388 275856
rect 100168 275816 100174 275828
rect 161382 275816 161388 275828
rect 161440 275816 161446 275868
rect 161566 275816 161572 275868
rect 161624 275816 161630 275868
rect 161750 275816 161756 275868
rect 161808 275856 161814 275868
rect 166994 275856 167000 275868
rect 161808 275828 167000 275856
rect 161808 275816 161814 275828
rect 166994 275816 167000 275828
rect 167052 275816 167058 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 217134 275816 217140 275868
rect 217192 275856 217198 275868
rect 224034 275856 224040 275868
rect 217192 275828 224040 275856
rect 217192 275816 217198 275828
rect 224034 275816 224040 275828
rect 224092 275816 224098 275868
rect 232498 275816 232504 275868
rect 232556 275856 232562 275868
rect 239858 275856 239864 275868
rect 232556 275828 239864 275856
rect 232556 275816 232562 275828
rect 239858 275816 239864 275828
rect 239916 275816 239922 275868
rect 284570 275816 284576 275868
rect 284628 275856 284634 275868
rect 290090 275856 290096 275868
rect 284628 275828 290096 275856
rect 284628 275816 284634 275828
rect 290090 275816 290096 275828
rect 290148 275816 290154 275868
rect 445018 275816 445024 275868
rect 445076 275856 445082 275868
rect 454696 275856 454724 275964
rect 457438 275952 457444 276004
rect 457496 275992 457502 276004
rect 509050 275992 509056 276004
rect 457496 275964 509056 275992
rect 457496 275952 457502 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 517146 275952 517152 276004
rect 517204 275992 517210 276004
rect 608410 275992 608416 276004
rect 517204 275964 608416 275992
rect 517204 275952 517210 275964
rect 608410 275952 608416 275964
rect 608468 275952 608474 276004
rect 475378 275856 475384 275868
rect 445076 275828 454632 275856
rect 454696 275828 475384 275856
rect 445076 275816 445082 275828
rect 93026 275680 93032 275732
rect 93084 275720 93090 275732
rect 155954 275720 155960 275732
rect 93084 275692 155960 275720
rect 93084 275680 93090 275692
rect 155954 275680 155960 275692
rect 156012 275680 156018 275732
rect 161584 275720 161612 275816
rect 163130 275720 163136 275732
rect 161584 275692 163136 275720
rect 163130 275680 163136 275692
rect 163188 275680 163194 275732
rect 164050 275680 164056 275732
rect 164108 275720 164114 275732
rect 164108 275692 166488 275720
rect 164108 275680 164114 275692
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 156874 275544 156880 275596
rect 156932 275584 156938 275596
rect 166460 275584 166488 275692
rect 171042 275680 171048 275732
rect 171100 275720 171106 275732
rect 211062 275720 211068 275732
rect 171100 275692 211068 275720
rect 171100 275680 171106 275692
rect 211062 275680 211068 275692
rect 211120 275680 211126 275732
rect 224218 275680 224224 275732
rect 224276 275720 224282 275732
rect 232774 275720 232780 275732
rect 224276 275692 232780 275720
rect 224276 275680 224282 275692
rect 232774 275680 232780 275692
rect 232832 275680 232838 275732
rect 236086 275680 236092 275732
rect 236144 275720 236150 275732
rect 253382 275720 253388 275732
rect 236144 275692 253388 275720
rect 236144 275680 236150 275692
rect 253382 275680 253388 275692
rect 253440 275680 253446 275732
rect 435634 275680 435640 275732
rect 435692 275720 435698 275732
rect 454402 275720 454408 275732
rect 435692 275692 454408 275720
rect 435692 275680 435698 275692
rect 454402 275680 454408 275692
rect 454460 275680 454466 275732
rect 454604 275720 454632 275828
rect 475378 275816 475384 275828
rect 475436 275816 475442 275868
rect 479518 275816 479524 275868
rect 479576 275856 479582 275868
rect 523310 275856 523316 275868
rect 479576 275828 523316 275856
rect 479576 275816 479582 275828
rect 523310 275816 523316 275828
rect 523368 275816 523374 275868
rect 524138 275816 524144 275868
rect 524196 275856 524202 275868
rect 615494 275856 615500 275868
rect 524196 275828 615500 275856
rect 524196 275816 524202 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 498470 275720 498476 275732
rect 454604 275692 498476 275720
rect 498470 275680 498476 275692
rect 498528 275680 498534 275732
rect 507854 275680 507860 275732
rect 507912 275720 507918 275732
rect 545758 275720 545764 275732
rect 507912 275692 545764 275720
rect 507912 275680 507918 275692
rect 545758 275680 545764 275692
rect 545816 275680 545822 275732
rect 277486 275612 277492 275664
rect 277544 275652 277550 275664
rect 284294 275652 284300 275664
rect 277544 275624 284300 275652
rect 277544 275612 277550 275624
rect 284294 275612 284300 275624
rect 284352 275612 284358 275664
rect 206370 275584 206376 275596
rect 156932 275556 166304 275584
rect 166460 275556 206376 275584
rect 156932 275544 156938 275556
rect 81250 275408 81256 275460
rect 81308 275448 81314 275460
rect 145558 275448 145564 275460
rect 81308 275420 145564 275448
rect 81308 275408 81314 275420
rect 145558 275408 145564 275420
rect 145616 275408 145622 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 161842 275448 161848 275460
rect 160520 275420 161848 275448
rect 160520 275408 160526 275420
rect 161842 275408 161848 275420
rect 161900 275408 161906 275460
rect 166276 275448 166304 275556
rect 206370 275544 206376 275556
rect 206428 275544 206434 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 239398 275584 239404 275596
rect 221976 275556 239404 275584
rect 221976 275544 221982 275556
rect 239398 275544 239404 275556
rect 239456 275544 239462 275596
rect 243170 275544 243176 275596
rect 243228 275584 243234 275596
rect 255314 275584 255320 275596
rect 243228 275556 255320 275584
rect 243228 275544 243234 275556
rect 255314 275544 255320 275556
rect 255372 275544 255378 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262858 275584 262864 275596
rect 257396 275556 262864 275584
rect 257396 275544 257402 275556
rect 262858 275544 262864 275556
rect 262916 275544 262922 275596
rect 286870 275544 286876 275596
rect 286928 275584 286934 275596
rect 291838 275584 291844 275596
rect 286928 275556 291844 275584
rect 286928 275544 286934 275556
rect 291838 275544 291844 275556
rect 291896 275544 291902 275596
rect 430206 275544 430212 275596
rect 430264 275584 430270 275596
rect 484302 275584 484308 275596
rect 430264 275556 484308 275584
rect 430264 275544 430270 275556
rect 484302 275544 484308 275556
rect 484360 275544 484366 275596
rect 501598 275544 501604 275596
rect 501656 275584 501662 275596
rect 512638 275584 512644 275596
rect 501656 275556 512644 275584
rect 501656 275544 501662 275556
rect 512638 275544 512644 275556
rect 512696 275544 512702 275596
rect 515398 275544 515404 275596
rect 515456 275584 515462 275596
rect 526806 275584 526812 275596
rect 515456 275556 526812 275584
rect 515456 275544 515462 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 528186 275544 528192 275596
rect 528244 275584 528250 275596
rect 622578 275584 622584 275596
rect 528244 275556 622584 275584
rect 528244 275544 528250 275556
rect 622578 275544 622584 275556
rect 622636 275544 622642 275596
rect 198734 275448 198740 275460
rect 166276 275420 198740 275448
rect 198734 275408 198740 275420
rect 198792 275408 198798 275460
rect 214834 275408 214840 275460
rect 214892 275448 214898 275460
rect 236638 275448 236644 275460
rect 214892 275420 236644 275448
rect 214892 275408 214898 275420
rect 236638 275408 236644 275420
rect 236696 275408 236702 275460
rect 239582 275408 239588 275460
rect 239640 275448 239646 275460
rect 251910 275448 251916 275460
rect 239640 275420 251916 275448
rect 239640 275408 239646 275420
rect 251910 275408 251916 275420
rect 251968 275408 251974 275460
rect 263226 275408 263232 275460
rect 263284 275448 263290 275460
rect 273254 275448 273260 275460
rect 263284 275420 273260 275448
rect 263284 275408 263290 275420
rect 273254 275408 273260 275420
rect 273312 275408 273318 275460
rect 285674 275408 285680 275460
rect 285732 275448 285738 275460
rect 291194 275448 291200 275460
rect 285732 275420 291200 275448
rect 285732 275408 285738 275420
rect 291194 275408 291200 275420
rect 291252 275408 291258 275460
rect 291654 275408 291660 275460
rect 291712 275448 291718 275460
rect 295426 275448 295432 275460
rect 291712 275420 295432 275448
rect 291712 275408 291718 275420
rect 295426 275408 295432 275420
rect 295484 275408 295490 275460
rect 386046 275408 386052 275460
rect 386104 275448 386110 275460
rect 420454 275448 420460 275460
rect 386104 275420 420460 275448
rect 386104 275408 386110 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 423398 275408 423404 275460
rect 423456 275448 423462 275460
rect 473354 275448 473360 275460
rect 423456 275420 473360 275448
rect 423456 275408 423462 275420
rect 473354 275408 473360 275420
rect 473412 275408 473418 275460
rect 475378 275408 475384 275460
rect 475436 275448 475442 275460
rect 485038 275448 485044 275460
rect 475436 275420 485044 275448
rect 475436 275408 475442 275420
rect 485038 275408 485044 275420
rect 485096 275408 485102 275460
rect 485222 275408 485228 275460
rect 485280 275448 485286 275460
rect 537478 275448 537484 275460
rect 485280 275420 537484 275448
rect 485280 275408 485286 275420
rect 537478 275408 537484 275420
rect 537536 275408 537542 275460
rect 636746 275448 636752 275460
rect 537772 275420 636752 275448
rect 297542 275340 297548 275392
rect 297600 275380 297606 275392
rect 299566 275380 299572 275392
rect 297600 275352 299572 275380
rect 297600 275340 297606 275352
rect 299566 275340 299572 275352
rect 299624 275340 299630 275392
rect 299934 275340 299940 275392
rect 299992 275380 299998 275392
rect 301130 275380 301136 275392
rect 299992 275352 301136 275380
rect 299992 275340 299998 275352
rect 301130 275340 301136 275352
rect 301188 275340 301194 275392
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 141050 275312 141056 275324
rect 71832 275284 141056 275312
rect 71832 275272 71838 275284
rect 141050 275272 141056 275284
rect 141108 275272 141114 275324
rect 146202 275272 146208 275324
rect 146260 275312 146266 275324
rect 189074 275312 189080 275324
rect 146260 275284 189080 275312
rect 146260 275272 146266 275284
rect 189074 275272 189080 275284
rect 189132 275272 189138 275324
rect 218330 275272 218336 275324
rect 218388 275312 218394 275324
rect 243078 275312 243084 275324
rect 218388 275284 243084 275312
rect 218388 275272 218394 275284
rect 243078 275272 243084 275284
rect 243136 275272 243142 275324
rect 256142 275272 256148 275324
rect 256200 275312 256206 275324
rect 268654 275312 268660 275324
rect 256200 275284 268660 275312
rect 256200 275272 256206 275284
rect 268654 275272 268660 275284
rect 268712 275272 268718 275324
rect 273898 275272 273904 275324
rect 273956 275312 273962 275324
rect 282914 275312 282920 275324
rect 273956 275284 282920 275312
rect 273956 275272 273962 275284
rect 282914 275272 282920 275284
rect 282972 275272 282978 275324
rect 361206 275272 361212 275324
rect 361264 275312 361270 275324
rect 385034 275312 385040 275324
rect 361264 275284 385040 275312
rect 361264 275272 361270 275284
rect 385034 275272 385040 275284
rect 385092 275272 385098 275324
rect 416406 275272 416412 275324
rect 416464 275312 416470 275324
rect 462958 275312 462964 275324
rect 416464 275284 462964 275312
rect 416464 275272 416470 275284
rect 462958 275272 462964 275284
rect 463016 275272 463022 275324
rect 463142 275272 463148 275324
rect 463200 275312 463206 275324
rect 530394 275312 530400 275324
rect 463200 275284 530400 275312
rect 463200 275272 463206 275284
rect 530394 275272 530400 275284
rect 530452 275272 530458 275324
rect 532326 275272 532332 275324
rect 532384 275312 532390 275324
rect 537294 275312 537300 275324
rect 532384 275284 537300 275312
rect 532384 275272 532390 275284
rect 537294 275272 537300 275284
rect 537352 275272 537358 275324
rect 537570 275272 537576 275324
rect 537628 275312 537634 275324
rect 537772 275312 537800 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 537628 275284 537800 275312
rect 537628 275272 537634 275284
rect 537938 275272 537944 275324
rect 537996 275312 538002 275324
rect 540974 275312 540980 275324
rect 537996 275284 540980 275312
rect 537996 275272 538002 275284
rect 540974 275272 540980 275284
rect 541032 275272 541038 275324
rect 542998 275272 543004 275324
rect 543056 275312 543062 275324
rect 629662 275312 629668 275324
rect 543056 275284 629668 275312
rect 543056 275272 543062 275284
rect 629662 275272 629668 275284
rect 629720 275272 629726 275324
rect 290458 275204 290464 275256
rect 290516 275244 290522 275256
rect 294138 275244 294144 275256
rect 290516 275216 294144 275244
rect 290516 275204 290522 275216
rect 294138 275204 294144 275216
rect 294196 275204 294202 275256
rect 298738 275204 298744 275256
rect 298796 275244 298802 275256
rect 300026 275244 300032 275256
rect 298796 275216 300032 275244
rect 298796 275204 298802 275216
rect 300026 275204 300032 275216
rect 300084 275204 300090 275256
rect 139118 275136 139124 275188
rect 139176 275176 139182 275188
rect 146938 275176 146944 275188
rect 139176 275148 146944 275176
rect 139176 275136 139182 275148
rect 146938 275136 146944 275148
rect 146996 275136 147002 275188
rect 149790 275136 149796 275188
rect 149848 275176 149854 275188
rect 191742 275176 191748 275188
rect 149848 275148 191748 275176
rect 149848 275136 149854 275148
rect 191742 275136 191748 275148
rect 191800 275136 191806 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 485038 275136 485044 275188
rect 485096 275176 485102 275188
rect 491386 275176 491392 275188
rect 485096 275148 491392 275176
rect 485096 275136 485102 275148
rect 491386 275136 491392 275148
rect 491444 275136 491450 275188
rect 493318 275136 493324 275188
rect 493376 275176 493382 275188
rect 493376 275148 495112 275176
rect 493376 275136 493382 275148
rect 269206 275068 269212 275120
rect 269264 275108 269270 275120
rect 274910 275108 274916 275120
rect 269264 275080 274916 275108
rect 269264 275068 269270 275080
rect 274910 275068 274916 275080
rect 274968 275068 274974 275120
rect 110782 275000 110788 275052
rect 110840 275040 110846 275052
rect 149698 275040 149704 275052
rect 110840 275012 149704 275040
rect 110840 275000 110846 275012
rect 149698 275000 149704 275012
rect 149756 275000 149762 275052
rect 153378 275000 153384 275052
rect 153436 275040 153442 275052
rect 154482 275040 154488 275052
rect 153436 275012 154488 275040
rect 153436 275000 153442 275012
rect 154482 275000 154488 275012
rect 154540 275000 154546 275052
rect 161658 275040 161664 275052
rect 161446 275012 161664 275040
rect 132034 274864 132040 274916
rect 132092 274904 132098 274916
rect 161446 274904 161474 275012
rect 161658 275000 161664 275012
rect 161716 275000 161722 275052
rect 161842 275000 161848 275052
rect 161900 275040 161906 275052
rect 175918 275040 175924 275052
rect 161900 275012 175924 275040
rect 161900 275000 161906 275012
rect 175918 275000 175924 275012
rect 175976 275000 175982 275052
rect 189994 275000 190000 275052
rect 190052 275040 190058 275052
rect 218698 275040 218704 275052
rect 190052 275012 218704 275040
rect 190052 275000 190058 275012
rect 218698 275000 218704 275012
rect 218756 275000 218762 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292666 275040 292672 275052
rect 288124 275012 292672 275040
rect 288124 275000 288130 275012
rect 292666 275000 292672 275012
rect 292724 275000 292730 275052
rect 420638 275000 420644 275052
rect 420696 275040 420702 275052
rect 470134 275040 470140 275052
rect 420696 275012 470140 275040
rect 420696 275000 420702 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 476114 275000 476120 275052
rect 476172 275040 476178 275052
rect 485222 275040 485228 275052
rect 476172 275012 485228 275040
rect 476172 275000 476178 275012
rect 485222 275000 485228 275012
rect 485280 275000 485286 275052
rect 492398 275000 492404 275052
rect 492456 275040 492462 275052
rect 494882 275040 494888 275052
rect 492456 275012 494888 275040
rect 492456 275000 492462 275012
rect 494882 275000 494888 275012
rect 494940 275000 494946 275052
rect 495084 275040 495112 275148
rect 497458 275136 497464 275188
rect 497516 275176 497522 275188
rect 505554 275176 505560 275188
rect 497516 275148 505560 275176
rect 497516 275136 497522 275148
rect 505554 275136 505560 275148
rect 505612 275136 505618 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 501966 275040 501972 275052
rect 495084 275012 501972 275040
rect 501966 275000 501972 275012
rect 502024 275000 502030 275052
rect 503438 275000 503444 275052
rect 503496 275040 503502 275052
rect 587066 275040 587072 275052
rect 503496 275012 587072 275040
rect 503496 275000 503502 275012
rect 587066 275000 587072 275012
rect 587124 275000 587130 275052
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 296806 274972 296812 274984
rect 294012 274944 296812 274972
rect 294012 274932 294018 274944
rect 296806 274932 296812 274944
rect 296864 274932 296870 274984
rect 132092 274876 161474 274904
rect 132092 274864 132098 274876
rect 167546 274864 167552 274916
rect 167604 274904 167610 274916
rect 169018 274904 169024 274916
rect 167604 274876 169024 274904
rect 167604 274864 167610 274876
rect 169018 274864 169024 274876
rect 169076 274864 169082 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 293402 274904 293408 274916
rect 289320 274876 293408 274904
rect 289320 274864 289326 274876
rect 293402 274864 293408 274876
rect 293460 274864 293466 274916
rect 413462 274864 413468 274916
rect 413520 274904 413526 274916
rect 459462 274904 459468 274916
rect 413520 274876 459468 274904
rect 413520 274864 413526 274876
rect 459462 274864 459468 274876
rect 459520 274864 459526 274916
rect 473354 274864 473360 274916
rect 473412 274904 473418 274916
rect 544562 274904 544568 274916
rect 473412 274876 544568 274904
rect 473412 274864 473418 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 122668 274808 122834 274836
rect 103698 274728 103704 274780
rect 103756 274768 103762 274780
rect 104802 274768 104808 274780
rect 103756 274740 104808 274768
rect 103756 274728 103762 274740
rect 104802 274728 104808 274740
rect 104860 274728 104866 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76742 274700 76748 274712
rect 74224 274672 76748 274700
rect 74224 274660 74230 274672
rect 76742 274660 76748 274672
rect 76800 274660 76806 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 117682 274632 117688 274644
rect 103486 274604 117688 274632
rect 96614 274524 96620 274576
rect 96672 274564 96678 274576
rect 103486 274564 103514 274604
rect 117682 274592 117688 274604
rect 117740 274592 117746 274644
rect 117866 274592 117872 274644
rect 117924 274632 117930 274644
rect 122668 274632 122696 274808
rect 117924 274604 122696 274632
rect 122806 274632 122834 274808
rect 174630 274796 174636 274848
rect 174688 274836 174694 274848
rect 182726 274836 182732 274848
rect 174688 274808 182732 274836
rect 174688 274796 174694 274808
rect 182726 274796 182732 274808
rect 182784 274796 182790 274848
rect 295150 274796 295156 274848
rect 295208 274836 295214 274848
rect 297450 274836 297456 274848
rect 295208 274808 297456 274836
rect 295208 274796 295214 274808
rect 297450 274796 297456 274808
rect 297508 274796 297514 274848
rect 136818 274728 136824 274780
rect 136876 274768 136882 274780
rect 137646 274768 137652 274780
rect 136876 274740 137652 274768
rect 136876 274728 136882 274740
rect 137646 274728 137652 274740
rect 137704 274728 137710 274780
rect 143902 274728 143908 274780
rect 143960 274768 143966 274780
rect 144362 274768 144368 274780
rect 143960 274740 144368 274768
rect 143960 274728 143966 274740
rect 144362 274728 144368 274740
rect 144420 274728 144426 274780
rect 146938 274728 146944 274780
rect 146996 274768 147002 274780
rect 174446 274768 174452 274780
rect 146996 274740 174452 274768
rect 146996 274728 147002 274740
rect 174446 274728 174452 274740
rect 174504 274728 174510 274780
rect 469858 274728 469864 274780
rect 469916 274768 469922 274780
rect 516226 274768 516232 274780
rect 469916 274740 516232 274768
rect 469916 274728 469922 274740
rect 516226 274728 516232 274740
rect 516284 274728 516290 274780
rect 526438 274728 526444 274780
rect 526496 274768 526502 274780
rect 533890 274768 533896 274780
rect 526496 274740 533896 274768
rect 526496 274728 526502 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 537938 274768 537944 274780
rect 534776 274740 537944 274768
rect 534776 274728 534782 274740
rect 537938 274728 537944 274740
rect 537996 274728 538002 274780
rect 538122 274728 538128 274780
rect 538180 274768 538186 274780
rect 542998 274768 543004 274780
rect 538180 274740 543004 274768
rect 538180 274728 538186 274740
rect 542998 274728 543004 274740
rect 543056 274728 543062 274780
rect 543182 274728 543188 274780
rect 543240 274768 543246 274780
rect 643830 274768 643836 274780
rect 543240 274740 643836 274768
rect 543240 274728 543246 274740
rect 643830 274728 643836 274740
rect 643888 274728 643894 274780
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 258350 274700 258356 274712
rect 253900 274672 258356 274700
rect 253900 274660 253906 274672
rect 258350 274660 258356 274672
rect 258408 274660 258414 274712
rect 268010 274660 268016 274712
rect 268068 274700 268074 274712
rect 272426 274700 272432 274712
rect 268068 274672 272432 274700
rect 268068 274660 268074 274672
rect 272426 274660 272432 274672
rect 272484 274660 272490 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 292850 274660 292856 274712
rect 292908 274700 292914 274712
rect 295794 274700 295800 274712
rect 292908 274672 295800 274700
rect 292908 274660 292914 274672
rect 295794 274660 295800 274672
rect 295852 274660 295858 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 350718 274660 350724 274712
rect 350776 274700 350782 274712
rect 353110 274700 353116 274712
rect 350776 274672 353116 274700
rect 350776 274660 350782 274672
rect 353110 274660 353116 274672
rect 353168 274660 353174 274712
rect 174170 274632 174176 274644
rect 122806 274604 174176 274632
rect 117924 274592 117930 274604
rect 174170 274592 174176 274604
rect 174228 274592 174234 274644
rect 182910 274592 182916 274644
rect 182968 274632 182974 274644
rect 214558 274632 214564 274644
rect 182968 274604 214564 274632
rect 182968 274592 182974 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 382918 274592 382924 274644
rect 382976 274632 382982 274644
rect 392118 274632 392124 274644
rect 382976 274604 392124 274632
rect 382976 274592 382982 274604
rect 392118 274592 392124 274604
rect 392176 274592 392182 274644
rect 404170 274592 404176 274644
rect 404228 274632 404234 274644
rect 446490 274632 446496 274644
rect 404228 274604 446496 274632
rect 404228 274592 404234 274604
rect 446490 274592 446496 274604
rect 446548 274592 446554 274644
rect 450538 274592 450544 274644
rect 450596 274632 450602 274644
rect 480714 274632 480720 274644
rect 450596 274604 480720 274632
rect 450596 274592 450602 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 488350 274592 488356 274644
rect 488408 274632 488414 274644
rect 567010 274632 567016 274644
rect 488408 274604 567016 274632
rect 488408 274592 488414 274604
rect 567010 274592 567016 274604
rect 567068 274592 567074 274644
rect 96672 274536 103514 274564
rect 96672 274524 96678 274536
rect 95878 274496 95884 274508
rect 84166 274468 95884 274496
rect 67082 274320 67088 274372
rect 67140 274360 67146 274372
rect 84166 274360 84194 274468
rect 95878 274456 95884 274468
rect 95936 274456 95942 274508
rect 105170 274456 105176 274508
rect 105228 274496 105234 274508
rect 163314 274496 163320 274508
rect 105228 274468 163320 274496
rect 105228 274456 105234 274468
rect 163314 274456 163320 274468
rect 163372 274456 163378 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208486 274496 208492 274508
rect 168800 274468 208492 274496
rect 168800 274456 168806 274468
rect 208486 274456 208492 274468
rect 208544 274456 208550 274508
rect 227806 274456 227812 274508
rect 227864 274496 227870 274508
rect 248874 274496 248880 274508
rect 227864 274468 248880 274496
rect 227864 274456 227870 274468
rect 248874 274456 248880 274468
rect 248932 274456 248938 274508
rect 358078 274456 358084 274508
rect 358136 274496 358142 274508
rect 369578 274496 369584 274508
rect 358136 274468 369584 274496
rect 358136 274456 358142 274468
rect 369578 274456 369584 274468
rect 369636 274456 369642 274508
rect 395614 274496 395620 274508
rect 369780 274468 395620 274496
rect 67140 274332 84194 274360
rect 67140 274320 67146 274332
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 166350 274320 166356 274372
rect 166408 274360 166414 274372
rect 207290 274360 207296 274372
rect 166408 274332 207296 274360
rect 166408 274320 166414 274332
rect 207290 274320 207296 274332
rect 207348 274320 207354 274372
rect 207750 274320 207756 274372
rect 207808 274360 207814 274372
rect 233878 274360 233884 274372
rect 207808 274332 233884 274360
rect 207808 274320 207814 274332
rect 233878 274320 233884 274332
rect 233936 274320 233942 274372
rect 249058 274320 249064 274372
rect 249116 274360 249122 274372
rect 265250 274360 265256 274372
rect 249116 274332 265256 274360
rect 249116 274320 249122 274332
rect 265250 274320 265256 274332
rect 265308 274320 265314 274372
rect 333790 274320 333796 274372
rect 333848 274360 333854 274372
rect 345934 274360 345940 274372
rect 333848 274332 345940 274360
rect 333848 274320 333854 274332
rect 345934 274320 345940 274332
rect 345992 274320 345998 274372
rect 347038 274320 347044 274372
rect 347096 274360 347102 274372
rect 358998 274360 359004 274372
rect 347096 274332 359004 274360
rect 347096 274320 347102 274332
rect 358998 274320 359004 274332
rect 359056 274320 359062 274372
rect 369302 274320 369308 274372
rect 369360 274360 369366 274372
rect 369780 274360 369808 274468
rect 395614 274456 395620 274468
rect 395672 274456 395678 274508
rect 409230 274456 409236 274508
rect 409288 274496 409294 274508
rect 453574 274496 453580 274508
rect 409288 274468 453580 274496
rect 409288 274456 409294 274468
rect 453574 274456 453580 274468
rect 453632 274456 453638 274508
rect 453758 274456 453764 274508
rect 453816 274496 453822 274508
rect 486602 274496 486608 274508
rect 453816 274468 486608 274496
rect 453816 274456 453822 274468
rect 486602 274456 486608 274468
rect 486660 274456 486666 274508
rect 536742 274456 536748 274508
rect 536800 274496 536806 274508
rect 634354 274496 634360 274508
rect 536800 274468 634360 274496
rect 536800 274456 536806 274468
rect 634354 274456 634360 274468
rect 634412 274456 634418 274508
rect 369360 274332 369808 274360
rect 369360 274320 369366 274332
rect 373258 274320 373264 274372
rect 373316 274360 373322 274372
rect 400306 274360 400312 274372
rect 373316 274332 400312 274360
rect 373316 274320 373322 274332
rect 400306 274320 400312 274332
rect 400364 274320 400370 274372
rect 413830 274320 413836 274372
rect 413888 274360 413894 274372
rect 460658 274360 460664 274372
rect 413888 274332 460664 274360
rect 413888 274320 413894 274332
rect 460658 274320 460664 274332
rect 460716 274320 460722 274372
rect 465718 274320 465724 274372
rect 465776 274360 465782 274372
rect 487798 274360 487804 274372
rect 465776 274332 487804 274360
rect 465776 274320 465782 274332
rect 487798 274320 487804 274332
rect 487856 274320 487862 274372
rect 508590 274320 508596 274372
rect 508648 274360 508654 274372
rect 595070 274360 595076 274372
rect 508648 274332 595076 274360
rect 508648 274320 508654 274332
rect 595070 274320 595076 274332
rect 595128 274320 595134 274372
rect 595438 274320 595444 274372
rect 595496 274360 595502 274372
rect 640334 274360 640340 274372
rect 595496 274332 640340 274360
rect 595496 274320 595502 274332
rect 640334 274320 640340 274332
rect 640392 274320 640398 274372
rect 282178 274252 282184 274304
rect 282236 274292 282242 274304
rect 287698 274292 287704 274304
rect 282236 274264 287704 274292
rect 282236 274252 282242 274264
rect 287698 274252 287704 274264
rect 287756 274252 287762 274304
rect 89438 274184 89444 274236
rect 89496 274224 89502 274236
rect 151998 274224 152004 274236
rect 89496 274196 152004 274224
rect 89496 274184 89502 274196
rect 151998 274184 152004 274196
rect 152056 274184 152062 274236
rect 155678 274184 155684 274236
rect 155736 274224 155742 274236
rect 200114 274224 200120 274236
rect 155736 274196 200120 274224
rect 155736 274184 155742 274196
rect 200114 274184 200120 274196
rect 200172 274184 200178 274236
rect 205358 274184 205364 274236
rect 205416 274224 205422 274236
rect 234706 274224 234712 274236
rect 205416 274196 234712 274224
rect 205416 274184 205422 274196
rect 234706 274184 234712 274196
rect 234764 274184 234770 274236
rect 237282 274184 237288 274236
rect 237340 274224 237346 274236
rect 256970 274224 256976 274236
rect 237340 274196 256976 274224
rect 237340 274184 237346 274196
rect 256970 274184 256976 274196
rect 257028 274184 257034 274236
rect 325326 274184 325332 274236
rect 325384 274224 325390 274236
rect 332962 274224 332968 274236
rect 325384 274196 332968 274224
rect 325384 274184 325390 274196
rect 332962 274184 332968 274196
rect 333020 274184 333026 274236
rect 343450 274184 343456 274236
rect 343508 274224 343514 274236
rect 360194 274224 360200 274236
rect 343508 274196 360200 274224
rect 343508 274184 343514 274196
rect 360194 274184 360200 274196
rect 360252 274184 360258 274236
rect 364978 274184 364984 274236
rect 365036 274224 365042 274236
rect 374362 274224 374368 274236
rect 365036 274196 374368 274224
rect 365036 274184 365042 274196
rect 374362 274184 374368 274196
rect 374420 274184 374426 274236
rect 379330 274184 379336 274236
rect 379388 274224 379394 274236
rect 410978 274224 410984 274236
rect 379388 274196 410984 274224
rect 379388 274184 379394 274196
rect 410978 274184 410984 274196
rect 411036 274184 411042 274236
rect 416590 274184 416596 274236
rect 416648 274224 416654 274236
rect 464154 274224 464160 274236
rect 416648 274196 464160 274224
rect 416648 274184 416654 274196
rect 464154 274184 464160 274196
rect 464212 274184 464218 274236
rect 474366 274184 474372 274236
rect 474424 274224 474430 274236
rect 507854 274224 507860 274236
rect 474424 274196 507860 274224
rect 474424 274184 474430 274196
rect 507854 274184 507860 274196
rect 507912 274184 507918 274236
rect 511810 274184 511816 274236
rect 511868 274224 511874 274236
rect 598934 274224 598940 274236
rect 511868 274196 598940 274224
rect 511868 274184 511874 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 77720 274060 142154 274088
rect 77720 274048 77726 274060
rect 65886 273912 65892 273964
rect 65944 273952 65950 273964
rect 136818 273952 136824 273964
rect 65944 273924 136824 273952
rect 65944 273912 65950 273924
rect 136818 273912 136824 273924
rect 136876 273912 136882 273964
rect 142126 273952 142154 274060
rect 145098 274048 145104 274100
rect 145156 274088 145162 274100
rect 192386 274088 192392 274100
rect 145156 274060 192392 274088
rect 145156 274048 145162 274060
rect 192386 274048 192392 274060
rect 192444 274048 192450 274100
rect 198274 274048 198280 274100
rect 198332 274088 198338 274100
rect 229186 274088 229192 274100
rect 198332 274060 229192 274088
rect 198332 274048 198338 274060
rect 229186 274048 229192 274060
rect 229244 274048 229250 274100
rect 234890 274048 234896 274100
rect 234948 274088 234954 274100
rect 234948 274060 251956 274088
rect 234948 274048 234954 274060
rect 145098 273952 145104 273964
rect 142126 273924 145104 273952
rect 145098 273912 145104 273924
rect 145156 273912 145162 273964
rect 147398 273912 147404 273964
rect 147456 273952 147462 273964
rect 193398 273952 193404 273964
rect 147456 273924 193404 273952
rect 147456 273912 147462 273924
rect 193398 273912 193404 273924
rect 193456 273912 193462 273964
rect 195882 273912 195888 273964
rect 195940 273952 195946 273964
rect 227898 273952 227904 273964
rect 195940 273924 227904 273952
rect 195940 273912 195946 273924
rect 227898 273912 227904 273924
rect 227956 273912 227962 273964
rect 229002 273912 229008 273964
rect 229060 273952 229066 273964
rect 250438 273952 250444 273964
rect 229060 273924 250444 273952
rect 229060 273912 229066 273924
rect 250438 273912 250444 273924
rect 250496 273912 250502 273964
rect 251928 273952 251956 274060
rect 255314 274048 255320 274100
rect 255372 274088 255378 274100
rect 261018 274088 261024 274100
rect 255372 274060 261024 274088
rect 255372 274048 255378 274060
rect 261018 274048 261024 274060
rect 261076 274048 261082 274100
rect 261202 274048 261208 274100
rect 261260 274088 261266 274100
rect 273530 274088 273536 274100
rect 261260 274060 273536 274088
rect 261260 274048 261266 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 275094 274048 275100 274100
rect 275152 274088 275158 274100
rect 283466 274088 283472 274100
rect 275152 274060 283472 274088
rect 275152 274048 275158 274060
rect 283466 274048 283472 274060
rect 283524 274048 283530 274100
rect 332318 274048 332324 274100
rect 332376 274088 332382 274100
rect 343634 274088 343640 274100
rect 332376 274060 343640 274088
rect 332376 274048 332382 274060
rect 343634 274048 343640 274060
rect 343692 274048 343698 274100
rect 350350 274048 350356 274100
rect 350408 274088 350414 274100
rect 368474 274088 368480 274100
rect 350408 274060 368480 274088
rect 350408 274048 350414 274060
rect 368474 274048 368480 274060
rect 368532 274048 368538 274100
rect 369118 274048 369124 274100
rect 369176 274088 369182 274100
rect 387334 274088 387340 274100
rect 369176 274060 387340 274088
rect 369176 274048 369182 274060
rect 387334 274048 387340 274060
rect 387392 274048 387398 274100
rect 394326 274048 394332 274100
rect 394384 274088 394390 274100
rect 432230 274088 432236 274100
rect 394384 274060 432236 274088
rect 394384 274048 394390 274060
rect 432230 274048 432236 274060
rect 432288 274048 432294 274100
rect 432598 274048 432604 274100
rect 432656 274088 432662 274100
rect 485498 274088 485504 274100
rect 432656 274060 485504 274088
rect 432656 274048 432662 274060
rect 485498 274048 485504 274060
rect 485556 274048 485562 274100
rect 491202 274048 491208 274100
rect 491260 274088 491266 274100
rect 569954 274088 569960 274100
rect 491260 274060 569960 274088
rect 491260 274048 491266 274060
rect 569954 274048 569960 274060
rect 570012 274048 570018 274100
rect 571978 274048 571984 274100
rect 572036 274088 572042 274100
rect 583570 274088 583576 274100
rect 572036 274060 583576 274088
rect 572036 274048 572042 274060
rect 583570 274048 583576 274060
rect 583628 274048 583634 274100
rect 255406 273952 255412 273964
rect 251928 273924 255412 273952
rect 255406 273912 255412 273924
rect 255464 273912 255470 273964
rect 258534 273912 258540 273964
rect 258592 273952 258598 273964
rect 272058 273952 272064 273964
rect 258592 273924 272064 273952
rect 258592 273912 258598 273924
rect 272058 273912 272064 273924
rect 272116 273912 272122 273964
rect 272702 273912 272708 273964
rect 272760 273952 272766 273964
rect 281810 273952 281816 273964
rect 272760 273924 281816 273952
rect 272760 273912 272766 273924
rect 281810 273912 281816 273924
rect 281868 273912 281874 273964
rect 324038 273912 324044 273964
rect 324096 273952 324102 273964
rect 331766 273952 331772 273964
rect 324096 273924 331772 273952
rect 324096 273912 324102 273924
rect 331766 273912 331772 273924
rect 331824 273912 331830 273964
rect 331950 273912 331956 273964
rect 332008 273952 332014 273964
rect 341242 273952 341248 273964
rect 332008 273924 341248 273952
rect 332008 273912 332014 273924
rect 341242 273912 341248 273924
rect 341300 273912 341306 273964
rect 342070 273912 342076 273964
rect 342128 273952 342134 273964
rect 357802 273952 357808 273964
rect 342128 273924 357808 273952
rect 342128 273912 342134 273924
rect 357802 273912 357808 273924
rect 357860 273912 357866 273964
rect 360102 273912 360108 273964
rect 360160 273952 360166 273964
rect 382642 273952 382648 273964
rect 360160 273924 382648 273952
rect 360160 273912 360166 273924
rect 382642 273912 382648 273924
rect 382700 273912 382706 273964
rect 387426 273912 387432 273964
rect 387484 273952 387490 273964
rect 421650 273952 421656 273964
rect 387484 273924 421656 273952
rect 387484 273912 387490 273924
rect 421650 273912 421656 273924
rect 421708 273912 421714 273964
rect 421834 273912 421840 273964
rect 421892 273952 421898 273964
rect 471238 273952 471244 273964
rect 421892 273924 471244 273952
rect 421892 273912 421898 273924
rect 471238 273912 471244 273924
rect 471296 273912 471302 273964
rect 475746 273912 475752 273964
rect 475804 273952 475810 273964
rect 547506 273952 547512 273964
rect 475804 273924 547512 273952
rect 475804 273912 475810 273924
rect 547506 273912 547512 273924
rect 547564 273912 547570 273964
rect 547690 273912 547696 273964
rect 547748 273952 547754 273964
rect 639138 273952 639144 273964
rect 547748 273924 639144 273952
rect 547748 273912 547754 273924
rect 639138 273912 639144 273924
rect 639196 273912 639202 273964
rect 113450 273776 113456 273828
rect 113508 273816 113514 273828
rect 169938 273816 169944 273828
rect 113508 273788 169944 273816
rect 113508 273776 113514 273788
rect 169938 273776 169944 273788
rect 169996 273776 170002 273828
rect 175918 273776 175924 273828
rect 175976 273816 175982 273828
rect 204254 273816 204260 273828
rect 175976 273788 204260 273816
rect 175976 273776 175982 273788
rect 204254 273776 204260 273788
rect 204312 273776 204318 273828
rect 206554 273776 206560 273828
rect 206612 273816 206618 273828
rect 235442 273816 235448 273828
rect 206612 273788 235448 273816
rect 206612 273776 206618 273788
rect 235442 273776 235448 273788
rect 235500 273776 235506 273828
rect 400122 273776 400128 273828
rect 400180 273816 400186 273828
rect 439314 273816 439320 273828
rect 400180 273788 439320 273816
rect 400180 273776 400186 273788
rect 439314 273776 439320 273788
rect 439372 273776 439378 273828
rect 442258 273776 442264 273828
rect 442316 273816 442322 273828
rect 481910 273816 481916 273828
rect 442316 273788 481916 273816
rect 442316 273776 442322 273788
rect 481910 273776 481916 273788
rect 481968 273776 481974 273828
rect 487062 273776 487068 273828
rect 487120 273816 487126 273828
rect 487120 273788 562456 273816
rect 487120 273776 487126 273788
rect 123754 273640 123760 273692
rect 123812 273680 123818 273692
rect 177482 273680 177488 273692
rect 123812 273652 177488 273680
rect 123812 273640 123818 273652
rect 177482 273640 177488 273652
rect 177540 273640 177546 273692
rect 392578 273640 392584 273692
rect 392636 273680 392642 273692
rect 409782 273680 409788 273692
rect 392636 273652 409788 273680
rect 392636 273640 392642 273652
rect 409782 273640 409788 273652
rect 409840 273640 409846 273692
rect 440878 273640 440884 273692
rect 440936 273680 440942 273692
rect 474826 273680 474832 273692
rect 440936 273652 474832 273680
rect 440936 273640 440942 273652
rect 474826 273640 474832 273652
rect 474884 273640 474890 273692
rect 484302 273640 484308 273692
rect 484360 273680 484366 273692
rect 552658 273680 552664 273692
rect 484360 273652 552664 273680
rect 484360 273640 484366 273652
rect 552658 273640 552664 273652
rect 552716 273640 552722 273692
rect 552842 273640 552848 273692
rect 552900 273680 552906 273692
rect 562226 273680 562232 273692
rect 552900 273652 562232 273680
rect 552900 273640 552906 273652
rect 562226 273640 562232 273652
rect 562284 273640 562290 273692
rect 562428 273680 562456 273788
rect 562594 273776 562600 273828
rect 562652 273816 562658 273828
rect 571978 273816 571984 273828
rect 562652 273788 571984 273816
rect 562652 273776 562658 273788
rect 571978 273776 571984 273788
rect 572036 273776 572042 273828
rect 597738 273816 597744 273828
rect 576826 273788 597744 273816
rect 563422 273680 563428 273692
rect 562428 273652 563428 273680
rect 563422 273640 563428 273652
rect 563480 273640 563486 273692
rect 563698 273640 563704 273692
rect 563756 273680 563762 273692
rect 576826 273680 576854 273788
rect 597738 273776 597744 273788
rect 597796 273776 597802 273828
rect 563756 273652 576854 273680
rect 563756 273640 563762 273652
rect 134426 273504 134432 273556
rect 134484 273544 134490 273556
rect 185118 273544 185124 273556
rect 134484 273516 185124 273544
rect 134484 273504 134490 273516
rect 185118 273504 185124 273516
rect 185176 273504 185182 273556
rect 446398 273504 446404 273556
rect 446456 273544 446462 273556
rect 475930 273544 475936 273556
rect 446456 273516 475936 273544
rect 446456 273504 446462 273516
rect 475930 273504 475936 273516
rect 475988 273504 475994 273556
rect 481358 273504 481364 273556
rect 481416 273544 481422 273556
rect 556338 273544 556344 273556
rect 481416 273516 556344 273544
rect 481416 273504 481422 273516
rect 556338 273504 556344 273516
rect 556396 273504 556402 273556
rect 556798 273504 556804 273556
rect 556856 273544 556862 273556
rect 590654 273544 590660 273556
rect 556856 273516 590660 273544
rect 556856 273504 556862 273516
rect 590654 273504 590660 273516
rect 590712 273504 590718 273556
rect 135622 273368 135628 273420
rect 135680 273408 135686 273420
rect 146938 273408 146944 273420
rect 135680 273380 146944 273408
rect 135680 273368 135686 273380
rect 146938 273368 146944 273380
rect 146996 273368 147002 273420
rect 460014 273368 460020 273420
rect 460072 273408 460078 273420
rect 465718 273408 465724 273420
rect 460072 273380 465724 273408
rect 460072 273368 460078 273380
rect 465718 273368 465724 273380
rect 465776 273368 465782 273420
rect 467558 273368 467564 273420
rect 467616 273408 467622 273420
rect 476114 273408 476120 273420
rect 467616 273380 476120 273408
rect 467616 273368 467622 273380
rect 476114 273368 476120 273380
rect 476172 273368 476178 273420
rect 478690 273368 478696 273420
rect 478748 273408 478754 273420
rect 552474 273408 552480 273420
rect 478748 273380 552480 273408
rect 478748 273368 478754 273380
rect 552474 273368 552480 273380
rect 552532 273368 552538 273420
rect 552658 273368 552664 273420
rect 552716 273408 552722 273420
rect 559926 273408 559932 273420
rect 552716 273380 559932 273408
rect 552716 273368 552722 273380
rect 559926 273368 559932 273380
rect 559984 273368 559990 273420
rect 374638 273300 374644 273352
rect 374696 273340 374702 273352
rect 377858 273340 377864 273352
rect 374696 273312 377864 273340
rect 374696 273300 374702 273312
rect 377858 273300 377864 273312
rect 377916 273300 377922 273352
rect 453298 273300 453304 273352
rect 453356 273340 453362 273352
rect 453758 273340 453764 273352
rect 453356 273312 453764 273340
rect 453356 273300 453362 273312
rect 453758 273300 453764 273312
rect 453816 273300 453822 273352
rect 318702 273232 318708 273284
rect 318760 273272 318766 273284
rect 324682 273272 324688 273284
rect 318760 273244 324688 273272
rect 318760 273232 318766 273244
rect 324682 273232 324688 273244
rect 324740 273232 324746 273284
rect 327534 273232 327540 273284
rect 327592 273272 327598 273284
rect 329466 273272 329472 273284
rect 327592 273244 329472 273272
rect 327592 273232 327598 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 114370 273164 114376 273216
rect 114428 273204 114434 273216
rect 171594 273204 171600 273216
rect 114428 273176 171600 273204
rect 114428 273164 114434 273176
rect 171594 273164 171600 273176
rect 171652 273164 171658 273216
rect 184106 273164 184112 273216
rect 184164 273204 184170 273216
rect 218882 273204 218888 273216
rect 184164 273176 218888 273204
rect 184164 273164 184170 273176
rect 218882 273164 218888 273176
rect 218940 273164 218946 273216
rect 366358 273164 366364 273216
rect 366416 273204 366422 273216
rect 383838 273204 383844 273216
rect 366416 273176 383844 273204
rect 366416 273164 366422 273176
rect 383838 273164 383844 273176
rect 383896 273164 383902 273216
rect 401502 273164 401508 273216
rect 401560 273204 401566 273216
rect 442902 273204 442908 273216
rect 401560 273176 442908 273204
rect 401560 273164 401566 273176
rect 442902 273164 442908 273176
rect 442960 273164 442966 273216
rect 452286 273164 452292 273216
rect 452344 273204 452350 273216
rect 515030 273204 515036 273216
rect 452344 273176 515036 273204
rect 452344 273164 452350 273176
rect 515030 273164 515036 273176
rect 515088 273164 515094 273216
rect 515214 273164 515220 273216
rect 515272 273204 515278 273216
rect 519722 273204 519728 273216
rect 515272 273176 519728 273204
rect 515272 273164 515278 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 278590 273096 278596 273148
rect 278648 273136 278654 273148
rect 285858 273136 285864 273148
rect 278648 273108 285864 273136
rect 278648 273096 278654 273108
rect 285858 273096 285864 273108
rect 285916 273096 285922 273148
rect 101306 273028 101312 273080
rect 101364 273068 101370 273080
rect 160186 273068 160192 273080
rect 101364 273040 160192 273068
rect 101364 273028 101370 273040
rect 160186 273028 160192 273040
rect 160244 273028 160250 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 210602 273068 210608 273080
rect 172296 273040 210608 273068
rect 172296 273028 172302 273040
rect 210602 273028 210608 273040
rect 210660 273028 210666 273080
rect 224034 273028 224040 273080
rect 224092 273068 224098 273080
rect 243262 273068 243268 273080
rect 224092 273040 243268 273068
rect 224092 273028 224098 273040
rect 243262 273028 243268 273040
rect 243320 273028 243326 273080
rect 329466 273028 329472 273080
rect 329524 273068 329530 273080
rect 338850 273068 338856 273080
rect 329524 273040 338856 273068
rect 329524 273028 329530 273040
rect 338850 273028 338856 273040
rect 338908 273028 338914 273080
rect 349798 273028 349804 273080
rect 349856 273068 349862 273080
rect 366082 273068 366088 273080
rect 349856 273040 366088 273068
rect 349856 273028 349862 273040
rect 366082 273028 366088 273040
rect 366140 273028 366146 273080
rect 377398 273028 377404 273080
rect 377456 273068 377462 273080
rect 399202 273068 399208 273080
rect 377456 273040 399208 273068
rect 377456 273028 377462 273040
rect 399202 273028 399208 273040
rect 399260 273028 399266 273080
rect 408218 273028 408224 273080
rect 408276 273068 408282 273080
rect 450814 273068 450820 273080
rect 408276 273040 450820 273068
rect 408276 273028 408282 273040
rect 450814 273028 450820 273040
rect 450872 273028 450878 273080
rect 451182 273028 451188 273080
rect 451240 273068 451246 273080
rect 513834 273068 513840 273080
rect 451240 273040 513840 273068
rect 451240 273028 451246 273040
rect 513834 273028 513840 273040
rect 513892 273028 513898 273080
rect 526806 273028 526812 273080
rect 526864 273068 526870 273080
rect 621382 273068 621388 273080
rect 526864 273040 621388 273068
rect 526864 273028 526870 273040
rect 621382 273028 621388 273040
rect 621440 273028 621446 273080
rect 99006 272892 99012 272944
rect 99064 272932 99070 272944
rect 160370 272932 160376 272944
rect 99064 272904 160376 272932
rect 99064 272892 99070 272904
rect 160370 272892 160376 272904
rect 160428 272892 160434 272944
rect 162762 272892 162768 272944
rect 162820 272932 162826 272944
rect 204714 272932 204720 272944
rect 162820 272904 204720 272932
rect 162820 272892 162826 272904
rect 204714 272892 204720 272904
rect 204772 272892 204778 272944
rect 219526 272892 219532 272944
rect 219584 272932 219590 272944
rect 244458 272932 244464 272944
rect 219584 272904 244464 272932
rect 219584 272892 219590 272904
rect 244458 272892 244464 272904
rect 244516 272892 244522 272944
rect 251450 272892 251456 272944
rect 251508 272932 251514 272944
rect 266998 272932 267004 272944
rect 251508 272904 267004 272932
rect 251508 272892 251514 272904
rect 266998 272892 267004 272904
rect 267056 272892 267062 272944
rect 335262 272892 335268 272944
rect 335320 272932 335326 272944
rect 346854 272932 346860 272944
rect 335320 272904 346860 272932
rect 335320 272892 335326 272904
rect 346854 272892 346860 272904
rect 346912 272892 346918 272944
rect 362770 272892 362776 272944
rect 362828 272932 362834 272944
rect 385862 272932 385868 272944
rect 362828 272904 385868 272932
rect 362828 272892 362834 272904
rect 385862 272892 385868 272904
rect 385920 272892 385926 272944
rect 406838 272892 406844 272944
rect 406896 272932 406902 272944
rect 449986 272932 449992 272944
rect 406896 272904 449992 272932
rect 406896 272892 406902 272904
rect 449986 272892 449992 272904
rect 450044 272892 450050 272944
rect 455230 272892 455236 272944
rect 455288 272932 455294 272944
rect 455288 272904 457300 272932
rect 455288 272892 455294 272904
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 158070 272756 158076 272808
rect 158128 272796 158134 272808
rect 200666 272796 200672 272808
rect 158128 272768 200672 272796
rect 158128 272756 158134 272768
rect 200666 272756 200672 272768
rect 200724 272756 200730 272808
rect 208854 272756 208860 272808
rect 208912 272796 208918 272808
rect 237374 272796 237380 272808
rect 208912 272768 237380 272796
rect 208912 272756 208918 272768
rect 237374 272756 237380 272768
rect 237432 272756 237438 272808
rect 252646 272756 252652 272808
rect 252704 272796 252710 272808
rect 252704 272768 262260 272796
rect 252704 272756 252710 272768
rect 72970 272620 72976 272672
rect 73028 272660 73034 272672
rect 142154 272660 142160 272672
rect 73028 272632 142160 272660
rect 73028 272620 73034 272632
rect 142154 272620 142160 272632
rect 142212 272620 142218 272672
rect 152182 272620 152188 272672
rect 152240 272660 152246 272672
rect 197538 272660 197544 272672
rect 152240 272632 197544 272660
rect 152240 272620 152246 272632
rect 197538 272620 197544 272632
rect 197596 272620 197602 272672
rect 199470 272620 199476 272672
rect 199528 272660 199534 272672
rect 230566 272660 230572 272672
rect 199528 272632 230572 272660
rect 199528 272620 199534 272632
rect 230566 272620 230572 272632
rect 230624 272620 230630 272672
rect 233694 272620 233700 272672
rect 233752 272660 233758 272672
rect 253934 272660 253940 272672
rect 233752 272632 253940 272660
rect 233752 272620 233758 272632
rect 253934 272620 253940 272632
rect 253992 272620 253998 272672
rect 69382 272484 69388 272536
rect 69440 272524 69446 272536
rect 139394 272524 139400 272536
rect 69440 272496 139400 272524
rect 69440 272484 69446 272496
rect 139394 272484 139400 272496
rect 139452 272484 139458 272536
rect 141510 272484 141516 272536
rect 141568 272524 141574 272536
rect 141568 272496 180794 272524
rect 141568 272484 141574 272496
rect 120258 272348 120264 272400
rect 120316 272388 120322 272400
rect 175274 272388 175280 272400
rect 120316 272360 175280 272388
rect 120316 272348 120322 272360
rect 175274 272348 175280 272360
rect 175332 272348 175338 272400
rect 180766 272388 180794 272496
rect 189074 272484 189080 272536
rect 189132 272524 189138 272536
rect 194042 272524 194048 272536
rect 189132 272496 194048 272524
rect 189132 272484 189138 272496
rect 194042 272484 194048 272496
rect 194100 272484 194106 272536
rect 194686 272484 194692 272536
rect 194744 272524 194750 272536
rect 227162 272524 227168 272536
rect 194744 272496 227168 272524
rect 194744 272484 194750 272496
rect 227162 272484 227168 272496
rect 227220 272484 227226 272536
rect 238478 272484 238484 272536
rect 238536 272524 238542 272536
rect 258074 272524 258080 272536
rect 238536 272496 258080 272524
rect 238536 272484 238542 272496
rect 258074 272484 258080 272496
rect 258132 272484 258138 272536
rect 262232 272524 262260 272768
rect 271506 272756 271512 272808
rect 271564 272796 271570 272808
rect 280338 272796 280344 272808
rect 271564 272768 280344 272796
rect 271564 272756 271570 272768
rect 280338 272756 280344 272768
rect 280396 272756 280402 272808
rect 336366 272756 336372 272808
rect 336424 272796 336430 272808
rect 349522 272796 349528 272808
rect 336424 272768 349528 272796
rect 336424 272756 336430 272768
rect 349522 272756 349528 272768
rect 349580 272756 349586 272808
rect 352558 272756 352564 272808
rect 352616 272796 352622 272808
rect 370774 272796 370780 272808
rect 352616 272768 370780 272796
rect 352616 272756 352622 272768
rect 370774 272756 370780 272768
rect 370832 272756 370838 272808
rect 375190 272756 375196 272808
rect 375248 272796 375254 272808
rect 403894 272796 403900 272808
rect 375248 272768 403900 272796
rect 375248 272756 375254 272768
rect 403894 272756 403900 272768
rect 403952 272756 403958 272808
rect 412266 272756 412272 272808
rect 412324 272796 412330 272808
rect 457070 272796 457076 272808
rect 412324 272768 457076 272796
rect 412324 272756 412330 272768
rect 457070 272756 457076 272768
rect 457128 272756 457134 272808
rect 457272 272796 457300 272904
rect 458082 272892 458088 272944
rect 458140 272932 458146 272944
rect 463326 272932 463332 272944
rect 458140 272904 463332 272932
rect 458140 272892 458146 272904
rect 463326 272892 463332 272904
rect 463384 272892 463390 272944
rect 518526 272932 518532 272944
rect 463712 272904 518532 272932
rect 463712 272796 463740 272904
rect 518526 272892 518532 272904
rect 518584 272892 518590 272944
rect 529842 272892 529848 272944
rect 529900 272932 529906 272944
rect 624970 272932 624976 272944
rect 529900 272904 624976 272932
rect 529900 272892 529906 272904
rect 624970 272892 624976 272904
rect 625028 272892 625034 272944
rect 457272 272768 463740 272796
rect 463878 272756 463884 272808
rect 463936 272796 463942 272808
rect 522114 272796 522120 272808
rect 463936 272768 522120 272796
rect 463936 272756 463942 272768
rect 522114 272756 522120 272768
rect 522172 272756 522178 272808
rect 522758 272756 522764 272808
rect 522816 272796 522822 272808
rect 524138 272796 524144 272808
rect 522816 272768 524144 272796
rect 522816 272756 522822 272768
rect 524138 272756 524144 272768
rect 524196 272756 524202 272808
rect 532510 272756 532516 272808
rect 532568 272796 532574 272808
rect 628466 272796 628472 272808
rect 532568 272768 628472 272796
rect 532568 272756 532574 272768
rect 628466 272756 628472 272768
rect 628524 272756 628530 272808
rect 266814 272620 266820 272672
rect 266872 272660 266878 272672
rect 277578 272660 277584 272672
rect 266872 272632 277584 272660
rect 266872 272620 266878 272632
rect 277578 272620 277584 272632
rect 277636 272620 277642 272672
rect 280982 272620 280988 272672
rect 281040 272660 281046 272672
rect 286318 272660 286324 272672
rect 281040 272632 286324 272660
rect 281040 272620 281046 272632
rect 286318 272620 286324 272632
rect 286376 272620 286382 272672
rect 322750 272620 322756 272672
rect 322808 272660 322814 272672
rect 330570 272660 330576 272672
rect 322808 272632 330576 272660
rect 322808 272620 322814 272632
rect 330570 272620 330576 272632
rect 330628 272620 330634 272672
rect 338022 272620 338028 272672
rect 338080 272660 338086 272672
rect 351914 272660 351920 272672
rect 338080 272632 351920 272660
rect 338080 272620 338086 272632
rect 351914 272620 351920 272632
rect 351972 272620 351978 272672
rect 354490 272620 354496 272672
rect 354548 272660 354554 272672
rect 375558 272660 375564 272672
rect 354548 272632 375564 272660
rect 354548 272620 354554 272632
rect 375558 272620 375564 272632
rect 375616 272620 375622 272672
rect 381998 272620 382004 272672
rect 382056 272660 382062 272672
rect 414566 272660 414572 272672
rect 382056 272632 414572 272660
rect 382056 272620 382062 272632
rect 414566 272620 414572 272632
rect 414624 272620 414630 272672
rect 419166 272620 419172 272672
rect 419224 272660 419230 272672
rect 467374 272660 467380 272672
rect 419224 272632 467380 272660
rect 419224 272620 419230 272632
rect 467374 272620 467380 272632
rect 467432 272620 467438 272672
rect 467742 272620 467748 272672
rect 467800 272660 467806 272672
rect 470410 272660 470416 272672
rect 467800 272632 470416 272660
rect 467800 272620 467806 272632
rect 470410 272620 470416 272632
rect 470468 272620 470474 272672
rect 470594 272620 470600 272672
rect 470652 272660 470658 272672
rect 536282 272660 536288 272672
rect 470652 272632 536288 272660
rect 470652 272620 470658 272632
rect 536282 272620 536288 272632
rect 536340 272620 536346 272672
rect 536558 272620 536564 272672
rect 536616 272660 536622 272672
rect 635550 272660 635556 272672
rect 536616 272632 635556 272660
rect 536616 272620 536622 272632
rect 635550 272620 635556 272632
rect 635608 272620 635614 272672
rect 267918 272524 267924 272536
rect 262232 272496 267924 272524
rect 267918 272484 267924 272496
rect 267976 272484 267982 272536
rect 325510 272484 325516 272536
rect 325568 272524 325574 272536
rect 334158 272524 334164 272536
rect 325568 272496 334164 272524
rect 325568 272484 325574 272496
rect 334158 272484 334164 272496
rect 334216 272484 334222 272536
rect 344646 272484 344652 272536
rect 344704 272524 344710 272536
rect 361390 272524 361396 272536
rect 344704 272496 361396 272524
rect 344704 272484 344710 272496
rect 361390 272484 361396 272496
rect 361448 272484 361454 272536
rect 363782 272484 363788 272536
rect 363840 272524 363846 272536
rect 388530 272524 388536 272536
rect 363840 272496 388536 272524
rect 363840 272484 363846 272496
rect 388530 272484 388536 272496
rect 388588 272484 388594 272536
rect 397270 272484 397276 272536
rect 397328 272524 397334 272536
rect 435818 272524 435824 272536
rect 397328 272496 435824 272524
rect 397328 272484 397334 272496
rect 435818 272484 435824 272496
rect 435876 272484 435882 272536
rect 438762 272484 438768 272536
rect 438820 272524 438826 272536
rect 489868 272524 489874 272536
rect 438820 272496 489874 272524
rect 438820 272484 438826 272496
rect 489868 272484 489874 272496
rect 489926 272484 489932 272536
rect 490006 272484 490012 272536
rect 490064 272524 490070 272536
rect 529198 272524 529204 272536
rect 490064 272496 529204 272524
rect 490064 272484 490070 272496
rect 529198 272484 529204 272496
rect 529256 272484 529262 272536
rect 533706 272484 533712 272536
rect 533764 272524 533770 272536
rect 632054 272524 632060 272536
rect 533764 272496 632060 272524
rect 533764 272484 533770 272496
rect 632054 272484 632060 272496
rect 632112 272484 632118 272536
rect 189166 272388 189172 272400
rect 180766 272360 189172 272388
rect 189166 272348 189172 272360
rect 189224 272348 189230 272400
rect 193582 272348 193588 272400
rect 193640 272388 193646 272400
rect 224218 272388 224224 272400
rect 193640 272360 224224 272388
rect 193640 272348 193646 272360
rect 224218 272348 224224 272360
rect 224276 272348 224282 272400
rect 264422 272348 264428 272400
rect 264480 272388 264486 272400
rect 276014 272388 276020 272400
rect 264480 272360 276020 272388
rect 264480 272348 264486 272360
rect 276014 272348 276020 272360
rect 276072 272348 276078 272400
rect 388990 272348 388996 272400
rect 389048 272388 389054 272400
rect 425146 272388 425152 272400
rect 389048 272360 425152 272388
rect 389048 272348 389054 272360
rect 425146 272348 425152 272360
rect 425204 272348 425210 272400
rect 449710 272348 449716 272400
rect 449768 272388 449774 272400
rect 511442 272388 511448 272400
rect 449768 272360 511448 272388
rect 449768 272348 449774 272360
rect 511442 272348 511448 272360
rect 511500 272348 511506 272400
rect 512638 272348 512644 272400
rect 512696 272388 512702 272400
rect 515214 272388 515220 272400
rect 512696 272360 515220 272388
rect 512696 272348 512702 272360
rect 515214 272348 515220 272360
rect 515272 272348 515278 272400
rect 517330 272348 517336 272400
rect 517388 272388 517394 272400
rect 607214 272388 607220 272400
rect 517388 272360 607220 272388
rect 517388 272348 517394 272360
rect 607214 272348 607220 272360
rect 607272 272348 607278 272400
rect 119062 272212 119068 272264
rect 119120 272252 119126 272264
rect 173250 272252 173256 272264
rect 119120 272224 173256 272252
rect 119120 272212 119126 272224
rect 173250 272212 173256 272224
rect 173308 272212 173314 272264
rect 174446 272212 174452 272264
rect 174504 272252 174510 272264
rect 189350 272252 189356 272264
rect 174504 272224 189356 272252
rect 174504 272212 174510 272224
rect 189350 272212 189356 272224
rect 189408 272212 189414 272264
rect 446950 272212 446956 272264
rect 447008 272252 447014 272264
rect 508038 272252 508044 272264
rect 447008 272224 508044 272252
rect 447008 272212 447014 272224
rect 508038 272212 508044 272224
rect 508096 272212 508102 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 130838 272076 130844 272128
rect 130896 272116 130902 272128
rect 182450 272116 182456 272128
rect 130896 272088 182456 272116
rect 130896 272076 130902 272088
rect 182450 272076 182456 272088
rect 182508 272076 182514 272128
rect 426342 272076 426348 272128
rect 426400 272116 426406 272128
rect 470548 272116 470554 272128
rect 426400 272088 470554 272116
rect 426400 272076 426406 272088
rect 470548 272076 470554 272088
rect 470606 272076 470612 272128
rect 470778 272076 470784 272128
rect 470836 272116 470842 272128
rect 489868 272116 489874 272128
rect 470836 272088 489874 272116
rect 470836 272076 470842 272088
rect 489868 272076 489874 272088
rect 489926 272076 489932 272128
rect 490006 272076 490012 272128
rect 490064 272116 490070 272128
rect 558730 272116 558736 272128
rect 490064 272088 558736 272116
rect 490064 272076 490070 272088
rect 558730 272076 558736 272088
rect 558788 272076 558794 272128
rect 191466 271940 191472 271992
rect 191524 271980 191530 271992
rect 191524 271952 192800 271980
rect 191524 271940 191530 271952
rect 108390 271804 108396 271856
rect 108448 271844 108454 271856
rect 165890 271844 165896 271856
rect 108448 271816 165896 271844
rect 108448 271804 108454 271816
rect 165890 271804 165896 271816
rect 165948 271804 165954 271856
rect 188798 271804 188804 271856
rect 188856 271844 188862 271856
rect 192570 271844 192576 271856
rect 188856 271816 192576 271844
rect 188856 271804 188862 271816
rect 192570 271804 192576 271816
rect 192628 271804 192634 271856
rect 192772 271844 192800 271952
rect 447778 271940 447784 271992
rect 447836 271980 447842 271992
rect 506750 271980 506756 271992
rect 447836 271952 506756 271980
rect 447836 271940 447842 271952
rect 506750 271940 506756 271952
rect 506808 271940 506814 271992
rect 507118 271940 507124 271992
rect 507176 271980 507182 271992
rect 569402 271980 569408 271992
rect 507176 271952 569408 271980
rect 507176 271940 507182 271952
rect 569402 271940 569408 271952
rect 569460 271940 569466 271992
rect 268654 271872 268660 271924
rect 268712 271912 268718 271924
rect 270494 271912 270500 271924
rect 268712 271884 270500 271912
rect 268712 271872 268718 271884
rect 270494 271872 270500 271884
rect 270552 271872 270558 271924
rect 225046 271844 225052 271856
rect 192772 271816 225052 271844
rect 225046 271804 225052 271816
rect 225104 271804 225110 271856
rect 225414 271804 225420 271856
rect 225472 271844 225478 271856
rect 228358 271844 228364 271856
rect 225472 271816 228364 271844
rect 225472 271804 225478 271816
rect 228358 271804 228364 271816
rect 228416 271804 228422 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 376570 271804 376576 271856
rect 376628 271844 376634 271856
rect 407482 271844 407488 271856
rect 376628 271816 407488 271844
rect 376628 271804 376634 271816
rect 407482 271804 407488 271816
rect 407540 271804 407546 271856
rect 407758 271804 407764 271856
rect 407816 271844 407822 271856
rect 437014 271844 437020 271856
rect 407816 271816 437020 271844
rect 407816 271804 407822 271816
rect 437014 271804 437020 271816
rect 437072 271804 437078 271856
rect 437198 271804 437204 271856
rect 437256 271844 437262 271856
rect 493686 271844 493692 271856
rect 437256 271816 493692 271844
rect 437256 271804 437262 271816
rect 493686 271804 493692 271816
rect 493744 271804 493750 271856
rect 496538 271804 496544 271856
rect 496596 271844 496602 271856
rect 578510 271844 578516 271856
rect 496596 271816 578516 271844
rect 496596 271804 496602 271816
rect 578510 271804 578516 271816
rect 578568 271804 578574 271856
rect 578878 271804 578884 271856
rect 578936 271844 578942 271856
rect 611906 271844 611912 271856
rect 578936 271816 611912 271844
rect 578936 271804 578942 271816
rect 611906 271804 611912 271816
rect 611964 271804 611970 271856
rect 106090 271668 106096 271720
rect 106148 271708 106154 271720
rect 164970 271708 164976 271720
rect 106148 271680 164976 271708
rect 106148 271668 106154 271680
rect 164970 271668 164976 271680
rect 165028 271668 165034 271720
rect 175734 271668 175740 271720
rect 175792 271708 175798 271720
rect 212994 271708 213000 271720
rect 175792 271680 213000 271708
rect 175792 271668 175798 271680
rect 212994 271668 213000 271680
rect 213052 271668 213058 271720
rect 239858 271668 239864 271720
rect 239916 271708 239922 271720
rect 254118 271708 254124 271720
rect 239916 271680 254124 271708
rect 239916 271668 239922 271680
rect 254118 271668 254124 271680
rect 254176 271668 254182 271720
rect 353938 271668 353944 271720
rect 353996 271708 354002 271720
rect 372798 271708 372804 271720
rect 353996 271680 372804 271708
rect 353996 271668 354002 271680
rect 372798 271668 372804 271680
rect 372856 271668 372862 271720
rect 384942 271668 384948 271720
rect 385000 271708 385006 271720
rect 418062 271708 418068 271720
rect 385000 271680 418068 271708
rect 385000 271668 385006 271680
rect 418062 271668 418068 271680
rect 418120 271668 418126 271720
rect 420178 271668 420184 271720
rect 420236 271708 420242 271720
rect 431126 271708 431132 271720
rect 420236 271680 431132 271708
rect 420236 271668 420242 271680
rect 431126 271668 431132 271680
rect 431184 271668 431190 271720
rect 434622 271668 434628 271720
rect 434680 271708 434686 271720
rect 485222 271708 485228 271720
rect 434680 271680 485228 271708
rect 434680 271668 434686 271680
rect 485222 271668 485228 271680
rect 485280 271668 485286 271720
rect 485406 271668 485412 271720
rect 485464 271708 485470 271720
rect 490006 271708 490012 271720
rect 485464 271680 490012 271708
rect 485464 271668 485470 271680
rect 490006 271668 490012 271680
rect 490064 271668 490070 271720
rect 501966 271668 501972 271720
rect 502024 271708 502030 271720
rect 585962 271708 585968 271720
rect 502024 271680 585968 271708
rect 502024 271668 502030 271680
rect 585962 271668 585968 271680
rect 586020 271668 586026 271720
rect 94222 271532 94228 271584
rect 94280 271572 94286 271584
rect 156138 271572 156144 271584
rect 94280 271544 156144 271572
rect 94280 271532 94286 271544
rect 156138 271532 156144 271544
rect 156196 271532 156202 271584
rect 170122 271532 170128 271584
rect 170180 271572 170186 271584
rect 209774 271572 209780 271584
rect 170180 271544 209780 271572
rect 170180 271532 170186 271544
rect 209774 271532 209780 271544
rect 209832 271532 209838 271584
rect 223114 271532 223120 271584
rect 223172 271572 223178 271584
rect 247218 271572 247224 271584
rect 223172 271544 247224 271572
rect 223172 271532 223178 271544
rect 247218 271532 247224 271544
rect 247276 271532 247282 271584
rect 357158 271532 357164 271584
rect 357216 271572 357222 271584
rect 379054 271572 379060 271584
rect 357216 271544 379060 271572
rect 357216 271532 357222 271544
rect 379054 271532 379060 271544
rect 379112 271532 379118 271584
rect 387610 271532 387616 271584
rect 387668 271572 387674 271584
rect 422846 271572 422852 271584
rect 387668 271544 422852 271572
rect 387668 271532 387674 271544
rect 422846 271532 422852 271544
rect 422904 271532 422910 271584
rect 439958 271532 439964 271584
rect 440016 271572 440022 271584
rect 497274 271572 497280 271584
rect 440016 271544 497280 271572
rect 440016 271532 440022 271544
rect 497274 271532 497280 271544
rect 497332 271532 497338 271584
rect 499298 271532 499304 271584
rect 499356 271572 499362 271584
rect 582374 271572 582380 271584
rect 499356 271544 582380 271572
rect 499356 271532 499362 271544
rect 582374 271532 582380 271544
rect 582432 271532 582438 271584
rect 585778 271532 585784 271584
rect 585836 271572 585842 271584
rect 626074 271572 626080 271584
rect 585836 271544 626080 271572
rect 585836 271532 585842 271544
rect 626074 271532 626080 271544
rect 626132 271532 626138 271584
rect 87138 271396 87144 271448
rect 87196 271436 87202 271448
rect 152182 271436 152188 271448
rect 87196 271408 152188 271436
rect 87196 271396 87202 271408
rect 152182 271396 152188 271408
rect 152240 271396 152246 271448
rect 159266 271396 159272 271448
rect 159324 271436 159330 271448
rect 202322 271436 202328 271448
rect 159324 271408 202328 271436
rect 159324 271396 159330 271408
rect 202322 271396 202328 271408
rect 202380 271396 202386 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 250254 271396 250260 271448
rect 250312 271436 250318 271448
rect 250312 271408 262444 271436
rect 250312 271396 250318 271408
rect 75362 271260 75368 271312
rect 75420 271300 75426 271312
rect 75420 271272 142154 271300
rect 75420 271260 75426 271272
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 142126 271164 142154 271272
rect 142706 271260 142712 271312
rect 142764 271300 142770 271312
rect 144178 271300 144184 271312
rect 142764 271272 144184 271300
rect 142764 271260 142770 271272
rect 144178 271260 144184 271272
rect 144236 271260 144242 271312
rect 154298 271260 154304 271312
rect 154356 271300 154362 271312
rect 198090 271300 198096 271312
rect 154356 271272 198096 271300
rect 154356 271260 154362 271272
rect 198090 271260 198096 271272
rect 198148 271260 198154 271312
rect 212258 271260 212264 271312
rect 212316 271300 212322 271312
rect 239306 271300 239312 271312
rect 212316 271272 239312 271300
rect 212316 271260 212322 271272
rect 239306 271260 239312 271272
rect 239364 271260 239370 271312
rect 244642 271260 244648 271312
rect 244700 271300 244706 271312
rect 262214 271300 262220 271312
rect 244700 271272 262220 271300
rect 244700 271260 244706 271272
rect 262214 271260 262220 271272
rect 262272 271260 262278 271312
rect 262416 271300 262444 271408
rect 265618 271396 265624 271448
rect 265676 271436 265682 271448
rect 276842 271436 276848 271448
rect 265676 271408 276848 271436
rect 265676 271396 265682 271408
rect 276842 271396 276848 271408
rect 276900 271396 276906 271448
rect 329650 271396 329656 271448
rect 329708 271436 329714 271448
rect 340046 271436 340052 271448
rect 329708 271408 340052 271436
rect 329708 271396 329714 271408
rect 340046 271396 340052 271408
rect 340104 271396 340110 271448
rect 340598 271396 340604 271448
rect 340656 271436 340662 271448
rect 355134 271436 355140 271448
rect 340656 271408 355140 271436
rect 340656 271396 340662 271408
rect 355134 271396 355140 271408
rect 355192 271396 355198 271448
rect 358722 271396 358728 271448
rect 358780 271436 358786 271448
rect 381446 271436 381452 271448
rect 358780 271408 381452 271436
rect 358780 271396 358786 271408
rect 381446 271396 381452 271408
rect 381504 271396 381510 271448
rect 393958 271396 393964 271448
rect 394016 271436 394022 271448
rect 429930 271436 429936 271448
rect 394016 271408 429936 271436
rect 394016 271396 394022 271408
rect 429930 271396 429936 271408
rect 429988 271396 429994 271448
rect 442902 271396 442908 271448
rect 442960 271436 442966 271448
rect 500862 271436 500868 271448
rect 442960 271408 500868 271436
rect 442960 271396 442966 271408
rect 500862 271396 500868 271408
rect 500920 271396 500926 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 266446 271300 266452 271312
rect 262416 271272 266452 271300
rect 266446 271260 266452 271272
rect 266504 271260 266510 271312
rect 276658 271260 276664 271312
rect 276716 271300 276722 271312
rect 284478 271300 284484 271312
rect 276716 271272 284484 271300
rect 276716 271260 276722 271272
rect 284478 271260 284484 271272
rect 284536 271260 284542 271312
rect 326430 271260 326436 271312
rect 326488 271300 326494 271312
rect 335078 271300 335084 271312
rect 326488 271272 335084 271300
rect 326488 271260 326494 271272
rect 335078 271260 335084 271272
rect 335136 271260 335142 271312
rect 339402 271260 339408 271312
rect 339460 271300 339466 271312
rect 354214 271300 354220 271312
rect 339460 271272 354220 271300
rect 339460 271260 339466 271272
rect 354214 271260 354220 271272
rect 354272 271260 354278 271312
rect 365438 271260 365444 271312
rect 365496 271300 365502 271312
rect 390922 271300 390928 271312
rect 365496 271272 390928 271300
rect 365496 271260 365502 271272
rect 390922 271260 390928 271272
rect 390980 271260 390986 271312
rect 391842 271260 391848 271312
rect 391900 271300 391906 271312
rect 428734 271300 428740 271312
rect 391900 271272 428740 271300
rect 391900 271260 391906 271272
rect 428734 271260 428740 271272
rect 428792 271260 428798 271312
rect 445662 271260 445668 271312
rect 445720 271300 445726 271312
rect 504358 271300 504364 271312
rect 445720 271272 504364 271300
rect 445720 271260 445726 271272
rect 504358 271260 504364 271272
rect 504416 271260 504422 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 611998 271260 612004 271312
rect 612056 271300 612062 271312
rect 618622 271300 618628 271312
rect 612056 271272 618628 271300
rect 612056 271260 612062 271272
rect 618622 271260 618628 271272
rect 618680 271260 618686 271312
rect 618898 271260 618904 271312
rect 618956 271300 618962 271312
rect 633250 271300 633256 271312
rect 618956 271272 633256 271300
rect 618956 271260 618962 271272
rect 633250 271260 633256 271272
rect 633308 271260 633314 271312
rect 142706 271164 142712 271176
rect 142126 271136 142712 271164
rect 142706 271124 142712 271136
rect 142764 271124 142770 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 197078 271124 197084 271176
rect 197136 271164 197142 271176
rect 229278 271164 229284 271176
rect 197136 271136 229284 271164
rect 197136 271124 197142 271136
rect 229278 271124 229284 271136
rect 229336 271124 229342 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 251726 271164 251732 271176
rect 230256 271136 251732 271164
rect 230256 271124 230262 271136
rect 251726 271124 251732 271136
rect 251784 271124 251790 271176
rect 254946 271124 254952 271176
rect 255004 271164 255010 271176
rect 269298 271164 269304 271176
rect 255004 271136 269304 271164
rect 255004 271124 255010 271136
rect 269298 271124 269304 271136
rect 269356 271124 269362 271176
rect 270310 271124 270316 271176
rect 270368 271164 270374 271176
rect 280522 271164 280528 271176
rect 270368 271136 280528 271164
rect 270368 271124 270374 271136
rect 280522 271124 280528 271136
rect 280580 271124 280586 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 347590 271124 347596 271176
rect 347648 271164 347654 271176
rect 364518 271164 364524 271176
rect 347648 271136 364524 271164
rect 347648 271124 347654 271136
rect 364518 271124 364524 271136
rect 364576 271124 364582 271176
rect 366910 271124 366916 271176
rect 366968 271164 366974 271176
rect 393314 271164 393320 271176
rect 366968 271136 393320 271164
rect 366968 271124 366974 271136
rect 393314 271124 393320 271136
rect 393372 271124 393378 271176
rect 402606 271124 402612 271176
rect 402664 271164 402670 271176
rect 444098 271164 444104 271176
rect 402664 271136 444104 271164
rect 402664 271124 402670 271136
rect 444098 271124 444104 271136
rect 444156 271124 444162 271176
rect 459462 271124 459468 271176
rect 459520 271164 459526 271176
rect 523862 271164 523868 271176
rect 459520 271136 523868 271164
rect 459520 271124 459526 271136
rect 523862 271124 523868 271136
rect 523920 271124 523926 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617794 271164 617800 271176
rect 524104 271136 617800 271164
rect 524104 271124 524110 271136
rect 617794 271124 617800 271136
rect 617852 271124 617858 271176
rect 625798 271124 625804 271176
rect 625856 271164 625862 271176
rect 645026 271164 645032 271176
rect 625856 271136 645032 271164
rect 625856 271124 625862 271136
rect 645026 271124 645032 271136
rect 645084 271124 645090 271176
rect 116670 270988 116676 271040
rect 116728 271028 116734 271040
rect 172514 271028 172520 271040
rect 116728 271000 172520 271028
rect 116728 270988 116734 271000
rect 172514 270988 172520 271000
rect 172572 270988 172578 271040
rect 192754 270988 192760 271040
rect 192812 271028 192818 271040
rect 225506 271028 225512 271040
rect 192812 271000 225512 271028
rect 192812 270988 192818 271000
rect 225506 270988 225512 271000
rect 225564 270988 225570 271040
rect 381538 270988 381544 271040
rect 381596 271028 381602 271040
rect 411806 271028 411812 271040
rect 381596 271000 411812 271028
rect 381596 270988 381602 271000
rect 411806 270988 411812 271000
rect 411864 270988 411870 271040
rect 414474 270988 414480 271040
rect 414532 271028 414538 271040
rect 438118 271028 438124 271040
rect 414532 271000 438124 271028
rect 414532 270988 414538 271000
rect 438118 270988 438124 271000
rect 438176 270988 438182 271040
rect 438302 270988 438308 271040
rect 438360 271028 438366 271040
rect 438360 271000 485084 271028
rect 438360 270988 438366 271000
rect 124950 270852 124956 270904
rect 125008 270892 125014 270904
rect 178678 270892 178684 270904
rect 125008 270864 178684 270892
rect 125008 270852 125014 270864
rect 178678 270852 178684 270864
rect 178736 270852 178742 270904
rect 417418 270852 417424 270904
rect 417476 270892 417482 270904
rect 427538 270892 427544 270904
rect 417476 270864 427544 270892
rect 417476 270852 417482 270864
rect 427538 270852 427544 270864
rect 427596 270852 427602 270904
rect 430390 270852 430396 270904
rect 430448 270892 430454 270904
rect 483106 270892 483112 270904
rect 430448 270864 483112 270892
rect 430448 270852 430454 270864
rect 483106 270852 483112 270864
rect 483164 270852 483170 270904
rect 485056 270892 485084 271000
rect 485222 270988 485228 271040
rect 485280 271028 485286 271040
rect 490190 271028 490196 271040
rect 485280 271000 490196 271028
rect 485280 270988 485286 271000
rect 490190 270988 490196 271000
rect 490248 270988 490254 271040
rect 495250 270988 495256 271040
rect 495308 271028 495314 271040
rect 575290 271028 575296 271040
rect 495308 271000 575296 271028
rect 495308 270988 495314 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 492398 270892 492404 270904
rect 485056 270864 492404 270892
rect 492398 270852 492404 270864
rect 492456 270852 492462 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571702 270892 571708 270904
rect 492640 270864 571708 270892
rect 492640 270852 492646 270864
rect 571702 270852 571708 270864
rect 571760 270852 571766 270904
rect 571978 270852 571984 270904
rect 572036 270892 572042 270904
rect 604822 270892 604828 270904
rect 572036 270864 604828 270892
rect 572036 270852 572042 270864
rect 604822 270852 604828 270864
rect 604880 270852 604886 270904
rect 127342 270716 127348 270768
rect 127400 270756 127406 270768
rect 179874 270756 179880 270768
rect 127400 270728 179880 270756
rect 127400 270716 127406 270728
rect 179874 270716 179880 270728
rect 179932 270716 179938 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 427446 270716 427452 270768
rect 427504 270756 427510 270768
rect 479150 270756 479156 270768
rect 427504 270728 479156 270756
rect 427504 270716 427510 270728
rect 479150 270716 479156 270728
rect 479208 270716 479214 270768
rect 486878 270716 486884 270768
rect 486936 270756 486942 270768
rect 564618 270756 564624 270768
rect 486936 270728 564624 270756
rect 486936 270716 486942 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 137922 270580 137928 270632
rect 137980 270620 137986 270632
rect 187694 270620 187700 270632
rect 137980 270592 187700 270620
rect 137980 270580 137986 270592
rect 187694 270580 187700 270592
rect 187752 270580 187758 270632
rect 422938 270580 422944 270632
rect 422996 270620 423002 270632
rect 445294 270620 445300 270632
rect 422996 270592 445300 270620
rect 422996 270580 423002 270592
rect 445294 270580 445300 270592
rect 445352 270580 445358 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 129458 270444 129464 270496
rect 129516 270484 129522 270496
rect 181162 270484 181168 270496
rect 129516 270456 181168 270484
rect 129516 270444 129522 270456
rect 181162 270444 181168 270456
rect 181220 270444 181226 270496
rect 191742 270444 191748 270496
rect 191800 270484 191806 270496
rect 196894 270484 196900 270496
rect 191800 270456 196900 270484
rect 191800 270444 191806 270456
rect 196894 270444 196900 270456
rect 196952 270444 196958 270496
rect 201770 270444 201776 270496
rect 201828 270484 201834 270496
rect 232222 270484 232228 270496
rect 201828 270456 232228 270484
rect 201828 270444 201834 270456
rect 232222 270444 232228 270456
rect 232280 270444 232286 270496
rect 395614 270444 395620 270496
rect 395672 270484 395678 270496
rect 433610 270484 433616 270496
rect 395672 270456 433616 270484
rect 395672 270444 395678 270456
rect 433610 270444 433616 270456
rect 433668 270444 433674 270496
rect 453574 270444 453580 270496
rect 453632 270484 453638 270496
rect 516778 270484 516784 270496
rect 453632 270456 516784 270484
rect 453632 270444 453638 270456
rect 516778 270444 516784 270456
rect 516836 270444 516842 270496
rect 517514 270444 517520 270496
rect 517572 270484 517578 270496
rect 579614 270484 579620 270496
rect 517572 270456 579620 270484
rect 517572 270444 517578 270456
rect 579614 270444 579620 270456
rect 579672 270444 579678 270496
rect 581638 270444 581644 270496
rect 581696 270484 581702 270496
rect 620278 270484 620284 270496
rect 581696 270456 620284 270484
rect 581696 270444 581702 270456
rect 620278 270444 620284 270456
rect 620336 270444 620342 270496
rect 88334 270308 88340 270360
rect 88392 270348 88398 270360
rect 121454 270348 121460 270360
rect 88392 270320 121460 270348
rect 88392 270308 88398 270320
rect 121454 270308 121460 270320
rect 121512 270308 121518 270360
rect 122466 270308 122472 270360
rect 122524 270348 122530 270360
rect 176194 270348 176200 270360
rect 122524 270320 176200 270348
rect 122524 270308 122530 270320
rect 176194 270308 176200 270320
rect 176252 270308 176258 270360
rect 180702 270308 180708 270360
rect 180760 270348 180766 270360
rect 215294 270348 215300 270360
rect 180760 270320 215300 270348
rect 180760 270308 180766 270320
rect 215294 270308 215300 270320
rect 215352 270308 215358 270360
rect 232774 270308 232780 270360
rect 232832 270348 232838 270360
rect 247862 270348 247868 270360
rect 232832 270320 247868 270348
rect 232832 270308 232838 270320
rect 247862 270308 247868 270320
rect 247920 270308 247926 270360
rect 262858 270308 262864 270360
rect 262916 270348 262922 270360
rect 262916 270320 267734 270348
rect 262916 270308 262922 270320
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 179322 270172 179328 270224
rect 179380 270212 179386 270224
rect 214098 270212 214104 270224
rect 179380 270184 214104 270212
rect 179380 270172 179386 270184
rect 214098 270172 214104 270184
rect 214156 270172 214162 270224
rect 226610 270172 226616 270224
rect 226668 270212 226674 270224
rect 249886 270212 249892 270224
rect 226668 270184 249892 270212
rect 226668 270172 226674 270184
rect 249886 270172 249892 270184
rect 249944 270172 249950 270224
rect 259730 270172 259736 270224
rect 259788 270212 259794 270224
rect 267706 270212 267734 270320
rect 367462 270308 367468 270360
rect 367520 270348 367526 270360
rect 393498 270348 393504 270360
rect 367520 270320 393504 270348
rect 367520 270308 367526 270320
rect 393498 270308 393504 270320
rect 393556 270308 393562 270360
rect 400858 270308 400864 270360
rect 400916 270348 400922 270360
rect 441614 270348 441620 270360
rect 400916 270320 441620 270348
rect 400916 270308 400922 270320
rect 441614 270308 441620 270320
rect 441672 270308 441678 270360
rect 456058 270308 456064 270360
rect 456116 270348 456122 270360
rect 520274 270348 520280 270360
rect 456116 270320 520280 270348
rect 456116 270308 456122 270320
rect 520274 270308 520280 270320
rect 520332 270308 520338 270360
rect 524414 270348 524420 270360
rect 521672 270320 524420 270348
rect 271414 270212 271420 270224
rect 259788 270184 265020 270212
rect 267706 270184 271420 270212
rect 259788 270172 259794 270184
rect 85482 270036 85488 270088
rect 85540 270076 85546 270088
rect 149422 270076 149428 270088
rect 85540 270048 149428 270076
rect 85540 270036 85546 270048
rect 149422 270036 149428 270048
rect 149480 270036 149486 270088
rect 173710 270036 173716 270088
rect 173768 270076 173774 270088
rect 212626 270076 212632 270088
rect 173768 270048 212632 270076
rect 173768 270036 173774 270048
rect 212626 270036 212632 270048
rect 212684 270036 212690 270088
rect 216490 270036 216496 270088
rect 216548 270076 216554 270088
rect 242434 270076 242440 270088
rect 216548 270048 242440 270076
rect 216548 270036 216554 270048
rect 242434 270036 242440 270048
rect 242492 270036 242498 270088
rect 248322 270036 248328 270088
rect 248380 270076 248386 270088
rect 264790 270076 264796 270088
rect 248380 270048 264796 270076
rect 248380 270036 248386 270048
rect 264790 270036 264796 270048
rect 264848 270036 264854 270088
rect 70578 269900 70584 269952
rect 70636 269940 70642 269952
rect 79962 269940 79968 269952
rect 70636 269912 79968 269940
rect 70636 269900 70642 269912
rect 79962 269900 79968 269912
rect 80020 269900 80026 269952
rect 80146 269900 80152 269952
rect 80204 269940 80210 269952
rect 146386 269940 146392 269952
rect 80204 269912 146392 269940
rect 80204 269900 80210 269912
rect 146386 269900 146392 269912
rect 146444 269900 146450 269952
rect 165430 269900 165436 269952
rect 165488 269940 165494 269952
rect 206002 269940 206008 269952
rect 165488 269912 206008 269940
rect 165488 269900 165494 269912
rect 206002 269900 206008 269912
rect 206060 269900 206066 269952
rect 210050 269900 210056 269952
rect 210108 269940 210114 269952
rect 238294 269940 238300 269952
rect 210108 269912 238300 269940
rect 210108 269900 210114 269912
rect 238294 269900 238300 269912
rect 238352 269900 238358 269952
rect 241974 269900 241980 269952
rect 242032 269940 242038 269952
rect 260374 269940 260380 269952
rect 242032 269912 260380 269940
rect 242032 269900 242038 269912
rect 260374 269900 260380 269912
rect 260432 269900 260438 269952
rect 264992 269940 265020 270184
rect 271414 270172 271420 270184
rect 271472 270172 271478 270224
rect 345106 270172 345112 270224
rect 345164 270212 345170 270224
rect 361574 270212 361580 270224
rect 345164 270184 361580 270212
rect 345164 270172 345170 270184
rect 361574 270172 361580 270184
rect 361632 270172 361638 270224
rect 364150 270172 364156 270224
rect 364208 270212 364214 270224
rect 389174 270212 389180 270224
rect 364208 270184 389180 270212
rect 364208 270172 364214 270184
rect 389174 270172 389180 270184
rect 389232 270172 389238 270224
rect 390094 270172 390100 270224
rect 390152 270212 390158 270224
rect 405734 270212 405740 270224
rect 390152 270184 405740 270212
rect 390152 270172 390158 270184
rect 405734 270172 405740 270184
rect 405792 270172 405798 270224
rect 409690 270172 409696 270224
rect 409748 270212 409754 270224
rect 454034 270212 454040 270224
rect 409748 270184 454040 270212
rect 409748 270172 409754 270184
rect 454034 270172 454040 270184
rect 454092 270172 454098 270224
rect 458542 270172 458548 270224
rect 458600 270212 458606 270224
rect 521672 270212 521700 270320
rect 524414 270308 524420 270320
rect 524472 270308 524478 270360
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 525668 270320 533384 270348
rect 525668 270308 525674 270320
rect 458600 270184 521700 270212
rect 458600 270172 458606 270184
rect 523126 270172 523132 270224
rect 523184 270212 523190 270224
rect 533154 270212 533160 270224
rect 523184 270184 533160 270212
rect 523184 270172 523190 270184
rect 533154 270172 533160 270184
rect 533212 270172 533218 270224
rect 533356 270212 533384 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 619634 270212 619640 270224
rect 533356 270184 619640 270212
rect 619634 270172 619640 270184
rect 619692 270172 619698 270224
rect 623958 270212 623964 270224
rect 619836 270184 623964 270212
rect 327718 270036 327724 270088
rect 327776 270076 327782 270088
rect 336734 270076 336740 270088
rect 327776 270048 336740 270076
rect 327776 270036 327782 270048
rect 336734 270036 336740 270048
rect 336792 270036 336798 270088
rect 345934 270036 345940 270088
rect 345992 270076 345998 270088
rect 362954 270076 362960 270088
rect 345992 270048 362960 270076
rect 345992 270036 345998 270048
rect 362954 270036 362960 270048
rect 363012 270036 363018 270088
rect 369946 270036 369952 270088
rect 370004 270076 370010 270088
rect 396074 270076 396080 270088
rect 370004 270048 396080 270076
rect 370004 270036 370010 270048
rect 396074 270036 396080 270048
rect 396132 270036 396138 270088
rect 399938 270036 399944 270088
rect 399996 270076 400002 270088
rect 412634 270076 412640 270088
rect 399996 270048 412640 270076
rect 399996 270036 400002 270048
rect 412634 270036 412640 270048
rect 412692 270036 412698 270088
rect 414658 270036 414664 270088
rect 414716 270076 414722 270088
rect 460934 270076 460940 270088
rect 414716 270048 460940 270076
rect 414716 270036 414722 270048
rect 460934 270036 460940 270048
rect 460992 270036 460998 270088
rect 461394 270036 461400 270088
rect 461452 270076 461458 270088
rect 527174 270076 527180 270088
rect 461452 270048 527180 270076
rect 461452 270036 461458 270048
rect 527174 270036 527180 270048
rect 527232 270036 527238 270088
rect 528370 270036 528376 270088
rect 528428 270076 528434 270088
rect 619836 270076 619864 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 528428 270048 619864 270076
rect 528428 270036 528434 270048
rect 620278 270036 620284 270088
rect 620336 270076 620342 270088
rect 630674 270076 630680 270088
rect 620336 270048 630680 270076
rect 620336 270036 620342 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 273070 269940 273076 269952
rect 264992 269912 273076 269940
rect 273070 269900 273076 269912
rect 273128 269900 273134 269952
rect 335078 269900 335084 269952
rect 335136 269940 335142 269952
rect 347774 269940 347780 269952
rect 335136 269912 347780 269940
rect 335136 269900 335142 269912
rect 347774 269900 347780 269912
rect 347832 269900 347838 269952
rect 351730 269900 351736 269952
rect 351788 269940 351794 269952
rect 371234 269940 371240 269952
rect 351788 269912 371240 269940
rect 351788 269900 351794 269912
rect 371234 269900 371240 269912
rect 371292 269900 371298 269952
rect 372430 269900 372436 269952
rect 372488 269940 372494 269952
rect 400490 269940 400496 269952
rect 372488 269912 400496 269940
rect 372488 269900 372494 269912
rect 400490 269900 400496 269912
rect 400548 269900 400554 269952
rect 401870 269900 401876 269952
rect 401928 269940 401934 269952
rect 416774 269940 416780 269952
rect 401928 269912 416780 269940
rect 401928 269900 401934 269912
rect 416774 269900 416780 269912
rect 416832 269900 416838 269952
rect 417142 269900 417148 269952
rect 417200 269940 417206 269952
rect 465074 269940 465080 269952
rect 417200 269912 465080 269940
rect 417200 269900 417206 269912
rect 465074 269900 465080 269912
rect 465132 269900 465138 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 468536 269912 531820 269940
rect 468536 269900 468542 269912
rect 76742 269764 76748 269816
rect 76800 269804 76806 269816
rect 143902 269804 143908 269816
rect 76800 269776 143908 269804
rect 76800 269764 76806 269776
rect 143902 269764 143908 269776
rect 143960 269764 143966 269816
rect 144362 269764 144368 269816
rect 144420 269804 144426 269816
rect 190822 269804 190828 269816
rect 144420 269776 190828 269804
rect 144420 269764 144426 269776
rect 190822 269764 190828 269776
rect 190880 269764 190886 269816
rect 202966 269764 202972 269816
rect 203024 269804 203030 269816
rect 233326 269804 233332 269816
rect 203024 269776 233332 269804
rect 203024 269764 203030 269776
rect 233326 269764 233332 269776
rect 233384 269764 233390 269816
rect 241422 269764 241428 269816
rect 241480 269804 241486 269816
rect 259822 269804 259828 269816
rect 241480 269776 259828 269804
rect 241480 269764 241486 269776
rect 259822 269764 259828 269776
rect 259880 269764 259886 269816
rect 261938 269764 261944 269816
rect 261996 269804 262002 269816
rect 274726 269804 274732 269816
rect 261996 269776 274732 269804
rect 261996 269764 262002 269776
rect 274726 269764 274732 269776
rect 274784 269764 274790 269816
rect 280062 269764 280068 269816
rect 280120 269804 280126 269816
rect 287146 269804 287152 269816
rect 280120 269776 287152 269804
rect 280120 269764 280126 269776
rect 287146 269764 287152 269776
rect 287204 269764 287210 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 336826 269764 336832 269816
rect 336884 269804 336890 269816
rect 350534 269804 350540 269816
rect 336884 269776 350540 269804
rect 336884 269764 336890 269776
rect 350534 269764 350540 269776
rect 350592 269764 350598 269816
rect 355042 269764 355048 269816
rect 355100 269804 355106 269816
rect 376938 269804 376944 269816
rect 355100 269776 376944 269804
rect 355100 269764 355106 269776
rect 376938 269764 376944 269776
rect 376996 269764 377002 269816
rect 377674 269764 377680 269816
rect 377732 269804 377738 269816
rect 408494 269804 408500 269816
rect 377732 269776 408500 269804
rect 377732 269764 377738 269776
rect 408494 269764 408500 269776
rect 408552 269764 408558 269816
rect 412450 269764 412456 269816
rect 412508 269804 412514 269816
rect 458266 269804 458272 269816
rect 412508 269776 458272 269804
rect 412508 269764 412514 269776
rect 458266 269764 458272 269776
rect 458324 269764 458330 269816
rect 463510 269764 463516 269816
rect 463568 269804 463574 269816
rect 531314 269804 531320 269816
rect 463568 269776 531320 269804
rect 463568 269764 463574 269776
rect 531314 269764 531320 269776
rect 531372 269764 531378 269816
rect 531792 269804 531820 269912
rect 531958 269900 531964 269952
rect 532016 269940 532022 269952
rect 533522 269940 533528 269952
rect 532016 269912 533528 269940
rect 532016 269900 532022 269912
rect 533522 269900 533528 269912
rect 533580 269900 533586 269952
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 537754 269940 537760 269952
rect 534040 269912 537760 269940
rect 534040 269900 534046 269912
rect 537754 269900 537760 269912
rect 537812 269900 537818 269952
rect 537938 269900 537944 269952
rect 537996 269940 538002 269952
rect 537996 269912 543044 269940
rect 537996 269900 538002 269912
rect 538490 269804 538496 269816
rect 531792 269776 538496 269804
rect 538490 269764 538496 269776
rect 538548 269764 538554 269816
rect 538674 269764 538680 269816
rect 538732 269804 538738 269816
rect 542814 269804 542820 269816
rect 538732 269776 542820 269804
rect 538732 269764 538738 269776
rect 542814 269764 542820 269776
rect 542872 269764 542878 269816
rect 543016 269804 543044 269912
rect 543182 269900 543188 269952
rect 543240 269940 543246 269952
rect 640518 269940 640524 269952
rect 543240 269912 640524 269940
rect 543240 269900 543246 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 637574 269804 637580 269816
rect 543016 269776 637580 269804
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 126882 269628 126888 269680
rect 126940 269668 126946 269680
rect 178310 269668 178316 269680
rect 126940 269640 178316 269668
rect 126940 269628 126946 269640
rect 178310 269628 178316 269640
rect 178368 269628 178374 269680
rect 200482 269628 200488 269680
rect 200540 269668 200546 269680
rect 226886 269668 226892 269680
rect 200540 269640 226892 269668
rect 200540 269628 200546 269640
rect 226886 269628 226892 269640
rect 226944 269628 226950 269680
rect 384758 269628 384764 269680
rect 384816 269668 384822 269680
rect 418246 269668 418252 269680
rect 384816 269640 418252 269668
rect 384816 269628 384822 269640
rect 418246 269628 418252 269640
rect 418304 269628 418310 269680
rect 422110 269628 422116 269680
rect 422168 269668 422174 269680
rect 471974 269668 471980 269680
rect 422168 269640 471980 269668
rect 422168 269628 422174 269640
rect 471974 269628 471980 269640
rect 472032 269628 472038 269680
rect 472618 269628 472624 269680
rect 472676 269668 472682 269680
rect 473354 269668 473360 269680
rect 472676 269640 473360 269668
rect 472676 269628 472682 269640
rect 473354 269628 473360 269640
rect 473412 269628 473418 269680
rect 530394 269668 530400 269680
rect 480226 269640 530400 269668
rect 78858 269492 78864 269544
rect 78916 269532 78922 269544
rect 130378 269532 130384 269544
rect 78916 269504 130384 269532
rect 78916 269492 78922 269504
rect 130378 269492 130384 269504
rect 130436 269492 130442 269544
rect 133782 269492 133788 269544
rect 133840 269532 133846 269544
rect 183646 269532 183652 269544
rect 133840 269504 183652 269532
rect 133840 269492 133846 269504
rect 183646 269492 183652 269504
rect 183704 269492 183710 269544
rect 186406 269492 186412 269544
rect 186464 269532 186470 269544
rect 204070 269532 204076 269544
rect 186464 269504 204076 269532
rect 186464 269492 186470 269504
rect 204070 269492 204076 269504
rect 204128 269492 204134 269544
rect 392026 269492 392032 269544
rect 392084 269532 392090 269544
rect 401686 269532 401692 269544
rect 392084 269504 401692 269532
rect 392084 269492 392090 269504
rect 401686 269492 401692 269504
rect 401744 269492 401750 269544
rect 404538 269492 404544 269544
rect 404596 269532 404602 269544
rect 423674 269532 423680 269544
rect 404596 269504 423680 269532
rect 404596 269492 404602 269504
rect 423674 269492 423680 269504
rect 423732 269492 423738 269544
rect 432230 269492 432236 269544
rect 432288 269532 432294 269544
rect 466454 269532 466460 269544
rect 432288 269504 466460 269532
rect 432288 269492 432294 269504
rect 466454 269492 466460 269504
rect 466512 269492 466518 269544
rect 480226 269532 480254 269640
rect 530394 269628 530400 269640
rect 530452 269628 530458 269680
rect 530578 269628 530584 269680
rect 530636 269668 530642 269680
rect 531958 269668 531964 269680
rect 530636 269640 531964 269668
rect 530636 269628 530642 269640
rect 531958 269628 531964 269640
rect 532016 269628 532022 269680
rect 533154 269628 533160 269680
rect 533212 269668 533218 269680
rect 616138 269668 616144 269680
rect 533212 269640 616144 269668
rect 533212 269628 533218 269640
rect 616138 269628 616144 269640
rect 616196 269628 616202 269680
rect 470566 269504 480254 269532
rect 140682 269356 140688 269408
rect 140740 269396 140746 269408
rect 188614 269396 188620 269408
rect 140740 269368 188620 269396
rect 140740 269356 140746 269368
rect 188614 269356 188620 269368
rect 188672 269356 188678 269408
rect 429102 269356 429108 269408
rect 429160 269396 429166 269408
rect 455414 269396 455420 269408
rect 429160 269368 455420 269396
rect 429160 269356 429166 269368
rect 455414 269356 455420 269368
rect 455472 269356 455478 269408
rect 465994 269356 466000 269408
rect 466052 269396 466058 269408
rect 470566 269396 470594 269504
rect 509050 269492 509056 269544
rect 509108 269532 509114 269544
rect 596174 269532 596180 269544
rect 509108 269504 596180 269532
rect 509108 269492 509114 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 466052 269368 470594 269396
rect 466052 269356 466058 269368
rect 474642 269356 474648 269408
rect 474700 269396 474706 269408
rect 538122 269396 538128 269408
rect 474700 269368 538128 269396
rect 474700 269356 474706 269368
rect 538122 269356 538128 269368
rect 538180 269356 538186 269408
rect 538306 269356 538312 269408
rect 538364 269396 538370 269408
rect 581638 269396 581644 269408
rect 538364 269368 581644 269396
rect 538364 269356 538370 269368
rect 581638 269356 581644 269368
rect 581696 269356 581702 269408
rect 121638 269220 121644 269272
rect 121696 269260 121702 269272
rect 167822 269260 167828 269272
rect 121696 269232 167828 269260
rect 121696 269220 121702 269232
rect 167822 269220 167828 269232
rect 167880 269220 167886 269272
rect 272426 269220 272432 269272
rect 272484 269260 272490 269272
rect 278866 269260 278872 269272
rect 272484 269232 278872 269260
rect 272484 269220 272490 269232
rect 278866 269220 278872 269232
rect 278924 269220 278930 269272
rect 423950 269220 423956 269272
rect 424008 269260 424014 269272
rect 448514 269260 448520 269272
rect 424008 269232 448520 269260
rect 424008 269220 424014 269232
rect 448514 269220 448520 269232
rect 448572 269220 448578 269272
rect 470962 269220 470968 269272
rect 471020 269260 471026 269272
rect 540606 269260 540612 269272
rect 471020 269232 540612 269260
rect 471020 269220 471026 269232
rect 540606 269220 540612 269232
rect 540664 269220 540670 269272
rect 540790 269220 540796 269272
rect 540848 269260 540854 269272
rect 543182 269260 543188 269272
rect 540848 269232 543188 269260
rect 540848 269220 540854 269232
rect 543182 269220 543188 269232
rect 543240 269220 543246 269272
rect 543366 269152 543372 269204
rect 543424 269192 543430 269204
rect 546494 269192 546500 269204
rect 543424 269164 546500 269192
rect 543424 269152 543430 269164
rect 546494 269152 546500 269164
rect 546552 269152 546558 269204
rect 274910 269084 274916 269136
rect 274968 269124 274974 269136
rect 279694 269124 279700 269136
rect 274968 269096 279700 269124
rect 274968 269084 274974 269096
rect 279694 269084 279700 269096
rect 279752 269084 279758 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 42150 269016 42156 269068
rect 42208 269056 42214 269068
rect 43162 269056 43168 269068
rect 42208 269028 43168 269056
rect 42208 269016 42214 269028
rect 43162 269016 43168 269028
rect 43220 269016 43226 269068
rect 84102 269016 84108 269068
rect 84160 269056 84166 269068
rect 137462 269056 137468 269068
rect 84160 269028 137468 269056
rect 84160 269016 84166 269028
rect 137462 269016 137468 269028
rect 137520 269016 137526 269068
rect 137646 269016 137652 269068
rect 137704 269056 137710 269068
rect 186130 269056 186136 269068
rect 137704 269028 186136 269056
rect 137704 269016 137710 269028
rect 186130 269016 186136 269028
rect 186188 269016 186194 269068
rect 379698 269016 379704 269068
rect 379756 269056 379762 269068
rect 404354 269056 404360 269068
rect 379756 269028 404360 269056
rect 379756 269016 379762 269028
rect 404354 269016 404360 269028
rect 404412 269016 404418 269068
rect 436186 269016 436192 269068
rect 436244 269056 436250 269068
rect 491754 269056 491760 269068
rect 436244 269028 491760 269056
rect 436244 269016 436250 269028
rect 491754 269016 491760 269028
rect 491812 269016 491818 269068
rect 498286 269016 498292 269068
rect 498344 269056 498350 269068
rect 580994 269056 581000 269068
rect 498344 269028 581000 269056
rect 498344 269016 498350 269028
rect 580994 269016 581000 269028
rect 581052 269016 581058 269068
rect 273254 268948 273260 269000
rect 273312 268988 273318 269000
rect 275554 268988 275560 269000
rect 273312 268960 275560 268988
rect 273312 268948 273318 268960
rect 275554 268948 275560 268960
rect 275612 268948 275618 269000
rect 111978 268880 111984 268932
rect 112036 268920 112042 268932
rect 168742 268920 168748 268932
rect 112036 268892 168748 268920
rect 112036 268880 112042 268892
rect 168742 268880 168748 268892
rect 168800 268880 168806 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415394 268920 415400 268932
rect 382424 268892 415400 268920
rect 382424 268880 382430 268892
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 433702 268880 433708 268932
rect 433760 268920 433766 268932
rect 488534 268920 488540 268932
rect 433760 268892 488540 268920
rect 433760 268880 433766 268892
rect 488534 268880 488540 268892
rect 488592 268880 488598 268932
rect 500770 268880 500776 268932
rect 500828 268920 500834 268932
rect 583754 268920 583760 268932
rect 500828 268892 583760 268920
rect 500828 268880 500834 268892
rect 583754 268880 583760 268892
rect 583812 268880 583818 268932
rect 115842 268744 115848 268796
rect 115900 268784 115906 268796
rect 115900 268756 166304 268784
rect 115900 268744 115906 268756
rect 110230 268608 110236 268660
rect 110288 268648 110294 268660
rect 110288 268620 164648 268648
rect 110288 268608 110294 268620
rect 102502 268472 102508 268524
rect 102560 268512 102566 268524
rect 162946 268512 162952 268524
rect 102560 268484 162952 268512
rect 102560 268472 102566 268484
rect 162946 268472 162952 268484
rect 163004 268472 163010 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 164620 268376 164648 268620
rect 166276 268512 166304 268756
rect 211338 268744 211344 268796
rect 211396 268784 211402 268796
rect 223482 268784 223488 268796
rect 211396 268756 223488 268784
rect 211396 268744 211402 268756
rect 223482 268744 223488 268756
rect 223540 268744 223546 268796
rect 389818 268744 389824 268796
rect 389876 268784 389882 268796
rect 425330 268784 425336 268796
rect 389876 268756 425336 268784
rect 389876 268744 389882 268756
rect 425330 268744 425336 268756
rect 425388 268744 425394 268796
rect 441154 268744 441160 268796
rect 441212 268784 441218 268796
rect 499574 268784 499580 268796
rect 441212 268756 499580 268784
rect 441212 268744 441218 268756
rect 499574 268744 499580 268756
rect 499632 268744 499638 268796
rect 505738 268744 505744 268796
rect 505796 268784 505802 268796
rect 590838 268784 590844 268796
rect 505796 268756 590844 268784
rect 505796 268744 505802 268756
rect 590838 268744 590844 268756
rect 590896 268744 590902 268796
rect 166994 268608 167000 268660
rect 167052 268648 167058 268660
rect 184474 268648 184480 268660
rect 167052 268620 184480 268648
rect 167052 268608 167058 268620
rect 184474 268608 184480 268620
rect 184532 268608 184538 268660
rect 187326 268608 187332 268660
rect 187384 268648 187390 268660
rect 219434 268648 219440 268660
rect 187384 268620 219440 268648
rect 187384 268608 187390 268620
rect 219434 268608 219440 268620
rect 219492 268608 219498 268660
rect 245562 268608 245568 268660
rect 245620 268648 245626 268660
rect 263134 268648 263140 268660
rect 245620 268620 263140 268648
rect 245620 268608 245626 268620
rect 263134 268608 263140 268620
rect 263192 268608 263198 268660
rect 396166 268608 396172 268660
rect 396224 268648 396230 268660
rect 433334 268648 433340 268660
rect 396224 268620 433340 268648
rect 396224 268608 396230 268620
rect 433334 268608 433340 268620
rect 433392 268608 433398 268660
rect 443638 268608 443644 268660
rect 443696 268648 443702 268660
rect 502334 268648 502340 268660
rect 443696 268620 502340 268648
rect 443696 268608 443702 268620
rect 502334 268608 502340 268620
rect 502392 268608 502398 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 171226 268512 171232 268524
rect 166276 268484 171232 268512
rect 171226 268472 171232 268484
rect 171284 268472 171290 268524
rect 176930 268472 176936 268524
rect 176988 268512 176994 268524
rect 215110 268512 215116 268524
rect 176988 268484 215116 268512
rect 176988 268472 176994 268484
rect 215110 268472 215116 268484
rect 215168 268472 215174 268524
rect 220446 268472 220452 268524
rect 220504 268512 220510 268524
rect 245746 268512 245752 268524
rect 220504 268484 245752 268512
rect 220504 268472 220510 268484
rect 245746 268472 245752 268484
rect 245804 268472 245810 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 350718 268512 350724 268524
rect 338540 268484 350724 268512
rect 338540 268472 338546 268484
rect 350718 268472 350724 268484
rect 350776 268472 350782 268524
rect 359826 268472 359832 268524
rect 359884 268512 359890 268524
rect 379514 268512 379520 268524
rect 359884 268484 379520 268512
rect 359884 268472 359890 268484
rect 379514 268472 379520 268484
rect 379572 268472 379578 268524
rect 403250 268472 403256 268524
rect 403308 268512 403314 268524
rect 440234 268512 440240 268524
rect 403308 268484 440240 268512
rect 403308 268472 403314 268484
rect 440234 268472 440240 268484
rect 440292 268472 440298 268524
rect 448606 268472 448612 268524
rect 448664 268512 448670 268524
rect 509234 268512 509240 268524
rect 448664 268484 509240 268512
rect 448664 268472 448670 268484
rect 509234 268472 509240 268484
rect 509292 268472 509298 268524
rect 513190 268472 513196 268524
rect 513248 268512 513254 268524
rect 601694 268512 601700 268524
rect 513248 268484 601700 268512
rect 513248 268472 513254 268484
rect 601694 268472 601700 268484
rect 601752 268472 601758 268524
rect 167638 268376 167644 268388
rect 164620 268348 167644 268376
rect 167638 268336 167644 268348
rect 167696 268336 167702 268388
rect 168006 268336 168012 268388
rect 168064 268376 168070 268388
rect 203518 268376 203524 268388
rect 168064 268348 203524 268376
rect 168064 268336 168070 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 203886 268336 203892 268388
rect 203944 268376 203950 268388
rect 230750 268376 230756 268388
rect 203944 268348 230756 268376
rect 203944 268336 203950 268348
rect 230750 268336 230756 268348
rect 230808 268336 230814 268388
rect 231670 268336 231676 268388
rect 231728 268376 231734 268388
rect 253198 268376 253204 268388
rect 231728 268348 253204 268376
rect 231728 268336 231734 268348
rect 253198 268336 253204 268348
rect 253256 268336 253262 268388
rect 258350 268336 258356 268388
rect 258408 268376 258414 268388
rect 268930 268376 268936 268388
rect 258408 268348 268936 268376
rect 258408 268336 258414 268348
rect 268930 268336 268936 268348
rect 268988 268336 268994 268388
rect 348418 268336 348424 268388
rect 348476 268376 348482 268388
rect 367094 268376 367100 268388
rect 348476 268348 367100 268376
rect 348476 268336 348482 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372154 268336 372160 268388
rect 372212 268376 372218 268388
rect 397454 268376 397460 268388
rect 372212 268348 397460 268376
rect 372212 268336 372218 268348
rect 397454 268336 397460 268348
rect 397512 268336 397518 268388
rect 408034 268336 408040 268388
rect 408092 268376 408098 268388
rect 451366 268376 451372 268388
rect 408092 268348 451372 268376
rect 408092 268336 408098 268348
rect 451366 268336 451372 268348
rect 451424 268336 451430 268388
rect 464338 268336 464344 268388
rect 464396 268376 464402 268388
rect 532694 268376 532700 268388
rect 464396 268348 532700 268376
rect 464396 268336 464402 268348
rect 532694 268336 532700 268348
rect 532752 268336 532758 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 128538 268200 128544 268252
rect 128596 268240 128602 268252
rect 150434 268240 150440 268252
rect 128596 268212 150440 268240
rect 128596 268200 128602 268212
rect 150434 268200 150440 268212
rect 150492 268200 150498 268252
rect 151722 268200 151728 268252
rect 151780 268240 151786 268252
rect 196066 268240 196072 268252
rect 151780 268212 196072 268240
rect 151780 268200 151786 268212
rect 196066 268200 196072 268212
rect 196124 268200 196130 268252
rect 419626 268200 419632 268252
rect 419684 268240 419690 268252
rect 467926 268240 467932 268252
rect 419684 268212 467932 268240
rect 419684 268200 419690 268212
rect 467926 268200 467932 268212
rect 467984 268200 467990 268252
rect 493594 268200 493600 268252
rect 493652 268240 493658 268252
rect 574094 268240 574100 268252
rect 493652 268212 574100 268240
rect 493652 268200 493658 268212
rect 574094 268200 574100 268212
rect 574152 268200 574158 268252
rect 163130 268064 163136 268116
rect 163188 268104 163194 268116
rect 168006 268104 168012 268116
rect 163188 268076 168012 268104
rect 163188 268064 163194 268076
rect 168006 268064 168012 268076
rect 168064 268064 168070 268116
rect 412634 268064 412640 268116
rect 412692 268104 412698 268116
rect 447134 268104 447140 268116
rect 412692 268076 447140 268104
rect 412692 268064 412698 268076
rect 447134 268064 447140 268076
rect 447192 268064 447198 268116
rect 495802 268064 495808 268116
rect 495860 268104 495866 268116
rect 576854 268104 576860 268116
rect 495860 268076 576860 268104
rect 495860 268064 495866 268076
rect 576854 268064 576860 268076
rect 576912 268064 576918 268116
rect 198734 267792 198740 267844
rect 198792 267832 198798 267844
rect 201862 267832 201868 267844
rect 198792 267804 201868 267832
rect 198792 267792 198798 267804
rect 201862 267792 201868 267804
rect 201920 267792 201926 267844
rect 117682 267656 117688 267708
rect 117740 267696 117746 267708
rect 159634 267696 159640 267708
rect 117740 267668 159640 267696
rect 117740 267656 117746 267668
rect 159634 267656 159640 267668
rect 159692 267656 159698 267708
rect 167822 267656 167828 267708
rect 167880 267696 167886 267708
rect 177022 267696 177028 267708
rect 167880 267668 177028 267696
rect 167880 267656 167886 267668
rect 177022 267656 177028 267668
rect 177080 267656 177086 267708
rect 181990 267656 181996 267708
rect 182048 267696 182054 267708
rect 182048 267668 182312 267696
rect 182048 267656 182054 267668
rect 95878 267520 95884 267572
rect 95936 267560 95942 267572
rect 138106 267560 138112 267572
rect 95936 267532 138112 267560
rect 95936 267520 95942 267532
rect 138106 267520 138112 267532
rect 138164 267520 138170 267572
rect 150434 267520 150440 267572
rect 150492 267560 150498 267572
rect 181990 267560 181996 267572
rect 150492 267532 181996 267560
rect 150492 267520 150498 267532
rect 181990 267520 181996 267532
rect 182048 267520 182054 267572
rect 182284 267560 182312 267668
rect 182726 267656 182732 267708
rect 182784 267696 182790 267708
rect 214282 267696 214288 267708
rect 182784 267668 214288 267696
rect 182784 267656 182790 267668
rect 214282 267656 214288 267668
rect 214340 267656 214346 267708
rect 378226 267656 378232 267708
rect 378284 267696 378290 267708
rect 392578 267696 392584 267708
rect 378284 267668 392584 267696
rect 378284 267656 378290 267668
rect 392578 267656 392584 267668
rect 392636 267656 392642 267708
rect 398098 267656 398104 267708
rect 398156 267696 398162 267708
rect 414474 267696 414480 267708
rect 398156 267668 414480 267696
rect 398156 267656 398162 267668
rect 414474 267656 414480 267668
rect 414532 267656 414538 267708
rect 423766 267656 423772 267708
rect 423824 267696 423830 267708
rect 440878 267696 440884 267708
rect 423824 267668 440884 267696
rect 423824 267656 423830 267668
rect 440878 267656 440884 267668
rect 440936 267656 440942 267708
rect 450262 267656 450268 267708
rect 450320 267696 450326 267708
rect 501598 267696 501604 267708
rect 450320 267668 501604 267696
rect 450320 267656 450326 267668
rect 501598 267656 501604 267668
rect 501656 267656 501662 267708
rect 514846 267656 514852 267708
rect 514904 267696 514910 267708
rect 571978 267696 571984 267708
rect 514904 267668 571984 267696
rect 514904 267656 514910 267668
rect 571978 267656 571984 267668
rect 572036 267656 572042 267708
rect 219250 267560 219256 267572
rect 182284 267532 219256 267560
rect 219250 267520 219256 267532
rect 219308 267520 219314 267572
rect 340966 267520 340972 267572
rect 341024 267560 341030 267572
rect 355318 267560 355324 267572
rect 341024 267532 355324 267560
rect 341024 267520 341030 267532
rect 355318 267520 355324 267532
rect 355376 267520 355382 267572
rect 362494 267520 362500 267572
rect 362552 267560 362558 267572
rect 369118 267560 369124 267572
rect 362552 267532 369124 267560
rect 362552 267520 362558 267532
rect 369118 267520 369124 267532
rect 369176 267520 369182 267572
rect 370774 267520 370780 267572
rect 370832 267560 370838 267572
rect 377398 267560 377404 267572
rect 370832 267532 377404 267560
rect 370832 267520 370838 267532
rect 377398 267520 377404 267532
rect 377456 267520 377462 267572
rect 380710 267520 380716 267572
rect 380768 267560 380774 267572
rect 399938 267560 399944 267572
rect 380768 267532 399944 267560
rect 380768 267520 380774 267532
rect 399938 267520 399944 267532
rect 399996 267520 400002 267572
rect 410518 267520 410524 267572
rect 410576 267560 410582 267572
rect 429102 267560 429108 267572
rect 410576 267532 429108 267560
rect 410576 267520 410582 267532
rect 429102 267520 429108 267532
rect 429160 267520 429166 267572
rect 445294 267520 445300 267572
rect 445352 267560 445358 267572
rect 497458 267560 497464 267572
rect 445352 267532 497464 267560
rect 445352 267520 445358 267532
rect 497458 267520 497464 267532
rect 497516 267520 497522 267572
rect 504818 267520 504824 267572
rect 504876 267560 504882 267572
rect 517514 267560 517520 267572
rect 504876 267532 517520 267560
rect 504876 267520 504882 267532
rect 517514 267520 517520 267532
rect 517572 267520 517578 267572
rect 529658 267520 529664 267572
rect 529716 267560 529722 267572
rect 585778 267560 585784 267572
rect 529716 267532 585784 267560
rect 529716 267520 529722 267532
rect 585778 267520 585784 267532
rect 585836 267520 585842 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 146938 267384 146944 267436
rect 146996 267424 147002 267436
rect 186958 267424 186964 267436
rect 146996 267396 186964 267424
rect 146996 267384 147002 267396
rect 186958 267384 186964 267396
rect 187016 267384 187022 267436
rect 236638 267384 236644 267436
rect 236696 267424 236702 267436
rect 241606 267424 241612 267436
rect 236696 267396 241612 267424
rect 236696 267384 236702 267396
rect 241606 267384 241612 267396
rect 241664 267384 241670 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 319162 267424 319168 267436
rect 315356 267396 319168 267424
rect 315356 267384 315362 267396
rect 319162 267384 319168 267396
rect 319220 267384 319226 267436
rect 350074 267384 350080 267436
rect 350132 267424 350138 267436
rect 358078 267424 358084 267436
rect 350132 267396 358084 267424
rect 350132 267384 350138 267396
rect 358078 267384 358084 267396
rect 358136 267384 358142 267436
rect 371602 267384 371608 267436
rect 371660 267424 371666 267436
rect 373258 267424 373264 267436
rect 371660 267396 373264 267424
rect 371660 267384 371666 267396
rect 373258 267384 373264 267396
rect 373316 267384 373322 267436
rect 383194 267384 383200 267436
rect 383252 267424 383258 267436
rect 401870 267424 401876 267436
rect 383252 267396 401876 267424
rect 383252 267384 383258 267396
rect 401870 267384 401876 267396
rect 401928 267384 401934 267436
rect 405550 267384 405556 267436
rect 405608 267424 405614 267436
rect 423950 267424 423956 267436
rect 405608 267396 423956 267424
rect 405608 267384 405614 267396
rect 423950 267384 423956 267396
rect 424008 267384 424014 267436
rect 432046 267384 432052 267436
rect 432104 267424 432110 267436
rect 453298 267424 453304 267436
rect 432104 267396 453304 267424
rect 432104 267384 432110 267396
rect 453298 267384 453304 267396
rect 453356 267384 453362 267436
rect 460198 267384 460204 267436
rect 460256 267424 460262 267436
rect 515398 267424 515404 267436
rect 460256 267396 515404 267424
rect 460256 267384 460262 267396
rect 515398 267384 515404 267396
rect 515456 267384 515462 267436
rect 519814 267384 519820 267436
rect 519872 267424 519878 267436
rect 578878 267424 578884 267436
rect 519872 267396 578884 267424
rect 519872 267384 519878 267396
rect 578878 267384 578884 267396
rect 578936 267384 578942 267436
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 169018 267248 169024 267300
rect 169076 267288 169082 267300
rect 209314 267288 209320 267300
rect 169076 267260 209320 267288
rect 169076 267248 169082 267260
rect 209314 267248 209320 267260
rect 209372 267248 209378 267300
rect 218698 267248 218704 267300
rect 218756 267288 218762 267300
rect 223022 267288 223028 267300
rect 218756 267260 223028 267288
rect 218756 267248 218762 267260
rect 223022 267248 223028 267260
rect 223080 267248 223086 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 239122 267288 239128 267300
rect 223540 267260 239128 267288
rect 223540 267248 223546 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 353386 267248 353392 267300
rect 353444 267288 353450 267300
rect 364978 267288 364984 267300
rect 353444 267260 364984 267288
rect 353444 267248 353450 267260
rect 364978 267248 364984 267260
rect 365036 267248 365042 267300
rect 373258 267248 373264 267300
rect 373316 267288 373322 267300
rect 392026 267288 392032 267300
rect 373316 267260 392032 267288
rect 373316 267248 373322 267260
rect 392026 267248 392032 267260
rect 392084 267248 392090 267300
rect 403066 267248 403072 267300
rect 403124 267288 403130 267300
rect 422938 267288 422944 267300
rect 403124 267260 422944 267288
rect 403124 267248 403130 267260
rect 422938 267248 422944 267260
rect 422996 267248 423002 267300
rect 424594 267248 424600 267300
rect 424652 267288 424658 267300
rect 446398 267288 446404 267300
rect 424652 267260 446404 267288
rect 424652 267248 424658 267260
rect 446398 267248 446404 267260
rect 446456 267248 446462 267300
rect 448146 267248 448152 267300
rect 448204 267288 448210 267300
rect 457438 267288 457444 267300
rect 448204 267260 457444 267288
rect 448204 267248 448210 267260
rect 457438 267248 457444 267260
rect 457496 267248 457502 267300
rect 470134 267248 470140 267300
rect 470192 267288 470198 267300
rect 534718 267288 534724 267300
rect 470192 267260 534724 267288
rect 470192 267248 470198 267260
rect 534718 267248 534724 267260
rect 534776 267248 534782 267300
rect 542998 267248 543004 267300
rect 543056 267288 543062 267300
rect 625798 267288 625804 267300
rect 543056 267260 625804 267288
rect 543056 267248 543062 267260
rect 625798 267248 625804 267260
rect 625856 267248 625862 267300
rect 79962 267112 79968 267164
rect 80020 267152 80026 267164
rect 140590 267152 140596 267164
rect 80020 267124 140596 267152
rect 80020 267112 80026 267124
rect 140590 267112 140596 267124
rect 140648 267112 140654 267164
rect 144178 267112 144184 267164
rect 144236 267152 144242 267164
rect 191926 267152 191932 267164
rect 144236 267124 191932 267152
rect 144236 267112 144242 267124
rect 191926 267112 191932 267124
rect 191984 267112 191990 267164
rect 192570 267112 192576 267164
rect 192628 267152 192634 267164
rect 223942 267152 223948 267164
rect 192628 267124 223948 267152
rect 192628 267112 192634 267124
rect 223942 267112 223948 267124
rect 224000 267112 224006 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 317782 267112 317788 267164
rect 317840 267152 317846 267164
rect 322934 267152 322940 267164
rect 317840 267124 322940 267152
rect 317840 267112 317846 267124
rect 322934 267112 322940 267124
rect 322992 267112 322998 267164
rect 365806 267112 365812 267164
rect 365864 267152 365870 267164
rect 382918 267152 382924 267164
rect 365864 267124 382924 267152
rect 365864 267112 365870 267124
rect 382918 267112 382924 267124
rect 382976 267112 382982 267164
rect 390646 267112 390652 267164
rect 390704 267152 390710 267164
rect 417418 267152 417424 267164
rect 390704 267124 417424 267152
rect 390704 267112 390710 267124
rect 417418 267112 417424 267124
rect 417476 267112 417482 267164
rect 417970 267112 417976 267164
rect 418028 267152 418034 267164
rect 432230 267152 432236 267164
rect 418028 267124 432236 267152
rect 418028 267112 418034 267124
rect 432230 267112 432236 267124
rect 432288 267112 432294 267164
rect 432874 267112 432880 267164
rect 432932 267152 432938 267164
rect 460014 267152 460020 267164
rect 432932 267124 460020 267152
rect 432932 267112 432938 267124
rect 460014 267112 460020 267124
rect 460072 267112 460078 267164
rect 465166 267112 465172 267164
rect 465224 267152 465230 267164
rect 526438 267152 526444 267164
rect 465224 267124 526444 267152
rect 465224 267112 465230 267124
rect 526438 267112 526444 267124
rect 526496 267112 526502 267164
rect 534718 267112 534724 267164
rect 534776 267152 534782 267164
rect 618898 267152 618904 267164
rect 534776 267124 618904 267152
rect 534776 267112 534782 267124
rect 618898 267112 618904 267124
rect 618956 267112 618962 267164
rect 90358 266976 90364 267028
rect 90416 267016 90422 267028
rect 151354 267016 151360 267028
rect 90416 266988 151360 267016
rect 90416 266976 90422 266988
rect 151354 266976 151360 266988
rect 151412 266976 151418 267028
rect 154482 266976 154488 267028
rect 154540 267016 154546 267028
rect 199378 267016 199384 267028
rect 154540 266988 199384 267016
rect 154540 266976 154546 266988
rect 199378 266976 199384 266988
rect 199436 266976 199442 267028
rect 218882 266976 218888 267028
rect 218940 267016 218946 267028
rect 220078 267016 220084 267028
rect 218940 266988 220084 267016
rect 218940 266976 218946 266988
rect 220078 266976 220084 266988
rect 220136 266976 220142 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 228416 266988 238754 267016
rect 228416 266976 228422 266988
rect 121454 266840 121460 266892
rect 121512 266880 121518 266892
rect 144914 266880 144920 266892
rect 121512 266852 144920 266880
rect 121512 266840 121518 266852
rect 144914 266840 144920 266852
rect 144972 266840 144978 266892
rect 145374 266840 145380 266892
rect 145432 266880 145438 266892
rect 150526 266880 150532 266892
rect 145432 266852 150532 266880
rect 145432 266840 145438 266852
rect 150526 266840 150532 266852
rect 150584 266840 150590 266892
rect 204070 266840 204076 266892
rect 204128 266880 204134 266892
rect 220906 266880 220912 266892
rect 204128 266852 220912 266880
rect 204128 266840 204134 266852
rect 220906 266840 220912 266852
rect 220964 266840 220970 266892
rect 238726 266880 238754 266988
rect 314470 266976 314476 267028
rect 314528 267016 314534 267028
rect 318978 267016 318984 267028
rect 314528 266988 318984 267016
rect 314528 266976 314534 266988
rect 318978 266976 318984 266988
rect 319036 266976 319042 267028
rect 355870 266976 355876 267028
rect 355928 267016 355934 267028
rect 374638 267016 374644 267028
rect 355928 266988 374644 267016
rect 355928 266976 355934 266988
rect 374638 266976 374644 266988
rect 374696 266976 374702 267028
rect 375742 266976 375748 267028
rect 375800 267016 375806 267028
rect 390094 267016 390100 267028
rect 375800 266988 390100 267016
rect 375800 266976 375806 266988
rect 390094 266976 390100 266988
rect 390152 266976 390158 267028
rect 393130 266976 393136 267028
rect 393188 267016 393194 267028
rect 420178 267016 420184 267028
rect 393188 266988 420184 267016
rect 393188 266976 393194 266988
rect 420178 266976 420184 266988
rect 420236 266976 420242 267028
rect 431218 266976 431224 267028
rect 431276 267016 431282 267028
rect 432598 267016 432604 267028
rect 431276 266988 432604 267016
rect 431276 266976 431282 266988
rect 432598 266976 432604 266988
rect 432656 266976 432662 267028
rect 450538 267016 450544 267028
rect 441586 266988 450544 267016
rect 249058 266880 249064 266892
rect 238726 266852 249064 266880
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 286318 266840 286324 266892
rect 286376 266880 286382 266892
rect 287974 266880 287980 266892
rect 286376 266852 287980 266880
rect 286376 266840 286382 266852
rect 287974 266840 287980 266852
rect 288032 266840 288038 266892
rect 313642 266840 313648 266892
rect 313700 266880 313706 266892
rect 317414 266880 317420 266892
rect 313700 266852 317420 266880
rect 313700 266840 313706 266852
rect 317414 266840 317420 266852
rect 317472 266840 317478 266892
rect 321922 266840 321928 266892
rect 321980 266880 321986 266892
rect 327534 266880 327540 266892
rect 321980 266852 327540 266880
rect 321980 266840 321986 266852
rect 327534 266840 327540 266852
rect 327592 266840 327598 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 392302 266840 392308 266892
rect 392360 266880 392366 266892
rect 393958 266880 393964 266892
rect 392360 266852 393964 266880
rect 392360 266840 392366 266852
rect 393958 266840 393964 266852
rect 394016 266840 394022 266892
rect 427906 266840 427912 266892
rect 427964 266880 427970 266892
rect 441586 266880 441614 266988
rect 450538 266976 450544 266988
rect 450596 266976 450602 267028
rect 455046 266976 455052 267028
rect 455104 267016 455110 267028
rect 512638 267016 512644 267028
rect 455104 266988 512644 267016
rect 455104 266976 455110 266988
rect 512638 266976 512644 266988
rect 512696 266976 512702 267028
rect 524782 266976 524788 267028
rect 524840 267016 524846 267028
rect 611998 267016 612004 267028
rect 524840 266988 612004 267016
rect 524840 266976 524846 266988
rect 611998 266976 612004 266988
rect 612056 266976 612062 267028
rect 427964 266852 441614 266880
rect 427964 266840 427970 266852
rect 442718 266840 442724 266892
rect 442776 266880 442782 266892
rect 493318 266880 493324 266892
rect 442776 266852 493324 266880
rect 442776 266840 442782 266852
rect 493318 266840 493324 266852
rect 493376 266840 493382 266892
rect 497458 266840 497464 266892
rect 497516 266880 497522 266892
rect 517698 266880 517704 266892
rect 497516 266852 517704 266880
rect 497516 266840 497522 266852
rect 517698 266840 517704 266852
rect 517756 266840 517762 266892
rect 518986 266840 518992 266892
rect 519044 266880 519050 266892
rect 520090 266880 520096 266892
rect 519044 266852 520096 266880
rect 519044 266840 519050 266852
rect 520090 266840 520096 266852
rect 520148 266840 520154 266892
rect 527266 266840 527272 266892
rect 527324 266880 527330 266892
rect 528186 266880 528192 266892
rect 527324 266852 528192 266880
rect 527324 266840 527330 266852
rect 528186 266840 528192 266852
rect 528244 266840 528250 266892
rect 528922 266840 528928 266892
rect 528980 266880 528986 266892
rect 529842 266880 529848 266892
rect 528980 266852 529848 266880
rect 528980 266840 528986 266852
rect 529842 266840 529848 266852
rect 529900 266840 529906 266892
rect 531406 266840 531412 266892
rect 531464 266880 531470 266892
rect 532510 266880 532516 266892
rect 531464 266852 532516 266880
rect 531464 266840 531470 266852
rect 532510 266840 532516 266852
rect 532568 266840 532574 266892
rect 533062 266840 533068 266892
rect 533120 266880 533126 266892
rect 533982 266880 533988 266892
rect 533120 266852 533988 266880
rect 533120 266840 533126 266852
rect 533982 266840 533988 266852
rect 534040 266840 534046 266892
rect 535546 266840 535552 266892
rect 535604 266880 535610 266892
rect 536742 266880 536748 266892
rect 535604 266852 536748 266880
rect 535604 266840 535610 266852
rect 536742 266840 536748 266852
rect 536800 266840 536806 266892
rect 539686 266840 539692 266892
rect 539744 266880 539750 266892
rect 595438 266880 595444 266892
rect 539744 266852 595444 266880
rect 539744 266840 539750 266852
rect 595438 266840 595444 266852
rect 595496 266840 595502 266892
rect 130378 266704 130384 266756
rect 130436 266744 130442 266756
rect 147214 266744 147220 266756
rect 130436 266716 147220 266744
rect 130436 266704 130442 266716
rect 147214 266704 147220 266716
rect 147272 266704 147278 266756
rect 149698 266704 149704 266756
rect 149756 266744 149762 266756
rect 169570 266744 169576 266756
rect 149756 266716 169576 266744
rect 149756 266704 149762 266716
rect 169570 266704 169576 266716
rect 169628 266704 169634 266756
rect 230750 266704 230756 266756
rect 230808 266744 230814 266756
rect 234154 266744 234160 266756
rect 230808 266716 234160 266744
rect 230808 266704 230814 266716
rect 234154 266704 234160 266716
rect 234212 266704 234218 266756
rect 252002 266704 252008 266756
rect 252060 266744 252066 266756
rect 258994 266744 259000 266756
rect 252060 266716 259000 266744
rect 252060 266704 252066 266716
rect 258994 266704 259000 266716
rect 259052 266704 259058 266756
rect 359642 266704 359648 266756
rect 359700 266744 359706 266756
rect 366358 266744 366364 266756
rect 359700 266716 366364 266744
rect 359700 266704 359706 266716
rect 366358 266704 366364 266716
rect 366416 266704 366422 266756
rect 388162 266704 388168 266756
rect 388220 266744 388226 266756
rect 388220 266716 393314 266744
rect 388220 266704 388226 266716
rect 214558 266636 214564 266688
rect 214616 266676 214622 266688
rect 218422 266676 218428 266688
rect 214616 266648 218428 266676
rect 214616 266636 214622 266648
rect 218422 266636 218428 266648
rect 218480 266636 218486 266688
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310606 266676 310612 266688
rect 308732 266648 310612 266676
rect 308732 266636 308738 266648
rect 310606 266636 310612 266648
rect 310664 266636 310670 266688
rect 312354 266636 312360 266688
rect 312412 266676 312418 266688
rect 314654 266676 314660 266688
rect 312412 266648 314660 266676
rect 312412 266636 312418 266648
rect 314654 266636 314660 266648
rect 314712 266636 314718 266688
rect 316954 266636 316960 266688
rect 317012 266676 317018 266688
rect 321554 266676 321560 266688
rect 317012 266648 321560 266676
rect 317012 266636 317018 266648
rect 321554 266636 321560 266648
rect 321612 266636 321618 266688
rect 342622 266636 342628 266688
rect 342680 266676 342686 266688
rect 347038 266676 347044 266688
rect 342680 266648 347044 266676
rect 342680 266636 342686 266648
rect 347038 266636 347044 266648
rect 347096 266636 347102 266688
rect 137462 266568 137468 266620
rect 137520 266608 137526 266620
rect 145374 266608 145380 266620
rect 137520 266580 145380 266608
rect 137520 266568 137526 266580
rect 145374 266568 145380 266580
rect 145432 266568 145438 266620
rect 145558 266568 145564 266620
rect 145616 266608 145622 266620
rect 148042 266608 148048 266620
rect 145616 266580 148048 266608
rect 145616 266568 145622 266580
rect 148042 266568 148048 266580
rect 148100 266568 148106 266620
rect 226886 266568 226892 266620
rect 226944 266608 226950 266620
rect 231670 266608 231676 266620
rect 226944 266580 231676 266608
rect 226944 266568 226950 266580
rect 231670 266568 231676 266580
rect 231728 266568 231734 266620
rect 393286 266608 393314 266716
rect 397086 266704 397092 266756
rect 397144 266744 397150 266756
rect 407758 266744 407764 266756
rect 397144 266716 407764 266744
rect 397144 266704 397150 266716
rect 407758 266704 407764 266716
rect 407816 266704 407822 266756
rect 428734 266704 428740 266756
rect 428792 266744 428798 266756
rect 442258 266744 442264 266756
rect 428792 266716 442264 266744
rect 428792 266704 428798 266716
rect 442258 266704 442264 266716
rect 442316 266704 442322 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 479518 266744 479524 266756
rect 457772 266716 479524 266744
rect 457772 266704 457778 266716
rect 479518 266704 479524 266716
rect 479576 266704 479582 266756
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 507118 266744 507124 266756
rect 490064 266716 507124 266744
rect 490064 266704 490070 266716
rect 507118 266704 507124 266716
rect 507176 266704 507182 266756
rect 509878 266704 509884 266756
rect 509936 266744 509942 266756
rect 563698 266744 563704 266756
rect 509936 266716 563704 266744
rect 509936 266704 509942 266716
rect 563698 266704 563704 266716
rect 563756 266704 563762 266756
rect 404538 266608 404544 266620
rect 393286 266580 404544 266608
rect 404538 266568 404544 266580
rect 404596 266568 404602 266620
rect 404722 266568 404728 266620
rect 404780 266608 404786 266620
rect 412634 266608 412640 266620
rect 404780 266580 412640 266608
rect 404780 266568 404786 266580
rect 412634 266568 412640 266580
rect 412692 266568 412698 266620
rect 440326 266568 440332 266620
rect 440384 266608 440390 266620
rect 445018 266608 445024 266620
rect 440384 266580 445024 266608
rect 440384 266568 440390 266580
rect 445018 266568 445024 266580
rect 445076 266568 445082 266620
rect 452746 266568 452752 266620
rect 452804 266608 452810 266620
rect 469858 266608 469864 266620
rect 452804 266580 469864 266608
rect 452804 266568 452810 266580
rect 469858 266568 469864 266580
rect 469916 266568 469922 266620
rect 499942 266568 499948 266620
rect 500000 266608 500006 266620
rect 500000 266580 509234 266608
rect 500000 266568 500006 266580
rect 214098 266500 214104 266552
rect 214156 266540 214162 266552
rect 215938 266540 215944 266552
rect 214156 266512 215944 266540
rect 214156 266500 214162 266512
rect 215938 266500 215944 266512
rect 215996 266500 216002 266552
rect 248874 266500 248880 266552
rect 248932 266540 248938 266552
rect 250714 266540 250720 266552
rect 248932 266512 250720 266540
rect 248932 266500 248938 266512
rect 250714 266500 250720 266512
rect 250772 266500 250778 266552
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312814 266500 312820 266552
rect 312872 266540 312878 266552
rect 316034 266540 316040 266552
rect 312872 266512 316040 266540
rect 312872 266500 312878 266512
rect 316034 266500 316040 266512
rect 316092 266500 316098 266552
rect 316402 266500 316408 266552
rect 316460 266540 316466 266552
rect 320174 266540 320180 266552
rect 316460 266512 320180 266540
rect 316460 266500 316466 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 347406 266500 347412 266552
rect 347464 266540 347470 266552
rect 349798 266540 349804 266552
rect 347464 266512 349804 266540
rect 347464 266500 347470 266512
rect 349798 266500 349804 266512
rect 349856 266500 349862 266552
rect 350902 266500 350908 266552
rect 350960 266540 350966 266552
rect 352558 266540 352564 266552
rect 350960 266512 352564 266540
rect 350960 266500 350966 266512
rect 352558 266500 352564 266512
rect 352616 266500 352622 266552
rect 357526 266500 357532 266552
rect 357584 266540 357590 266552
rect 359826 266540 359832 266552
rect 357584 266512 359832 266540
rect 357584 266500 357590 266512
rect 359826 266500 359832 266512
rect 359884 266500 359890 266552
rect 369118 266500 369124 266552
rect 369176 266540 369182 266552
rect 369946 266540 369952 266552
rect 369176 266512 369952 266540
rect 369176 266500 369182 266512
rect 369946 266500 369952 266512
rect 370004 266500 370010 266552
rect 374914 266500 374920 266552
rect 374972 266540 374978 266552
rect 379698 266540 379704 266552
rect 374972 266512 379704 266540
rect 374972 266500 374978 266512
rect 379698 266500 379704 266512
rect 379756 266500 379762 266552
rect 482554 266500 482560 266552
rect 482612 266540 482618 266552
rect 485038 266540 485044 266552
rect 482612 266512 485044 266540
rect 482612 266500 482618 266512
rect 485038 266500 485044 266512
rect 485096 266500 485102 266552
rect 144914 266432 144920 266484
rect 144972 266472 144978 266484
rect 153838 266472 153844 266484
rect 144972 266444 153844 266472
rect 144972 266432 144978 266444
rect 153838 266432 153844 266444
rect 153896 266432 153902 266484
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492582 266472 492588 266484
rect 491720 266444 492588 266472
rect 491720 266432 491726 266444
rect 492582 266432 492588 266444
rect 492640 266432 492646 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495250 266472 495256 266484
rect 494204 266444 495256 266472
rect 494204 266432 494210 266444
rect 495250 266432 495256 266444
rect 495308 266432 495314 266484
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503438 266472 503444 266484
rect 502484 266444 503444 266472
rect 502484 266432 502490 266444
rect 503438 266432 503444 266444
rect 503496 266432 503502 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 509206 266472 509234 266580
rect 510706 266568 510712 266620
rect 510764 266608 510770 266620
rect 511810 266608 511816 266620
rect 510764 266580 511816 266608
rect 510764 266568 510770 266580
rect 511810 266568 511816 266580
rect 511868 266568 511874 266620
rect 516502 266568 516508 266620
rect 516560 266608 516566 266620
rect 517330 266608 517336 266620
rect 516560 266580 517336 266608
rect 516560 266568 516566 266580
rect 517330 266568 517336 266580
rect 517388 266568 517394 266620
rect 517514 266568 517520 266620
rect 517572 266608 517578 266620
rect 556798 266608 556804 266620
rect 517572 266580 556804 266608
rect 517572 266568 517578 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 549898 266472 549904 266484
rect 509206 266444 549904 266472
rect 549898 266432 549904 266444
rect 549956 266432 549962 266484
rect 162118 266364 162124 266416
rect 162176 266404 162182 266416
rect 167086 266404 167092 266416
rect 162176 266376 167092 266404
rect 162176 266364 162182 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 178678 266364 178684 266416
rect 178736 266404 178742 266416
rect 179506 266404 179512 266416
rect 178736 266376 179512 266404
rect 178736 266364 178742 266376
rect 179506 266364 179512 266376
rect 179564 266364 179570 266416
rect 215294 266364 215300 266416
rect 215352 266404 215358 266416
rect 217594 266404 217600 266416
rect 215352 266376 217600 266404
rect 215352 266364 215358 266376
rect 217594 266364 217600 266376
rect 217652 266364 217658 266416
rect 219434 266364 219440 266416
rect 219492 266404 219498 266416
rect 222562 266404 222568 266416
rect 219492 266376 222568 266404
rect 219492 266364 219498 266376
rect 222562 266364 222568 266376
rect 222620 266364 222626 266416
rect 224218 266364 224224 266416
rect 224276 266404 224282 266416
rect 226702 266404 226708 266416
rect 224276 266376 226708 266404
rect 224276 266364 224282 266376
rect 226702 266364 226708 266376
rect 226760 266364 226766 266416
rect 233878 266364 233884 266416
rect 233936 266404 233942 266416
rect 236638 266404 236644 266416
rect 233936 266376 236644 266404
rect 233936 266364 233942 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 239582 266364 239588 266416
rect 239640 266404 239646 266416
rect 246574 266404 246580 266416
rect 239640 266376 246580 266404
rect 239640 266364 239646 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 250438 266364 250444 266416
rect 250496 266404 250502 266416
rect 251542 266404 251548 266416
rect 250496 266376 251548 266404
rect 250496 266364 250502 266376
rect 251542 266364 251548 266376
rect 251600 266364 251606 266416
rect 253382 266364 253388 266416
rect 253440 266404 253446 266416
rect 256510 266404 256516 266416
rect 253440 266376 256516 266404
rect 253440 266364 253446 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 287698 266364 287704 266416
rect 287756 266404 287762 266416
rect 288802 266404 288808 266416
rect 287756 266376 288808 266404
rect 287756 266364 287762 266376
rect 288802 266364 288808 266376
rect 288860 266364 288866 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302050 266404 302056 266416
rect 301004 266376 302056 266404
rect 301004 266364 301010 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310974 266404 310980 266416
rect 309560 266376 310980 266404
rect 309560 266364 309566 266376
rect 310974 266364 310980 266376
rect 311032 266364 311038 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329466 266404 329472 266416
rect 328604 266376 329472 266404
rect 328604 266364 328610 266376
rect 329466 266364 329472 266376
rect 329524 266364 329530 266416
rect 330202 266364 330208 266416
rect 330260 266404 330266 266416
rect 331950 266404 331956 266416
rect 330260 266376 331956 266404
rect 330260 266364 330266 266376
rect 331950 266364 331956 266376
rect 332008 266364 332014 266416
rect 334342 266364 334348 266416
rect 334400 266404 334406 266416
rect 335262 266404 335268 266416
rect 334400 266376 335268 266404
rect 334400 266364 334406 266376
rect 335262 266364 335268 266376
rect 335320 266364 335326 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347590 266404 347596 266416
rect 346820 266376 347596 266404
rect 346820 266364 346826 266376
rect 347590 266364 347596 266376
rect 347648 266364 347654 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 352558 266364 352564 266416
rect 352616 266404 352622 266416
rect 353938 266404 353944 266416
rect 352616 266376 353944 266404
rect 352616 266364 352622 266376
rect 353938 266364 353944 266376
rect 353996 266364 354002 266416
rect 359182 266364 359188 266416
rect 359240 266404 359246 266416
rect 360102 266404 360108 266416
rect 359240 266376 360108 266404
rect 359240 266364 359246 266376
rect 360102 266364 360108 266376
rect 360160 266364 360166 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 368290 266364 368296 266416
rect 368348 266404 368354 266416
rect 369302 266404 369308 266416
rect 368348 266376 369308 266404
rect 368348 266364 368354 266376
rect 369302 266364 369308 266376
rect 369360 266364 369366 266416
rect 369946 266364 369952 266416
rect 370004 266404 370010 266416
rect 372154 266404 372160 266416
rect 370004 266376 372160 266404
rect 370004 266364 370010 266376
rect 372154 266364 372160 266376
rect 372212 266364 372218 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375190 266404 375196 266416
rect 374144 266376 375196 266404
rect 374144 266364 374150 266376
rect 375190 266364 375196 266376
rect 375248 266364 375254 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 381538 266404 381544 266416
rect 379940 266376 381544 266404
rect 379940 266364 379946 266376
rect 381538 266364 381544 266376
rect 381596 266364 381602 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387426 266404 387432 266416
rect 386564 266376 387432 266404
rect 386564 266364 386570 266376
rect 387426 266364 387432 266376
rect 387484 266364 387490 266416
rect 394786 266364 394792 266416
rect 394844 266404 394850 266416
rect 396166 266404 396172 266416
rect 394844 266376 396172 266404
rect 394844 266364 394850 266376
rect 396166 266364 396172 266376
rect 396224 266364 396230 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 403250 266404 403256 266416
rect 400324 266376 403256 266404
rect 400122 266228 400128 266280
rect 400180 266268 400186 266280
rect 400324 266268 400352 266376
rect 403250 266364 403256 266376
rect 403308 266364 403314 266416
rect 407206 266364 407212 266416
rect 407264 266404 407270 266416
rect 408218 266404 408224 266416
rect 407264 266376 408224 266404
rect 407264 266364 407270 266376
rect 408218 266364 408224 266376
rect 408276 266364 408282 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 446122 266364 446128 266416
rect 446180 266404 446186 266416
rect 447778 266404 447784 266416
rect 446180 266376 447784 266404
rect 446180 266364 446186 266376
rect 447778 266364 447784 266376
rect 447836 266364 447842 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455230 266404 455236 266416
rect 454460 266376 455236 266404
rect 454460 266364 454466 266376
rect 455230 266364 455236 266376
rect 455288 266364 455294 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 458082 266404 458088 266416
rect 456944 266376 458088 266404
rect 456944 266364 456950 266376
rect 458082 266364 458088 266376
rect 458140 266364 458146 266416
rect 466822 266364 466828 266416
rect 466880 266404 466886 266416
rect 467742 266404 467748 266416
rect 466880 266376 467748 266404
rect 466880 266364 466886 266376
rect 467742 266364 467748 266376
rect 467800 266364 467806 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474366 266404 474372 266416
rect 473504 266376 474372 266404
rect 473504 266364 473510 266376
rect 474366 266364 474372 266376
rect 474424 266364 474430 266416
rect 477586 266364 477592 266416
rect 477644 266404 477650 266416
rect 478506 266404 478512 266416
rect 477644 266376 478512 266404
rect 477644 266364 477650 266376
rect 478506 266364 478512 266376
rect 478564 266364 478570 266416
rect 481726 266364 481732 266416
rect 481784 266404 481790 266416
rect 482830 266404 482836 266416
rect 481784 266376 482836 266404
rect 481784 266364 481790 266376
rect 482830 266364 482836 266376
rect 482888 266364 482894 266416
rect 483382 266364 483388 266416
rect 483440 266404 483446 266416
rect 484302 266404 484308 266416
rect 483440 266376 484308 266404
rect 483440 266364 483446 266376
rect 484302 266364 484308 266376
rect 484360 266364 484366 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 487062 266404 487068 266416
rect 485924 266376 487068 266404
rect 485924 266364 485930 266376
rect 487062 266364 487068 266376
rect 487120 266364 487126 266416
rect 560478 266336 560484 266348
rect 487264 266308 560484 266336
rect 400180 266240 400352 266268
rect 400180 266228 400186 266240
rect 484210 266228 484216 266280
rect 484268 266268 484274 266280
rect 487264 266268 487292 266308
rect 560478 266296 560484 266308
rect 560536 266296 560542 266348
rect 484268 266240 487292 266268
rect 484268 266228 484274 266240
rect 487522 266160 487528 266212
rect 487580 266200 487586 266212
rect 565814 266200 565820 266212
rect 487580 266172 565820 266200
rect 487580 266160 487586 266172
rect 565814 266160 565820 266172
rect 565872 266160 565878 266212
rect 492490 266024 492496 266076
rect 492548 266064 492554 266076
rect 572714 266064 572720 266076
rect 492548 266036 572720 266064
rect 492548 266024 492554 266036
rect 572714 266024 572720 266036
rect 572772 266024 572778 266076
rect 674466 265956 674472 266008
rect 674524 265996 674530 266008
rect 675478 265996 675484 266008
rect 674524 265968 675484 265996
rect 674524 265956 674530 265968
rect 675478 265956 675484 265968
rect 675536 265956 675542 266008
rect 512362 265888 512368 265940
rect 512420 265928 512426 265940
rect 600314 265928 600320 265940
rect 512420 265900 600320 265928
rect 512420 265888 512426 265900
rect 600314 265888 600320 265900
rect 600372 265888 600378 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 151998 265616 152004 265668
rect 152056 265656 152062 265668
rect 152734 265656 152740 265668
rect 152056 265628 152740 265656
rect 152056 265616 152062 265628
rect 152734 265616 152740 265628
rect 152792 265616 152798 265668
rect 155954 265616 155960 265668
rect 156012 265656 156018 265668
rect 156782 265656 156788 265668
rect 156012 265628 156788 265656
rect 156012 265616 156018 265628
rect 156782 265616 156788 265628
rect 156840 265616 156846 265668
rect 160186 265616 160192 265668
rect 160244 265656 160250 265668
rect 161014 265656 161020 265668
rect 160244 265628 161020 265656
rect 160244 265616 160250 265628
rect 161014 265616 161020 265628
rect 161072 265616 161078 265668
rect 189166 265616 189172 265668
rect 189224 265656 189230 265668
rect 189902 265656 189908 265668
rect 189224 265628 189908 265656
rect 189224 265616 189230 265628
rect 189902 265616 189908 265628
rect 189960 265616 189966 265668
rect 229094 265616 229100 265668
rect 229152 265656 229158 265668
rect 229646 265656 229652 265668
rect 229152 265628 229652 265656
rect 229152 265616 229158 265628
rect 229646 265616 229652 265628
rect 229704 265616 229710 265668
rect 243078 265616 243084 265668
rect 243136 265656 243142 265668
rect 243814 265656 243820 265668
rect 243136 265628 243820 265656
rect 243136 265616 243142 265628
rect 243814 265616 243820 265628
rect 243872 265616 243878 265668
rect 253934 265616 253940 265668
rect 253992 265656 253998 265668
rect 254486 265656 254492 265668
rect 253992 265628 254492 265656
rect 253992 265616 253998 265628
rect 254486 265616 254492 265628
rect 254544 265616 254550 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 520642 265616 520648 265668
rect 520700 265656 520706 265668
rect 612734 265656 612740 265668
rect 520700 265628 612740 265656
rect 520700 265616 520706 265628
rect 612734 265616 612740 265628
rect 612792 265616 612798 265668
rect 480070 265480 480076 265532
rect 480128 265520 480134 265532
rect 554774 265520 554780 265532
rect 480128 265492 554780 265520
rect 480128 265480 480134 265492
rect 554774 265480 554780 265492
rect 554832 265480 554838 265532
rect 479242 265344 479248 265396
rect 479300 265384 479306 265396
rect 553394 265384 553400 265396
rect 479300 265356 553400 265384
rect 479300 265344 479306 265356
rect 553394 265344 553400 265356
rect 553452 265344 553458 265396
rect 475102 265208 475108 265260
rect 475160 265248 475166 265260
rect 547874 265248 547880 265260
rect 475160 265220 547880 265248
rect 475160 265208 475166 265220
rect 547874 265208 547880 265220
rect 547932 265208 547938 265260
rect 469306 265072 469312 265124
rect 469364 265112 469370 265124
rect 539962 265112 539968 265124
rect 469364 265084 539968 265112
rect 469364 265072 469370 265084
rect 539962 265072 539968 265084
rect 540020 265072 540026 265124
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 675846 259564 675852 259616
rect 675904 259604 675910 259616
rect 676214 259604 676220 259616
rect 675904 259576 676220 259604
rect 675904 259564 675910 259576
rect 676214 259564 676220 259576
rect 676272 259564 676278 259616
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 560938 259468 560944 259480
rect 554372 259440 560944 259468
rect 554372 259428 554378 259440
rect 560938 259428 560944 259440
rect 560996 259428 561002 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 563698 256748 563704 256760
rect 554004 256720 563704 256748
rect 554004 256708 554010 256720
rect 563698 256708 563704 256720
rect 563756 256708 563762 256760
rect 553486 255552 553492 255604
rect 553544 255592 553550 255604
rect 555418 255592 555424 255604
rect 553544 255564 555424 255592
rect 553544 255552 553550 255564
rect 555418 255552 555424 255564
rect 555476 255552 555482 255604
rect 35802 255348 35808 255400
rect 35860 255388 35866 255400
rect 39758 255388 39764 255400
rect 35860 255360 39764 255388
rect 35860 255348 35866 255360
rect 39758 255348 39764 255360
rect 39816 255348 39822 255400
rect 675846 254668 675852 254720
rect 675904 254708 675910 254720
rect 683022 254708 683028 254720
rect 675904 254680 683028 254708
rect 675904 254668 675910 254680
rect 683022 254668 683028 254680
rect 683080 254668 683086 254720
rect 35802 254056 35808 254108
rect 35860 254096 35866 254108
rect 39206 254096 39212 254108
rect 35860 254068 39212 254096
rect 35860 254056 35866 254068
rect 39206 254056 39212 254068
rect 39264 254056 39270 254108
rect 675846 253852 675852 253904
rect 675904 253892 675910 253904
rect 680998 253892 681004 253904
rect 675904 253864 681004 253892
rect 675904 253852 675910 253864
rect 680998 253852 681004 253864
rect 681056 253852 681062 253904
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41414 252736 41420 252748
rect 35860 252708 41420 252736
rect 35860 252696 35866 252708
rect 41414 252696 41420 252708
rect 41472 252696 41478 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 40310 252600 40316 252612
rect 35676 252572 40316 252600
rect 35676 252560 35682 252572
rect 40310 252560 40316 252572
rect 40368 252560 40374 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251336 35808 251388
rect 35860 251376 35866 251388
rect 41690 251376 41696 251388
rect 35860 251348 41696 251376
rect 35860 251336 35866 251348
rect 41690 251336 41696 251348
rect 41748 251336 41754 251388
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 35802 249908 35808 249960
rect 35860 249948 35866 249960
rect 39666 249948 39672 249960
rect 35860 249920 39672 249948
rect 35860 249908 35866 249920
rect 39666 249908 39672 249920
rect 39724 249908 39730 249960
rect 35802 248616 35808 248668
rect 35860 248656 35866 248668
rect 41506 248656 41512 248668
rect 35860 248628 41512 248656
rect 35860 248616 35866 248628
rect 41506 248616 41512 248628
rect 41564 248616 41570 248668
rect 674834 248072 674840 248124
rect 674892 248072 674898 248124
rect 674852 247976 674880 248072
rect 675294 247976 675300 247988
rect 674852 247948 675300 247976
rect 675294 247936 675300 247948
rect 675352 247936 675358 247988
rect 35802 247188 35808 247240
rect 35860 247228 35866 247240
rect 41690 247228 41696 247240
rect 35860 247200 41696 247228
rect 35860 247188 35866 247200
rect 41690 247188 41696 247200
rect 41748 247188 41754 247240
rect 35618 247052 35624 247104
rect 35676 247092 35682 247104
rect 39850 247092 39856 247104
rect 35676 247064 39856 247092
rect 35676 247052 35682 247064
rect 39850 247052 39856 247064
rect 39908 247052 39914 247104
rect 558178 246304 558184 246356
rect 558236 246344 558242 246356
rect 647234 246344 647240 246356
rect 558236 246316 647240 246344
rect 558236 246304 558242 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 573358 244304 573364 244316
rect 554556 244276 573364 244304
rect 554556 244264 554562 244276
rect 573358 244264 573364 244276
rect 573416 244264 573422 244316
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 674834 239912 674840 239964
rect 674892 239952 674898 239964
rect 675202 239952 675208 239964
rect 674892 239924 675208 239952
rect 674892 239912 674898 239924
rect 675202 239912 675208 239924
rect 675260 239912 675266 239964
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 668762 237396 668768 237448
rect 668820 237436 668826 237448
rect 671614 237436 671620 237448
rect 668820 237408 671620 237436
rect 668820 237396 668826 237408
rect 671614 237396 671620 237408
rect 671672 237396 671678 237448
rect 672756 236892 672784 237082
rect 672736 236864 672784 236892
rect 672166 236784 672172 236836
rect 672224 236824 672230 236836
rect 672736 236824 672764 236864
rect 672224 236796 672764 236824
rect 672224 236784 672230 236796
rect 672874 236756 672902 236878
rect 672828 236728 672902 236756
rect 671614 236580 671620 236632
rect 671672 236620 671678 236632
rect 672828 236620 672856 236728
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 671672 236592 672856 236620
rect 671672 236580 671678 236592
rect 672966 236456 673118 236484
rect 671798 236376 671804 236428
rect 671856 236416 671862 236428
rect 672966 236416 672994 236456
rect 671856 236388 672994 236416
rect 671856 236376 671862 236388
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 672368 236048 673330 236076
rect 670142 235900 670148 235952
rect 670200 235940 670206 235952
rect 672166 235940 672172 235952
rect 670200 235912 672172 235940
rect 670200 235900 670206 235912
rect 672166 235900 672172 235912
rect 672224 235900 672230 235952
rect 670970 235764 670976 235816
rect 671028 235804 671034 235816
rect 672368 235804 672396 236048
rect 673270 235900 673276 235952
rect 673328 235940 673334 235952
rect 673328 235912 673440 235940
rect 673328 235900 673334 235912
rect 671028 235776 672396 235804
rect 671028 235764 671034 235776
rect 672994 235696 673000 235748
rect 673052 235736 673058 235748
rect 673052 235708 673554 235736
rect 673052 235696 673058 235708
rect 673086 235492 673092 235544
rect 673144 235532 673150 235544
rect 673144 235504 673670 235532
rect 673144 235492 673150 235504
rect 669590 235288 669596 235340
rect 669648 235328 669654 235340
rect 669648 235300 673778 235328
rect 669648 235288 669654 235300
rect 673886 234988 673914 235110
rect 673764 234960 673914 234988
rect 668210 234880 668216 234932
rect 668268 234920 668274 234932
rect 673764 234920 673792 234960
rect 668268 234892 673792 234920
rect 668268 234880 668274 234892
rect 673978 234852 674006 234906
rect 673886 234824 674006 234852
rect 673638 234784 673644 234796
rect 669286 234756 673644 234784
rect 661678 234608 661684 234660
rect 661736 234648 661742 234660
rect 669286 234648 669314 234756
rect 673638 234744 673644 234756
rect 673696 234744 673702 234796
rect 673886 234716 673914 234824
rect 661736 234620 669314 234648
rect 673764 234688 673914 234716
rect 661736 234608 661742 234620
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 668394 234472 668400 234524
rect 668452 234512 668458 234524
rect 673764 234512 673792 234688
rect 674100 234648 674128 234702
rect 674100 234620 674144 234648
rect 674116 234512 674144 234620
rect 668452 234484 673792 234512
rect 673886 234484 674144 234512
rect 668452 234472 668458 234484
rect 671154 234376 671160 234388
rect 670988 234348 671160 234376
rect 670988 234104 671016 234348
rect 671154 234336 671160 234348
rect 671212 234336 671218 234388
rect 671154 234200 671160 234252
rect 671212 234240 671218 234252
rect 673886 234240 673914 234484
rect 674208 234252 674236 234498
rect 671212 234212 673914 234240
rect 671212 234200 671218 234212
rect 674190 234200 674196 234252
rect 674248 234200 674254 234252
rect 675110 234104 675116 234116
rect 670988 234076 675116 234104
rect 675110 234064 675116 234076
rect 675168 234064 675174 234116
rect 683390 234036 683396 234048
rect 678946 234008 683396 234036
rect 675846 233928 675852 233980
rect 675904 233968 675910 233980
rect 678946 233968 678974 234008
rect 683390 233996 683396 234008
rect 683448 233996 683454 234048
rect 675904 233940 678974 233968
rect 675904 233928 675910 233940
rect 652202 233860 652208 233912
rect 652260 233900 652266 233912
rect 672166 233900 672172 233912
rect 652260 233872 672172 233900
rect 652260 233860 652266 233872
rect 672166 233860 672172 233872
rect 672224 233860 672230 233912
rect 675846 233724 675852 233776
rect 675904 233764 675910 233776
rect 678238 233764 678244 233776
rect 675904 233736 678244 233764
rect 675904 233724 675910 233736
rect 678238 233724 678244 233736
rect 678296 233724 678302 233776
rect 672258 233248 672264 233300
rect 672316 233288 672322 233300
rect 673086 233288 673092 233300
rect 672316 233260 673092 233288
rect 672316 233248 672322 233260
rect 673086 233248 673092 233260
rect 673144 233248 673150 233300
rect 670326 233044 670332 233096
rect 670384 233084 670390 233096
rect 672994 233084 673000 233096
rect 670384 233056 673000 233084
rect 670384 233044 670390 233056
rect 672994 233044 673000 233056
rect 673052 233044 673058 233096
rect 669406 232908 669412 232960
rect 669464 232948 669470 232960
rect 674190 232948 674196 232960
rect 669464 232920 674196 232948
rect 669464 232908 669470 232920
rect 674190 232908 674196 232920
rect 674248 232908 674254 232960
rect 639598 232500 639604 232552
rect 639656 232540 639662 232552
rect 654778 232540 654784 232552
rect 639656 232512 654784 232540
rect 639656 232500 639662 232512
rect 654778 232500 654784 232512
rect 654836 232500 654842 232552
rect 660298 232500 660304 232552
rect 660356 232540 660362 232552
rect 660356 232512 663794 232540
rect 660356 232500 660362 232512
rect 663766 232472 663794 232512
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 683206 232540 683212 232552
rect 675904 232512 683212 232540
rect 675904 232500 675910 232512
rect 683206 232500 683212 232512
rect 683264 232500 683270 232552
rect 670786 232472 670792 232484
rect 663766 232444 670792 232472
rect 670786 232432 670792 232444
rect 670844 232432 670850 232484
rect 665450 231616 665456 231668
rect 665508 231656 665514 231668
rect 674926 231656 674932 231668
rect 665508 231628 674932 231656
rect 665508 231616 665514 231628
rect 674926 231616 674932 231628
rect 674984 231616 674990 231668
rect 146202 231548 146208 231600
rect 146260 231588 146266 231600
rect 150526 231588 150532 231600
rect 146260 231560 150532 231588
rect 146260 231548 146266 231560
rect 150526 231548 150532 231560
rect 150584 231548 150590 231600
rect 155494 231548 155500 231600
rect 155552 231588 155558 231600
rect 156966 231588 156972 231600
rect 155552 231560 156972 231588
rect 155552 231548 155558 231560
rect 156966 231548 156972 231560
rect 157024 231548 157030 231600
rect 663058 231480 663064 231532
rect 663116 231520 663122 231532
rect 670786 231520 670792 231532
rect 663116 231492 670792 231520
rect 663116 231480 663122 231492
rect 670786 231480 670792 231492
rect 670844 231480 670850 231532
rect 675846 231480 675852 231532
rect 675904 231520 675910 231532
rect 683574 231520 683580 231532
rect 675904 231492 683580 231520
rect 675904 231480 675910 231492
rect 683574 231480 683580 231492
rect 683632 231480 683638 231532
rect 146754 231412 146760 231464
rect 146812 231452 146818 231464
rect 147214 231452 147220 231464
rect 146812 231424 147220 231452
rect 146812 231412 146818 231424
rect 147214 231412 147220 231424
rect 147272 231412 147278 231464
rect 156598 231412 156604 231464
rect 156656 231452 156662 231464
rect 163682 231452 163688 231464
rect 156656 231424 163688 231452
rect 156656 231412 156662 231424
rect 163682 231412 163688 231424
rect 163740 231412 163746 231464
rect 662322 231344 662328 231396
rect 662380 231384 662386 231396
rect 675110 231384 675116 231396
rect 662380 231356 675116 231384
rect 662380 231344 662386 231356
rect 675110 231344 675116 231356
rect 675168 231344 675174 231396
rect 137922 231276 137928 231328
rect 137980 231316 137986 231328
rect 152458 231316 152464 231328
rect 137980 231288 152464 231316
rect 137980 231276 137986 231288
rect 152458 231276 152464 231288
rect 152516 231276 152522 231328
rect 155770 231276 155776 231328
rect 155828 231316 155834 231328
rect 161750 231316 161756 231328
rect 155828 231288 161756 231316
rect 155828 231276 155834 231288
rect 161750 231276 161756 231288
rect 161808 231276 161814 231328
rect 91738 231140 91744 231192
rect 91796 231180 91802 231192
rect 168834 231180 168840 231192
rect 91796 231152 168840 231180
rect 91796 231140 91802 231152
rect 168834 231140 168840 231152
rect 168892 231140 168898 231192
rect 664990 231140 664996 231192
rect 665048 231180 665054 231192
rect 665048 231152 675326 231180
rect 665048 231140 665054 231152
rect 596818 231072 596824 231124
rect 596876 231112 596882 231124
rect 633618 231112 633624 231124
rect 596876 231084 633624 231112
rect 596876 231072 596882 231084
rect 633618 231072 633624 231084
rect 633676 231072 633682 231124
rect 636838 231072 636844 231124
rect 636896 231112 636902 231124
rect 650638 231112 650644 231124
rect 636896 231084 650644 231112
rect 636896 231072 636902 231084
rect 650638 231072 650644 231084
rect 650696 231072 650702 231124
rect 675116 231056 675168 231062
rect 128262 231004 128268 231056
rect 128320 231044 128326 231056
rect 195882 231044 195888 231056
rect 128320 231016 195888 231044
rect 128320 231004 128326 231016
rect 195882 231004 195888 231016
rect 195940 231004 195946 231056
rect 675116 230998 675168 231004
rect 97902 230868 97908 230920
rect 97960 230908 97966 230920
rect 173986 230908 173992 230920
rect 97960 230880 173992 230908
rect 97960 230868 97966 230880
rect 173986 230868 173992 230880
rect 174044 230868 174050 230920
rect 674956 230852 675008 230858
rect 674956 230794 675008 230800
rect 110322 230732 110328 230784
rect 110380 230772 110386 230784
rect 184290 230772 184296 230784
rect 110380 230744 184296 230772
rect 110380 230732 110386 230744
rect 184290 230732 184296 230744
rect 184348 230732 184354 230784
rect 118602 230596 118608 230648
rect 118660 230636 118666 230648
rect 188154 230636 188160 230648
rect 118660 230608 188160 230636
rect 118660 230596 118666 230608
rect 188154 230596 188160 230608
rect 188212 230596 188218 230648
rect 195054 230596 195060 230648
rect 195112 230636 195118 230648
rect 196894 230636 196900 230648
rect 195112 230608 196900 230636
rect 195112 230596 195118 230608
rect 196894 230596 196900 230608
rect 196952 230596 196958 230648
rect 672166 230596 672172 230648
rect 672224 230636 672230 230648
rect 672224 230608 674820 230636
rect 672224 230596 672230 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 152458 230460 152464 230512
rect 152516 230500 152522 230512
rect 203610 230500 203616 230512
rect 152516 230472 203616 230500
rect 152516 230460 152522 230472
rect 203610 230460 203616 230472
rect 203668 230460 203674 230512
rect 42426 230392 42432 230444
rect 42484 230432 42490 230444
rect 43162 230432 43168 230444
rect 42484 230404 43168 230432
rect 42484 230392 42490 230404
rect 43162 230392 43168 230404
rect 43220 230392 43226 230444
rect 130378 230392 130384 230444
rect 130436 230432 130442 230444
rect 142430 230432 142436 230444
rect 130436 230404 142436 230432
rect 130436 230392 130442 230404
rect 142430 230392 142436 230404
rect 142488 230392 142494 230444
rect 142614 230392 142620 230444
rect 142672 230432 142678 230444
rect 146202 230432 146208 230444
rect 142672 230404 146208 230432
rect 142672 230392 142678 230404
rect 146202 230392 146208 230404
rect 146260 230392 146266 230444
rect 147628 230392 147634 230444
rect 147686 230432 147692 230444
rect 149514 230432 149520 230444
rect 147686 230404 149520 230432
rect 147686 230392 147692 230404
rect 149514 230392 149520 230404
rect 149572 230392 149578 230444
rect 206278 230392 206284 230444
rect 206336 230432 206342 230444
rect 256418 230432 256424 230444
rect 206336 230404 256424 230432
rect 206336 230392 206342 230404
rect 256418 230392 256424 230404
rect 256476 230392 256482 230444
rect 287054 230392 287060 230444
rect 287112 230432 287118 230444
rect 307938 230432 307944 230444
rect 287112 230404 307944 230432
rect 287112 230392 287118 230404
rect 307938 230392 307944 230404
rect 307996 230392 308002 230444
rect 308398 230392 308404 230444
rect 308456 230432 308462 230444
rect 334986 230432 334992 230444
rect 308456 230404 334992 230432
rect 308456 230392 308462 230404
rect 334986 230392 334992 230404
rect 335044 230392 335050 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 444466 230392 444472 230444
rect 444524 230432 444530 230444
rect 447594 230432 447600 230444
rect 444524 230404 447600 230432
rect 444524 230392 444530 230404
rect 447594 230392 447600 230404
rect 447652 230392 447658 230444
rect 526898 230392 526904 230444
rect 526956 230432 526962 230444
rect 536098 230432 536104 230444
rect 526956 230404 536104 230432
rect 526956 230392 526962 230404
rect 536098 230392 536104 230404
rect 536156 230392 536162 230444
rect 673454 230392 673460 230444
rect 673512 230432 673518 230444
rect 673512 230404 674702 230432
rect 673512 230392 673518 230404
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 487614 230324 487620 230376
rect 487672 230364 487678 230376
rect 488442 230364 488448 230376
rect 487672 230336 488448 230364
rect 487672 230324 487678 230336
rect 488442 230324 488448 230336
rect 488500 230324 488506 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 511442 230324 511448 230376
rect 511500 230364 511506 230376
rect 517514 230364 517520 230376
rect 511500 230336 517520 230364
rect 511500 230324 511506 230336
rect 517514 230324 517520 230336
rect 517572 230324 517578 230376
rect 133782 230256 133788 230308
rect 133840 230296 133846 230308
rect 202322 230296 202328 230308
rect 133840 230268 202328 230296
rect 133840 230256 133846 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 210418 230256 210424 230308
rect 210476 230296 210482 230308
rect 261570 230296 261576 230308
rect 210476 230268 261576 230296
rect 210476 230256 210482 230268
rect 261570 230256 261576 230268
rect 261628 230256 261634 230308
rect 275646 230256 275652 230308
rect 275704 230296 275710 230308
rect 313090 230296 313096 230308
rect 275704 230268 313096 230296
rect 275704 230256 275710 230268
rect 313090 230256 313096 230268
rect 313148 230256 313154 230308
rect 436094 230256 436100 230308
rect 436152 230296 436158 230308
rect 436830 230296 436836 230308
rect 436152 230268 436836 230296
rect 436152 230256 436158 230268
rect 436830 230256 436836 230268
rect 436888 230256 436894 230308
rect 528830 230256 528836 230308
rect 528888 230296 528894 230308
rect 539594 230296 539600 230308
rect 528888 230268 539600 230296
rect 528888 230256 528894 230268
rect 539594 230256 539600 230268
rect 539652 230256 539658 230308
rect 388438 230188 388444 230240
rect 388496 230228 388502 230240
rect 391658 230228 391664 230240
rect 388496 230200 391664 230228
rect 388496 230188 388502 230200
rect 391658 230188 391664 230200
rect 391716 230188 391722 230240
rect 443822 230188 443828 230240
rect 443880 230228 443886 230240
rect 444650 230228 444656 230240
rect 443880 230200 444656 230228
rect 443880 230188 443886 230200
rect 444650 230188 444656 230200
rect 444708 230188 444714 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 453482 230188 453488 230240
rect 453540 230228 453546 230240
rect 455782 230228 455788 230240
rect 453540 230200 455788 230228
rect 453540 230188 453546 230200
rect 455782 230188 455788 230200
rect 455840 230188 455846 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 674374 230188 674380 230240
rect 674432 230228 674438 230240
rect 674432 230200 674590 230228
rect 674432 230188 674438 230200
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 157288 230160 157294 230172
rect 95292 230132 157294 230160
rect 95292 230120 95298 230132
rect 157288 230120 157294 230132
rect 157346 230120 157352 230172
rect 157426 230120 157432 230172
rect 157484 230160 157490 230172
rect 161106 230160 161112 230172
rect 157484 230132 161112 230160
rect 157484 230120 157490 230132
rect 161106 230120 161112 230132
rect 161164 230120 161170 230172
rect 176746 230120 176752 230172
rect 176804 230160 176810 230172
rect 235810 230160 235816 230172
rect 176804 230132 235816 230160
rect 176804 230120 176810 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 264238 230120 264244 230172
rect 264296 230160 264302 230172
rect 302786 230160 302792 230172
rect 264296 230132 302792 230160
rect 264296 230120 264302 230132
rect 302786 230120 302792 230132
rect 302844 230120 302850 230172
rect 312630 230120 312636 230172
rect 312688 230160 312694 230172
rect 340138 230160 340144 230172
rect 312688 230132 340144 230160
rect 312688 230120 312694 230132
rect 340138 230120 340144 230132
rect 340196 230120 340202 230172
rect 521102 230120 521108 230172
rect 521160 230160 521166 230172
rect 529198 230160 529204 230172
rect 521160 230132 529204 230160
rect 521160 230120 521166 230132
rect 529198 230120 529204 230132
rect 529256 230120 529262 230172
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 126882 229984 126888 230036
rect 126940 230024 126946 230036
rect 195054 230024 195060 230036
rect 126940 229996 195060 230024
rect 126940 229984 126946 229996
rect 195054 229984 195060 229996
rect 195112 229984 195118 230036
rect 195422 229984 195428 230036
rect 195480 230024 195486 230036
rect 214742 230024 214748 230036
rect 195480 229996 214748 230024
rect 195480 229984 195486 229996
rect 214742 229984 214748 229996
rect 214800 229984 214806 230036
rect 220078 229984 220084 230036
rect 220136 230024 220142 230036
rect 230658 230024 230664 230036
rect 220136 229996 230664 230024
rect 220136 229984 220142 229996
rect 230658 229984 230664 229996
rect 230716 229984 230722 230036
rect 242526 229984 242532 230036
rect 242584 230024 242590 230036
rect 287330 230024 287336 230036
rect 242584 229996 287336 230024
rect 242584 229984 242590 229996
rect 287330 229984 287336 229996
rect 287388 229984 287394 230036
rect 302878 229984 302884 230036
rect 302936 230024 302942 230036
rect 329834 230024 329840 230036
rect 302936 229996 329840 230024
rect 302936 229984 302942 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 334250 229984 334256 230036
rect 334308 230024 334314 230036
rect 355594 230024 355600 230036
rect 334308 229996 355600 230024
rect 334308 229984 334314 229996
rect 355594 229984 355600 229996
rect 355652 229984 355658 230036
rect 355778 229984 355784 230036
rect 355836 230024 355842 230036
rect 371050 230024 371056 230036
rect 355836 229996 371056 230024
rect 355836 229984 355842 229996
rect 371050 229984 371056 229996
rect 371108 229984 371114 230036
rect 457346 229984 457352 230036
rect 457404 230024 457410 230036
rect 463878 230024 463884 230036
rect 457404 229996 463884 230024
rect 457404 229984 457410 229996
rect 463878 229984 463884 229996
rect 463936 229984 463942 230036
rect 476666 229984 476672 230036
rect 476724 230024 476730 230036
rect 481634 230024 481640 230036
rect 476724 229996 481640 230024
rect 476724 229984 476730 229996
rect 481634 229984 481640 229996
rect 481692 229984 481698 230036
rect 517238 229984 517244 230036
rect 517296 230024 517302 230036
rect 526438 230024 526444 230036
rect 517296 229996 526444 230024
rect 517296 229984 517302 229996
rect 526438 229984 526444 229996
rect 526496 229984 526502 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 549254 230024 549260 230036
rect 534684 229996 549260 230024
rect 534684 229984 534690 229996
rect 549254 229984 549260 229996
rect 549312 229984 549318 230036
rect 674190 229984 674196 230036
rect 674248 229984 674254 230036
rect 86218 229848 86224 229900
rect 86276 229888 86282 229900
rect 156782 229888 156788 229900
rect 86276 229860 156788 229888
rect 86276 229848 86282 229860
rect 156782 229848 156788 229860
rect 156840 229848 156846 229900
rect 158530 229888 158536 229900
rect 157168 229860 158536 229888
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 142614 229752 142620 229764
rect 68336 229724 142620 229752
rect 68336 229712 68342 229724
rect 142614 229712 142620 229724
rect 142672 229712 142678 229764
rect 147766 229752 147772 229764
rect 147646 229724 147772 229752
rect 147646 229684 147674 229724
rect 147766 229712 147772 229724
rect 147824 229712 147830 229764
rect 157168 229752 157196 229860
rect 158530 229848 158536 229860
rect 158588 229848 158594 229900
rect 163958 229848 163964 229900
rect 164016 229888 164022 229900
rect 225506 229888 225512 229900
rect 164016 229860 225512 229888
rect 164016 229848 164022 229860
rect 225506 229848 225512 229860
rect 225564 229848 225570 229900
rect 230474 229848 230480 229900
rect 230532 229888 230538 229900
rect 277026 229888 277032 229900
rect 230532 229860 277032 229888
rect 230532 229848 230538 229860
rect 277026 229848 277032 229860
rect 277084 229848 277090 229900
rect 282546 229848 282552 229900
rect 282604 229888 282610 229900
rect 318242 229888 318248 229900
rect 282604 229860 318248 229888
rect 282604 229848 282610 229860
rect 318242 229848 318248 229860
rect 318300 229848 318306 229900
rect 324222 229848 324228 229900
rect 324280 229888 324286 229900
rect 350442 229888 350448 229900
rect 324280 229860 350448 229888
rect 324280 229848 324286 229860
rect 350442 229848 350448 229860
rect 350500 229848 350506 229900
rect 366726 229848 366732 229900
rect 366784 229888 366790 229900
rect 383930 229888 383936 229900
rect 366784 229860 383936 229888
rect 366784 229848 366790 229860
rect 383930 229848 383936 229860
rect 383988 229848 383994 229900
rect 449618 229848 449624 229900
rect 449676 229888 449682 229900
rect 450538 229888 450544 229900
rect 449676 229860 450544 229888
rect 449676 229848 449682 229860
rect 450538 229848 450544 229860
rect 450596 229848 450602 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 479242 229848 479248 229900
rect 479300 229888 479306 229900
rect 488074 229888 488080 229900
rect 479300 229860 488080 229888
rect 479300 229848 479306 229860
rect 488074 229848 488080 229860
rect 488132 229848 488138 229900
rect 492122 229848 492128 229900
rect 492180 229888 492186 229900
rect 492180 229860 495848 229888
rect 492180 229848 492186 229860
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 476022 229780 476028 229832
rect 476080 229820 476086 229832
rect 478598 229820 478604 229832
rect 476080 229792 478604 229820
rect 476080 229780 476086 229792
rect 478598 229780 478604 229792
rect 478656 229780 478662 229832
rect 147968 229724 157196 229752
rect 142816 229656 147674 229684
rect 82078 229576 82084 229628
rect 82136 229616 82142 229628
rect 142816 229616 142844 229656
rect 82136 229588 142844 229616
rect 82136 229576 82142 229588
rect 147122 229508 147128 229560
rect 147180 229548 147186 229560
rect 147968 229548 147996 229724
rect 171042 229712 171048 229764
rect 171100 229752 171106 229764
rect 220078 229752 220084 229764
rect 171100 229724 220084 229752
rect 171100 229712 171106 229724
rect 220078 229712 220084 229724
rect 220136 229712 220142 229764
rect 246114 229752 246120 229764
rect 224926 229724 246120 229752
rect 148134 229576 148140 229628
rect 148192 229616 148198 229628
rect 155954 229616 155960 229628
rect 148192 229588 155960 229616
rect 148192 229576 148198 229588
rect 155954 229576 155960 229588
rect 156012 229576 156018 229628
rect 157334 229576 157340 229628
rect 157392 229616 157398 229628
rect 157392 229588 214604 229616
rect 157392 229576 157398 229588
rect 147180 229520 147996 229548
rect 156800 229520 157012 229548
rect 147180 229508 147186 229520
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 143994 229480 144000 229492
rect 102192 229452 144000 229480
rect 102192 229440 102198 229452
rect 143994 229440 144000 229452
rect 144052 229440 144058 229492
rect 144178 229440 144184 229492
rect 144236 229480 144242 229492
rect 146938 229480 146944 229492
rect 144236 229452 146944 229480
rect 144236 229440 144242 229452
rect 146938 229440 146944 229452
rect 146996 229440 147002 229492
rect 156800 229480 156828 229520
rect 148060 229452 156828 229480
rect 156984 229480 157012 229520
rect 210050 229480 210056 229492
rect 156984 229452 210056 229480
rect 111058 229304 111064 229356
rect 111116 229344 111122 229356
rect 147582 229344 147588 229356
rect 111116 229316 147588 229344
rect 111116 229304 111122 229316
rect 147582 229304 147588 229316
rect 147640 229304 147646 229356
rect 147766 229304 147772 229356
rect 147824 229344 147830 229356
rect 148060 229344 148088 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 214576 229480 214604 229588
rect 214742 229576 214748 229628
rect 214800 229616 214806 229628
rect 224926 229616 224954 229724
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 256510 229712 256516 229764
rect 256568 229752 256574 229764
rect 297634 229752 297640 229764
rect 256568 229724 297640 229752
rect 256568 229712 256574 229724
rect 297634 229712 297640 229724
rect 297692 229712 297698 229764
rect 318058 229712 318064 229764
rect 318116 229752 318122 229764
rect 318116 229724 335354 229752
rect 318116 229712 318122 229724
rect 266722 229616 266728 229628
rect 214800 229588 224954 229616
rect 229066 229588 266728 229616
rect 214800 229576 214806 229588
rect 220354 229480 220360 229492
rect 214576 229452 220360 229480
rect 220354 229440 220360 229452
rect 220412 229440 220418 229492
rect 220630 229440 220636 229492
rect 220688 229480 220694 229492
rect 229066 229480 229094 229588
rect 266722 229576 266728 229588
rect 266780 229576 266786 229628
rect 276290 229576 276296 229628
rect 276348 229616 276354 229628
rect 292482 229616 292488 229628
rect 276348 229588 292488 229616
rect 276348 229576 276354 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 296990 229576 296996 229628
rect 297048 229616 297054 229628
rect 323394 229616 323400 229628
rect 297048 229588 323400 229616
rect 297048 229576 297054 229588
rect 323394 229576 323400 229588
rect 323452 229576 323458 229628
rect 335326 229616 335354 229724
rect 345014 229712 345020 229764
rect 345072 229752 345078 229764
rect 360746 229752 360752 229764
rect 345072 229724 360752 229752
rect 345072 229712 345078 229724
rect 360746 229712 360752 229724
rect 360804 229712 360810 229764
rect 361206 229712 361212 229764
rect 361264 229752 361270 229764
rect 378778 229752 378784 229764
rect 361264 229724 378784 229752
rect 361264 229712 361270 229724
rect 378778 229712 378784 229724
rect 378836 229712 378842 229764
rect 391198 229712 391204 229764
rect 391256 229752 391262 229764
rect 398742 229752 398748 229764
rect 391256 229724 398748 229752
rect 391256 229712 391262 229724
rect 398742 229712 398748 229724
rect 398800 229712 398806 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 410886 229712 410892 229764
rect 410944 229752 410950 229764
rect 417418 229752 417424 229764
rect 410944 229724 417424 229752
rect 410944 229712 410950 229724
rect 417418 229712 417424 229724
rect 417476 229712 417482 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 469640 229724 470594 229752
rect 469640 229712 469646 229724
rect 470566 229684 470594 229724
rect 481818 229712 481824 229764
rect 481876 229752 481882 229764
rect 489914 229752 489920 229764
rect 481876 229724 489920 229752
rect 481876 229712 481882 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 490190 229712 490196 229764
rect 490248 229752 490254 229764
rect 493594 229752 493600 229764
rect 490248 229724 493600 229752
rect 490248 229712 490254 229724
rect 493594 229712 493600 229724
rect 493652 229712 493658 229764
rect 495820 229752 495848 229860
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 507118 229888 507124 229900
rect 496044 229860 507124 229888
rect 496044 229848 496050 229860
rect 507118 229848 507124 229860
rect 507176 229848 507182 229900
rect 510798 229848 510804 229900
rect 510856 229888 510862 229900
rect 511902 229888 511908 229900
rect 510856 229860 511908 229888
rect 510856 229848 510862 229860
rect 511902 229848 511908 229860
rect 511960 229848 511966 229900
rect 515306 229848 515312 229900
rect 515364 229888 515370 229900
rect 525702 229888 525708 229900
rect 515364 229860 525708 229888
rect 515364 229848 515370 229860
rect 525702 229848 525708 229860
rect 525760 229848 525766 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 674208 229888 674236 229984
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674116 229860 674236 229888
rect 505186 229752 505192 229764
rect 495820 229724 505192 229752
rect 505186 229712 505192 229724
rect 505244 229712 505250 229764
rect 507578 229712 507584 229764
rect 507636 229752 507642 229764
rect 516778 229752 516784 229764
rect 507636 229724 516784 229752
rect 507636 229712 507642 229724
rect 516778 229712 516784 229724
rect 516836 229712 516842 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534810 229752 534816 229764
rect 523092 229724 534816 229752
rect 523092 229712 523098 229724
rect 534810 229712 534816 229724
rect 534868 229712 534874 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566458 229752 566464 229764
rect 538548 229724 566464 229752
rect 538548 229712 538554 229724
rect 566458 229712 566464 229724
rect 566516 229712 566522 229764
rect 476758 229684 476764 229696
rect 470566 229656 476764 229684
rect 476758 229644 476764 229656
rect 476816 229644 476822 229696
rect 345290 229616 345296 229628
rect 335326 229588 345296 229616
rect 345290 229576 345296 229588
rect 345348 229576 345354 229628
rect 509510 229576 509516 229628
rect 509568 229616 509574 229628
rect 515398 229616 515404 229628
rect 509568 229588 515404 229616
rect 509568 229576 509574 229588
rect 515398 229576 515404 229588
rect 515456 229576 515462 229628
rect 530118 229576 530124 229628
rect 530176 229616 530182 229628
rect 531130 229616 531136 229628
rect 530176 229588 531136 229616
rect 530176 229576 530182 229588
rect 531130 229576 531136 229588
rect 531188 229576 531194 229628
rect 538306 229616 538312 229628
rect 538186 229588 538312 229616
rect 384298 229508 384304 229560
rect 384356 229548 384362 229560
rect 389082 229548 389088 229560
rect 384356 229520 389088 229548
rect 384356 229508 384362 229520
rect 389082 229508 389088 229520
rect 389140 229508 389146 229560
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451366 229548 451372 229560
rect 449032 229520 451372 229548
rect 449032 229508 449038 229520
rect 451366 229508 451372 229520
rect 451424 229508 451430 229560
rect 220688 229452 229094 229480
rect 220688 229440 220694 229452
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 271874 229480 271880 229492
rect 231176 229452 271880 229480
rect 231176 229440 231182 229452
rect 271874 229440 271880 229452
rect 271932 229440 271938 229492
rect 530762 229440 530768 229492
rect 530820 229480 530826 229492
rect 538186 229480 538214 229588
rect 538306 229576 538312 229588
rect 538364 229576 538370 229628
rect 674116 229616 674144 229860
rect 674334 229764 674386 229770
rect 674334 229706 674386 229712
rect 674116 229588 674268 229616
rect 530820 229452 538214 229480
rect 530820 229440 530826 229452
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448790 229412 448796 229424
rect 446456 229384 448796 229412
rect 446456 229372 446462 229384
rect 448790 229372 448796 229384
rect 448848 229372 448854 229424
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 453022 229412 453028 229424
rect 450964 229384 453028 229412
rect 450964 229372 450970 229384
rect 453022 229372 453028 229384
rect 453080 229372 453086 229424
rect 673178 229372 673184 229424
rect 673236 229412 673242 229424
rect 673236 229384 674130 229412
rect 673236 229372 673242 229384
rect 147824 229316 148088 229344
rect 147824 229304 147830 229316
rect 151170 229304 151176 229356
rect 151228 229344 151234 229356
rect 151228 229316 153608 229344
rect 151228 229304 151234 229316
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 153378 229208 153384 229220
rect 123536 229180 153384 229208
rect 123536 229168 123542 229180
rect 153378 229168 153384 229180
rect 153436 229168 153442 229220
rect 153580 229208 153608 229316
rect 153838 229304 153844 229356
rect 153896 229344 153902 229356
rect 156598 229344 156604 229356
rect 153896 229316 156604 229344
rect 153896 229304 153902 229316
rect 156598 229304 156604 229316
rect 156656 229304 156662 229356
rect 159358 229304 159364 229356
rect 159416 229344 159422 229356
rect 215202 229344 215208 229356
rect 159416 229316 215208 229344
rect 159416 229304 159422 229316
rect 215202 229304 215208 229316
rect 215260 229304 215266 229356
rect 246482 229304 246488 229356
rect 246540 229344 246546 229356
rect 282178 229344 282184 229356
rect 246540 229316 282184 229344
rect 246540 229304 246546 229316
rect 282178 229304 282184 229316
rect 282236 229304 282242 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 472158 229304 472164 229356
rect 472216 229344 472222 229356
rect 472986 229344 472992 229356
rect 472216 229316 472992 229344
rect 472216 229304 472222 229316
rect 472986 229304 472992 229316
rect 473044 229304 473050 229356
rect 488258 229304 488264 229356
rect 488316 229344 488322 229356
rect 490374 229344 490380 229356
rect 488316 229316 490380 229344
rect 488316 229304 488322 229316
rect 490374 229304 490380 229316
rect 490432 229304 490438 229356
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451826 229276 451832 229288
rect 450320 229248 451832 229276
rect 450320 229236 450326 229248
rect 451826 229236 451832 229248
rect 451884 229236 451890 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 505646 229236 505652 229288
rect 505704 229276 505710 229288
rect 510614 229276 510620 229288
rect 505704 229248 510620 229276
rect 505704 229236 505710 229248
rect 510614 229236 510620 229248
rect 510672 229236 510678 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519354 229276 519360 229288
rect 513432 229248 519360 229276
rect 513432 229236 513438 229248
rect 519354 229236 519360 229248
rect 519412 229236 519418 229288
rect 155770 229208 155776 229220
rect 153580 229180 155776 229208
rect 155770 229168 155776 229180
rect 155828 229168 155834 229220
rect 157610 229168 157616 229220
rect 157668 229208 157674 229220
rect 166258 229208 166264 229220
rect 157668 229180 166264 229208
rect 157668 229168 157674 229180
rect 166258 229168 166264 229180
rect 166316 229168 166322 229220
rect 167362 229168 167368 229220
rect 167420 229208 167426 229220
rect 174262 229208 174268 229220
rect 167420 229180 174268 229208
rect 167420 229168 167426 229180
rect 174262 229168 174268 229180
rect 174320 229168 174326 229220
rect 184658 229168 184664 229220
rect 184716 229208 184722 229220
rect 240962 229208 240968 229220
rect 184716 229180 240968 229208
rect 184716 229168 184722 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 166920 229112 167132 229140
rect 100662 229032 100668 229084
rect 100720 229072 100726 229084
rect 100720 229044 103514 229072
rect 100720 229032 100726 229044
rect 103486 228936 103514 229044
rect 106182 229032 106188 229084
rect 106240 229072 106246 229084
rect 142982 229072 142988 229084
rect 106240 229044 142988 229072
rect 106240 229032 106246 229044
rect 142982 229032 142988 229044
rect 143040 229032 143046 229084
rect 143442 229032 143448 229084
rect 143500 229072 143506 229084
rect 146202 229072 146208 229084
rect 143500 229044 146208 229072
rect 143500 229032 143506 229044
rect 146202 229032 146208 229044
rect 146260 229032 146266 229084
rect 146386 229032 146392 229084
rect 146444 229072 146450 229084
rect 156874 229072 156880 229084
rect 146444 229044 156880 229072
rect 146444 229032 146450 229044
rect 156874 229032 156880 229044
rect 156932 229032 156938 229084
rect 157518 229032 157524 229084
rect 157576 229072 157582 229084
rect 166920 229072 166948 229112
rect 157576 229044 166948 229072
rect 167104 229072 167132 229112
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 519170 229100 519176 229152
rect 519228 229140 519234 229152
rect 519228 229112 521654 229140
rect 519228 229100 519234 229112
rect 202874 229072 202880 229084
rect 167104 229044 202880 229072
rect 157576 229032 157582 229044
rect 202874 229032 202880 229044
rect 202932 229032 202938 229084
rect 204714 229032 204720 229084
rect 204772 229072 204778 229084
rect 212350 229072 212356 229084
rect 204772 229044 212356 229072
rect 204772 229032 204778 229044
rect 212350 229032 212356 229044
rect 212408 229032 212414 229084
rect 213914 229032 213920 229084
rect 213972 229072 213978 229084
rect 214558 229072 214564 229084
rect 213972 229044 214564 229072
rect 213972 229032 213978 229044
rect 214558 229032 214564 229044
rect 214616 229032 214622 229084
rect 214742 229032 214748 229084
rect 214800 229072 214806 229084
rect 257062 229072 257068 229084
rect 214800 229044 257068 229072
rect 214800 229032 214806 229044
rect 257062 229032 257068 229044
rect 257120 229032 257126 229084
rect 257890 229032 257896 229084
rect 257948 229072 257954 229084
rect 296346 229072 296352 229084
rect 257948 229044 296352 229072
rect 257948 229032 257954 229044
rect 296346 229032 296352 229044
rect 296404 229032 296410 229084
rect 302142 229032 302148 229084
rect 302200 229072 302206 229084
rect 331122 229072 331128 229084
rect 302200 229044 331128 229072
rect 302200 229032 302206 229044
rect 331122 229032 331128 229044
rect 331180 229032 331186 229084
rect 521626 229004 521654 229112
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 660942 229100 660948 229152
rect 661000 229140 661006 229152
rect 665450 229140 665456 229152
rect 661000 229112 665456 229140
rect 661000 229100 661006 229112
rect 665450 229100 665456 229112
rect 665508 229100 665514 229152
rect 673362 229100 673368 229152
rect 673420 229140 673426 229152
rect 673420 229112 674038 229140
rect 673420 229100 673426 229112
rect 521626 228976 528554 229004
rect 166994 228936 167000 228948
rect 103486 228908 167000 228936
rect 166994 228896 167000 228908
rect 167052 228896 167058 228948
rect 167362 228896 167368 228948
rect 167420 228936 167426 228948
rect 169478 228936 169484 228948
rect 167420 228908 169484 228936
rect 167420 228896 167426 228908
rect 169478 228896 169484 228908
rect 169536 228896 169542 228948
rect 179690 228936 179696 228948
rect 171980 228908 179696 228936
rect 171980 228868 172008 228908
rect 179690 228896 179696 228908
rect 179748 228896 179754 228948
rect 180058 228896 180064 228948
rect 180116 228936 180122 228948
rect 219894 228936 219900 228948
rect 180116 228908 219900 228936
rect 180116 228896 180122 228908
rect 219894 228896 219900 228908
rect 219952 228896 219958 228948
rect 246758 228936 246764 228948
rect 224926 228908 246764 228936
rect 171888 228840 172008 228868
rect 93762 228760 93768 228812
rect 93820 228800 93826 228812
rect 166810 228800 166816 228812
rect 93820 228772 166816 228800
rect 93820 228760 93826 228772
rect 166810 228760 166816 228772
rect 166868 228760 166874 228812
rect 166948 228760 166954 228812
rect 167006 228800 167012 228812
rect 171888 228800 171916 228840
rect 167006 228772 171916 228800
rect 167006 228760 167012 228772
rect 174814 228760 174820 228812
rect 174872 228800 174878 228812
rect 218146 228800 218152 228812
rect 174872 228772 218152 228800
rect 174872 228760 174878 228772
rect 218146 228760 218152 228772
rect 218204 228760 218210 228812
rect 224926 228800 224954 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 257706 228896 257712 228948
rect 257764 228936 257770 228948
rect 299566 228936 299572 228948
rect 257764 228908 299572 228936
rect 257764 228896 257770 228908
rect 299566 228896 299572 228908
rect 299624 228896 299630 228948
rect 300670 228896 300676 228948
rect 300728 228936 300734 228948
rect 330478 228936 330484 228948
rect 300728 228908 330484 228936
rect 300728 228896 300734 228908
rect 330478 228896 330484 228908
rect 330536 228896 330542 228948
rect 502426 228896 502432 228948
rect 502484 228936 502490 228948
rect 521010 228936 521016 228948
rect 502484 228908 521016 228936
rect 502484 228896 502490 228908
rect 521010 228896 521016 228908
rect 521068 228896 521074 228948
rect 528526 228936 528554 228976
rect 542446 228936 542452 228948
rect 528526 228908 542452 228936
rect 542446 228896 542452 228908
rect 542504 228896 542510 228948
rect 219912 228772 224954 228800
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 67600 228636 142844 228664
rect 67600 228624 67606 228636
rect 61654 228488 61660 228540
rect 61712 228528 61718 228540
rect 142614 228528 142620 228540
rect 61712 228500 142620 228528
rect 61712 228488 61718 228500
rect 142614 228488 142620 228500
rect 142672 228488 142678 228540
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 141142 228392 141148 228404
rect 57296 228364 141148 228392
rect 57296 228352 57302 228364
rect 141142 228352 141148 228364
rect 141200 228352 141206 228404
rect 142816 228392 142844 228636
rect 142982 228624 142988 228676
rect 143040 228664 143046 228676
rect 152458 228664 152464 228676
rect 143040 228636 152464 228664
rect 143040 228624 143046 228636
rect 152458 228624 152464 228636
rect 152516 228624 152522 228676
rect 153102 228624 153108 228676
rect 153160 228664 153166 228676
rect 153160 228636 212212 228664
rect 153160 228624 153166 228636
rect 142982 228488 142988 228540
rect 143040 228528 143046 228540
rect 145926 228528 145932 228540
rect 143040 228500 145932 228528
rect 143040 228488 143046 228500
rect 145926 228488 145932 228500
rect 145984 228488 145990 228540
rect 146110 228488 146116 228540
rect 146168 228528 146174 228540
rect 210694 228528 210700 228540
rect 146168 228500 210700 228528
rect 146168 228488 146174 228500
rect 210694 228488 210700 228500
rect 210752 228488 210758 228540
rect 212184 228528 212212 228636
rect 212350 228624 212356 228676
rect 212408 228664 212414 228676
rect 219912 228664 219940 228772
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 282822 228800 282828 228812
rect 238628 228772 282828 228800
rect 238628 228760 238634 228772
rect 282822 228760 282828 228772
rect 282880 228760 282886 228812
rect 296622 228760 296628 228812
rect 296680 228800 296686 228812
rect 329190 228800 329196 228812
rect 296680 228772 329196 228800
rect 296680 228760 296686 228772
rect 329190 228760 329196 228772
rect 329248 228760 329254 228812
rect 336458 228760 336464 228812
rect 336516 228800 336522 228812
rect 358814 228800 358820 228812
rect 336516 228772 358820 228800
rect 336516 228760 336522 228772
rect 358814 228760 358820 228772
rect 358872 228760 358878 228812
rect 359918 228760 359924 228812
rect 359976 228800 359982 228812
rect 376846 228800 376852 228812
rect 359976 228772 376852 228800
rect 359976 228760 359982 228772
rect 376846 228760 376852 228772
rect 376904 228760 376910 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490190 228800 490196 228812
rect 478932 228772 490196 228800
rect 478932 228760 478938 228772
rect 490190 228760 490196 228772
rect 490248 228760 490254 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541618 228800 541624 228812
rect 518584 228772 541624 228800
rect 518584 228760 518590 228772
rect 541618 228760 541624 228772
rect 541676 228760 541682 228812
rect 264790 228664 264796 228676
rect 212408 228636 219940 228664
rect 220004 228636 264796 228664
rect 212408 228624 212414 228636
rect 215846 228528 215852 228540
rect 212184 228500 215852 228528
rect 215846 228488 215852 228500
rect 215904 228488 215910 228540
rect 216214 228488 216220 228540
rect 216272 228528 216278 228540
rect 220004 228528 220032 228636
rect 264790 228624 264796 228636
rect 264848 228624 264854 228676
rect 285490 228624 285496 228676
rect 285548 228664 285554 228676
rect 318886 228664 318892 228676
rect 285548 228636 318892 228664
rect 285548 228624 285554 228636
rect 318886 228624 318892 228636
rect 318944 228624 318950 228676
rect 326890 228624 326896 228676
rect 326948 228664 326954 228676
rect 351086 228664 351092 228676
rect 326948 228636 351092 228664
rect 326948 228624 326954 228636
rect 351086 228624 351092 228636
rect 351144 228624 351150 228676
rect 354582 228624 354588 228676
rect 354640 228664 354646 228676
rect 372338 228664 372344 228676
rect 354640 228636 372344 228664
rect 354640 228624 354646 228636
rect 372338 228624 372344 228636
rect 372396 228624 372402 228676
rect 377766 228624 377772 228676
rect 377824 228664 377830 228676
rect 390370 228664 390376 228676
rect 377824 228636 390376 228664
rect 377824 228624 377830 228636
rect 390370 228624 390376 228636
rect 390428 228624 390434 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 515766 228664 515772 228676
rect 498620 228636 515772 228664
rect 498620 228624 498626 228636
rect 515766 228624 515772 228636
rect 515824 228624 515830 228676
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 554958 228664 554964 228676
rect 539652 228636 554964 228664
rect 539652 228624 539658 228636
rect 554958 228624 554964 228636
rect 555016 228624 555022 228676
rect 216272 228500 220032 228528
rect 216272 228488 216278 228500
rect 220170 228488 220176 228540
rect 220228 228528 220234 228540
rect 260282 228528 260288 228540
rect 220228 228500 260288 228528
rect 220228 228488 220234 228500
rect 260282 228488 260288 228500
rect 260340 228488 260346 228540
rect 268930 228488 268936 228540
rect 268988 228528 268994 228540
rect 306006 228528 306012 228540
rect 268988 228500 306012 228528
rect 268988 228488 268994 228500
rect 306006 228488 306012 228500
rect 306064 228488 306070 228540
rect 313918 228488 313924 228540
rect 313976 228528 313982 228540
rect 320818 228528 320824 228540
rect 313976 228500 320824 228528
rect 313976 228488 313982 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 325510 228488 325516 228540
rect 325568 228528 325574 228540
rect 349154 228528 349160 228540
rect 325568 228500 349160 228528
rect 325568 228488 325574 228500
rect 349154 228488 349160 228500
rect 349212 228488 349218 228540
rect 350442 228488 350448 228540
rect 350500 228528 350506 228540
rect 369118 228528 369124 228540
rect 350500 228500 369124 228528
rect 350500 228488 350506 228500
rect 369118 228488 369124 228500
rect 369176 228488 369182 228540
rect 373442 228488 373448 228540
rect 373500 228528 373506 228540
rect 387150 228528 387156 228540
rect 373500 228500 387156 228528
rect 373500 228488 373506 228500
rect 387150 228488 387156 228500
rect 387208 228488 387214 228540
rect 390462 228488 390468 228540
rect 390520 228528 390526 228540
rect 400030 228528 400036 228540
rect 390520 228500 400036 228528
rect 390520 228488 390526 228500
rect 400030 228488 400036 228500
rect 400088 228488 400094 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 148870 228392 148876 228404
rect 142816 228364 148876 228392
rect 148870 228352 148876 228364
rect 148928 228352 148934 228404
rect 152458 228352 152464 228404
rect 152516 228392 152522 228404
rect 166810 228392 166816 228404
rect 152516 228364 166816 228392
rect 152516 228352 152522 228364
rect 166810 228352 166816 228364
rect 166868 228352 166874 228404
rect 166948 228352 166954 228404
rect 167006 228392 167012 228404
rect 214558 228392 214564 228404
rect 167006 228364 214564 228392
rect 167006 228352 167012 228364
rect 214558 228352 214564 228364
rect 214616 228352 214622 228404
rect 218146 228352 218152 228404
rect 218204 228392 218210 228404
rect 231302 228392 231308 228404
rect 218204 228364 231308 228392
rect 218204 228352 218210 228364
rect 231302 228352 231308 228364
rect 231360 228352 231366 228404
rect 233878 228352 233884 228404
rect 233936 228392 233942 228404
rect 273806 228392 273812 228404
rect 233936 228364 273812 228392
rect 233936 228352 233942 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 274266 228352 274272 228404
rect 274324 228392 274330 228404
rect 312446 228392 312452 228404
rect 274324 228364 312452 228392
rect 274324 228352 274330 228364
rect 312446 228352 312452 228364
rect 312504 228352 312510 228404
rect 320082 228352 320088 228404
rect 320140 228392 320146 228404
rect 346854 228392 346860 228404
rect 320140 228364 346860 228392
rect 320140 228352 320146 228364
rect 346854 228352 346860 228364
rect 346912 228352 346918 228404
rect 347038 228352 347044 228404
rect 347096 228392 347102 228404
rect 365898 228392 365904 228404
rect 347096 228364 365904 228392
rect 347096 228352 347102 228364
rect 365898 228352 365904 228364
rect 365956 228352 365962 228404
rect 371142 228352 371148 228404
rect 371200 228392 371206 228404
rect 385218 228392 385224 228404
rect 371200 228364 385224 228392
rect 371200 228352 371206 228364
rect 385218 228352 385224 228364
rect 385276 228352 385282 228404
rect 386230 228352 386236 228404
rect 386288 228392 386294 228404
rect 397454 228392 397460 228404
rect 386288 228364 397460 228392
rect 386288 228352 386294 228364
rect 397454 228352 397460 228364
rect 397512 228352 397518 228404
rect 112806 228216 112812 228268
rect 112864 228256 112870 228268
rect 184934 228256 184940 228268
rect 112864 228228 184940 228256
rect 112864 228216 112870 228228
rect 184934 228216 184940 228228
rect 184992 228216 184998 228268
rect 189718 228216 189724 228268
rect 189776 228256 189782 228268
rect 239030 228256 239036 228268
rect 189776 228228 239036 228256
rect 189776 228216 189782 228228
rect 239030 228216 239036 228228
rect 239088 228216 239094 228268
rect 254946 228216 254952 228268
rect 255004 228256 255010 228268
rect 295702 228256 295708 228268
rect 255004 228228 295708 228256
rect 255004 228216 255010 228228
rect 295702 228216 295708 228228
rect 295760 228216 295766 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485682 228488 485688 228540
rect 485740 228528 485746 228540
rect 498286 228528 498292 228540
rect 485740 228500 498292 228528
rect 485740 228488 485746 228500
rect 498286 228488 498292 228500
rect 498344 228488 498350 228540
rect 499850 228488 499856 228540
rect 499908 228528 499914 228540
rect 517698 228528 517704 228540
rect 499908 228500 517704 228528
rect 499908 228488 499914 228500
rect 517698 228488 517704 228500
rect 517756 228488 517762 228540
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553210 228528 553216 228540
rect 527600 228500 553216 228528
rect 527600 228488 527606 228500
rect 553210 228488 553216 228500
rect 553268 228488 553274 228540
rect 555418 228488 555424 228540
rect 555476 228528 555482 228540
rect 571334 228528 571340 228540
rect 555476 228500 571340 228528
rect 555476 228488 555482 228500
rect 571334 228488 571340 228500
rect 571392 228488 571398 228540
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484578 228392 484584 228404
rect 474516 228364 484584 228392
rect 474516 228352 474522 228364
rect 484578 228352 484584 228364
rect 484636 228352 484642 228404
rect 485038 228352 485044 228404
rect 485096 228392 485102 228404
rect 498562 228392 498568 228404
rect 485096 228364 498568 228392
rect 485096 228352 485102 228364
rect 498562 228352 498568 228364
rect 498620 228352 498626 228404
rect 507118 228352 507124 228404
rect 507176 228392 507182 228404
rect 507176 228364 509234 228392
rect 507176 228352 507182 228364
rect 400140 228228 400260 228256
rect 509206 228256 509234 228364
rect 512086 228352 512092 228404
rect 512144 228392 512150 228404
rect 532970 228392 532976 228404
rect 512144 228364 532976 228392
rect 512144 228352 512150 228364
rect 532970 228352 532976 228364
rect 533028 228352 533034 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 663518 228352 663524 228404
rect 663576 228392 663582 228404
rect 672166 228392 672172 228404
rect 663576 228364 672172 228392
rect 663576 228352 663582 228364
rect 672166 228352 672172 228364
rect 672224 228352 672230 228404
rect 512730 228256 512736 228268
rect 509206 228228 512736 228256
rect 400140 228132 400168 228228
rect 512730 228216 512736 228228
rect 512788 228216 512794 228268
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540882 228256 540888 228268
rect 539468 228228 540888 228256
rect 539468 228216 539474 228228
rect 540882 228216 540888 228228
rect 540940 228216 540946 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 190086 228120 190092 228132
rect 120040 228092 190092 228120
rect 120040 228080 120046 228092
rect 190086 228080 190092 228092
rect 190144 228080 190150 228132
rect 192938 228080 192944 228132
rect 192996 228120 193002 228132
rect 204714 228120 204720 228132
rect 192996 228092 204720 228120
rect 192996 228080 193002 228092
rect 204714 228080 204720 228092
rect 204772 228080 204778 228132
rect 214558 228080 214564 228132
rect 214616 228120 214622 228132
rect 214616 228092 215294 228120
rect 214616 228080 214622 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 195146 227984 195152 227996
rect 126756 227956 195152 227984
rect 126756 227944 126762 227956
rect 195146 227944 195152 227956
rect 195204 227944 195210 227996
rect 205450 227944 205456 227996
rect 205508 227984 205514 227996
rect 214742 227984 214748 227996
rect 205508 227956 214748 227984
rect 205508 227944 205514 227956
rect 214742 227944 214748 227956
rect 214800 227944 214806 227996
rect 215266 227984 215294 228092
rect 217502 228080 217508 228132
rect 217560 228120 217566 228132
rect 219434 228120 219440 228132
rect 217560 228092 219440 228120
rect 217560 228080 217566 228092
rect 219434 228080 219440 228092
rect 219492 228080 219498 228132
rect 219894 228080 219900 228132
rect 219952 228120 219958 228132
rect 225782 228120 225788 228132
rect 219952 228092 225788 228120
rect 219952 228080 219958 228092
rect 225782 228080 225788 228092
rect 225840 228080 225846 228132
rect 225966 228080 225972 228132
rect 226024 228120 226030 228132
rect 272518 228120 272524 228132
rect 226024 228092 272524 228120
rect 226024 228080 226030 228092
rect 272518 228080 272524 228092
rect 272576 228080 272582 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 220998 227984 221004 227996
rect 215266 227956 221004 227984
rect 220998 227944 221004 227956
rect 221056 227944 221062 227996
rect 251266 227984 251272 227996
rect 221200 227956 251272 227984
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 200390 227848 200396 227860
rect 133564 227820 200396 227848
rect 133564 227808 133570 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 203518 227808 203524 227860
rect 203576 227848 203582 227860
rect 203576 227820 205128 227848
rect 203576 227808 203582 227820
rect 42426 227672 42432 227724
rect 42484 227712 42490 227724
rect 42978 227712 42984 227724
rect 42484 227684 42984 227712
rect 42484 227672 42490 227684
rect 42978 227672 42984 227684
rect 43036 227672 43042 227724
rect 64782 227672 64788 227724
rect 64840 227712 64846 227724
rect 111058 227712 111064 227724
rect 64840 227684 111064 227712
rect 64840 227672 64846 227684
rect 111058 227672 111064 227684
rect 111116 227672 111122 227724
rect 117222 227672 117228 227724
rect 117280 227712 117286 227724
rect 187510 227712 187516 227724
rect 117280 227684 187516 227712
rect 117280 227672 117286 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 187694 227672 187700 227724
rect 187752 227712 187758 227724
rect 187752 227684 193076 227712
rect 187752 227672 187758 227684
rect 110138 227536 110144 227588
rect 110196 227576 110202 227588
rect 182358 227576 182364 227588
rect 110196 227548 182364 227576
rect 110196 227536 110202 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 185394 227536 185400 227588
rect 185452 227576 185458 227588
rect 192662 227576 192668 227588
rect 185452 227548 192668 227576
rect 185452 227536 185458 227548
rect 192662 227536 192668 227548
rect 192720 227536 192726 227588
rect 193048 227576 193076 227684
rect 200022 227672 200028 227724
rect 200080 227712 200086 227724
rect 204898 227712 204904 227724
rect 200080 227684 204904 227712
rect 200080 227672 200086 227684
rect 204898 227672 204904 227684
rect 204956 227672 204962 227724
rect 205100 227712 205128 227820
rect 210970 227808 210976 227860
rect 211028 227848 211034 227860
rect 220078 227848 220084 227860
rect 211028 227820 220084 227848
rect 211028 227808 211034 227820
rect 220078 227808 220084 227820
rect 220136 227808 220142 227860
rect 221200 227848 221228 227956
rect 251266 227944 251272 227956
rect 251324 227944 251330 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 233878 227848 233884 227860
rect 220280 227820 221228 227848
rect 226352 227820 233884 227848
rect 217778 227712 217784 227724
rect 205100 227684 217784 227712
rect 217778 227672 217784 227684
rect 217836 227672 217842 227724
rect 219434 227672 219440 227724
rect 219492 227712 219498 227724
rect 220280 227712 220308 227820
rect 224586 227740 224592 227792
rect 224644 227780 224650 227792
rect 224644 227752 224954 227780
rect 224644 227740 224650 227752
rect 219492 227684 220308 227712
rect 219492 227672 219498 227684
rect 220446 227672 220452 227724
rect 220504 227712 220510 227724
rect 223574 227712 223580 227724
rect 220504 227684 223580 227712
rect 220504 227672 220510 227684
rect 223574 227672 223580 227684
rect 223632 227672 223638 227724
rect 224926 227712 224954 227752
rect 226352 227712 226380 227820
rect 233878 227808 233884 227820
rect 233936 227808 233942 227860
rect 239306 227808 239312 227860
rect 239364 227848 239370 227860
rect 243538 227848 243544 227860
rect 239364 227820 243544 227848
rect 239364 227808 239370 227820
rect 243538 227808 243544 227820
rect 243596 227808 243602 227860
rect 246298 227808 246304 227860
rect 246356 227848 246362 227860
rect 248690 227848 248696 227860
rect 246356 227820 248696 227848
rect 246356 227808 246362 227820
rect 248690 227808 248696 227820
rect 248748 227808 248754 227860
rect 249058 227808 249064 227860
rect 249116 227848 249122 227860
rect 253842 227848 253848 227860
rect 249116 227820 253848 227848
rect 249116 227808 249122 227820
rect 253842 227808 253848 227820
rect 253900 227808 253906 227860
rect 331030 227740 331036 227792
rect 331088 227780 331094 227792
rect 334250 227780 334256 227792
rect 331088 227752 334256 227780
rect 331088 227740 331094 227752
rect 334250 227740 334256 227752
rect 334308 227740 334314 227792
rect 351086 227740 351092 227792
rect 351144 227780 351150 227792
rect 353018 227780 353024 227792
rect 351144 227752 353024 227780
rect 351144 227740 351150 227752
rect 353018 227740 353024 227752
rect 353076 227740 353082 227792
rect 371786 227740 371792 227792
rect 371844 227780 371850 227792
rect 373626 227780 373632 227792
rect 371844 227752 373632 227780
rect 371844 227740 371850 227752
rect 373626 227740 373632 227752
rect 373684 227740 373690 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 489914 227740 489920 227792
rect 489972 227780 489978 227792
rect 494514 227780 494520 227792
rect 489972 227752 494520 227780
rect 489972 227740 489978 227752
rect 494514 227740 494520 227752
rect 494572 227740 494578 227792
rect 660482 227740 660488 227792
rect 660540 227780 660546 227792
rect 665266 227780 665272 227792
rect 660540 227752 665272 227780
rect 660540 227740 660546 227752
rect 665266 227740 665272 227752
rect 665324 227740 665330 227792
rect 669038 227740 669044 227792
rect 669096 227780 669102 227792
rect 672902 227780 672908 227792
rect 669096 227752 672908 227780
rect 669096 227740 669102 227752
rect 672902 227740 672908 227752
rect 672960 227740 672966 227792
rect 224926 227684 226380 227712
rect 226702 227672 226708 227724
rect 226760 227712 226766 227724
rect 268010 227712 268016 227724
rect 226760 227684 268016 227712
rect 226760 227672 226766 227684
rect 268010 227672 268016 227684
rect 268068 227672 268074 227724
rect 293770 227672 293776 227724
rect 293828 227712 293834 227724
rect 325326 227712 325332 227724
rect 293828 227684 325332 227712
rect 293828 227672 293834 227684
rect 325326 227672 325332 227684
rect 325384 227672 325390 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 214742 227576 214748 227588
rect 193048 227548 214748 227576
rect 214742 227536 214748 227548
rect 214800 227536 214806 227588
rect 214926 227536 214932 227588
rect 214984 227576 214990 227588
rect 262214 227576 262220 227588
rect 214984 227548 262220 227576
rect 214984 227536 214990 227548
rect 262214 227536 262220 227548
rect 262272 227536 262278 227588
rect 264790 227536 264796 227588
rect 264848 227576 264854 227588
rect 304718 227576 304724 227588
rect 264848 227548 304724 227576
rect 264848 227536 264854 227548
rect 304718 227536 304724 227548
rect 304776 227536 304782 227588
rect 315482 227536 315488 227588
rect 315540 227576 315546 227588
rect 341426 227576 341432 227588
rect 315540 227548 341432 227576
rect 315540 227536 315546 227548
rect 341426 227536 341432 227548
rect 341484 227536 341490 227588
rect 525702 227536 525708 227588
rect 525760 227576 525766 227588
rect 537478 227576 537484 227588
rect 525760 227548 537484 227576
rect 525760 227536 525766 227548
rect 537478 227536 537484 227548
rect 537536 227536 537542 227588
rect 60642 227400 60648 227452
rect 60700 227440 60706 227452
rect 102134 227440 102140 227452
rect 60700 227412 102140 227440
rect 60700 227400 60706 227412
rect 102134 227400 102140 227412
rect 102192 227400 102198 227452
rect 103422 227400 103428 227452
rect 103480 227440 103486 227452
rect 171226 227440 171232 227452
rect 103480 227412 171232 227440
rect 103480 227400 103486 227412
rect 171226 227400 171232 227412
rect 171284 227400 171290 227452
rect 172146 227400 172152 227452
rect 172204 227440 172210 227452
rect 177206 227440 177212 227452
rect 172204 227412 177212 227440
rect 172204 227400 172210 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 181346 227400 181352 227452
rect 181404 227440 181410 227452
rect 181404 227412 185900 227440
rect 181404 227400 181410 227412
rect 96430 227264 96436 227316
rect 96488 227304 96494 227316
rect 169478 227304 169484 227316
rect 96488 227276 157196 227304
rect 96488 227264 96494 227276
rect 89622 227128 89628 227180
rect 89680 227168 89686 227180
rect 156874 227168 156880 227180
rect 89680 227140 156880 227168
rect 89680 227128 89686 227140
rect 156874 227128 156880 227140
rect 156932 227128 156938 227180
rect 157168 227168 157196 227276
rect 157444 227276 169484 227304
rect 157444 227168 157472 227276
rect 169478 227264 169484 227276
rect 169536 227264 169542 227316
rect 185578 227304 185584 227316
rect 171336 227276 185584 227304
rect 157168 227140 157472 227168
rect 160186 227128 160192 227180
rect 160244 227168 160250 227180
rect 171336 227168 171364 227276
rect 185578 227264 185584 227276
rect 185636 227264 185642 227316
rect 185872 227304 185900 227412
rect 186130 227400 186136 227452
rect 186188 227440 186194 227452
rect 187694 227440 187700 227452
rect 186188 227412 187700 227440
rect 186188 227400 186194 227412
rect 187694 227400 187700 227412
rect 187752 227400 187758 227452
rect 189902 227400 189908 227452
rect 189960 227440 189966 227452
rect 204714 227440 204720 227452
rect 189960 227412 204720 227440
rect 189960 227400 189966 227412
rect 204714 227400 204720 227412
rect 204772 227400 204778 227452
rect 204898 227400 204904 227452
rect 204956 227440 204962 227452
rect 251910 227440 251916 227452
rect 204956 227412 251916 227440
rect 204956 227400 204962 227412
rect 251910 227400 251916 227412
rect 251968 227400 251974 227452
rect 259362 227400 259368 227452
rect 259420 227440 259426 227452
rect 298278 227440 298284 227452
rect 259420 227412 298284 227440
rect 259420 227400 259426 227412
rect 298278 227400 298284 227412
rect 298336 227400 298342 227452
rect 306190 227400 306196 227452
rect 306248 227440 306254 227452
rect 336918 227440 336924 227452
rect 306248 227412 336924 227440
rect 306248 227400 306254 227412
rect 336918 227400 336924 227412
rect 336976 227400 336982 227452
rect 337746 227400 337752 227452
rect 337804 227440 337810 227452
rect 345014 227440 345020 227452
rect 337804 227412 345020 227440
rect 337804 227400 337810 227412
rect 345014 227400 345020 227412
rect 345072 227400 345078 227452
rect 352558 227400 352564 227452
rect 352616 227440 352622 227452
rect 363230 227440 363236 227452
rect 352616 227412 363236 227440
rect 352616 227400 352622 227412
rect 363230 227400 363236 227412
rect 363288 227400 363294 227452
rect 494698 227400 494704 227452
rect 494756 227440 494762 227452
rect 511074 227440 511080 227452
rect 494756 227412 511080 227440
rect 494756 227400 494762 227412
rect 511074 227400 511080 227412
rect 511132 227400 511138 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 536098 227400 536104 227452
rect 536156 227440 536162 227452
rect 552474 227440 552480 227452
rect 536156 227412 552480 227440
rect 536156 227400 536162 227412
rect 552474 227400 552480 227412
rect 552532 227400 552538 227452
rect 219434 227304 219440 227316
rect 185872 227276 219440 227304
rect 219434 227264 219440 227276
rect 219492 227264 219498 227316
rect 219802 227264 219808 227316
rect 219860 227304 219866 227316
rect 241606 227304 241612 227316
rect 219860 227276 241612 227304
rect 219860 227264 219866 227276
rect 241606 227264 241612 227276
rect 241664 227264 241670 227316
rect 249242 227264 249248 227316
rect 249300 227304 249306 227316
rect 290550 227304 290556 227316
rect 249300 227276 290556 227304
rect 249300 227264 249306 227276
rect 290550 227264 290556 227276
rect 290608 227264 290614 227316
rect 291010 227264 291016 227316
rect 291068 227304 291074 227316
rect 322106 227304 322112 227316
rect 291068 227276 322112 227304
rect 291068 227264 291074 227276
rect 322106 227264 322112 227276
rect 322164 227264 322170 227316
rect 340690 227264 340696 227316
rect 340748 227304 340754 227316
rect 361390 227304 361396 227316
rect 340748 227276 361396 227304
rect 340748 227264 340754 227276
rect 361390 227264 361396 227276
rect 361448 227264 361454 227316
rect 363598 227264 363604 227316
rect 363656 227304 363662 227316
rect 368474 227304 368480 227316
rect 363656 227276 368480 227304
rect 363656 227264 363662 227276
rect 368474 227264 368480 227276
rect 368532 227264 368538 227316
rect 382090 227264 382096 227316
rect 382148 227304 382154 227316
rect 392946 227304 392952 227316
rect 382148 227276 392952 227304
rect 382148 227264 382154 227276
rect 392946 227264 392952 227276
rect 393004 227264 393010 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 160244 227140 171364 227168
rect 160244 227128 160250 227140
rect 171594 227128 171600 227180
rect 171652 227168 171658 227180
rect 171652 227140 220124 227168
rect 171652 227128 171658 227140
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142154 227032 142160 227044
rect 56560 227004 142160 227032
rect 56560 226992 56566 227004
rect 142154 226992 142160 227004
rect 142212 226992 142218 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 204070 227032 204076 227044
rect 143316 227004 204076 227032
rect 143316 226992 143322 227004
rect 204070 226992 204076 227004
rect 204128 226992 204134 227044
rect 214098 227032 214104 227044
rect 204916 227004 214104 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 204916 226896 204944 227004
rect 214098 226992 214104 227004
rect 214156 226992 214162 227044
rect 220096 227032 220124 227140
rect 220262 227128 220268 227180
rect 220320 227168 220326 227180
rect 233694 227168 233700 227180
rect 220320 227140 233700 227168
rect 220320 227128 220326 227140
rect 233694 227128 233700 227140
rect 233752 227128 233758 227180
rect 235810 227128 235816 227180
rect 235868 227168 235874 227180
rect 280246 227168 280252 227180
rect 235868 227140 280252 227168
rect 235868 227128 235874 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 281350 227128 281356 227180
rect 281408 227168 281414 227180
rect 317598 227168 317604 227180
rect 281408 227140 317604 227168
rect 281408 227128 281414 227140
rect 317598 227128 317604 227140
rect 317656 227128 317662 227180
rect 322198 227128 322204 227180
rect 322256 227168 322262 227180
rect 332410 227168 332416 227180
rect 322256 227140 332416 227168
rect 322256 227128 322262 227140
rect 332410 227128 332416 227140
rect 332468 227128 332474 227180
rect 333882 227128 333888 227180
rect 333940 227168 333946 227180
rect 356238 227168 356244 227180
rect 333940 227140 356244 227168
rect 333940 227128 333946 227140
rect 356238 227128 356244 227140
rect 356296 227128 356302 227180
rect 357250 227128 357256 227180
rect 357308 227168 357314 227180
rect 374270 227168 374276 227180
rect 357308 227140 374276 227168
rect 357308 227128 357314 227140
rect 374270 227128 374276 227140
rect 374328 227128 374334 227180
rect 376662 227128 376668 227180
rect 376720 227168 376726 227180
rect 389726 227168 389732 227180
rect 376720 227140 389732 227168
rect 376720 227128 376726 227140
rect 389726 227128 389732 227140
rect 389784 227128 389790 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 510614 227264 510620 227316
rect 510672 227304 510678 227316
rect 524414 227304 524420 227316
rect 510672 227276 524420 227304
rect 510672 227264 510678 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 551554 227304 551560 227316
rect 526312 227276 551560 227304
rect 526312 227264 526318 227276
rect 551554 227264 551560 227276
rect 551612 227264 551618 227316
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 490374 227128 490380 227180
rect 490432 227168 490438 227180
rect 503162 227168 503168 227180
rect 490432 227140 503168 227168
rect 490432 227128 490438 227140
rect 503162 227128 503168 227140
rect 503220 227128 503226 227180
rect 505002 227128 505008 227180
rect 505060 227168 505066 227180
rect 523034 227168 523040 227180
rect 505060 227140 523040 227168
rect 505060 227128 505066 227140
rect 523034 227128 523040 227140
rect 523092 227128 523098 227180
rect 523678 227128 523684 227180
rect 523736 227168 523742 227180
rect 548150 227168 548156 227180
rect 523736 227140 548156 227168
rect 523736 227128 523742 227140
rect 548150 227128 548156 227140
rect 548208 227128 548214 227180
rect 556798 227128 556804 227180
rect 556856 227168 556862 227180
rect 570598 227168 570604 227180
rect 556856 227140 570604 227168
rect 556856 227128 556862 227140
rect 570598 227128 570604 227140
rect 570656 227128 570662 227180
rect 668578 227128 668584 227180
rect 668636 227168 668642 227180
rect 673546 227168 673552 227180
rect 668636 227140 673552 227168
rect 668636 227128 668642 227140
rect 673546 227128 673552 227140
rect 673604 227128 673610 227180
rect 228726 227032 228732 227044
rect 214576 227004 220032 227032
rect 220096 227004 228732 227032
rect 214576 226896 214604 227004
rect 185636 226868 204944 226896
rect 209746 226868 214604 226896
rect 185636 226856 185642 226868
rect 129550 226720 129556 226772
rect 129608 226760 129614 226772
rect 197446 226760 197452 226772
rect 129608 226732 197452 226760
rect 129608 226720 129614 226732
rect 197446 226720 197452 226732
rect 197504 226720 197510 226772
rect 204714 226720 204720 226772
rect 204772 226760 204778 226772
rect 209746 226760 209774 226868
rect 214742 226856 214748 226908
rect 214800 226896 214806 226908
rect 219802 226896 219808 226908
rect 214800 226868 219808 226896
rect 214800 226856 214806 226868
rect 219802 226856 219808 226868
rect 219860 226856 219866 226908
rect 220004 226896 220032 227004
rect 228726 226992 228732 227004
rect 228784 226992 228790 227044
rect 228910 226992 228916 227044
rect 228968 227032 228974 227044
rect 271230 227032 271236 227044
rect 228968 227004 271236 227032
rect 228968 226992 228974 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 310330 226992 310336 227044
rect 310388 227032 310394 227044
rect 338206 227032 338212 227044
rect 310388 227004 338212 227032
rect 310388 226992 310394 227004
rect 338206 226992 338212 227004
rect 338264 226992 338270 227044
rect 338666 226992 338672 227044
rect 338724 227032 338730 227044
rect 360102 227032 360108 227044
rect 338724 227004 360108 227032
rect 338724 226992 338730 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 362770 226992 362776 227044
rect 362828 227032 362834 227044
rect 379054 227032 379060 227044
rect 362828 227004 379060 227032
rect 362828 226992 362834 227004
rect 379054 226992 379060 227004
rect 379112 226992 379118 227044
rect 391750 226992 391756 227044
rect 391808 227032 391814 227044
rect 403526 227032 403532 227044
rect 391808 227004 403532 227032
rect 391808 226992 391814 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 506290 226992 506296 227044
rect 506348 227032 506354 227044
rect 526622 227032 526628 227044
rect 506348 227004 526628 227032
rect 506348 226992 506354 227004
rect 526622 226992 526628 227004
rect 526680 226992 526686 227044
rect 533338 226992 533344 227044
rect 533396 227032 533402 227044
rect 560754 227032 560760 227044
rect 533396 227004 560760 227032
rect 533396 226992 533402 227004
rect 560754 226992 560760 227004
rect 560812 226992 560818 227044
rect 652018 226992 652024 227044
rect 652076 227032 652082 227044
rect 673546 227032 673552 227044
rect 652076 227004 673552 227032
rect 652076 226992 652082 227004
rect 673546 226992 673552 227004
rect 673604 226992 673610 227044
rect 426434 226924 426440 226976
rect 426492 226964 426498 226976
rect 426986 226964 426992 226976
rect 426492 226936 426992 226964
rect 426492 226924 426498 226936
rect 426986 226924 426992 226936
rect 427044 226924 427050 226976
rect 220262 226896 220268 226908
rect 220004 226868 220268 226896
rect 220262 226856 220268 226868
rect 220320 226856 220326 226908
rect 267366 226896 267372 226908
rect 224926 226868 267372 226896
rect 204772 226732 209774 226760
rect 204772 226720 204778 226732
rect 214098 226720 214104 226772
rect 214156 226760 214162 226772
rect 218422 226760 218428 226772
rect 214156 226732 218428 226760
rect 214156 226720 214162 226732
rect 218422 226720 218428 226732
rect 218480 226720 218486 226772
rect 219342 226720 219348 226772
rect 219400 226760 219406 226772
rect 224926 226760 224954 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 378778 226788 378784 226840
rect 378836 226828 378842 226840
rect 385862 226828 385868 226840
rect 378836 226800 385868 226828
rect 378836 226788 378842 226800
rect 385862 226788 385868 226800
rect 385920 226788 385926 226840
rect 219400 226732 224954 226760
rect 219400 226720 219406 226732
rect 225598 226720 225604 226772
rect 225656 226760 225662 226772
rect 238386 226760 238392 226772
rect 225656 226732 238392 226760
rect 225656 226720 225662 226732
rect 238386 226720 238392 226732
rect 238444 226720 238450 226772
rect 241146 226720 241152 226772
rect 241204 226760 241210 226772
rect 286686 226760 286692 226772
rect 241204 226732 286692 226760
rect 241204 226720 241210 226732
rect 286686 226720 286692 226732
rect 286744 226720 286750 226772
rect 136542 226584 136548 226636
rect 136600 226624 136606 226636
rect 203150 226624 203156 226636
rect 136600 226596 203156 226624
rect 136600 226584 136606 226596
rect 203150 226584 203156 226596
rect 203208 226584 203214 226636
rect 204070 226584 204076 226636
rect 204128 226624 204134 226636
rect 208118 226624 208124 226636
rect 204128 226596 208124 226624
rect 204128 226584 204134 226596
rect 208118 226584 208124 226596
rect 208176 226584 208182 226636
rect 212166 226584 212172 226636
rect 212224 226624 212230 226636
rect 214926 226624 214932 226636
rect 212224 226596 214932 226624
rect 212224 226584 212230 226596
rect 214926 226584 214932 226596
rect 214984 226584 214990 226636
rect 220446 226584 220452 226636
rect 220504 226624 220510 226636
rect 226702 226624 226708 226636
rect 220504 226596 226708 226624
rect 220504 226584 220510 226596
rect 226702 226584 226708 226596
rect 226760 226584 226766 226636
rect 670786 226516 670792 226568
rect 670844 226556 670850 226568
rect 672994 226556 673000 226568
rect 670844 226528 672644 226556
rect 672842 226528 673000 226556
rect 670844 226516 670850 226528
rect 106918 226448 106924 226500
rect 106976 226488 106982 226500
rect 146570 226488 146576 226500
rect 106976 226460 146576 226488
rect 106976 226448 106982 226460
rect 146570 226448 146576 226460
rect 146628 226448 146634 226500
rect 150066 226448 150072 226500
rect 150124 226488 150130 226500
rect 213270 226488 213276 226500
rect 150124 226460 213276 226488
rect 150124 226448 150130 226460
rect 213270 226448 213276 226460
rect 213328 226448 213334 226500
rect 216398 226448 216404 226500
rect 216456 226488 216462 226500
rect 220630 226488 220636 226500
rect 216456 226460 220636 226488
rect 216456 226448 216462 226460
rect 220630 226448 220636 226460
rect 220688 226448 220694 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 228910 226488 228916 226500
rect 221884 226460 228916 226488
rect 221884 226448 221890 226460
rect 228910 226448 228916 226460
rect 228968 226448 228974 226500
rect 369118 226448 369124 226500
rect 369176 226488 369182 226500
rect 376202 226488 376208 226500
rect 369176 226460 376208 226488
rect 369176 226448 369182 226460
rect 376202 226448 376208 226460
rect 376260 226448 376266 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672616 226488 672644 226528
rect 672994 226516 673000 226528
rect 673052 226516 673058 226568
rect 672616 226460 672750 226488
rect 386046 226380 386052 226432
rect 386104 226420 386110 226432
rect 391198 226420 391204 226432
rect 386104 226392 391204 226420
rect 386104 226380 386110 226392
rect 391198 226380 391204 226392
rect 391256 226380 391262 226432
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 488074 226312 488080 226364
rect 488132 226352 488138 226364
rect 490006 226352 490012 226364
rect 488132 226324 490012 226352
rect 488132 226312 488138 226324
rect 490006 226312 490012 226324
rect 490064 226312 490070 226364
rect 672150 226312 672156 226364
rect 672208 226352 672214 226364
rect 672208 226324 672304 226352
rect 672208 226312 672214 226324
rect 122558 226244 122564 226296
rect 122616 226284 122622 226296
rect 193950 226284 193956 226296
rect 122616 226256 193956 226284
rect 122616 226244 122622 226256
rect 193950 226244 193956 226256
rect 194008 226244 194014 226296
rect 194134 226244 194140 226296
rect 194192 226284 194198 226296
rect 204898 226284 204904 226296
rect 194192 226256 204904 226284
rect 194192 226244 194198 226256
rect 204898 226244 204904 226256
rect 204956 226244 204962 226296
rect 205082 226244 205088 226296
rect 205140 226284 205146 226296
rect 255130 226284 255136 226296
rect 205140 226256 255136 226284
rect 205140 226244 205146 226256
rect 255130 226244 255136 226256
rect 255188 226244 255194 226296
rect 260650 226244 260656 226296
rect 260708 226284 260714 226296
rect 298922 226284 298928 226296
rect 260708 226256 298928 226284
rect 260708 226244 260714 226256
rect 298922 226244 298928 226256
rect 298980 226244 298986 226296
rect 308214 226244 308220 226296
rect 308272 226284 308278 226296
rect 336274 226284 336280 226296
rect 308272 226256 336280 226284
rect 308272 226244 308278 226256
rect 336274 226244 336280 226256
rect 336332 226244 336338 226296
rect 388622 226244 388628 226296
rect 388680 226284 388686 226296
rect 394234 226284 394240 226296
rect 388680 226256 394240 226284
rect 388680 226244 388686 226256
rect 394234 226244 394240 226256
rect 394292 226244 394298 226296
rect 539962 226284 539968 226296
rect 528526 226256 539968 226284
rect 72418 226108 72424 226160
rect 72476 226148 72482 226160
rect 141142 226148 141148 226160
rect 72476 226120 141148 226148
rect 72476 226108 72482 226120
rect 141142 226108 141148 226120
rect 141200 226108 141206 226160
rect 141510 226108 141516 226160
rect 141568 226148 141574 226160
rect 145006 226148 145012 226160
rect 141568 226120 145012 226148
rect 141568 226108 141574 226120
rect 145006 226108 145012 226120
rect 145064 226108 145070 226160
rect 145190 226108 145196 226160
rect 145248 226148 145254 226160
rect 146754 226148 146760 226160
rect 145248 226120 146760 226148
rect 145248 226108 145254 226120
rect 146754 226108 146760 226120
rect 146812 226108 146818 226160
rect 148962 226108 148968 226160
rect 149020 226148 149026 226160
rect 213454 226148 213460 226160
rect 149020 226120 213460 226148
rect 149020 226108 149026 226120
rect 213454 226108 213460 226120
rect 213512 226108 213518 226160
rect 213638 226108 213644 226160
rect 213696 226148 213702 226160
rect 220078 226148 220084 226160
rect 213696 226120 220084 226148
rect 213696 226108 213702 226120
rect 220078 226108 220084 226120
rect 220136 226108 220142 226160
rect 222010 226108 222016 226160
rect 222068 226148 222074 226160
rect 269942 226148 269948 226160
rect 222068 226120 269948 226148
rect 222068 226108 222074 226120
rect 269942 226108 269948 226120
rect 270000 226108 270006 226160
rect 270218 226108 270224 226160
rect 270276 226148 270282 226160
rect 287054 226148 287060 226160
rect 270276 226120 287060 226148
rect 270276 226108 270282 226120
rect 287054 226108 287060 226120
rect 287112 226108 287118 226160
rect 288066 226108 288072 226160
rect 288124 226148 288130 226160
rect 322750 226148 322756 226160
rect 288124 226120 322756 226148
rect 288124 226108 288130 226120
rect 322750 226108 322756 226120
rect 322808 226108 322814 226160
rect 526438 226108 526444 226160
rect 526496 226148 526502 226160
rect 528526 226148 528554 226256
rect 539962 226244 539968 226256
rect 540020 226244 540026 226296
rect 563698 226244 563704 226296
rect 563756 226284 563762 226296
rect 568114 226284 568120 226296
rect 563756 226256 568120 226284
rect 563756 226244 563762 226256
rect 568114 226244 568120 226256
rect 568172 226244 568178 226296
rect 672276 226284 672304 226324
rect 672276 226256 672630 226284
rect 538490 226148 538496 226160
rect 526496 226120 528554 226148
rect 538186 226120 538496 226148
rect 526496 226108 526502 226120
rect 83458 225972 83464 226024
rect 83516 226012 83522 226024
rect 163038 226012 163044 226024
rect 83516 225984 163044 226012
rect 83516 225972 83522 225984
rect 163038 225972 163044 225984
rect 163096 225972 163102 226024
rect 196342 225972 196348 226024
rect 196400 226012 196406 226024
rect 236454 226012 236460 226024
rect 196400 225984 236460 226012
rect 196400 225972 196406 225984
rect 236454 225972 236460 225984
rect 236512 225972 236518 226024
rect 252462 225972 252468 226024
rect 252520 226012 252526 226024
rect 293126 226012 293132 226024
rect 252520 225984 293132 226012
rect 252520 225972 252526 225984
rect 293126 225972 293132 225984
rect 293184 225972 293190 226024
rect 299382 225972 299388 226024
rect 299440 226012 299446 226024
rect 328546 226012 328552 226024
rect 299440 225984 328552 226012
rect 299440 225972 299446 225984
rect 328546 225972 328552 225984
rect 328604 225972 328610 226024
rect 335170 225972 335176 226024
rect 335228 226012 335234 226024
rect 356882 226012 356888 226024
rect 335228 225984 356888 226012
rect 335228 225972 335234 225984
rect 356882 225972 356888 225984
rect 356940 225972 356946 226024
rect 361206 225972 361212 226024
rect 361264 226012 361270 226024
rect 377490 226012 377496 226024
rect 361264 225984 377496 226012
rect 361264 225972 361270 225984
rect 377490 225972 377496 225984
rect 377548 225972 377554 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538186 226012 538214 226120
rect 538490 226108 538496 226120
rect 538548 226108 538554 226160
rect 670786 226040 670792 226092
rect 670844 226080 670850 226092
rect 670844 226052 672520 226080
rect 670844 226040 670850 226052
rect 516652 225984 538214 226012
rect 516652 225972 516658 225984
rect 538306 225972 538312 226024
rect 538364 226012 538370 226024
rect 556154 226012 556160 226024
rect 538364 225984 556160 226012
rect 538364 225972 538370 225984
rect 556154 225972 556160 225984
rect 556212 225972 556218 226024
rect 76558 225836 76564 225888
rect 76616 225876 76622 225888
rect 157886 225876 157892 225888
rect 76616 225848 157892 225876
rect 76616 225836 76622 225848
rect 157886 225836 157892 225848
rect 157944 225836 157950 225888
rect 169662 225836 169668 225888
rect 169720 225876 169726 225888
rect 171594 225876 171600 225888
rect 169720 225848 171600 225876
rect 169720 225836 169726 225848
rect 171594 225836 171600 225848
rect 171652 225836 171658 225888
rect 171778 225836 171784 225888
rect 171836 225876 171842 225888
rect 204530 225876 204536 225888
rect 171836 225848 204536 225876
rect 171836 225836 171842 225848
rect 204530 225836 204536 225848
rect 204588 225836 204594 225888
rect 204898 225836 204904 225888
rect 204956 225876 204962 225888
rect 213638 225876 213644 225888
rect 204956 225848 213644 225876
rect 204956 225836 204962 225848
rect 213638 225836 213644 225848
rect 213696 225836 213702 225888
rect 220078 225836 220084 225888
rect 220136 225876 220142 225888
rect 244182 225876 244188 225888
rect 220136 225848 244188 225876
rect 220136 225836 220142 225848
rect 244182 225836 244188 225848
rect 244240 225836 244246 225888
rect 261846 225836 261852 225888
rect 261904 225876 261910 225888
rect 300854 225876 300860 225888
rect 261904 225848 300860 225876
rect 261904 225836 261910 225848
rect 300854 225836 300860 225848
rect 300912 225836 300918 225888
rect 312906 225836 312912 225888
rect 312964 225876 312970 225888
rect 341702 225876 341708 225888
rect 312964 225848 341708 225876
rect 312964 225836 312970 225848
rect 341702 225836 341708 225848
rect 341760 225836 341766 225888
rect 341978 225836 341984 225888
rect 342036 225876 342042 225888
rect 365254 225876 365260 225888
rect 342036 225848 365260 225876
rect 342036 225836 342042 225848
rect 365254 225836 365260 225848
rect 365312 225836 365318 225888
rect 375006 225836 375012 225888
rect 375064 225876 375070 225888
rect 387794 225876 387800 225888
rect 375064 225848 387800 225876
rect 375064 225836 375070 225848
rect 387794 225836 387800 225848
rect 387852 225836 387858 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519170 225876 519176 225888
rect 501196 225848 519176 225876
rect 501196 225836 501202 225848
rect 519170 225836 519176 225848
rect 519228 225836 519234 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 672258 225836 672264 225888
rect 672316 225876 672322 225888
rect 672316 225848 672406 225876
rect 672316 225836 672322 225848
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 66162 225700 66168 225752
rect 66220 225740 66226 225752
rect 149790 225740 149796 225752
rect 66220 225712 149796 225740
rect 66220 225700 66226 225712
rect 149790 225700 149796 225712
rect 149848 225700 149854 225752
rect 151262 225700 151268 225752
rect 151320 225740 151326 225752
rect 151320 225712 203380 225740
rect 151320 225700 151326 225712
rect 58986 225564 58992 225616
rect 59044 225604 59050 225616
rect 141510 225604 141516 225616
rect 59044 225576 141516 225604
rect 59044 225564 59050 225576
rect 141510 225564 141516 225576
rect 141568 225564 141574 225616
rect 141786 225564 141792 225616
rect 141844 225604 141850 225616
rect 203150 225604 203156 225616
rect 141844 225576 203156 225604
rect 141844 225564 141850 225576
rect 203150 225564 203156 225576
rect 203208 225564 203214 225616
rect 203352 225604 203380 225712
rect 203886 225700 203892 225752
rect 203944 225740 203950 225752
rect 204714 225740 204720 225752
rect 203944 225712 204720 225740
rect 203944 225700 203950 225712
rect 204714 225700 204720 225712
rect 204772 225700 204778 225752
rect 204898 225700 204904 225752
rect 204956 225740 204962 225752
rect 248874 225740 248880 225752
rect 204956 225712 248880 225740
rect 204956 225700 204962 225712
rect 248874 225700 248880 225712
rect 248932 225700 248938 225752
rect 251082 225700 251088 225752
rect 251140 225740 251146 225752
rect 294414 225740 294420 225752
rect 251140 225712 294420 225740
rect 251140 225700 251146 225712
rect 294414 225700 294420 225712
rect 294472 225700 294478 225752
rect 296438 225700 296444 225752
rect 296496 225740 296502 225752
rect 327902 225740 327908 225752
rect 296496 225712 327908 225740
rect 296496 225700 296502 225712
rect 327902 225700 327908 225712
rect 327960 225700 327966 225752
rect 329742 225700 329748 225752
rect 329800 225740 329806 225752
rect 353662 225740 353668 225752
rect 329800 225712 353668 225740
rect 329800 225700 329806 225712
rect 353662 225700 353668 225712
rect 353720 225700 353726 225752
rect 365346 225700 365352 225752
rect 365404 225740 365410 225752
rect 383286 225740 383292 225752
rect 365404 225712 383292 225740
rect 365404 225700 365410 225712
rect 383286 225700 383292 225712
rect 383344 225700 383350 225752
rect 387702 225700 387708 225752
rect 387760 225740 387766 225752
rect 397822 225740 397828 225752
rect 387760 225712 397828 225740
rect 387760 225700 387766 225712
rect 397822 225700 397828 225712
rect 397880 225700 397886 225752
rect 481174 225700 481180 225752
rect 481232 225740 481238 225752
rect 492674 225740 492680 225752
rect 481232 225712 492680 225740
rect 481232 225700 481238 225712
rect 492674 225700 492680 225712
rect 492732 225700 492738 225752
rect 493594 225700 493600 225752
rect 493652 225740 493658 225752
rect 505370 225740 505376 225752
rect 493652 225712 505376 225740
rect 493652 225700 493658 225712
rect 505370 225700 505376 225712
rect 505428 225700 505434 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563054 225740 563060 225752
rect 535972 225712 563060 225740
rect 535972 225700 535978 225712
rect 563054 225700 563060 225712
rect 563112 225700 563118 225752
rect 217134 225604 217140 225616
rect 203352 225576 217140 225604
rect 217134 225564 217140 225576
rect 217192 225564 217198 225616
rect 220078 225564 220084 225616
rect 220136 225604 220142 225616
rect 266078 225604 266084 225616
rect 220136 225576 266084 225604
rect 220136 225564 220142 225576
rect 266078 225564 266084 225576
rect 266136 225564 266142 225616
rect 266998 225564 267004 225616
rect 267056 225604 267062 225616
rect 274450 225604 274456 225616
rect 267056 225576 274456 225604
rect 267056 225564 267062 225576
rect 274450 225564 274456 225576
rect 274508 225564 274514 225616
rect 278406 225564 278412 225616
rect 278464 225604 278470 225616
rect 313274 225604 313280 225616
rect 278464 225576 313280 225604
rect 278464 225564 278470 225576
rect 313274 225564 313280 225576
rect 313332 225564 313338 225616
rect 327718 225564 327724 225616
rect 327776 225604 327782 225616
rect 352374 225604 352380 225616
rect 327776 225576 352380 225604
rect 327776 225564 327782 225576
rect 352374 225564 352380 225576
rect 352432 225564 352438 225616
rect 352926 225564 352932 225616
rect 352984 225604 352990 225616
rect 371602 225604 371608 225616
rect 352984 225576 371608 225604
rect 352984 225564 352990 225576
rect 371602 225564 371608 225576
rect 371660 225564 371666 225616
rect 382918 225564 382924 225616
rect 382976 225604 382982 225616
rect 396166 225604 396172 225616
rect 382976 225576 396172 225604
rect 382976 225564 382982 225576
rect 396166 225564 396172 225576
rect 396224 225564 396230 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488718 225604 488724 225616
rect 477368 225576 488724 225604
rect 477368 225564 477374 225576
rect 488718 225564 488724 225576
rect 488776 225564 488782 225616
rect 489362 225564 489368 225616
rect 489420 225604 489426 225616
rect 502978 225604 502984 225616
rect 489420 225576 502984 225604
rect 489420 225564 489426 225576
rect 502978 225564 502984 225576
rect 503036 225564 503042 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530578 225604 530584 225616
rect 510212 225576 530584 225604
rect 510212 225564 510218 225576
rect 530578 225564 530584 225576
rect 530636 225564 530642 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558178 225604 558184 225616
rect 531464 225576 558184 225604
rect 531464 225564 531470 225576
rect 558178 225564 558184 225576
rect 558236 225564 558242 225616
rect 672264 225548 672316 225554
rect 672264 225490 672316 225496
rect 125226 225428 125232 225480
rect 125284 225468 125290 225480
rect 196158 225468 196164 225480
rect 125284 225440 196164 225468
rect 125284 225428 125290 225440
rect 196158 225428 196164 225440
rect 196216 225428 196222 225480
rect 197998 225428 198004 225480
rect 198056 225468 198062 225480
rect 204898 225468 204904 225480
rect 198056 225440 204904 225468
rect 198056 225428 198062 225440
rect 204898 225428 204904 225440
rect 204956 225428 204962 225480
rect 209590 225428 209596 225480
rect 209648 225468 209654 225480
rect 259638 225468 259644 225480
rect 209648 225440 259644 225468
rect 209648 225428 209654 225440
rect 259638 225428 259644 225440
rect 259696 225428 259702 225480
rect 297358 225428 297364 225480
rect 297416 225468 297422 225480
rect 310514 225468 310520 225480
rect 297416 225440 310520 225468
rect 297416 225428 297422 225440
rect 310514 225428 310520 225440
rect 310572 225428 310578 225480
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 672156 225344 672208 225350
rect 129366 225292 129372 225344
rect 129424 225332 129430 225344
rect 199102 225332 199108 225344
rect 129424 225304 199108 225332
rect 129424 225292 129430 225304
rect 199102 225292 199108 225304
rect 199160 225292 199166 225344
rect 203150 225292 203156 225344
rect 203208 225332 203214 225344
rect 209406 225332 209412 225344
rect 203208 225304 209412 225332
rect 203208 225292 203214 225304
rect 209406 225292 209412 225304
rect 209464 225292 209470 225344
rect 222930 225332 222936 225344
rect 209746 225304 222936 225332
rect 62022 225156 62028 225208
rect 62080 225196 62086 225208
rect 130378 225196 130384 225208
rect 62080 225168 130384 225196
rect 62080 225156 62086 225168
rect 130378 225156 130384 225168
rect 130436 225156 130442 225208
rect 135070 225156 135076 225208
rect 135128 225196 135134 225208
rect 204254 225196 204260 225208
rect 135128 225168 204260 225196
rect 135128 225156 135134 225168
rect 204254 225156 204260 225168
rect 204312 225156 204318 225208
rect 204530 225156 204536 225208
rect 204588 225196 204594 225208
rect 209746 225196 209774 225304
rect 222930 225292 222936 225304
rect 222988 225292 222994 225344
rect 242894 225292 242900 225344
rect 242952 225332 242958 225344
rect 285030 225332 285036 225344
rect 242952 225304 285036 225332
rect 242952 225292 242958 225304
rect 285030 225292 285036 225304
rect 285088 225292 285094 225344
rect 672156 225286 672208 225292
rect 671246 225224 671252 225276
rect 671304 225264 671310 225276
rect 671304 225236 672060 225264
rect 671304 225224 671310 225236
rect 204588 225168 209774 225196
rect 204588 225156 204594 225168
rect 215202 225156 215208 225208
rect 215260 225196 215266 225208
rect 220078 225196 220084 225208
rect 215260 225168 220084 225196
rect 215260 225156 215266 225168
rect 220078 225156 220084 225168
rect 220136 225156 220142 225208
rect 132402 225020 132408 225072
rect 132460 225060 132466 225072
rect 201678 225060 201684 225072
rect 132460 225032 201684 225060
rect 132460 225020 132466 225032
rect 201678 225020 201684 225032
rect 201736 225020 201742 225072
rect 202598 225020 202604 225072
rect 202656 225060 202662 225072
rect 254486 225060 254492 225072
rect 202656 225032 254492 225060
rect 202656 225020 202662 225032
rect 254486 225020 254492 225032
rect 254544 225020 254550 225072
rect 554958 225020 554964 225072
rect 555016 225060 555022 225072
rect 559098 225060 559104 225072
rect 555016 225032 559104 225060
rect 555016 225020 555022 225032
rect 559098 225020 559104 225032
rect 559156 225020 559162 225072
rect 666462 225020 666468 225072
rect 666520 225060 666526 225072
rect 666520 225032 671968 225060
rect 666520 225020 666526 225032
rect 355226 224952 355232 225004
rect 355284 224992 355290 225004
rect 358170 224992 358176 225004
rect 355284 224964 358176 224992
rect 355284 224952 355290 224964
rect 358170 224952 358176 224964
rect 358228 224952 358234 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 172974 224924 172980 224936
rect 96304 224896 172980 224924
rect 96304 224884 96310 224896
rect 172974 224884 172980 224896
rect 173032 224884 173038 224936
rect 177482 224884 177488 224936
rect 177540 224924 177546 224936
rect 199746 224924 199752 224936
rect 177540 224896 199752 224924
rect 177540 224884 177546 224896
rect 199746 224884 199752 224896
rect 199804 224884 199810 224936
rect 199930 224884 199936 224936
rect 199988 224924 199994 224936
rect 248046 224924 248052 224936
rect 199988 224896 248052 224924
rect 199988 224884 199994 224896
rect 248046 224884 248052 224896
rect 248104 224884 248110 224936
rect 266262 224884 266268 224936
rect 266320 224924 266326 224936
rect 303430 224924 303436 224936
rect 266320 224896 303436 224924
rect 266320 224884 266326 224896
rect 303430 224884 303436 224896
rect 303488 224884 303494 224936
rect 304258 224884 304264 224936
rect 304316 224924 304322 224936
rect 315298 224924 315304 224936
rect 304316 224896 315304 224924
rect 304316 224884 304322 224896
rect 315298 224884 315304 224896
rect 315356 224884 315362 224936
rect 319806 224884 319812 224936
rect 319864 224924 319870 224936
rect 345934 224924 345940 224936
rect 319864 224896 345940 224924
rect 319864 224884 319870 224896
rect 345934 224884 345940 224896
rect 345992 224884 345998 224936
rect 460566 224884 460572 224936
rect 460624 224924 460630 224936
rect 463142 224924 463148 224936
rect 460624 224896 463148 224924
rect 460624 224884 460630 224896
rect 463142 224884 463148 224896
rect 463200 224884 463206 224936
rect 519354 224884 519360 224936
rect 519412 224924 519418 224936
rect 534994 224924 535000 224936
rect 519412 224896 535000 224924
rect 519412 224884 519418 224896
rect 534994 224884 535000 224896
rect 535052 224924 535058 224936
rect 621014 224924 621020 224936
rect 535052 224896 621020 224924
rect 535052 224884 535058 224896
rect 621014 224884 621020 224896
rect 621072 224884 621078 224936
rect 350258 224816 350264 224868
rect 350316 224856 350322 224868
rect 355778 224856 355784 224868
rect 350316 224828 355784 224856
rect 350316 224816 350322 224828
rect 355778 224816 355784 224828
rect 355836 224816 355842 224868
rect 670786 224816 670792 224868
rect 670844 224856 670850 224868
rect 670844 224828 671846 224856
rect 670844 224816 670850 224828
rect 89438 224748 89444 224800
rect 89496 224788 89502 224800
rect 168190 224788 168196 224800
rect 89496 224760 168196 224788
rect 89496 224748 89502 224760
rect 168190 224748 168196 224760
rect 168248 224748 168254 224800
rect 171962 224788 171968 224800
rect 169496 224760 171968 224788
rect 79962 224612 79968 224664
rect 80020 224652 80026 224664
rect 160462 224652 160468 224664
rect 80020 224624 160468 224652
rect 80020 224612 80026 224624
rect 160462 224612 160468 224624
rect 160520 224612 160526 224664
rect 165154 224612 165160 224664
rect 165212 224652 165218 224664
rect 169496 224652 169524 224760
rect 171962 224748 171968 224760
rect 172020 224748 172026 224800
rect 172146 224748 172152 224800
rect 172204 224788 172210 224800
rect 178954 224788 178960 224800
rect 172204 224760 178960 224788
rect 172204 224748 172210 224760
rect 178954 224748 178960 224760
rect 179012 224748 179018 224800
rect 179322 224748 179328 224800
rect 179380 224788 179386 224800
rect 237742 224788 237748 224800
rect 179380 224760 237748 224788
rect 179380 224748 179386 224760
rect 237742 224748 237748 224760
rect 237800 224748 237806 224800
rect 248322 224748 248328 224800
rect 248380 224788 248386 224800
rect 291838 224788 291844 224800
rect 248380 224760 291844 224788
rect 248380 224748 248386 224760
rect 291838 224748 291844 224760
rect 291896 224748 291902 224800
rect 294874 224748 294880 224800
rect 294932 224788 294938 224800
rect 325970 224788 325976 224800
rect 294932 224760 325976 224788
rect 294932 224748 294938 224760
rect 325970 224748 325976 224760
rect 326028 224748 326034 224800
rect 331858 224748 331864 224800
rect 331916 224788 331922 224800
rect 337562 224788 337568 224800
rect 331916 224760 337568 224788
rect 331916 224748 331922 224760
rect 337562 224748 337568 224760
rect 337620 224748 337626 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526346 224788 526352 224800
rect 506992 224760 526352 224788
rect 506992 224748 506998 224760
rect 526346 224748 526352 224760
rect 526404 224748 526410 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 529992 224760 547874 224788
rect 529992 224748 529998 224760
rect 224862 224652 224868 224664
rect 165212 224624 169524 224652
rect 169588 224624 224868 224652
rect 165212 224612 165218 224624
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 169588 224516 169616 224624
rect 224862 224612 224868 224624
rect 224920 224612 224926 224664
rect 227530 224612 227536 224664
rect 227588 224652 227594 224664
rect 272334 224652 272340 224664
rect 227588 224624 272340 224652
rect 227588 224612 227594 224624
rect 272334 224612 272340 224624
rect 272392 224612 272398 224664
rect 272518 224612 272524 224664
rect 272576 224652 272582 224664
rect 309870 224652 309876 224664
rect 272576 224624 309876 224652
rect 272576 224612 272582 224624
rect 309870 224612 309876 224624
rect 309928 224612 309934 224664
rect 311526 224612 311532 224664
rect 311584 224652 311590 224664
rect 338850 224652 338856 224664
rect 311584 224624 338856 224652
rect 311584 224612 311590 224624
rect 338850 224612 338856 224624
rect 338908 224612 338914 224664
rect 346302 224612 346308 224664
rect 346360 224652 346366 224664
rect 366542 224652 366548 224664
rect 346360 224624 366548 224652
rect 346360 224612 346366 224624
rect 366542 224612 366548 224624
rect 366600 224612 366606 224664
rect 494054 224612 494060 224664
rect 494112 224652 494118 224664
rect 510154 224652 510160 224664
rect 494112 224624 510160 224652
rect 494112 224612 494118 224624
rect 510154 224612 510160 224624
rect 510212 224612 510218 224664
rect 520458 224612 520464 224664
rect 520516 224652 520522 224664
rect 544102 224652 544108 224664
rect 520516 224624 544108 224652
rect 520516 224612 520522 224624
rect 544102 224612 544108 224624
rect 544160 224612 544166 224664
rect 547846 224652 547874 224760
rect 548334 224748 548340 224800
rect 548392 224788 548398 224800
rect 550818 224788 550824 224800
rect 548392 224760 550824 224788
rect 548392 224748 548398 224760
rect 550818 224748 550824 224760
rect 550876 224748 550882 224800
rect 555786 224788 555792 224800
rect 553366 224760 555792 224788
rect 549070 224652 549076 224664
rect 547846 224624 549076 224652
rect 549070 224612 549076 224624
rect 549128 224612 549134 224664
rect 549254 224612 549260 224664
rect 549312 224652 549318 224664
rect 553366 224652 553394 224760
rect 555786 224748 555792 224760
rect 555844 224748 555850 224800
rect 556154 224748 556160 224800
rect 556212 224788 556218 224800
rect 557350 224788 557356 224800
rect 556212 224760 557356 224788
rect 556212 224748 556218 224760
rect 557350 224748 557356 224760
rect 557408 224788 557414 224800
rect 558822 224788 558828 224800
rect 557408 224760 558828 224788
rect 557408 224748 557414 224760
rect 558822 224748 558828 224760
rect 558880 224748 558886 224800
rect 559098 224748 559104 224800
rect 559156 224788 559162 224800
rect 559156 224760 562456 224788
rect 559156 224748 559162 224760
rect 562428 224720 562456 224760
rect 562686 224748 562692 224800
rect 562744 224788 562750 224800
rect 571518 224788 571524 224800
rect 562744 224760 571524 224788
rect 562744 224748 562750 224760
rect 571518 224748 571524 224760
rect 571576 224748 571582 224800
rect 610986 224788 610992 224800
rect 605806 224760 610992 224788
rect 562428 224692 562548 224720
rect 549312 224624 553394 224652
rect 549312 224612 549318 224624
rect 557810 224612 557816 224664
rect 557868 224652 557874 224664
rect 562134 224652 562140 224664
rect 557868 224624 562140 224652
rect 557868 224612 557874 224624
rect 562134 224612 562140 224624
rect 562192 224612 562198 224664
rect 562520 224652 562548 224692
rect 605806 224652 605834 224760
rect 610986 224748 610992 224760
rect 611044 224748 611050 224800
rect 562520 224624 605834 224652
rect 610618 224612 610624 224664
rect 610676 224652 610682 224664
rect 617058 224652 617064 224664
rect 610676 224624 617064 224652
rect 610676 224612 610682 224624
rect 617058 224612 617064 224624
rect 617116 224612 617122 224664
rect 671712 224528 671764 224534
rect 165770 224488 169616 224516
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 155310 224380 155316 224392
rect 73764 224352 155316 224380
rect 73764 224340 73770 224352
rect 155310 224340 155316 224352
rect 155368 224340 155374 224392
rect 156690 224340 156696 224392
rect 156748 224380 156754 224392
rect 157334 224380 157340 224392
rect 156748 224352 157340 224380
rect 156748 224340 156754 224352
rect 157334 224340 157340 224352
rect 157392 224340 157398 224392
rect 161658 224340 161664 224392
rect 161716 224380 161722 224392
rect 165770 224380 165798 224488
rect 171594 224476 171600 224528
rect 171652 224516 171658 224528
rect 178494 224516 178500 224528
rect 171652 224488 178500 224516
rect 171652 224476 171658 224488
rect 178494 224476 178500 224488
rect 178552 224476 178558 224528
rect 178954 224476 178960 224528
rect 179012 224516 179018 224528
rect 232590 224516 232596 224528
rect 179012 224488 232596 224516
rect 179012 224476 179018 224488
rect 232590 224476 232596 224488
rect 232648 224476 232654 224528
rect 233142 224476 233148 224528
rect 233200 224516 233206 224528
rect 272334 224516 272340 224528
rect 233200 224488 272340 224516
rect 233200 224476 233206 224488
rect 272334 224476 272340 224488
rect 272392 224476 272398 224528
rect 275094 224516 275100 224528
rect 272628 224488 275100 224516
rect 161716 224352 165798 224380
rect 161716 224340 161722 224352
rect 165982 224340 165988 224392
rect 166040 224380 166046 224392
rect 171778 224380 171784 224392
rect 166040 224352 171784 224380
rect 166040 224340 166046 224352
rect 171778 224340 171784 224352
rect 171836 224340 171842 224392
rect 171962 224340 171968 224392
rect 172020 224380 172026 224392
rect 227070 224380 227076 224392
rect 172020 224352 227076 224380
rect 172020 224340 172026 224352
rect 227070 224340 227076 224352
rect 227128 224340 227134 224392
rect 228726 224340 228732 224392
rect 228784 224380 228790 224392
rect 272628 224380 272656 224488
rect 275094 224476 275100 224488
rect 275152 224476 275158 224528
rect 286318 224476 286324 224528
rect 286376 224516 286382 224528
rect 289906 224516 289912 224528
rect 286376 224488 289912 224516
rect 286376 224476 286382 224488
rect 289906 224476 289912 224488
rect 289964 224476 289970 224528
rect 290826 224476 290832 224528
rect 290884 224516 290890 224528
rect 324038 224516 324044 224528
rect 290884 224488 324044 224516
rect 290884 224476 290890 224488
rect 324038 224476 324044 224488
rect 324096 224476 324102 224528
rect 342162 224476 342168 224528
rect 342220 224516 342226 224528
rect 362034 224516 362040 224528
rect 342220 224488 362040 224516
rect 342220 224476 342226 224488
rect 362034 224476 362040 224488
rect 362092 224476 362098 224528
rect 366726 224476 366732 224528
rect 366784 224516 366790 224528
rect 381630 224516 381636 224528
rect 366784 224488 381636 224516
rect 366784 224476 366790 224488
rect 381630 224476 381636 224488
rect 381688 224476 381694 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506014 224516 506020 224528
rect 491352 224488 506020 224516
rect 491352 224476 491358 224488
rect 506014 224476 506020 224488
rect 506072 224476 506078 224528
rect 535270 224476 535276 224528
rect 535328 224516 535334 224528
rect 562134 224516 562140 224528
rect 535328 224488 562140 224516
rect 535328 224476 535334 224488
rect 562134 224476 562140 224488
rect 562192 224476 562198 224528
rect 562318 224476 562324 224528
rect 562376 224516 562382 224528
rect 610802 224516 610808 224528
rect 562376 224488 610808 224516
rect 562376 224476 562382 224488
rect 610802 224476 610808 224488
rect 610860 224476 610866 224528
rect 671712 224470 671764 224476
rect 670602 224408 670608 224460
rect 670660 224448 670666 224460
rect 670660 224420 671622 224448
rect 670660 224408 670666 224420
rect 228784 224352 272656 224380
rect 228784 224340 228790 224352
rect 275094 224340 275100 224392
rect 275152 224380 275158 224392
rect 311158 224380 311164 224392
rect 275152 224352 311164 224380
rect 275152 224340 275158 224352
rect 311158 224340 311164 224352
rect 311216 224340 311222 224392
rect 322842 224340 322848 224392
rect 322900 224380 322906 224392
rect 349798 224380 349804 224392
rect 322900 224352 349804 224380
rect 322900 224340 322906 224352
rect 349798 224340 349804 224352
rect 349856 224340 349862 224392
rect 359458 224340 359464 224392
rect 359516 224380 359522 224392
rect 378134 224380 378140 224392
rect 359516 224352 378140 224380
rect 359516 224340 359522 224352
rect 378134 224340 378140 224352
rect 378192 224340 378198 224392
rect 379238 224340 379244 224392
rect 379296 224380 379302 224392
rect 393590 224380 393596 224392
rect 379296 224352 393596 224380
rect 379296 224340 379302 224352
rect 393590 224340 393596 224352
rect 393648 224340 393654 224392
rect 394510 224340 394516 224392
rect 394568 224380 394574 224392
rect 404538 224380 404544 224392
rect 394568 224352 404544 224380
rect 394568 224340 394574 224352
rect 404538 224340 404544 224352
rect 404596 224340 404602 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492858 224380 492864 224392
rect 480588 224352 492864 224380
rect 480588 224340 480594 224352
rect 492858 224340 492864 224352
rect 492916 224340 492922 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516594 224380 516600 224392
rect 499264 224352 516600 224380
rect 499264 224340 499270 224352
rect 516594 224340 516600 224352
rect 516652 224340 516658 224392
rect 525518 224340 525524 224392
rect 525576 224380 525582 224392
rect 548334 224380 548340 224392
rect 525576 224352 548340 224380
rect 525576 224340 525582 224352
rect 548334 224340 548340 224352
rect 548392 224340 548398 224392
rect 548518 224340 548524 224392
rect 548576 224380 548582 224392
rect 558178 224380 558184 224392
rect 548576 224352 558184 224380
rect 548576 224340 548582 224352
rect 558178 224340 558184 224352
rect 558236 224340 558242 224392
rect 558822 224340 558828 224392
rect 558880 224380 558886 224392
rect 626534 224380 626540 224392
rect 558880 224352 626540 224380
rect 558880 224340 558886 224352
rect 626534 224340 626540 224352
rect 626592 224340 626598 224392
rect 68922 224204 68928 224256
rect 68980 224244 68986 224256
rect 152734 224244 152740 224256
rect 68980 224216 152740 224244
rect 68980 224204 68986 224216
rect 152734 224204 152740 224216
rect 152792 224204 152798 224256
rect 155770 224204 155776 224256
rect 155828 224244 155834 224256
rect 160186 224244 160192 224256
rect 155828 224216 160192 224244
rect 155828 224204 155834 224216
rect 160186 224204 160192 224216
rect 160244 224204 160250 224256
rect 168282 224204 168288 224256
rect 168340 224244 168346 224256
rect 230014 224244 230020 224256
rect 168340 224216 230020 224244
rect 168340 224204 168346 224216
rect 230014 224204 230020 224216
rect 230072 224204 230078 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 231728 224216 258074 224244
rect 231728 224204 231734 224216
rect 102042 224068 102048 224120
rect 102100 224108 102106 224120
rect 171594 224108 171600 224120
rect 102100 224080 171600 224108
rect 102100 224068 102106 224080
rect 171594 224068 171600 224080
rect 171652 224068 171658 224120
rect 171778 224068 171784 224120
rect 171836 224108 171842 224120
rect 194594 224108 194600 224120
rect 171836 224080 194600 224108
rect 171836 224068 171842 224080
rect 194594 224068 194600 224080
rect 194652 224068 194658 224120
rect 194778 224068 194784 224120
rect 194836 224108 194842 224120
rect 250622 224108 250628 224120
rect 194836 224080 250628 224108
rect 194836 224068 194842 224080
rect 250622 224068 250628 224080
rect 250680 224068 250686 224120
rect 258046 224108 258074 224216
rect 272334 224204 272340 224256
rect 272392 224244 272398 224256
rect 277670 224244 277676 224256
rect 272392 224216 277676 224244
rect 272392 224204 272398 224216
rect 277670 224204 277676 224216
rect 277728 224204 277734 224256
rect 289722 224204 289728 224256
rect 289780 224244 289786 224256
rect 296990 224244 296996 224256
rect 289780 224216 296996 224244
rect 289780 224204 289786 224216
rect 296990 224204 296996 224216
rect 297048 224204 297054 224256
rect 299106 224204 299112 224256
rect 299164 224244 299170 224256
rect 331398 224244 331404 224256
rect 299164 224216 331404 224244
rect 299164 224204 299170 224216
rect 331398 224204 331404 224216
rect 331456 224204 331462 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 362310 224244 362316 224256
rect 339460 224216 362316 224244
rect 339460 224204 339466 224216
rect 362310 224204 362316 224216
rect 362368 224204 362374 224256
rect 372522 224204 372528 224256
rect 372580 224244 372586 224256
rect 387426 224244 387432 224256
rect 372580 224216 387432 224244
rect 372580 224204 372586 224216
rect 387426 224204 387432 224216
rect 387484 224204 387490 224256
rect 390186 224204 390192 224256
rect 390244 224244 390250 224256
rect 401962 224244 401968 224256
rect 390244 224216 401968 224244
rect 390244 224204 390250 224216
rect 401962 224204 401968 224216
rect 402020 224204 402026 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 427906 224204 427912 224256
rect 427964 224244 427970 224256
rect 428734 224244 428740 224256
rect 427964 224216 428740 224244
rect 427964 224204 427970 224216
rect 428734 224204 428740 224216
rect 428792 224204 428798 224256
rect 451366 224204 451372 224256
rect 451424 224244 451430 224256
rect 452194 224244 452200 224256
rect 451424 224216 452200 224244
rect 451424 224204 451430 224216
rect 452194 224204 452200 224216
rect 452252 224204 452258 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480346 224244 480352 224256
rect 470284 224216 480352 224244
rect 470284 224204 470290 224216
rect 480346 224204 480352 224216
rect 480404 224204 480410 224256
rect 483750 224204 483756 224256
rect 483808 224244 483814 224256
rect 496906 224244 496912 224256
rect 483808 224216 496912 224244
rect 483808 224204 483814 224216
rect 496906 224204 496912 224216
rect 496964 224204 496970 224256
rect 523494 224244 523500 224256
rect 505066 224216 523500 224244
rect 278958 224108 278964 224120
rect 258046 224080 278964 224108
rect 278958 224068 278964 224080
rect 279016 224068 279022 224120
rect 504358 224068 504364 224120
rect 504416 224108 504422 224120
rect 505066 224108 505094 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 524414 224204 524420 224256
rect 524472 224244 524478 224256
rect 525058 224244 525064 224256
rect 524472 224216 525064 224244
rect 524472 224204 524478 224216
rect 525058 224204 525064 224216
rect 525116 224244 525122 224256
rect 619634 224244 619640 224256
rect 525116 224216 619640 224244
rect 525116 224204 525122 224216
rect 619634 224204 619640 224216
rect 619692 224204 619698 224256
rect 651282 224204 651288 224256
rect 651340 224244 651346 224256
rect 666462 224244 666468 224256
rect 651340 224216 666468 224244
rect 651340 224204 651346 224216
rect 666462 224204 666468 224216
rect 666520 224204 666526 224256
rect 668026 224204 668032 224256
rect 668084 224244 668090 224256
rect 668084 224216 671508 224244
rect 668084 224204 668090 224216
rect 620186 224136 620192 224188
rect 620244 224176 620250 224188
rect 625430 224176 625436 224188
rect 620244 224148 625436 224176
rect 620244 224136 620250 224148
rect 625430 224136 625436 224148
rect 625488 224136 625494 224188
rect 504416 224080 505094 224108
rect 504416 224068 504422 224080
rect 667842 224068 667848 224120
rect 667900 224108 667906 224120
rect 667900 224080 670740 224108
rect 667900 224068 667906 224080
rect 279418 224000 279424 224052
rect 279476 224040 279482 224052
rect 284754 224040 284760 224052
rect 279476 224012 284760 224040
rect 279476 224000 279482 224012
rect 284754 224000 284760 224012
rect 284812 224000 284818 224052
rect 517698 224000 517704 224052
rect 517756 224040 517762 224052
rect 610618 224040 610624 224052
rect 517756 224012 610624 224040
rect 517756 224000 517762 224012
rect 610618 224000 610624 224012
rect 610676 224000 610682 224052
rect 610986 224000 610992 224052
rect 611044 224040 611050 224052
rect 670712 224040 670740 224080
rect 611044 224012 620416 224040
rect 670712 224012 671398 224040
rect 611044 224000 611050 224012
rect 105998 223932 106004 223984
rect 106056 223972 106062 223984
rect 181070 223972 181076 223984
rect 106056 223944 181076 223972
rect 106056 223932 106062 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 191558 223932 191564 223984
rect 191616 223972 191622 223984
rect 199838 223972 199844 223984
rect 191616 223944 199844 223972
rect 191616 223932 191622 223944
rect 199838 223932 199844 223944
rect 199896 223932 199902 223984
rect 201402 223932 201408 223984
rect 201460 223972 201466 223984
rect 255774 223972 255780 223984
rect 201460 223944 255780 223972
rect 201460 223932 201466 223944
rect 255774 223932 255780 223944
rect 255832 223932 255838 223984
rect 515950 223864 515956 223916
rect 516008 223904 516014 223916
rect 538490 223904 538496 223916
rect 516008 223876 538496 223904
rect 516008 223864 516014 223876
rect 538490 223864 538496 223876
rect 538548 223904 538554 223916
rect 539502 223904 539508 223916
rect 538548 223876 539508 223904
rect 538548 223864 538554 223876
rect 539502 223864 539508 223876
rect 539560 223864 539566 223916
rect 542446 223864 542452 223916
rect 542504 223904 542510 223916
rect 548518 223904 548524 223916
rect 542504 223876 548524 223904
rect 542504 223864 542510 223876
rect 548518 223864 548524 223876
rect 548576 223864 548582 223916
rect 549254 223864 549260 223916
rect 549312 223904 549318 223916
rect 549898 223904 549904 223916
rect 549312 223876 549904 223904
rect 549312 223864 549318 223876
rect 549898 223864 549904 223876
rect 549956 223904 549962 223916
rect 557810 223904 557816 223916
rect 549956 223876 557816 223904
rect 549956 223864 549962 223876
rect 557810 223864 557816 223876
rect 557868 223864 557874 223916
rect 558178 223864 558184 223916
rect 558236 223904 558242 223916
rect 610618 223904 610624 223916
rect 558236 223876 610624 223904
rect 558236 223864 558242 223876
rect 610618 223864 610624 223876
rect 610676 223864 610682 223916
rect 610802 223864 610808 223916
rect 610860 223904 610866 223916
rect 620186 223904 620192 223916
rect 610860 223876 620192 223904
rect 610860 223864 610866 223876
rect 620186 223864 620192 223876
rect 620244 223864 620250 223916
rect 620388 223904 620416 224012
rect 625246 223904 625252 223916
rect 620388 223876 625252 223904
rect 625246 223864 625252 223876
rect 625304 223864 625310 223916
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183646 223836 183652 223848
rect 108724 223808 183652 223836
rect 108724 223796 108730 223808
rect 183646 223796 183652 223808
rect 183704 223796 183710 223848
rect 184382 223796 184388 223848
rect 184440 223836 184446 223848
rect 207474 223836 207480 223848
rect 184440 223808 207480 223836
rect 184440 223796 184446 223808
rect 207474 223796 207480 223808
rect 207532 223796 207538 223848
rect 207658 223796 207664 223848
rect 207716 223836 207722 223848
rect 228082 223836 228088 223848
rect 207716 223808 228088 223836
rect 207716 223796 207722 223808
rect 228082 223796 228088 223808
rect 228140 223796 228146 223848
rect 245470 223796 245476 223848
rect 245528 223836 245534 223848
rect 287606 223836 287612 223848
rect 245528 223808 287612 223836
rect 245528 223796 245534 223808
rect 287606 223796 287612 223808
rect 287664 223796 287670 223848
rect 670712 223808 671278 223836
rect 505186 223728 505192 223780
rect 505244 223768 505250 223780
rect 507670 223768 507676 223780
rect 505244 223740 507676 223768
rect 505244 223728 505250 223740
rect 507670 223728 507676 223740
rect 507728 223728 507734 223780
rect 539962 223728 539968 223780
rect 540020 223768 540026 223780
rect 622670 223768 622676 223780
rect 540020 223740 622676 223768
rect 540020 223728 540026 223740
rect 622670 223728 622676 223740
rect 622728 223728 622734 223780
rect 670712 223768 670740 223808
rect 670620 223740 670740 223768
rect 115290 223660 115296 223712
rect 115348 223700 115354 223712
rect 188798 223700 188804 223712
rect 115348 223672 188804 223700
rect 115348 223660 115354 223672
rect 188798 223660 188804 223672
rect 188856 223660 188862 223712
rect 505370 223592 505376 223644
rect 505428 223632 505434 223644
rect 505428 223604 610480 223632
rect 505428 223592 505434 223604
rect 99282 223524 99288 223576
rect 99340 223564 99346 223576
rect 175734 223564 175740 223576
rect 99340 223536 175740 223564
rect 99340 223524 99346 223536
rect 175734 223524 175740 223536
rect 175792 223524 175798 223576
rect 183186 223524 183192 223576
rect 183244 223564 183250 223576
rect 184658 223564 184664 223576
rect 183244 223536 184664 223564
rect 183244 223524 183250 223536
rect 184658 223524 184664 223536
rect 184716 223524 184722 223576
rect 187326 223524 187332 223576
rect 187384 223564 187390 223576
rect 242250 223564 242256 223576
rect 187384 223536 242256 223564
rect 187384 223524 187390 223536
rect 242250 223524 242256 223536
rect 242308 223524 242314 223576
rect 249426 223524 249432 223576
rect 249484 223564 249490 223576
rect 276290 223564 276296 223576
rect 249484 223536 276296 223564
rect 249484 223524 249490 223536
rect 276290 223524 276296 223536
rect 276348 223524 276354 223576
rect 278590 223524 278596 223576
rect 278648 223564 278654 223576
rect 315022 223564 315028 223576
rect 278648 223536 315028 223564
rect 278648 223524 278654 223536
rect 315022 223524 315028 223536
rect 315080 223524 315086 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 610452 223496 610480 223604
rect 610618 223592 610624 223644
rect 610676 223632 610682 223644
rect 622486 223632 622492 223644
rect 610676 223604 622492 223632
rect 610676 223592 610682 223604
rect 622486 223592 622492 223604
rect 622544 223592 622550 223644
rect 614942 223496 614948 223508
rect 610452 223468 614948 223496
rect 614942 223456 614948 223468
rect 615000 223456 615006 223508
rect 81342 223388 81348 223440
rect 81400 223428 81406 223440
rect 157242 223428 157248 223440
rect 81400 223400 157248 223428
rect 81400 223388 81406 223400
rect 157242 223388 157248 223400
rect 157300 223388 157306 223440
rect 157426 223388 157432 223440
rect 157484 223428 157490 223440
rect 159818 223428 159824 223440
rect 157484 223400 159824 223428
rect 157484 223388 157490 223400
rect 159818 223388 159824 223400
rect 159876 223388 159882 223440
rect 162118 223388 162124 223440
rect 162176 223428 162182 223440
rect 162176 223400 166994 223428
rect 162176 223388 162182 223400
rect 85298 223252 85304 223304
rect 85356 223292 85362 223304
rect 162394 223292 162400 223304
rect 85356 223264 162400 223292
rect 85356 223252 85362 223264
rect 162394 223252 162400 223264
rect 162452 223252 162458 223304
rect 166966 223292 166994 223400
rect 171778 223388 171784 223440
rect 171836 223428 171842 223440
rect 181714 223428 181720 223440
rect 171836 223400 181720 223428
rect 171836 223388 171842 223400
rect 181714 223388 181720 223400
rect 181772 223388 181778 223440
rect 184842 223388 184848 223440
rect 184900 223428 184906 223440
rect 239674 223428 239680 223440
rect 184900 223400 239680 223428
rect 184900 223388 184906 223400
rect 239674 223388 239680 223400
rect 239732 223388 239738 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 291194 223428 291200 223440
rect 287026 223400 291200 223428
rect 186866 223292 186872 223304
rect 166966 223264 186872 223292
rect 186866 223252 186872 223264
rect 186924 223252 186930 223304
rect 188154 223252 188160 223304
rect 188212 223292 188218 223304
rect 245102 223292 245108 223304
rect 188212 223264 245108 223292
rect 188212 223252 188218 223264
rect 245102 223252 245108 223264
rect 245160 223252 245166 223304
rect 250898 223252 250904 223304
rect 250956 223292 250962 223304
rect 287026 223292 287054 223400
rect 291194 223388 291200 223400
rect 291252 223388 291258 223440
rect 316678 223388 316684 223440
rect 316736 223428 316742 223440
rect 327258 223428 327264 223440
rect 316736 223400 327264 223428
rect 316736 223388 316742 223400
rect 327258 223388 327264 223400
rect 327316 223388 327322 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 532510 223428 532516 223440
rect 517572 223400 532516 223428
rect 517572 223388 517578 223400
rect 532510 223388 532516 223400
rect 532568 223388 532574 223440
rect 534810 223388 534816 223440
rect 534868 223428 534874 223440
rect 547506 223428 547512 223440
rect 534868 223400 547512 223428
rect 534868 223388 534874 223400
rect 547506 223388 547512 223400
rect 547564 223388 547570 223440
rect 297542 223320 297548 223372
rect 297600 223360 297606 223372
rect 305362 223360 305368 223372
rect 297600 223332 305368 223360
rect 297600 223320 297606 223332
rect 305362 223320 305368 223332
rect 305420 223320 305426 223372
rect 250956 223264 287054 223292
rect 250956 223252 250962 223264
rect 288986 223252 288992 223304
rect 289044 223292 289050 223304
rect 295058 223292 295064 223304
rect 289044 223264 295064 223292
rect 289044 223252 289050 223264
rect 295058 223252 295064 223264
rect 295116 223252 295122 223304
rect 307662 223252 307668 223304
rect 307720 223292 307726 223304
rect 335630 223292 335636 223304
rect 307720 223264 335636 223292
rect 307720 223252 307726 223264
rect 335630 223252 335636 223264
rect 335688 223252 335694 223304
rect 337930 223252 337936 223304
rect 337988 223292 337994 223304
rect 359182 223292 359188 223304
rect 337988 223264 359188 223292
rect 337988 223252 337994 223264
rect 359182 223252 359188 223264
rect 359240 223252 359246 223304
rect 493042 223252 493048 223304
rect 493100 223292 493106 223304
rect 508498 223292 508504 223304
rect 493100 223264 508504 223292
rect 493100 223252 493106 223264
rect 508498 223252 508504 223264
rect 508556 223252 508562 223304
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 535454 223292 535460 223304
rect 514720 223264 535460 223292
rect 514720 223252 514726 223264
rect 535454 223252 535460 223264
rect 535512 223252 535518 223304
rect 68738 223116 68744 223168
rect 68796 223156 68802 223168
rect 146570 223156 146576 223168
rect 68796 223128 146576 223156
rect 68796 223116 68802 223128
rect 146570 223116 146576 223128
rect 146628 223116 146634 223168
rect 146754 223116 146760 223168
rect 146812 223156 146818 223168
rect 147628 223156 147634 223168
rect 146812 223128 147634 223156
rect 146812 223116 146818 223128
rect 147628 223116 147634 223128
rect 147686 223116 147692 223168
rect 147766 223116 147772 223168
rect 147824 223156 147830 223168
rect 176286 223156 176292 223168
rect 147824 223128 176292 223156
rect 147824 223116 147830 223128
rect 176286 223116 176292 223128
rect 176344 223116 176350 223168
rect 181990 223116 181996 223168
rect 182048 223156 182054 223168
rect 240318 223156 240324 223168
rect 182048 223128 240324 223156
rect 182048 223116 182054 223128
rect 240318 223116 240324 223128
rect 240376 223116 240382 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321462 223156 321468 223168
rect 288308 223128 321468 223156
rect 288308 223116 288314 223128
rect 321462 223116 321468 223128
rect 321520 223116 321526 223168
rect 323946 223116 323952 223168
rect 324004 223156 324010 223168
rect 348510 223156 348516 223168
rect 324004 223128 348516 223156
rect 324004 223116 324010 223128
rect 348510 223116 348516 223128
rect 348568 223116 348574 223168
rect 358538 223116 358544 223168
rect 358596 223156 358602 223168
rect 374638 223156 374644 223168
rect 358596 223128 374644 223156
rect 358596 223116 358602 223128
rect 374638 223116 374644 223128
rect 374696 223116 374702 223168
rect 483106 223116 483112 223168
rect 483164 223156 483170 223168
rect 496078 223156 496084 223168
rect 483164 223128 496084 223156
rect 483164 223116 483170 223128
rect 496078 223116 496084 223128
rect 496136 223116 496142 223168
rect 503346 223116 503352 223168
rect 503404 223156 503410 223168
rect 521746 223156 521752 223168
rect 503404 223128 521752 223156
rect 503404 223116 503410 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 529474 223116 529480 223168
rect 529532 223156 529538 223168
rect 555694 223156 555700 223168
rect 529532 223128 555700 223156
rect 529532 223116 529538 223128
rect 555694 223116 555700 223128
rect 555752 223116 555758 223168
rect 557534 223116 557540 223168
rect 557592 223156 557598 223168
rect 559926 223156 559932 223168
rect 557592 223128 559932 223156
rect 557592 223116 557598 223128
rect 559926 223116 559932 223128
rect 559984 223156 559990 223168
rect 562870 223156 562876 223168
rect 559984 223128 562876 223156
rect 559984 223116 559990 223128
rect 562870 223116 562876 223128
rect 562928 223116 562934 223168
rect 75822 222980 75828 223032
rect 75880 223020 75886 223032
rect 154942 223020 154948 223032
rect 75880 222992 154948 223020
rect 75880 222980 75886 222992
rect 154942 222980 154948 222992
rect 155000 222980 155006 223032
rect 155126 222980 155132 223032
rect 155184 223020 155190 223032
rect 155184 222992 157334 223020
rect 155184 222980 155190 222992
rect 71406 222844 71412 222896
rect 71464 222884 71470 222896
rect 152090 222884 152096 222896
rect 71464 222856 152096 222884
rect 71464 222844 71470 222856
rect 152090 222844 152096 222856
rect 152148 222844 152154 222896
rect 152274 222844 152280 222896
rect 152332 222884 152338 222896
rect 155494 222884 155500 222896
rect 152332 222856 155500 222884
rect 152332 222844 152338 222856
rect 155494 222844 155500 222856
rect 155552 222844 155558 222896
rect 157306 222884 157334 222992
rect 157518 222980 157524 223032
rect 157576 223020 157582 223032
rect 219066 223020 219072 223032
rect 157576 222992 219072 223020
rect 157576 222980 157582 222992
rect 219066 222980 219072 222992
rect 219124 222980 219130 223032
rect 245286 222980 245292 223032
rect 245344 223020 245350 223032
rect 289262 223020 289268 223032
rect 245344 222992 289268 223020
rect 245344 222980 245350 222992
rect 289262 222980 289268 222992
rect 289320 222980 289326 223032
rect 291470 222980 291476 223032
rect 291528 223020 291534 223032
rect 300210 223020 300216 223032
rect 291528 222992 300216 223020
rect 291528 222980 291534 222992
rect 300210 222980 300216 222992
rect 300268 222980 300274 223032
rect 315666 222980 315672 223032
rect 315724 223020 315730 223032
rect 344646 223020 344652 223032
rect 315724 222992 344652 223020
rect 315724 222980 315730 222992
rect 344646 222980 344652 222992
rect 344704 222980 344710 223032
rect 349062 222980 349068 223032
rect 349120 223020 349126 223032
rect 367186 223020 367192 223032
rect 349120 222992 367192 223020
rect 349120 222980 349126 222992
rect 367186 222980 367192 222992
rect 367244 222980 367250 223032
rect 368382 222980 368388 223032
rect 368440 223020 368446 223032
rect 382642 223020 382648 223032
rect 368440 222992 382648 223020
rect 368440 222980 368446 222992
rect 382642 222980 382648 222992
rect 382700 222980 382706 223032
rect 383562 222980 383568 223032
rect 383620 223020 383626 223032
rect 394878 223020 394884 223032
rect 383620 222992 394884 223020
rect 383620 222980 383626 222992
rect 394878 222980 394884 222992
rect 394936 222980 394942 223032
rect 486602 222980 486608 223032
rect 486660 223020 486666 223032
rect 500034 223020 500040 223032
rect 486660 222992 500040 223020
rect 486660 222980 486666 222992
rect 500034 222980 500040 222992
rect 500092 222980 500098 223032
rect 508222 222980 508228 223032
rect 508280 223020 508286 223032
rect 527174 223020 527180 223032
rect 508280 222992 527180 223020
rect 508280 222980 508286 222992
rect 527174 222980 527180 222992
rect 527232 222980 527238 223032
rect 532050 222980 532056 223032
rect 532108 223020 532114 223032
rect 559006 223020 559012 223032
rect 532108 222992 559012 223020
rect 532108 222980 532114 222992
rect 559006 222980 559012 222992
rect 559064 222980 559070 223032
rect 171778 222884 171784 222896
rect 157306 222856 171784 222884
rect 171778 222844 171784 222856
rect 171836 222844 171842 222896
rect 172882 222844 172888 222896
rect 172940 222884 172946 222896
rect 212626 222884 212632 222896
rect 172940 222856 212632 222884
rect 172940 222844 172946 222856
rect 212626 222844 212632 222856
rect 212684 222844 212690 222896
rect 213178 222844 213184 222896
rect 213236 222884 213242 222896
rect 233326 222884 233332 222896
rect 213236 222856 233332 222884
rect 213236 222844 213242 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282730 222844 282736 222896
rect 282788 222884 282794 222896
rect 316310 222884 316316 222896
rect 282788 222856 316316 222884
rect 282788 222844 282794 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 321462 222844 321468 222896
rect 321520 222884 321526 222896
rect 346578 222884 346584 222896
rect 321520 222856 346584 222884
rect 321520 222844 321526 222856
rect 346578 222844 346584 222856
rect 346636 222844 346642 222896
rect 347222 222844 347228 222896
rect 347280 222884 347286 222896
rect 367830 222884 367836 222896
rect 347280 222856 367836 222884
rect 347280 222844 347286 222856
rect 367830 222844 367836 222856
rect 367888 222844 367894 222896
rect 375190 222844 375196 222896
rect 375248 222884 375254 222896
rect 391014 222884 391020 222896
rect 375248 222856 391020 222884
rect 375248 222844 375254 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 492030 222884 492036 222896
rect 479944 222856 492036 222884
rect 479944 222844 479950 222856
rect 492030 222844 492036 222856
rect 492088 222844 492094 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 543366 222884 543372 222896
rect 519872 222856 543372 222884
rect 519872 222844 519878 222856
rect 543366 222844 543372 222856
rect 543424 222844 543430 222896
rect 554038 222844 554044 222896
rect 554096 222884 554102 222896
rect 632698 222884 632704 222896
rect 554096 222856 632704 222884
rect 554096 222844 554102 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 78582 222708 78588 222760
rect 78640 222748 78646 222760
rect 98546 222748 98552 222760
rect 78640 222720 98552 222748
rect 78640 222708 78646 222720
rect 98546 222708 98552 222720
rect 98604 222708 98610 222760
rect 164970 222748 164976 222760
rect 98748 222720 164976 222748
rect 87966 222572 87972 222624
rect 88024 222612 88030 222624
rect 98748 222612 98776 222720
rect 164970 222708 164976 222720
rect 165028 222708 165034 222760
rect 165614 222708 165620 222760
rect 165672 222748 165678 222760
rect 192018 222748 192024 222760
rect 165672 222720 192024 222748
rect 165672 222708 165678 222720
rect 192018 222708 192024 222720
rect 192076 222708 192082 222760
rect 193950 222708 193956 222760
rect 194008 222748 194014 222760
rect 247402 222748 247408 222760
rect 194008 222720 247408 222748
rect 194008 222708 194014 222720
rect 247402 222708 247408 222720
rect 247460 222708 247466 222760
rect 284202 222708 284208 222760
rect 284260 222748 284266 222760
rect 316954 222748 316960 222760
rect 284260 222720 316960 222748
rect 284260 222708 284266 222720
rect 316954 222708 316960 222720
rect 317012 222708 317018 222760
rect 345658 222708 345664 222760
rect 345716 222748 345722 222760
rect 347866 222748 347872 222760
rect 345716 222720 347872 222748
rect 345716 222708 345722 222720
rect 347866 222708 347872 222720
rect 347924 222708 347930 222760
rect 532510 222708 532516 222760
rect 532568 222748 532574 222760
rect 533522 222748 533528 222760
rect 532568 222720 533528 222748
rect 532568 222708 532574 222720
rect 533522 222708 533528 222720
rect 533580 222708 533586 222760
rect 558178 222708 558184 222760
rect 558236 222748 558242 222760
rect 558236 222720 596174 222748
rect 558236 222708 558242 222720
rect 126514 222612 126520 222624
rect 88024 222584 98776 222612
rect 103486 222584 126520 222612
rect 88024 222572 88030 222584
rect 98546 222436 98552 222488
rect 98604 222476 98610 222488
rect 103486 222476 103514 222584
rect 126514 222572 126520 222584
rect 126572 222572 126578 222624
rect 191374 222612 191380 222624
rect 127084 222584 191380 222612
rect 98604 222448 103514 222476
rect 98604 222436 98610 222448
rect 118418 222436 118424 222488
rect 118476 222476 118482 222488
rect 127084 222476 127112 222584
rect 191374 222572 191380 222584
rect 191432 222572 191438 222624
rect 197170 222572 197176 222624
rect 197228 222612 197234 222624
rect 249978 222612 249984 222624
rect 197228 222584 249984 222612
rect 197228 222572 197234 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 482738 222572 482744 222624
rect 482796 222612 482802 222624
rect 593966 222612 593972 222624
rect 482796 222584 593972 222612
rect 482796 222572 482802 222584
rect 593966 222572 593972 222584
rect 594024 222572 594030 222624
rect 596146 222612 596174 222720
rect 670620 222680 670648 223740
rect 670786 223592 670792 223644
rect 670844 223632 670850 223644
rect 670844 223604 671186 223632
rect 670844 223592 670850 223604
rect 671022 223372 671074 223378
rect 671022 223314 671074 223320
rect 670786 223116 670792 223168
rect 670844 223156 670850 223168
rect 670844 223128 670956 223156
rect 670844 223116 670850 223128
rect 670620 222652 670832 222680
rect 630674 222612 630680 222624
rect 596146 222584 630680 222612
rect 630674 222572 630680 222584
rect 630732 222572 630738 222624
rect 146754 222476 146760 222488
rect 118476 222448 127112 222476
rect 132466 222448 146760 222476
rect 118476 222436 118482 222448
rect 126514 222300 126520 222352
rect 126572 222340 126578 222352
rect 132466 222340 132494 222448
rect 146754 222436 146760 222448
rect 146812 222436 146818 222488
rect 206830 222476 206836 222488
rect 146956 222448 206836 222476
rect 126572 222312 132494 222340
rect 126572 222300 126578 222312
rect 139118 222300 139124 222352
rect 139176 222340 139182 222352
rect 146956 222340 146984 222448
rect 206830 222436 206836 222448
rect 206888 222436 206894 222488
rect 207842 222436 207848 222488
rect 207900 222476 207906 222488
rect 258350 222476 258356 222488
rect 207900 222448 258356 222476
rect 207900 222436 207906 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 500218 222436 500224 222488
rect 500276 222476 500282 222488
rect 533338 222476 533344 222488
rect 500276 222448 533344 222476
rect 500276 222436 500282 222448
rect 533338 222436 533344 222448
rect 533396 222436 533402 222488
rect 533522 222436 533528 222488
rect 533580 222476 533586 222488
rect 621198 222476 621204 222488
rect 533580 222448 621204 222476
rect 533580 222436 533586 222448
rect 621198 222436 621204 222448
rect 621256 222436 621262 222488
rect 670804 222420 670832 222652
rect 490006 222368 490012 222420
rect 490064 222408 490070 222420
rect 490064 222380 495434 222408
rect 490064 222368 490070 222380
rect 139176 222312 146984 222340
rect 139176 222300 139182 222312
rect 147122 222300 147128 222352
rect 147180 222340 147186 222352
rect 211982 222340 211988 222352
rect 147180 222312 211988 222340
rect 147180 222300 147186 222312
rect 211982 222300 211988 222312
rect 212040 222300 212046 222352
rect 237006 222300 237012 222352
rect 237064 222340 237070 222352
rect 280890 222340 280896 222352
rect 237064 222312 280896 222340
rect 237064 222300 237070 222312
rect 280890 222300 280896 222312
rect 280948 222300 280954 222352
rect 484578 222300 484584 222352
rect 484636 222340 484642 222352
rect 495406 222340 495434 222380
rect 670786 222368 670792 222420
rect 670844 222368 670850 222420
rect 629846 222340 629852 222352
rect 484636 222312 489914 222340
rect 495406 222312 629852 222340
rect 484636 222300 484642 222312
rect 489886 222204 489914 222312
rect 629846 222300 629852 222312
rect 629904 222300 629910 222352
rect 500218 222204 500224 222216
rect 489886 222176 500224 222204
rect 500218 222164 500224 222176
rect 500276 222164 500282 222216
rect 533338 222164 533344 222216
rect 533396 222204 533402 222216
rect 558178 222204 558184 222216
rect 533396 222176 558184 222204
rect 533396 222164 533402 222176
rect 558178 222164 558184 222176
rect 558236 222164 558242 222216
rect 562870 222164 562876 222216
rect 562928 222204 562934 222216
rect 627086 222204 627092 222216
rect 562928 222176 627092 222204
rect 562928 222164 562934 222176
rect 627086 222164 627092 222176
rect 627144 222164 627150 222216
rect 111978 222096 111984 222148
rect 112036 222136 112042 222148
rect 185854 222136 185860 222148
rect 112036 222108 185860 222136
rect 112036 222096 112042 222108
rect 185854 222096 185860 222108
rect 185912 222096 185918 222148
rect 200390 222096 200396 222148
rect 200448 222136 200454 222148
rect 252922 222136 252928 222148
rect 200448 222108 252928 222136
rect 200448 222096 200454 222108
rect 252922 222096 252928 222108
rect 252980 222096 252986 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263870 222136 263876 222148
rect 258132 222108 263876 222136
rect 258132 222096 258138 222108
rect 263870 222096 263876 222108
rect 263928 222096 263934 222148
rect 270034 222096 270040 222148
rect 270092 222136 270098 222148
rect 306374 222136 306380 222148
rect 270092 222108 306380 222136
rect 270092 222096 270098 222108
rect 306374 222096 306380 222108
rect 306432 222096 306438 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353938 222136 353944 222148
rect 331456 222108 353944 222136
rect 331456 222096 331462 222108
rect 353938 222096 353944 222108
rect 353996 222096 354002 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 560938 222096 560944 222148
rect 560996 222136 561002 222148
rect 562502 222136 562508 222148
rect 560996 222108 562508 222136
rect 560996 222096 561002 222108
rect 562502 222096 562508 222108
rect 562560 222096 562566 222148
rect 533154 222028 533160 222080
rect 533212 222068 533218 222080
rect 538766 222068 538772 222080
rect 533212 222040 538772 222068
rect 533212 222028 533218 222040
rect 538766 222028 538772 222040
rect 538824 222028 538830 222080
rect 539502 222028 539508 222080
rect 539560 222068 539566 222080
rect 543182 222068 543188 222080
rect 539560 222040 543188 222068
rect 539560 222028 539566 222040
rect 543182 222028 543188 222040
rect 543240 222028 543246 222080
rect 543366 222028 543372 222080
rect 543424 222068 543430 222080
rect 546954 222068 546960 222080
rect 543424 222040 546960 222068
rect 543424 222028 543430 222040
rect 546954 222028 546960 222040
rect 547012 222028 547018 222080
rect 547138 222028 547144 222080
rect 547196 222068 547202 222080
rect 547690 222068 547696 222080
rect 547196 222040 547696 222068
rect 547196 222028 547202 222040
rect 547690 222028 547696 222040
rect 547748 222028 547754 222080
rect 547874 222028 547880 222080
rect 547932 222068 547938 222080
rect 598566 222068 598572 222080
rect 547932 222040 556384 222068
rect 547932 222028 547938 222040
rect 91278 221960 91284 222012
rect 91336 222000 91342 222012
rect 167178 222000 167184 222012
rect 91336 221972 167184 222000
rect 91336 221960 91342 221972
rect 167178 221960 167184 221972
rect 167236 221960 167242 222012
rect 167454 221960 167460 222012
rect 167512 222000 167518 222012
rect 220630 222000 220636 222012
rect 167512 221972 220636 222000
rect 167512 221960 167518 221972
rect 220630 221960 220636 221972
rect 220688 221960 220694 222012
rect 220814 221960 220820 222012
rect 220872 222000 220878 222012
rect 222194 222000 222200 222012
rect 220872 221972 222200 222000
rect 220872 221960 220878 221972
rect 222194 221960 222200 221972
rect 222252 221960 222258 222012
rect 232130 221960 232136 222012
rect 232188 222000 232194 222012
rect 234706 222000 234712 222012
rect 232188 221972 234712 222000
rect 232188 221960 232194 221972
rect 234706 221960 234712 221972
rect 234764 221960 234770 222012
rect 261018 221960 261024 222012
rect 261076 222000 261082 222012
rect 301682 222000 301688 222012
rect 261076 221972 301688 222000
rect 261076 221960 261082 221972
rect 301682 221960 301688 221972
rect 301740 221960 301746 222012
rect 313182 221960 313188 222012
rect 313240 222000 313246 222012
rect 340414 222000 340420 222012
rect 313240 221972 340420 222000
rect 313240 221960 313246 221972
rect 340414 221960 340420 221972
rect 340472 221960 340478 222012
rect 516778 221960 516784 222012
rect 516836 222000 516842 222012
rect 527542 222000 527548 222012
rect 516836 221972 527548 222000
rect 516836 221960 516842 221972
rect 527542 221960 527548 221972
rect 527600 221960 527606 222012
rect 556356 222000 556384 222040
rect 563026 222040 598572 222068
rect 563026 222000 563054 222040
rect 598566 222028 598572 222040
rect 598624 222028 598630 222080
rect 556356 221972 563054 222000
rect 598750 221960 598756 222012
rect 598808 222000 598814 222012
rect 603074 222000 603080 222012
rect 598808 221972 603080 222000
rect 598808 221960 598814 221972
rect 603074 221960 603080 221972
rect 603132 221960 603138 222012
rect 533982 221892 533988 221944
rect 534040 221932 534046 221944
rect 534040 221904 553716 221932
rect 534040 221892 534046 221904
rect 94590 221824 94596 221876
rect 94648 221864 94654 221876
rect 169846 221864 169852 221876
rect 94648 221836 169852 221864
rect 94648 221824 94654 221836
rect 169846 221824 169852 221836
rect 169904 221824 169910 221876
rect 172698 221864 172704 221876
rect 170048 221836 172704 221864
rect 97718 221688 97724 221740
rect 97776 221728 97782 221740
rect 170048 221728 170076 221836
rect 172698 221824 172704 221836
rect 172756 221824 172762 221876
rect 174078 221824 174084 221876
rect 174136 221864 174142 221876
rect 231946 221864 231952 221876
rect 174136 221836 231952 221864
rect 174136 221824 174142 221836
rect 231946 221824 231952 221836
rect 232004 221824 232010 221876
rect 233694 221824 233700 221876
rect 233752 221864 233758 221876
rect 277946 221864 277952 221876
rect 233752 221836 277952 221864
rect 233752 221824 233758 221836
rect 277946 221824 277952 221836
rect 278004 221824 278010 221876
rect 280062 221824 280068 221876
rect 280120 221864 280126 221876
rect 313734 221864 313740 221876
rect 280120 221836 313740 221864
rect 280120 221824 280126 221836
rect 313734 221824 313740 221836
rect 313792 221824 313798 221876
rect 318242 221824 318248 221876
rect 318300 221864 318306 221876
rect 343818 221864 343824 221876
rect 318300 221836 343824 221864
rect 318300 221824 318306 221836
rect 343818 221824 343824 221836
rect 343876 221824 343882 221876
rect 353294 221824 353300 221876
rect 353352 221864 353358 221876
rect 372706 221864 372712 221876
rect 353352 221836 372712 221864
rect 353352 221824 353358 221836
rect 372706 221824 372712 221836
rect 372764 221824 372770 221876
rect 380342 221864 380348 221876
rect 373966 221836 380348 221864
rect 97776 221700 170076 221728
rect 97776 221688 97782 221700
rect 171594 221688 171600 221740
rect 171652 221728 171658 221740
rect 171652 221700 172008 221728
rect 171652 221688 171658 221700
rect 73890 221552 73896 221604
rect 73948 221592 73954 221604
rect 82078 221592 82084 221604
rect 73948 221564 82084 221592
rect 73948 221552 73954 221564
rect 82078 221552 82084 221564
rect 82136 221552 82142 221604
rect 86310 221552 86316 221604
rect 86368 221592 86374 221604
rect 164326 221592 164332 221604
rect 86368 221564 164332 221592
rect 86368 221552 86374 221564
rect 164326 221552 164332 221564
rect 164384 221552 164390 221604
rect 164510 221552 164516 221604
rect 164568 221592 164574 221604
rect 171778 221592 171784 221604
rect 164568 221564 171784 221592
rect 164568 221552 164574 221564
rect 171778 221552 171784 221564
rect 171836 221552 171842 221604
rect 171980 221592 172008 221700
rect 174906 221688 174912 221740
rect 174964 221728 174970 221740
rect 174964 221700 185348 221728
rect 174964 221688 174970 221700
rect 185320 221660 185348 221700
rect 185762 221688 185768 221740
rect 185820 221728 185826 221740
rect 243078 221728 243084 221740
rect 185820 221700 243084 221728
rect 185820 221688 185826 221700
rect 243078 221688 243084 221700
rect 243136 221688 243142 221740
rect 263134 221728 263140 221740
rect 243556 221700 263140 221728
rect 185320 221632 185440 221660
rect 182634 221592 182640 221604
rect 171980 221564 182640 221592
rect 182634 221552 182640 221564
rect 182692 221552 182698 221604
rect 185412 221592 185440 221632
rect 232130 221592 232136 221604
rect 185412 221564 232136 221592
rect 232130 221552 232136 221564
rect 232188 221552 232194 221604
rect 243556 221592 243584 221700
rect 263134 221688 263140 221700
rect 263192 221688 263198 221740
rect 263502 221688 263508 221740
rect 263560 221728 263566 221740
rect 301038 221728 301044 221740
rect 263560 221700 301044 221728
rect 263560 221688 263566 221700
rect 301038 221688 301044 221700
rect 301096 221688 301102 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332778 221728 332784 221740
rect 303304 221700 332784 221728
rect 303304 221688 303310 221700
rect 332778 221688 332784 221700
rect 332836 221688 332842 221740
rect 344646 221688 344652 221740
rect 344704 221728 344710 221740
rect 364518 221728 364524 221740
rect 344704 221700 364524 221728
rect 344704 221688 344710 221700
rect 364518 221688 364524 221700
rect 364576 221688 364582 221740
rect 370958 221688 370964 221740
rect 371016 221728 371022 221740
rect 373966 221728 373994 221836
rect 380342 221824 380348 221836
rect 380400 221824 380406 221876
rect 492490 221824 492496 221876
rect 492548 221864 492554 221876
rect 506842 221864 506848 221876
rect 492548 221836 506848 221864
rect 492548 221824 492554 221836
rect 506842 221824 506848 221836
rect 506900 221824 506906 221876
rect 523494 221824 523500 221876
rect 523552 221864 523558 221876
rect 533706 221864 533712 221876
rect 523552 221836 533712 221864
rect 523552 221824 523558 221836
rect 533706 221824 533712 221836
rect 533764 221824 533770 221876
rect 424962 221756 424968 221808
rect 425020 221796 425026 221808
rect 429194 221796 429200 221808
rect 425020 221768 429200 221796
rect 425020 221756 425026 221768
rect 429194 221756 429200 221768
rect 429252 221756 429258 221808
rect 547874 221756 547880 221808
rect 547932 221796 547938 221808
rect 553486 221796 553492 221808
rect 547932 221768 553492 221796
rect 547932 221756 547938 221768
rect 553486 221756 553492 221768
rect 553544 221756 553550 221808
rect 371016 221700 373994 221728
rect 371016 221688 371022 221700
rect 380066 221688 380072 221740
rect 380124 221728 380130 221740
rect 386506 221728 386512 221740
rect 380124 221700 386512 221728
rect 380124 221688 380130 221700
rect 386506 221688 386512 221700
rect 386564 221688 386570 221740
rect 475838 221688 475844 221740
rect 475896 221728 475902 221740
rect 486142 221728 486148 221740
rect 475896 221700 486148 221728
rect 475896 221688 475902 221700
rect 486142 221688 486148 221700
rect 486200 221688 486206 221740
rect 496262 221688 496268 221740
rect 496320 221728 496326 221740
rect 513558 221728 513564 221740
rect 496320 221700 513564 221728
rect 496320 221688 496326 221700
rect 513558 221688 513564 221700
rect 513616 221688 513622 221740
rect 524230 221688 524236 221740
rect 524288 221728 524294 221740
rect 547690 221728 547696 221740
rect 524288 221700 547696 221728
rect 524288 221688 524294 221700
rect 547690 221688 547696 221700
rect 547748 221688 547754 221740
rect 553688 221728 553716 221904
rect 553854 221824 553860 221876
rect 553912 221864 553918 221876
rect 598934 221864 598940 221876
rect 553912 221836 598940 221864
rect 553912 221824 553918 221836
rect 598934 221824 598940 221836
rect 598992 221824 598998 221876
rect 599118 221824 599124 221876
rect 599176 221864 599182 221876
rect 606110 221864 606116 221876
rect 599176 221836 606116 221864
rect 599176 221824 599182 221836
rect 606110 221824 606116 221836
rect 606168 221824 606174 221876
rect 559374 221728 559380 221740
rect 553688 221700 559380 221728
rect 559374 221688 559380 221700
rect 559432 221688 559438 221740
rect 559558 221688 559564 221740
rect 559616 221728 559622 221740
rect 562686 221728 562692 221740
rect 559616 221700 562692 221728
rect 559616 221688 559622 221700
rect 562686 221688 562692 221700
rect 562744 221688 562750 221740
rect 562870 221688 562876 221740
rect 562928 221728 562934 221740
rect 567010 221728 567016 221740
rect 562928 221700 567016 221728
rect 562928 221688 562934 221700
rect 567010 221688 567016 221700
rect 567068 221688 567074 221740
rect 567194 221688 567200 221740
rect 567252 221728 567258 221740
rect 609422 221728 609428 221740
rect 567252 221700 609428 221728
rect 567252 221688 567258 221700
rect 609422 221688 609428 221700
rect 609480 221688 609486 221740
rect 233896 221564 243584 221592
rect 59354 221416 59360 221468
rect 59412 221456 59418 221468
rect 141326 221456 141332 221468
rect 59412 221428 141332 221456
rect 59412 221416 59418 221428
rect 141326 221416 141332 221428
rect 141384 221416 141390 221468
rect 147582 221416 147588 221468
rect 147640 221456 147646 221468
rect 204898 221456 204904 221468
rect 147640 221428 204904 221456
rect 147640 221416 147646 221428
rect 204898 221416 204904 221428
rect 204956 221416 204962 221468
rect 205082 221416 205088 221468
rect 205140 221456 205146 221468
rect 220814 221456 220820 221468
rect 205140 221428 220820 221456
rect 205140 221416 205146 221428
rect 220814 221416 220820 221428
rect 220872 221416 220878 221468
rect 220998 221416 221004 221468
rect 221056 221456 221062 221468
rect 233896 221456 233924 221564
rect 243722 221552 243728 221604
rect 243780 221592 243786 221604
rect 283742 221592 283748 221604
rect 243780 221564 283748 221592
rect 243780 221552 243786 221564
rect 283742 221552 283748 221564
rect 283800 221552 283806 221604
rect 302418 221552 302424 221604
rect 302476 221592 302482 221604
rect 334066 221592 334072 221604
rect 302476 221564 334072 221592
rect 302476 221552 302482 221564
rect 334066 221552 334072 221564
rect 334124 221552 334130 221604
rect 348786 221552 348792 221604
rect 348844 221592 348850 221604
rect 370038 221592 370044 221604
rect 348844 221564 370044 221592
rect 348844 221552 348850 221564
rect 370038 221552 370044 221564
rect 370096 221552 370102 221604
rect 373718 221552 373724 221604
rect 373776 221592 373782 221604
rect 384298 221592 384304 221604
rect 373776 221564 384304 221592
rect 373776 221552 373782 221564
rect 384298 221552 384304 221564
rect 384356 221552 384362 221604
rect 391014 221552 391020 221604
rect 391072 221592 391078 221604
rect 400398 221592 400404 221604
rect 391072 221564 400404 221592
rect 391072 221552 391078 221564
rect 400398 221552 400404 221564
rect 400456 221552 400462 221604
rect 401318 221552 401324 221604
rect 401376 221592 401382 221604
rect 405826 221592 405832 221604
rect 401376 221564 405832 221592
rect 401376 221552 401382 221564
rect 405826 221552 405832 221564
rect 405884 221552 405890 221604
rect 484762 221552 484768 221604
rect 484820 221592 484826 221604
rect 498102 221592 498108 221604
rect 484820 221564 498108 221592
rect 484820 221552 484826 221564
rect 498102 221552 498108 221564
rect 498160 221552 498166 221604
rect 501322 221552 501328 221604
rect 501380 221592 501386 221604
rect 520182 221592 520188 221604
rect 501380 221564 520188 221592
rect 501380 221552 501386 221564
rect 520182 221552 520188 221564
rect 520240 221552 520246 221604
rect 522666 221552 522672 221604
rect 522724 221592 522730 221604
rect 522724 221564 533384 221592
rect 522724 221552 522730 221564
rect 221056 221428 233924 221456
rect 221056 221416 221062 221428
rect 234062 221416 234068 221468
rect 234120 221456 234126 221468
rect 276106 221456 276112 221468
rect 234120 221428 276112 221456
rect 234120 221416 234126 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 284018 221416 284024 221468
rect 284076 221456 284082 221468
rect 320358 221456 320364 221468
rect 284076 221428 320364 221456
rect 284076 221416 284082 221428
rect 320358 221416 320364 221428
rect 320416 221416 320422 221468
rect 333422 221416 333428 221468
rect 333480 221456 333486 221468
rect 357526 221456 357532 221468
rect 333480 221428 357532 221456
rect 333480 221416 333486 221428
rect 357526 221416 357532 221428
rect 357584 221416 357590 221468
rect 369486 221416 369492 221468
rect 369544 221456 369550 221468
rect 384114 221456 384120 221468
rect 369544 221428 384120 221456
rect 369544 221416 369550 221428
rect 384114 221416 384120 221428
rect 384172 221416 384178 221468
rect 384390 221416 384396 221468
rect 384448 221456 384454 221468
rect 395154 221456 395160 221468
rect 384448 221428 395160 221456
rect 384448 221416 384454 221428
rect 395154 221416 395160 221428
rect 395212 221416 395218 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 533154 221456 533160 221468
rect 483808 221428 533160 221456
rect 483808 221416 483814 221428
rect 533154 221416 533160 221428
rect 533212 221416 533218 221468
rect 533356 221456 533384 221564
rect 533522 221552 533528 221604
rect 533580 221592 533586 221604
rect 598750 221592 598756 221604
rect 533580 221564 598756 221592
rect 533580 221552 533586 221564
rect 598750 221552 598756 221564
rect 598808 221552 598814 221604
rect 598934 221552 598940 221604
rect 598992 221592 598998 221604
rect 605926 221592 605932 221604
rect 598992 221564 605932 221592
rect 598992 221552 598998 221564
rect 605926 221552 605932 221564
rect 605984 221552 605990 221604
rect 546586 221456 546592 221468
rect 533356 221428 546592 221456
rect 546586 221416 546592 221428
rect 546644 221416 546650 221468
rect 546770 221416 546776 221468
rect 546828 221456 546834 221468
rect 599118 221456 599124 221468
rect 546828 221428 599124 221456
rect 546828 221416 546834 221428
rect 599118 221416 599124 221428
rect 599176 221416 599182 221468
rect 599302 221348 599308 221400
rect 599360 221388 599366 221400
rect 605006 221388 605012 221400
rect 599360 221360 605012 221388
rect 599360 221348 599366 221360
rect 605006 221348 605012 221360
rect 605064 221348 605070 221400
rect 104526 221280 104532 221332
rect 104584 221320 104590 221332
rect 176470 221320 176476 221332
rect 104584 221292 176476 221320
rect 104584 221280 104590 221292
rect 176470 221280 176476 221292
rect 176528 221280 176534 221332
rect 176626 221292 185532 221320
rect 111150 221144 111156 221196
rect 111208 221184 111214 221196
rect 171594 221184 171600 221196
rect 111208 221156 171600 221184
rect 111208 221144 111214 221156
rect 171594 221144 171600 221156
rect 171652 221144 171658 221196
rect 171778 221144 171784 221196
rect 171836 221184 171842 221196
rect 176626 221184 176654 221292
rect 185504 221252 185532 221292
rect 185854 221280 185860 221332
rect 185912 221320 185918 221332
rect 234246 221320 234252 221332
rect 185912 221292 234252 221320
rect 185912 221280 185918 221292
rect 234246 221280 234252 221292
rect 234304 221280 234310 221332
rect 237834 221280 237840 221332
rect 237892 221320 237898 221332
rect 243722 221320 243728 221332
rect 237892 221292 243728 221320
rect 237892 221280 237898 221292
rect 243722 221280 243728 221292
rect 243780 221280 243786 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 527174 221280 527180 221332
rect 527232 221320 527238 221332
rect 528186 221320 528192 221332
rect 527232 221292 528192 221320
rect 527232 221280 527238 221292
rect 528186 221280 528192 221292
rect 528244 221320 528250 221332
rect 533522 221320 533528 221332
rect 528244 221292 533528 221320
rect 528244 221280 528250 221292
rect 533522 221280 533528 221292
rect 533580 221280 533586 221332
rect 185504 221224 185716 221252
rect 171836 221156 176654 221184
rect 171836 221144 171842 221156
rect 177298 221144 177304 221196
rect 177356 221184 177362 221196
rect 185302 221184 185308 221196
rect 177356 221156 185308 221184
rect 177356 221144 177362 221156
rect 185302 221144 185308 221156
rect 185360 221144 185366 221196
rect 185688 221184 185716 221224
rect 533706 221212 533712 221264
rect 533764 221252 533770 221264
rect 601694 221252 601700 221264
rect 533764 221224 601700 221252
rect 533764 221212 533770 221224
rect 601694 221212 601700 221224
rect 601752 221212 601758 221264
rect 185688 221156 200114 221184
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 193306 221048 193312 221060
rect 124456 221020 193312 221048
rect 124456 221008 124462 221020
rect 193306 221008 193312 221020
rect 193364 221008 193370 221060
rect 200086 221048 200114 221156
rect 204898 221144 204904 221196
rect 204956 221184 204962 221196
rect 211154 221184 211160 221196
rect 204956 221156 211160 221184
rect 204956 221144 204962 221156
rect 211154 221144 211160 221156
rect 211212 221144 211218 221196
rect 211522 221144 211528 221196
rect 211580 221184 211586 221196
rect 260834 221184 260840 221196
rect 211580 221156 260840 221184
rect 211580 221144 211586 221156
rect 260834 221144 260840 221156
rect 260892 221144 260898 221196
rect 521010 221076 521016 221128
rect 521068 221116 521074 221128
rect 601142 221116 601148 221128
rect 521068 221088 601148 221116
rect 521068 221076 521074 221088
rect 601142 221076 601148 221088
rect 601200 221076 601206 221128
rect 205082 221048 205088 221060
rect 200086 221020 205088 221048
rect 205082 221008 205088 221020
rect 205140 221008 205146 221060
rect 218054 221008 218060 221060
rect 218112 221048 218118 221060
rect 220998 221048 221004 221060
rect 218112 221020 221004 221048
rect 218112 221008 218118 221020
rect 220998 221008 221004 221020
rect 221056 221008 221062 221060
rect 226518 221048 226524 221060
rect 221200 221020 226524 221048
rect 82998 220940 83004 220992
rect 83056 220980 83062 220992
rect 83056 220952 93854 220980
rect 83056 220940 83062 220952
rect 93826 220912 93854 220952
rect 151078 220912 151084 220924
rect 93826 220884 151084 220912
rect 151078 220872 151084 220884
rect 151136 220872 151142 220924
rect 155034 220872 155040 220924
rect 155092 220912 155098 220924
rect 219618 220912 219624 220924
rect 155092 220884 219624 220912
rect 155092 220872 155098 220884
rect 219618 220872 219624 220884
rect 219676 220872 219682 220924
rect 220630 220872 220636 220924
rect 220688 220912 220694 220924
rect 221200 220912 221228 221020
rect 226518 221008 226524 221020
rect 226576 221008 226582 221060
rect 227898 221008 227904 221060
rect 227956 221048 227962 221060
rect 234062 221048 234068 221060
rect 227956 221020 234068 221048
rect 227956 221008 227962 221020
rect 234062 221008 234068 221020
rect 234120 221008 234126 221060
rect 268194 221048 268200 221060
rect 238726 221020 268200 221048
rect 220688 220884 221228 220912
rect 220688 220872 220694 220884
rect 223482 220872 223488 220924
rect 223540 220912 223546 220924
rect 238726 220912 238754 221020
rect 268194 221008 268200 221020
rect 268252 221008 268258 221060
rect 517514 220940 517520 220992
rect 517572 220980 517578 220992
rect 518434 220980 518440 220992
rect 517572 220952 518440 220980
rect 517572 220940 517578 220952
rect 518434 220940 518440 220952
rect 518492 220980 518498 220992
rect 600314 220980 600320 220992
rect 518492 220952 600320 220980
rect 518492 220940 518498 220952
rect 600314 220940 600320 220952
rect 600372 220940 600378 220992
rect 223540 220884 238754 220912
rect 223540 220872 223546 220884
rect 253842 220872 253848 220924
rect 253900 220912 253906 220924
rect 258626 220912 258632 220924
rect 253900 220884 258632 220912
rect 253900 220872 253906 220884
rect 258626 220872 258632 220884
rect 258684 220872 258690 220924
rect 80514 220804 80520 220856
rect 80572 220844 80578 220856
rect 86126 220844 86132 220856
rect 80572 220816 86132 220844
rect 80572 220804 80578 220816
rect 86126 220804 86132 220816
rect 86184 220804 86190 220856
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 456702 220804 456708 220856
rect 456760 220844 456766 220856
rect 462130 220844 462136 220856
rect 456760 220816 462136 220844
rect 456760 220804 456766 220816
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471422 220844 471428 220856
rect 466144 220816 471428 220844
rect 466144 220804 466150 220816
rect 471422 220804 471428 220816
rect 471480 220804 471486 220856
rect 515766 220804 515772 220856
rect 515824 220844 515830 220856
rect 600498 220844 600504 220856
rect 515824 220816 600504 220844
rect 515824 220804 515830 220816
rect 600498 220804 600504 220816
rect 600556 220804 600562 220856
rect 101214 220736 101220 220788
rect 101272 220776 101278 220788
rect 166948 220776 166954 220788
rect 101272 220748 166954 220776
rect 101272 220736 101278 220748
rect 166948 220736 166954 220748
rect 167006 220736 167012 220788
rect 167178 220736 167184 220788
rect 167236 220776 167242 220788
rect 176470 220776 176476 220788
rect 167236 220748 176476 220776
rect 167236 220736 167242 220748
rect 176470 220736 176476 220748
rect 176528 220736 176534 220788
rect 176608 220736 176614 220788
rect 176666 220776 176672 220788
rect 180518 220776 180524 220788
rect 176666 220748 180524 220776
rect 176666 220736 176672 220748
rect 180518 220736 180524 220748
rect 180576 220736 180582 220788
rect 180702 220736 180708 220788
rect 180760 220776 180766 220788
rect 236730 220776 236736 220788
rect 180760 220748 236736 220776
rect 180760 220736 180766 220748
rect 236730 220736 236736 220748
rect 236788 220736 236794 220788
rect 254394 220736 254400 220788
rect 254452 220776 254458 220788
rect 296806 220776 296812 220788
rect 254452 220748 296812 220776
rect 254452 220736 254458 220748
rect 296806 220736 296812 220748
rect 296864 220736 296870 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 455322 220668 455328 220720
rect 455380 220708 455386 220720
rect 458818 220708 458824 220720
rect 455380 220680 458824 220708
rect 455380 220668 455386 220680
rect 458818 220668 458824 220680
rect 458876 220668 458882 220720
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 511810 220668 511816 220720
rect 511868 220708 511874 220720
rect 511868 220680 518894 220708
rect 511868 220668 511874 220680
rect 76374 220600 76380 220652
rect 76432 220640 76438 220652
rect 149238 220640 149244 220652
rect 76432 220612 149244 220640
rect 76432 220600 76438 220612
rect 149238 220600 149244 220612
rect 149296 220600 149302 220652
rect 149422 220600 149428 220652
rect 149480 220640 149486 220652
rect 166350 220640 166356 220652
rect 149480 220612 166356 220640
rect 149480 220600 149486 220612
rect 166350 220600 166356 220612
rect 166408 220600 166414 220652
rect 166534 220600 166540 220652
rect 166592 220640 166598 220652
rect 221274 220640 221280 220652
rect 166592 220612 221280 220640
rect 166592 220600 166598 220612
rect 221274 220600 221280 220612
rect 221332 220600 221338 220652
rect 223758 220640 223764 220652
rect 221568 220612 223764 220640
rect 79686 220464 79692 220516
rect 79744 220504 79750 220516
rect 158898 220504 158904 220516
rect 79744 220476 158904 220504
rect 79744 220464 79750 220476
rect 158898 220464 158904 220476
rect 158956 220464 158962 220516
rect 164142 220464 164148 220516
rect 164200 220504 164206 220516
rect 166902 220504 166908 220516
rect 164200 220476 166908 220504
rect 164200 220464 164206 220476
rect 166902 220464 166908 220476
rect 166960 220464 166966 220516
rect 167086 220464 167092 220516
rect 167144 220504 167150 220516
rect 221568 220504 221596 220612
rect 223758 220600 223764 220612
rect 223816 220600 223822 220652
rect 236178 220600 236184 220652
rect 236236 220640 236242 220652
rect 246482 220640 246488 220652
rect 236236 220612 246488 220640
rect 236236 220600 236242 220612
rect 246482 220600 246488 220612
rect 246540 220600 246546 220652
rect 246942 220600 246948 220652
rect 247000 220640 247006 220652
rect 288618 220640 288624 220652
rect 247000 220612 288624 220640
rect 247000 220600 247006 220612
rect 288618 220600 288624 220612
rect 288676 220600 288682 220652
rect 304902 220600 304908 220652
rect 304960 220640 304966 220652
rect 333238 220640 333244 220652
rect 304960 220612 333244 220640
rect 304960 220600 304966 220612
rect 333238 220600 333244 220612
rect 333296 220600 333302 220652
rect 500402 220600 500408 220652
rect 500460 220640 500466 220652
rect 500460 220612 505094 220640
rect 500460 220600 500466 220612
rect 505066 220572 505094 220612
rect 511810 220572 511816 220584
rect 505066 220544 511816 220572
rect 511810 220532 511816 220544
rect 511868 220532 511874 220584
rect 167144 220476 221596 220504
rect 167144 220464 167150 220476
rect 223758 220464 223764 220516
rect 223816 220504 223822 220516
rect 270586 220504 270592 220516
rect 223816 220476 270592 220504
rect 223816 220464 223822 220476
rect 270586 220464 270592 220476
rect 270644 220464 270650 220516
rect 276750 220464 276756 220516
rect 276808 220504 276814 220516
rect 311342 220504 311348 220516
rect 276808 220476 311348 220504
rect 276808 220464 276814 220476
rect 311342 220464 311348 220476
rect 311400 220464 311406 220516
rect 328086 220464 328092 220516
rect 328144 220504 328150 220516
rect 351270 220504 351276 220516
rect 328144 220476 351276 220504
rect 328144 220464 328150 220476
rect 351270 220464 351276 220476
rect 351328 220464 351334 220516
rect 364518 220464 364524 220516
rect 364576 220504 364582 220516
rect 379698 220504 379704 220516
rect 364576 220476 379704 220504
rect 364576 220464 364582 220476
rect 379698 220464 379704 220476
rect 379756 220464 379762 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 518866 220504 518894 220680
rect 567010 220668 567016 220720
rect 567068 220708 567074 220720
rect 567194 220708 567200 220720
rect 567068 220680 567200 220708
rect 567068 220668 567074 220680
rect 567194 220668 567200 220680
rect 567252 220668 567258 220720
rect 529014 220600 529020 220652
rect 529072 220640 529078 220652
rect 544930 220640 544936 220652
rect 529072 220612 544936 220640
rect 529072 220600 529078 220612
rect 544930 220600 544936 220612
rect 544988 220600 544994 220652
rect 550818 220600 550824 220652
rect 550876 220640 550882 220652
rect 550876 220612 563054 220640
rect 550876 220600 550882 220612
rect 531682 220504 531688 220516
rect 518866 220476 531688 220504
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 548334 220464 548340 220516
rect 548392 220504 548398 220516
rect 551186 220504 551192 220516
rect 548392 220476 551192 220504
rect 548392 220464 548398 220476
rect 551186 220464 551192 220476
rect 551244 220464 551250 220516
rect 560754 220464 560760 220516
rect 560812 220504 560818 220516
rect 562870 220504 562876 220516
rect 560812 220476 562876 220504
rect 560812 220464 560818 220476
rect 562870 220464 562876 220476
rect 562928 220464 562934 220516
rect 563026 220504 563054 220612
rect 563238 220600 563244 220652
rect 563296 220640 563302 220652
rect 566826 220640 566832 220652
rect 563296 220612 566832 220640
rect 563296 220600 563302 220612
rect 566826 220600 566832 220612
rect 566884 220600 566890 220652
rect 567378 220600 567384 220652
rect 567436 220640 567442 220652
rect 611446 220640 611452 220652
rect 567436 220612 611452 220640
rect 567436 220600 567442 220612
rect 611446 220600 611452 220612
rect 611504 220600 611510 220652
rect 607306 220504 607312 220516
rect 563026 220476 607312 220504
rect 607306 220464 607312 220476
rect 607364 220464 607370 220516
rect 64598 220328 64604 220380
rect 64656 220368 64662 220380
rect 141970 220368 141976 220380
rect 64656 220340 141976 220368
rect 64656 220328 64662 220340
rect 141970 220328 141976 220340
rect 142028 220328 142034 220380
rect 144638 220368 144644 220380
rect 142126 220340 144644 220368
rect 69750 220192 69756 220244
rect 69808 220232 69814 220244
rect 142126 220232 142154 220340
rect 144638 220328 144644 220340
rect 144696 220328 144702 220380
rect 144822 220328 144828 220380
rect 144880 220368 144886 220380
rect 202414 220368 202420 220380
rect 144880 220340 202420 220368
rect 144880 220328 144886 220340
rect 202414 220328 202420 220340
rect 202472 220328 202478 220380
rect 202782 220328 202788 220380
rect 202840 220368 202846 220380
rect 214558 220368 214564 220380
rect 202840 220340 214564 220368
rect 202840 220328 202846 220340
rect 214558 220328 214564 220340
rect 214616 220328 214622 220380
rect 262398 220368 262404 220380
rect 214760 220340 262404 220368
rect 69808 220204 142154 220232
rect 69808 220192 69814 220204
rect 142246 220192 142252 220244
rect 142304 220232 142310 220244
rect 149422 220232 149428 220244
rect 142304 220204 149428 220232
rect 142304 220192 142310 220204
rect 149422 220192 149428 220204
rect 149480 220192 149486 220244
rect 150894 220192 150900 220244
rect 150952 220232 150958 220244
rect 150952 220204 211936 220232
rect 150952 220192 150958 220204
rect 73062 220056 73068 220108
rect 73120 220096 73126 220108
rect 153562 220096 153568 220108
rect 73120 220068 153568 220096
rect 73120 220056 73126 220068
rect 153562 220056 153568 220068
rect 153620 220056 153626 220108
rect 154206 220056 154212 220108
rect 154264 220096 154270 220108
rect 211706 220096 211712 220108
rect 154264 220068 211712 220096
rect 154264 220056 154270 220068
rect 211706 220056 211712 220068
rect 211764 220056 211770 220108
rect 211908 220096 211936 220204
rect 213822 220192 213828 220244
rect 213880 220232 213886 220244
rect 214760 220232 214788 220340
rect 262398 220328 262404 220340
rect 262456 220328 262462 220380
rect 262674 220328 262680 220380
rect 262732 220368 262738 220380
rect 264238 220368 264244 220380
rect 262732 220340 264244 220368
rect 262732 220328 262738 220340
rect 264238 220328 264244 220340
rect 264296 220328 264302 220380
rect 264606 220328 264612 220380
rect 264664 220368 264670 220380
rect 269298 220368 269304 220380
rect 264664 220340 269304 220368
rect 264664 220328 264670 220340
rect 269298 220328 269304 220340
rect 269356 220328 269362 220380
rect 273438 220328 273444 220380
rect 273496 220368 273502 220380
rect 309226 220368 309232 220380
rect 273496 220340 309232 220368
rect 273496 220328 273502 220340
rect 309226 220328 309232 220340
rect 309284 220328 309290 220380
rect 316494 220328 316500 220380
rect 316552 220368 316558 220380
rect 316552 220340 339908 220368
rect 316552 220328 316558 220340
rect 213880 220204 214788 220232
rect 213880 220192 213886 220204
rect 217134 220192 217140 220244
rect 217192 220232 217198 220244
rect 265158 220232 265164 220244
rect 217192 220204 265164 220232
rect 217192 220192 217198 220204
rect 265158 220192 265164 220204
rect 265216 220192 265222 220244
rect 267642 220192 267648 220244
rect 267700 220232 267706 220244
rect 306834 220232 306840 220244
rect 267700 220204 306840 220232
rect 267700 220192 267706 220204
rect 306834 220192 306840 220204
rect 306892 220192 306898 220244
rect 308950 220192 308956 220244
rect 309008 220232 309014 220244
rect 339678 220232 339684 220244
rect 309008 220204 339684 220232
rect 309008 220192 309014 220204
rect 339678 220192 339684 220204
rect 339736 220192 339742 220244
rect 339880 220232 339908 220340
rect 340322 220328 340328 220380
rect 340380 220368 340386 220380
rect 342438 220368 342444 220380
rect 340380 220340 342444 220368
rect 340380 220328 340386 220340
rect 342438 220328 342444 220340
rect 342496 220328 342502 220380
rect 342990 220368 342996 220380
rect 342640 220340 342996 220368
rect 342640 220232 342668 220340
rect 342990 220328 342996 220340
rect 343048 220328 343054 220380
rect 351270 220328 351276 220380
rect 351328 220368 351334 220380
rect 369302 220368 369308 220380
rect 351328 220340 369308 220368
rect 351328 220328 351334 220340
rect 369302 220328 369308 220340
rect 369360 220328 369366 220380
rect 376938 220328 376944 220380
rect 376996 220368 377002 220380
rect 388438 220368 388444 220380
rect 376996 220340 388444 220368
rect 376996 220328 377002 220340
rect 388438 220328 388444 220340
rect 388496 220328 388502 220380
rect 436278 220328 436284 220380
rect 436336 220368 436342 220380
rect 437014 220368 437020 220380
rect 436336 220340 437020 220368
rect 436336 220328 436342 220340
rect 437014 220328 437020 220340
rect 437072 220328 437078 220380
rect 472986 220328 472992 220380
rect 473044 220368 473050 220380
rect 481174 220368 481180 220380
rect 473044 220340 481180 220368
rect 473044 220328 473050 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 509878 220328 509884 220380
rect 509936 220368 509942 220380
rect 522574 220368 522580 220380
rect 509936 220340 522580 220368
rect 509936 220328 509942 220340
rect 522574 220328 522580 220340
rect 522632 220328 522638 220380
rect 528370 220328 528376 220380
rect 528428 220368 528434 220380
rect 553946 220368 553952 220380
rect 528428 220340 553952 220368
rect 528428 220328 528434 220340
rect 553946 220328 553952 220340
rect 554004 220328 554010 220380
rect 558178 220328 558184 220380
rect 558236 220368 558242 220380
rect 566458 220368 566464 220380
rect 558236 220340 566464 220368
rect 558236 220328 558242 220340
rect 566458 220328 566464 220340
rect 566516 220328 566522 220380
rect 567838 220328 567844 220380
rect 567896 220368 567902 220380
rect 610526 220368 610532 220380
rect 567896 220340 610532 220368
rect 567896 220328 567902 220340
rect 610526 220328 610532 220340
rect 610584 220328 610590 220380
rect 566642 220260 566648 220312
rect 566700 220300 566706 220312
rect 567148 220300 567154 220312
rect 566700 220272 567154 220300
rect 566700 220260 566706 220272
rect 567148 220260 567154 220272
rect 567206 220260 567212 220312
rect 339880 220204 342668 220232
rect 342990 220192 342996 220244
rect 343048 220232 343054 220244
rect 363322 220232 363328 220244
rect 343048 220204 363328 220232
rect 343048 220192 343054 220204
rect 363322 220192 363328 220204
rect 363380 220192 363386 220244
rect 363690 220192 363696 220244
rect 363748 220232 363754 220244
rect 381078 220232 381084 220244
rect 363748 220204 381084 220232
rect 363748 220192 363754 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388438 220192 388444 220244
rect 388496 220232 388502 220244
rect 400950 220232 400956 220244
rect 388496 220204 400956 220232
rect 388496 220192 388502 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 429562 220192 429568 220244
rect 429620 220232 429626 220244
rect 432046 220232 432052 220244
rect 429620 220204 432052 220232
rect 429620 220192 429626 220204
rect 432046 220192 432052 220204
rect 432104 220192 432110 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 473170 220192 473176 220244
rect 473228 220232 473234 220244
rect 482002 220232 482008 220244
rect 473228 220204 482008 220232
rect 473228 220192 473234 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495342 220232 495348 220244
rect 482980 220204 495348 220232
rect 482980 220192 482986 220204
rect 495342 220192 495348 220204
rect 495400 220192 495406 220244
rect 497458 220192 497464 220244
rect 497516 220232 497522 220244
rect 515214 220232 515220 220244
rect 497516 220204 515220 220232
rect 497516 220192 497522 220204
rect 515214 220192 515220 220204
rect 515272 220192 515278 220244
rect 515398 220192 515404 220244
rect 515456 220232 515462 220244
rect 530026 220232 530032 220244
rect 515456 220204 530032 220232
rect 515456 220192 515462 220204
rect 530026 220192 530032 220204
rect 530084 220192 530090 220244
rect 531130 220192 531136 220244
rect 531188 220232 531194 220244
rect 552290 220232 552296 220244
rect 531188 220204 552296 220232
rect 531188 220192 531194 220204
rect 552290 220192 552296 220204
rect 552348 220192 552354 220244
rect 552658 220192 552664 220244
rect 552716 220232 552722 220244
rect 552716 220204 563054 220232
rect 552716 220192 552722 220204
rect 563026 220164 563054 220204
rect 576762 220192 576768 220244
rect 576820 220232 576826 220244
rect 610066 220232 610072 220244
rect 576820 220204 610072 220232
rect 576820 220192 576826 220204
rect 610066 220192 610072 220204
rect 610124 220192 610130 220244
rect 576578 220164 576584 220176
rect 563026 220136 576584 220164
rect 576578 220124 576584 220136
rect 576636 220124 576642 220176
rect 214282 220096 214288 220108
rect 211908 220068 214288 220096
rect 214282 220056 214288 220068
rect 214340 220056 214346 220108
rect 214558 220056 214564 220108
rect 214616 220096 214622 220108
rect 229278 220096 229284 220108
rect 214616 220068 229284 220096
rect 214616 220056 214622 220068
rect 229278 220056 229284 220068
rect 229336 220056 229342 220108
rect 230198 220056 230204 220108
rect 230256 220096 230262 220108
rect 275278 220096 275284 220108
rect 230256 220068 275284 220096
rect 230256 220056 230262 220068
rect 275278 220056 275284 220068
rect 275336 220056 275342 220108
rect 292482 220056 292488 220108
rect 292540 220096 292546 220108
rect 326154 220096 326160 220108
rect 292540 220068 326160 220096
rect 292540 220056 292546 220068
rect 326154 220056 326160 220068
rect 326212 220056 326218 220108
rect 328914 220056 328920 220108
rect 328972 220096 328978 220108
rect 354766 220096 354772 220108
rect 328972 220068 354772 220096
rect 328972 220056 328978 220068
rect 354766 220056 354772 220068
rect 354824 220056 354830 220108
rect 355410 220056 355416 220108
rect 355468 220096 355474 220108
rect 375558 220096 375564 220108
rect 355468 220068 375564 220096
rect 355468 220056 355474 220068
rect 375558 220056 375564 220068
rect 375616 220056 375622 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426710 220096 426716 220108
rect 421708 220068 426716 220096
rect 421708 220056 421714 220068
rect 426710 220056 426716 220068
rect 426768 220056 426774 220108
rect 431954 220056 431960 220108
rect 432012 220096 432018 220108
rect 434806 220096 434812 220108
rect 432012 220068 434812 220096
rect 432012 220056 432018 220068
rect 434806 220056 434812 220068
rect 434864 220056 434870 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 489638 220056 489644 220108
rect 489696 220096 489702 220108
rect 504358 220096 504364 220108
rect 489696 220068 504364 220096
rect 489696 220056 489702 220068
rect 504358 220056 504364 220068
rect 504416 220056 504422 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 558178 220096 558184 220108
rect 538180 220068 558184 220096
rect 538180 220056 538186 220068
rect 558178 220056 558184 220068
rect 558236 220056 558242 220108
rect 582466 220056 582472 220108
rect 582524 220096 582530 220108
rect 633434 220096 633440 220108
rect 582524 220068 633440 220096
rect 582524 220056 582530 220068
rect 633434 220056 633440 220068
rect 633492 220056 633498 220108
rect 558362 219988 558368 220040
rect 558420 220028 558426 220040
rect 576762 220028 576768 220040
rect 558420 220000 576768 220028
rect 558420 219988 558426 220000
rect 576762 219988 576768 220000
rect 576820 219988 576826 220040
rect 576946 219988 576952 220040
rect 577004 220028 577010 220040
rect 581638 220028 581644 220040
rect 577004 220000 581644 220028
rect 577004 219988 577010 220000
rect 581638 219988 581644 220000
rect 581696 219988 581702 220040
rect 581822 219988 581828 220040
rect 581880 220028 581886 220040
rect 582328 220028 582334 220040
rect 581880 220000 582334 220028
rect 581880 219988 581886 220000
rect 582328 219988 582334 220000
rect 582386 219988 582392 220040
rect 107838 219920 107844 219972
rect 107896 219960 107902 219972
rect 127618 219960 127624 219972
rect 107896 219932 127624 219960
rect 107896 219920 107902 219932
rect 127618 219920 127624 219932
rect 127676 219920 127682 219972
rect 127802 219920 127808 219972
rect 127860 219960 127866 219972
rect 127860 219932 185348 219960
rect 127860 219920 127866 219932
rect 185320 219892 185348 219932
rect 185762 219920 185768 219972
rect 185820 219960 185826 219972
rect 185820 219932 190316 219960
rect 185820 219920 185826 219932
rect 185320 219864 185440 219892
rect 114462 219784 114468 219836
rect 114520 219824 114526 219836
rect 185118 219824 185124 219836
rect 114520 219796 185124 219824
rect 114520 219784 114526 219796
rect 185118 219784 185124 219796
rect 185176 219784 185182 219836
rect 185412 219824 185440 219864
rect 190086 219824 190092 219836
rect 185412 219796 190092 219824
rect 190086 219784 190092 219796
rect 190144 219784 190150 219836
rect 190288 219824 190316 219932
rect 190638 219920 190644 219972
rect 190696 219960 190702 219972
rect 244458 219960 244464 219972
rect 190696 219932 244464 219960
rect 190696 219920 190702 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 253566 219920 253572 219972
rect 253624 219960 253630 219972
rect 293310 219960 293316 219972
rect 253624 219932 293316 219960
rect 253624 219920 253630 219932
rect 293310 219920 293316 219932
rect 293368 219920 293374 219972
rect 527542 219852 527548 219904
rect 527600 219892 527606 219904
rect 527600 219864 528554 219892
rect 527600 219852 527606 219864
rect 202782 219824 202788 219836
rect 190288 219796 202788 219824
rect 202782 219784 202788 219796
rect 202840 219784 202846 219836
rect 252738 219824 252744 219836
rect 202984 219796 252744 219824
rect 121086 219648 121092 219700
rect 121144 219688 121150 219700
rect 121144 219660 122834 219688
rect 121144 219648 121150 219660
rect 122806 219552 122834 219660
rect 127618 219648 127624 219700
rect 127676 219688 127682 219700
rect 140774 219688 140780 219700
rect 127676 219660 140780 219688
rect 127676 219648 127682 219660
rect 140774 219648 140780 219660
rect 140832 219648 140838 219700
rect 140958 219648 140964 219700
rect 141016 219688 141022 219700
rect 141016 219660 200988 219688
rect 141016 219648 141022 219660
rect 127802 219552 127808 219564
rect 122806 219524 127808 219552
rect 127802 219512 127808 219524
rect 127860 219512 127866 219564
rect 134334 219512 134340 219564
rect 134392 219552 134398 219564
rect 200758 219552 200764 219564
rect 134392 219524 200764 219552
rect 134392 219512 134398 219524
rect 200758 219512 200764 219524
rect 200816 219512 200822 219564
rect 200960 219552 200988 219660
rect 201126 219648 201132 219700
rect 201184 219688 201190 219700
rect 202984 219688 203012 219796
rect 252738 219784 252744 219796
rect 252796 219784 252802 219836
rect 270770 219784 270776 219836
rect 270828 219824 270834 219836
rect 279142 219824 279148 219836
rect 270828 219796 279148 219824
rect 270828 219784 270834 219796
rect 279142 219784 279148 219796
rect 279200 219784 279206 219836
rect 286686 219784 286692 219836
rect 286744 219824 286750 219836
rect 319070 219824 319076 219836
rect 286744 219796 319076 219824
rect 286744 219784 286750 219796
rect 319070 219784 319076 219796
rect 319128 219784 319134 219836
rect 528526 219756 528554 219864
rect 530026 219852 530032 219904
rect 530084 219892 530090 219904
rect 552658 219892 552664 219904
rect 530084 219864 552664 219892
rect 530084 219852 530090 219864
rect 552658 219852 552664 219864
rect 552716 219852 552722 219904
rect 552842 219852 552848 219904
rect 552900 219892 552906 219904
rect 598382 219892 598388 219904
rect 552900 219864 598388 219892
rect 552900 219852 552906 219864
rect 598382 219852 598388 219864
rect 598440 219852 598446 219904
rect 598566 219852 598572 219904
rect 598624 219892 598630 219904
rect 598624 219864 615494 219892
rect 598624 219852 598630 219864
rect 558362 219756 558368 219768
rect 528526 219728 558368 219756
rect 558362 219716 558368 219728
rect 558420 219716 558426 219768
rect 558546 219716 558552 219768
rect 558604 219756 558610 219768
rect 608594 219756 608600 219768
rect 558604 219728 608600 219756
rect 558604 219716 558610 219728
rect 608594 219716 608600 219728
rect 608652 219716 608658 219768
rect 615466 219756 615494 219864
rect 620002 219756 620008 219768
rect 615466 219728 620008 219756
rect 620002 219716 620008 219728
rect 620060 219716 620066 219768
rect 201184 219660 203012 219688
rect 201184 219648 201190 219660
rect 203150 219648 203156 219700
rect 203208 219688 203214 219700
rect 203208 219660 206048 219688
rect 203208 219648 203214 219660
rect 205818 219552 205824 219564
rect 200960 219524 205824 219552
rect 205818 219512 205824 219524
rect 205876 219512 205882 219564
rect 206020 219552 206048 219660
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 506014 219580 506020 219632
rect 506072 219620 506078 219632
rect 576762 219620 576768 219632
rect 506072 219592 576768 219620
rect 506072 219580 506078 219592
rect 576762 219580 576768 219592
rect 576820 219580 576826 219632
rect 581638 219580 581644 219632
rect 581696 219620 581702 219632
rect 582328 219620 582334 219632
rect 581696 219592 582334 219620
rect 581696 219580 581702 219592
rect 582328 219580 582334 219592
rect 582386 219580 582392 219632
rect 582466 219580 582472 219632
rect 582524 219620 582530 219632
rect 598566 219620 598572 219632
rect 582524 219592 598572 219620
rect 582524 219580 582530 219592
rect 598566 219580 598572 219592
rect 598624 219580 598630 219632
rect 619818 219620 619824 219632
rect 598768 219592 619824 219620
rect 208578 219552 208584 219564
rect 206020 219524 208584 219552
rect 208578 219512 208584 219524
rect 208636 219512 208642 219564
rect 211706 219512 211712 219564
rect 211764 219552 211770 219564
rect 215938 219552 215944 219564
rect 211764 219524 215944 219552
rect 211764 219512 211770 219524
rect 215938 219512 215944 219524
rect 215996 219512 216002 219564
rect 366726 219512 366732 219564
rect 366784 219552 366790 219564
rect 366784 219524 367048 219552
rect 366784 219512 366790 219524
rect 105814 219444 105820 219496
rect 105872 219484 105878 219496
rect 105872 219456 106182 219484
rect 105872 219444 105878 219456
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 106154 219416 106182 219456
rect 289832 219456 291332 219484
rect 147122 219416 147128 219428
rect 106154 219388 147128 219416
rect 147122 219376 147128 219388
rect 147180 219376 147186 219428
rect 148410 219376 148416 219428
rect 148468 219416 148474 219428
rect 148962 219416 148968 219428
rect 148468 219388 148968 219416
rect 148468 219376 148474 219388
rect 148962 219376 148968 219388
rect 149020 219376 149026 219428
rect 149238 219376 149244 219428
rect 149296 219416 149302 219428
rect 149974 219416 149980 219428
rect 149296 219388 149980 219416
rect 149296 219376 149302 219388
rect 149974 219376 149980 219388
rect 150032 219376 150038 219428
rect 152550 219376 152556 219428
rect 152608 219416 152614 219428
rect 153102 219416 153108 219428
rect 152608 219388 153108 219416
rect 152608 219376 152614 219388
rect 153102 219376 153108 219388
rect 153160 219376 153166 219428
rect 159174 219376 159180 219428
rect 159232 219416 159238 219428
rect 160002 219416 160008 219428
rect 159232 219388 160008 219416
rect 159232 219376 159238 219388
rect 160002 219376 160008 219388
rect 160060 219376 160066 219428
rect 163314 219376 163320 219428
rect 163372 219416 163378 219428
rect 163958 219416 163964 219428
rect 163372 219388 163964 219416
rect 163372 219376 163378 219388
rect 163958 219376 163964 219388
rect 164016 219376 164022 219428
rect 204530 219416 204536 219428
rect 166966 219388 204536 219416
rect 106918 219280 106924 219292
rect 64846 219252 106924 219280
rect 63126 219104 63132 219156
rect 63184 219144 63190 219156
rect 64846 219144 64874 219252
rect 106918 219240 106924 219252
rect 106976 219240 106982 219292
rect 113634 219240 113640 219292
rect 113692 219280 113698 219292
rect 152366 219280 152372 219292
rect 113692 219252 152372 219280
rect 113692 219240 113698 219252
rect 152366 219240 152372 219252
rect 152424 219240 152430 219292
rect 153194 219240 153200 219292
rect 153252 219280 153258 219292
rect 153838 219280 153844 219292
rect 153252 219252 153844 219280
rect 153252 219240 153258 219252
rect 153838 219240 153844 219252
rect 153896 219240 153902 219292
rect 160002 219240 160008 219292
rect 160060 219280 160066 219292
rect 166966 219280 166994 219388
rect 204530 219376 204536 219388
rect 204588 219376 204594 219428
rect 209682 219376 209688 219428
rect 209740 219416 209746 219428
rect 210418 219416 210424 219428
rect 209740 219388 210424 219416
rect 209740 219376 209746 219388
rect 210418 219376 210424 219388
rect 210476 219376 210482 219428
rect 212994 219376 213000 219428
rect 213052 219416 213058 219428
rect 258074 219416 258080 219428
rect 213052 219388 258080 219416
rect 213052 219376 213058 219388
rect 258074 219376 258080 219388
rect 258132 219376 258138 219428
rect 272886 219376 272892 219428
rect 272944 219416 272950 219428
rect 289832 219416 289860 219456
rect 272944 219388 289860 219416
rect 291304 219416 291332 219456
rect 367020 219434 367048 219524
rect 576964 219524 579752 219552
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 297358 219416 297364 219428
rect 291304 219388 297364 219416
rect 272944 219376 272950 219388
rect 297358 219376 297364 219388
rect 297416 219376 297422 219428
rect 304074 219376 304080 219428
rect 304132 219416 304138 219428
rect 308398 219416 308404 219428
rect 304132 219388 308404 219416
rect 304132 219376 304138 219388
rect 308398 219376 308404 219388
rect 308456 219376 308462 219428
rect 310974 219376 310980 219428
rect 311032 219416 311038 219428
rect 322198 219416 322204 219428
rect 311032 219388 322204 219416
rect 311032 219376 311038 219388
rect 322198 219376 322204 219388
rect 322256 219376 322262 219428
rect 341334 219376 341340 219428
rect 341392 219416 341398 219428
rect 342254 219416 342260 219428
rect 341392 219388 342260 219416
rect 341392 219376 341398 219388
rect 342254 219376 342260 219388
rect 342312 219376 342318 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 349614 219376 349620 219428
rect 349672 219416 349678 219428
rect 350534 219416 350540 219428
rect 349672 219388 350540 219416
rect 349672 219376 349678 219388
rect 350534 219376 350540 219388
rect 350592 219376 350598 219428
rect 366174 219376 366180 219428
rect 366232 219416 366238 219428
rect 366928 219416 367048 219434
rect 366232 219406 367048 219416
rect 366232 219388 366956 219406
rect 366232 219376 366238 219388
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 501046 219444 501052 219496
rect 501104 219484 501110 219496
rect 576964 219484 576992 219524
rect 501104 219456 576992 219484
rect 579724 219484 579752 219524
rect 591574 219484 591580 219496
rect 579724 219456 591580 219484
rect 501104 219444 501110 219456
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 438210 219376 438216 219428
rect 438268 219416 438274 219428
rect 438854 219416 438860 219428
rect 438268 219388 438860 219416
rect 438268 219376 438274 219388
rect 438854 219376 438860 219388
rect 438912 219376 438918 219428
rect 439866 219376 439872 219428
rect 439924 219416 439930 219428
rect 440326 219416 440332 219428
rect 439924 219388 440332 219416
rect 439924 219376 439930 219388
rect 440326 219376 440332 219388
rect 440384 219376 440390 219428
rect 577130 219394 577136 219446
rect 577188 219434 577194 219446
rect 591574 219444 591580 219456
rect 591632 219444 591638 219496
rect 598768 219484 598796 219592
rect 619818 219580 619824 219592
rect 619876 219580 619882 219632
rect 591776 219456 598796 219484
rect 577188 219406 579614 219434
rect 577188 219394 577194 219406
rect 553210 219308 553216 219360
rect 553268 219348 553274 219360
rect 558546 219348 558552 219360
rect 553268 219320 558552 219348
rect 553268 219308 553274 219320
rect 558546 219308 558552 219320
rect 558604 219308 558610 219360
rect 572438 219308 572444 219360
rect 572496 219348 572502 219360
rect 574646 219348 574652 219360
rect 572496 219320 574652 219348
rect 572496 219308 572502 219320
rect 574646 219308 574652 219320
rect 574704 219308 574710 219360
rect 579586 219348 579614 219406
rect 582466 219348 582472 219360
rect 579586 219320 582472 219348
rect 582466 219308 582472 219320
rect 582524 219308 582530 219360
rect 582650 219308 582656 219360
rect 582708 219348 582714 219360
rect 591776 219348 591804 219456
rect 598934 219444 598940 219496
rect 598992 219484 598998 219496
rect 607490 219484 607496 219496
rect 598992 219456 607496 219484
rect 598992 219444 598998 219456
rect 607490 219444 607496 219456
rect 607548 219444 607554 219496
rect 672994 219376 673000 219428
rect 673052 219416 673058 219428
rect 673454 219416 673460 219428
rect 673052 219388 673460 219416
rect 673052 219376 673058 219388
rect 673454 219376 673460 219388
rect 673512 219376 673518 219428
rect 582708 219320 591804 219348
rect 582708 219308 582714 219320
rect 591942 219308 591948 219360
rect 592000 219348 592006 219360
rect 596818 219348 596824 219360
rect 592000 219320 596824 219348
rect 592000 219308 592006 219320
rect 596818 219308 596824 219320
rect 596876 219308 596882 219360
rect 160060 219252 166994 219280
rect 160060 219240 160066 219252
rect 169110 219240 169116 219292
rect 169168 219280 169174 219292
rect 169662 219280 169668 219292
rect 169168 219252 169668 219280
rect 169168 219240 169174 219252
rect 169662 219240 169668 219252
rect 169720 219240 169726 219292
rect 171594 219240 171600 219292
rect 171652 219280 171658 219292
rect 172146 219280 172152 219292
rect 171652 219252 172152 219280
rect 171652 219240 171658 219252
rect 172146 219240 172152 219252
rect 172204 219240 172210 219292
rect 172422 219240 172428 219292
rect 172480 219280 172486 219292
rect 173342 219280 173348 219292
rect 172480 219252 173348 219280
rect 172480 219240 172486 219252
rect 173342 219240 173348 219252
rect 173400 219240 173406 219292
rect 182358 219240 182364 219292
rect 182416 219280 182422 219292
rect 189718 219280 189724 219292
rect 182416 219252 189724 219280
rect 182416 219240 182422 219252
rect 189718 219240 189724 219252
rect 189776 219240 189782 219292
rect 192294 219240 192300 219292
rect 192352 219280 192358 219292
rect 192938 219280 192944 219292
rect 192352 219252 192944 219280
rect 192352 219240 192358 219252
rect 192938 219240 192944 219252
rect 192996 219240 193002 219292
rect 193122 219240 193128 219292
rect 193180 219280 193186 219292
rect 198182 219280 198188 219292
rect 193180 219252 198188 219280
rect 193180 219240 193186 219252
rect 198182 219240 198188 219252
rect 198240 219240 198246 219292
rect 198918 219240 198924 219292
rect 198976 219280 198982 219292
rect 200022 219280 200028 219292
rect 198976 219252 200028 219280
rect 198976 219240 198982 219252
rect 200022 219240 200028 219252
rect 200080 219240 200086 219292
rect 202598 219240 202604 219292
rect 202656 219280 202662 219292
rect 207658 219280 207664 219292
rect 202656 219252 207664 219280
rect 202656 219240 202662 219252
rect 207658 219240 207664 219252
rect 207716 219240 207722 219292
rect 211338 219240 211344 219292
rect 211396 219280 211402 219292
rect 218054 219280 218060 219292
rect 211396 219252 218060 219280
rect 211396 219240 211402 219252
rect 218054 219240 218060 219252
rect 218112 219240 218118 219292
rect 239490 219240 239496 219292
rect 239548 219280 239554 219292
rect 272702 219280 272708 219292
rect 239548 219252 272708 219280
rect 239548 219240 239554 219252
rect 272702 219240 272708 219252
rect 272760 219240 272766 219292
rect 279050 219240 279056 219292
rect 279108 219280 279114 219292
rect 286318 219280 286324 219292
rect 279108 219252 286324 219280
rect 279108 219240 279114 219252
rect 286318 219240 286324 219252
rect 286376 219240 286382 219292
rect 291654 219240 291660 219292
rect 291712 219280 291718 219292
rect 313918 219280 313924 219292
rect 291712 219252 313924 219280
rect 291712 219240 291718 219252
rect 313918 219240 313924 219252
rect 313976 219240 313982 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 561858 219240 561864 219292
rect 561916 219280 561922 219292
rect 565078 219280 565084 219292
rect 561916 219252 565084 219280
rect 561916 219240 561922 219252
rect 565078 219240 565084 219252
rect 565136 219240 565142 219292
rect 568390 219240 568396 219292
rect 568448 219280 568454 219292
rect 571978 219280 571984 219292
rect 568448 219252 571984 219280
rect 568448 219240 568454 219252
rect 571978 219240 571984 219252
rect 572036 219240 572042 219292
rect 355226 219212 355232 219224
rect 335326 219184 355232 219212
rect 63184 219116 64874 219144
rect 63184 219104 63190 219116
rect 70578 219104 70584 219156
rect 70636 219144 70642 219156
rect 117958 219144 117964 219156
rect 70636 219116 117964 219144
rect 70636 219104 70642 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 132586 219104 132592 219156
rect 132644 219144 132650 219156
rect 177482 219144 177488 219156
rect 132644 219116 177488 219144
rect 132644 219104 132650 219116
rect 177482 219104 177488 219116
rect 177540 219104 177546 219156
rect 179046 219104 179052 219156
rect 179104 219144 179110 219156
rect 195882 219144 195888 219156
rect 179104 219116 195888 219144
rect 179104 219104 179110 219116
rect 195882 219104 195888 219116
rect 195940 219104 195946 219156
rect 199746 219104 199752 219156
rect 199804 219144 199810 219156
rect 243538 219144 243544 219156
rect 199804 219116 243544 219144
rect 199804 219104 199810 219116
rect 243538 219104 243544 219116
rect 243596 219104 243602 219156
rect 272334 219104 272340 219156
rect 272392 219144 272398 219156
rect 272392 219116 291884 219144
rect 272392 219104 272398 219116
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 77202 218968 77208 219020
rect 77260 219008 77266 219020
rect 140038 219008 140044 219020
rect 77260 218980 140044 219008
rect 77260 218968 77266 218980
rect 140038 218968 140044 218980
rect 140096 218968 140102 219020
rect 153194 219008 153200 219020
rect 142126 218980 153200 219008
rect 50706 218832 50712 218884
rect 50764 218872 50770 218884
rect 62758 218872 62764 218884
rect 50764 218844 62764 218872
rect 50764 218832 50770 218844
rect 62758 218832 62764 218844
rect 62816 218832 62822 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 142126 218872 142154 218980
rect 153194 218968 153200 218980
rect 153252 218968 153258 219020
rect 153378 218968 153384 219020
rect 153436 219008 153442 219020
rect 203518 219008 203524 219020
rect 153436 218980 203524 219008
rect 153436 218968 153442 218980
rect 203518 218968 203524 218980
rect 203576 218968 203582 219020
rect 206370 218968 206376 219020
rect 206428 219008 206434 219020
rect 253842 219008 253848 219020
rect 206428 218980 253848 219008
rect 206428 218968 206434 218980
rect 253842 218968 253848 218980
rect 253900 218968 253906 219020
rect 259178 218968 259184 219020
rect 259236 219008 259242 219020
rect 291470 219008 291476 219020
rect 259236 218980 291476 219008
rect 259236 218968 259242 218980
rect 291470 218968 291476 218980
rect 291528 218968 291534 219020
rect 83884 218844 142154 218872
rect 83884 218832 83890 218844
rect 142430 218832 142436 218884
rect 142488 218872 142494 218884
rect 152182 218872 152188 218884
rect 142488 218844 152188 218872
rect 142488 218832 142494 218844
rect 152182 218832 152188 218844
rect 152240 218832 152246 218884
rect 152366 218832 152372 218884
rect 152424 218872 152430 218884
rect 162118 218872 162124 218884
rect 152424 218844 162124 218872
rect 152424 218832 152430 218844
rect 162118 218832 162124 218844
rect 162176 218832 162182 218884
rect 162486 218832 162492 218884
rect 162544 218872 162550 218884
rect 169754 218872 169760 218884
rect 162544 218844 169760 218872
rect 162544 218832 162550 218844
rect 169754 218832 169760 218844
rect 169812 218832 169818 218884
rect 169938 218832 169944 218884
rect 169996 218872 170002 218884
rect 171042 218872 171048 218884
rect 169996 218844 171048 218872
rect 169996 218832 170002 218844
rect 171042 218832 171048 218844
rect 171100 218832 171106 218884
rect 180058 218872 180064 218884
rect 171796 218844 180064 218872
rect 59814 218696 59820 218748
rect 59872 218736 59878 218748
rect 143718 218736 143724 218748
rect 59872 218708 143724 218736
rect 59872 218696 59878 218708
rect 143718 218696 143724 218708
rect 143776 218696 143782 218748
rect 146754 218696 146760 218748
rect 146812 218736 146818 218748
rect 161934 218736 161940 218748
rect 146812 218708 161940 218736
rect 146812 218696 146818 218708
rect 161934 218696 161940 218708
rect 161992 218696 161998 218748
rect 165798 218696 165804 218748
rect 165856 218736 165862 218748
rect 171796 218736 171824 218844
rect 180058 218832 180064 218844
rect 180116 218832 180122 218884
rect 180766 218844 184612 218872
rect 165856 218708 171824 218736
rect 165856 218696 165862 218708
rect 175734 218696 175740 218748
rect 175792 218736 175798 218748
rect 180766 218736 180794 218844
rect 175792 218708 180794 218736
rect 175792 218696 175798 218708
rect 181162 218696 181168 218748
rect 181220 218736 181226 218748
rect 184382 218736 184388 218748
rect 181220 218708 184388 218736
rect 181220 218696 181226 218708
rect 184382 218696 184388 218708
rect 184440 218696 184446 218748
rect 184584 218736 184612 218844
rect 188982 218832 188988 218884
rect 189040 218872 189046 218884
rect 194134 218872 194140 218884
rect 189040 218844 194140 218872
rect 189040 218832 189046 218844
rect 194134 218832 194140 218844
rect 194192 218832 194198 218884
rect 194318 218832 194324 218884
rect 194376 218872 194382 218884
rect 239306 218872 239312 218884
rect 194376 218844 239312 218872
rect 194376 218832 194382 218844
rect 239306 218832 239312 218844
rect 239364 218832 239370 218884
rect 246114 218832 246120 218884
rect 246172 218872 246178 218884
rect 279050 218872 279056 218884
rect 246172 218844 279056 218872
rect 246172 218832 246178 218844
rect 279050 218832 279056 218844
rect 279108 218832 279114 218884
rect 279234 218832 279240 218884
rect 279292 218872 279298 218884
rect 279292 218844 282316 218872
rect 279292 218832 279298 218844
rect 189626 218736 189632 218748
rect 184584 218708 189632 218736
rect 189626 218696 189632 218708
rect 189684 218696 189690 218748
rect 189810 218696 189816 218748
rect 189868 218736 189874 218748
rect 195330 218736 195336 218748
rect 189868 218708 195336 218736
rect 189868 218696 189874 218708
rect 195330 218696 195336 218708
rect 195388 218696 195394 218748
rect 195606 218696 195612 218748
rect 195664 218736 195670 218748
rect 197998 218736 198004 218748
rect 195664 218708 198004 218736
rect 195664 218696 195670 218708
rect 197998 218696 198004 218708
rect 198056 218696 198062 218748
rect 198182 218696 198188 218748
rect 198240 218736 198246 218748
rect 246298 218736 246304 218748
rect 198240 218708 246304 218736
rect 198240 218696 198246 218708
rect 246298 218696 246304 218708
rect 246356 218696 246362 218748
rect 252738 218696 252744 218748
rect 252796 218736 252802 218748
rect 252796 218708 282224 218736
rect 252796 218696 252802 218708
rect 100386 218560 100392 218612
rect 100444 218600 100450 218612
rect 105814 218600 105820 218612
rect 100444 218572 105820 218600
rect 100444 218560 100450 218572
rect 105814 218560 105820 218572
rect 105872 218560 105878 218612
rect 107010 218560 107016 218612
rect 107068 218600 107074 218612
rect 142430 218600 142436 218612
rect 107068 218572 142436 218600
rect 107068 218560 107074 218572
rect 142430 218560 142436 218572
rect 142488 218560 142494 218612
rect 142614 218560 142620 218612
rect 142672 218600 142678 218612
rect 143258 218600 143264 218612
rect 142672 218572 143264 218600
rect 142672 218560 142678 218572
rect 143258 218560 143264 218572
rect 143316 218560 143322 218612
rect 144270 218560 144276 218612
rect 144328 218600 144334 218612
rect 144822 218600 144828 218612
rect 144328 218572 144828 218600
rect 144328 218560 144334 218572
rect 144822 218560 144828 218572
rect 144880 218560 144886 218612
rect 145098 218560 145104 218612
rect 145156 218600 145162 218612
rect 145926 218600 145932 218612
rect 145156 218572 145932 218600
rect 145156 218560 145162 218572
rect 145926 218560 145932 218572
rect 145984 218560 145990 218612
rect 165614 218600 165620 218612
rect 157306 218572 165620 218600
rect 120258 218424 120264 218476
rect 120316 218464 120322 218476
rect 157306 218464 157334 218572
rect 165614 218560 165620 218572
rect 165672 218560 165678 218612
rect 166626 218560 166632 218612
rect 166684 218600 166690 218612
rect 202598 218600 202604 218612
rect 166684 218572 202604 218600
rect 166684 218560 166690 218572
rect 202598 218560 202604 218572
rect 202656 218560 202662 218612
rect 203058 218560 203064 218612
rect 203116 218600 203122 218612
rect 206186 218600 206192 218612
rect 203116 218572 206192 218600
rect 203116 218560 203122 218572
rect 206186 218560 206192 218572
rect 206244 218560 206250 218612
rect 208026 218560 208032 218612
rect 208084 218600 208090 218612
rect 208084 218572 209774 218600
rect 208084 218560 208090 218572
rect 120316 218436 157334 218464
rect 120316 218424 120322 218436
rect 161934 218424 161940 218476
rect 161992 218464 161998 218476
rect 169570 218464 169576 218476
rect 161992 218436 169576 218464
rect 161992 218424 161998 218436
rect 169570 218424 169576 218436
rect 169628 218424 169634 218476
rect 169754 218424 169760 218476
rect 169812 218464 169818 218476
rect 181346 218464 181352 218476
rect 169812 218436 181352 218464
rect 169812 218424 169818 218436
rect 181346 218424 181352 218436
rect 181404 218424 181410 218476
rect 186498 218424 186504 218476
rect 186556 218464 186562 218476
rect 194318 218464 194324 218476
rect 186556 218436 194324 218464
rect 186556 218424 186562 218436
rect 194318 218424 194324 218436
rect 194376 218424 194382 218476
rect 198090 218424 198096 218476
rect 198148 218464 198154 218476
rect 200390 218464 200396 218476
rect 198148 218436 200396 218464
rect 198148 218424 198154 218436
rect 200390 218424 200396 218436
rect 200448 218424 200454 218476
rect 202230 218424 202236 218476
rect 202288 218464 202294 218476
rect 202782 218464 202788 218476
rect 202288 218436 202788 218464
rect 202288 218424 202294 218436
rect 202782 218424 202788 218436
rect 202840 218424 202846 218476
rect 204714 218424 204720 218476
rect 204772 218464 204778 218476
rect 207842 218464 207848 218476
rect 204772 218436 207848 218464
rect 204772 218424 204778 218436
rect 207842 218424 207848 218436
rect 207900 218424 207906 218476
rect 208854 218424 208860 218476
rect 208912 218464 208918 218476
rect 209498 218464 209504 218476
rect 208912 218436 209504 218464
rect 208912 218424 208918 218436
rect 209498 218424 209504 218436
rect 209556 218424 209562 218476
rect 209746 218464 209774 218572
rect 210142 218560 210148 218612
rect 210200 218600 210206 218612
rect 217318 218600 217324 218612
rect 210200 218572 217324 218600
rect 210200 218560 210206 218572
rect 217318 218560 217324 218572
rect 217376 218560 217382 218612
rect 219618 218560 219624 218612
rect 219676 218600 219682 218612
rect 264606 218600 264612 218612
rect 219676 218572 264612 218600
rect 219676 218560 219682 218572
rect 264606 218560 264612 218572
rect 264664 218560 264670 218612
rect 265986 218560 265992 218612
rect 266044 218600 266050 218612
rect 272334 218600 272340 218612
rect 266044 218572 272340 218600
rect 266044 218560 266050 218572
rect 272334 218560 272340 218572
rect 272392 218560 272398 218612
rect 272702 218560 272708 218612
rect 272760 218600 272766 218612
rect 279418 218600 279424 218612
rect 272760 218572 279424 218600
rect 272760 218560 272766 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 211522 218464 211528 218476
rect 209746 218436 211528 218464
rect 211522 218424 211528 218436
rect 211580 218424 211586 218476
rect 217962 218424 217968 218476
rect 218020 218464 218026 218476
rect 223482 218464 223488 218476
rect 218020 218436 223488 218464
rect 218020 218424 218026 218436
rect 223482 218424 223488 218436
rect 223540 218424 223546 218476
rect 225966 218424 225972 218476
rect 226024 218464 226030 218476
rect 266998 218464 267004 218476
rect 226024 218436 267004 218464
rect 226024 218424 226030 218436
rect 266998 218424 267004 218436
rect 267056 218424 267062 218476
rect 282196 218464 282224 218708
rect 282288 218600 282316 218844
rect 285858 218832 285864 218884
rect 285916 218872 285922 218884
rect 291654 218872 291660 218884
rect 285916 218844 291660 218872
rect 285916 218832 285922 218844
rect 291654 218832 291660 218844
rect 291712 218832 291718 218884
rect 291856 218872 291884 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 307386 219104 307392 219156
rect 307444 219144 307450 219156
rect 331858 219144 331864 219156
rect 307444 219116 331864 219144
rect 307444 219104 307450 219116
rect 331858 219104 331864 219116
rect 331916 219104 331922 219156
rect 333698 219104 333704 219156
rect 333756 219144 333762 219156
rect 335326 219144 335354 219184
rect 355226 219172 355232 219184
rect 355284 219172 355290 219224
rect 333756 219116 335354 219144
rect 333756 219104 333762 219116
rect 362034 219104 362040 219156
rect 362092 219144 362098 219156
rect 370958 219144 370964 219156
rect 362092 219116 370964 219144
rect 362092 219104 362098 219116
rect 370958 219104 370964 219116
rect 371016 219104 371022 219156
rect 552658 219104 552664 219156
rect 552716 219144 552722 219156
rect 558178 219144 558184 219156
rect 552716 219116 558184 219144
rect 552716 219104 552722 219116
rect 558178 219104 558184 219116
rect 558236 219104 558242 219156
rect 563054 219104 563060 219156
rect 563112 219144 563118 219156
rect 563974 219144 563980 219156
rect 563112 219116 563980 219144
rect 563112 219104 563118 219116
rect 563974 219104 563980 219116
rect 564032 219104 564038 219156
rect 567286 219104 567292 219156
rect 567344 219144 567350 219156
rect 626350 219144 626356 219156
rect 567344 219116 626356 219144
rect 567344 219104 567350 219116
rect 626350 219104 626356 219116
rect 626408 219104 626414 219156
rect 294138 218968 294144 219020
rect 294196 219008 294202 219020
rect 311158 219008 311164 219020
rect 294196 218980 311164 219008
rect 294196 218968 294202 218980
rect 311158 218968 311164 218980
rect 311216 218968 311222 219020
rect 325326 218968 325332 219020
rect 325384 219008 325390 219020
rect 327718 219008 327724 219020
rect 325384 218980 327724 219008
rect 325384 218968 325390 218980
rect 327718 218968 327724 218980
rect 327776 218968 327782 219020
rect 330478 218968 330484 219020
rect 330536 219008 330542 219020
rect 330536 218980 345014 219008
rect 330536 218968 330542 218980
rect 297542 218872 297548 218884
rect 291856 218844 297548 218872
rect 297542 218832 297548 218844
rect 297600 218832 297606 218884
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 340322 218872 340328 218884
rect 314068 218844 340328 218872
rect 314068 218832 314074 218844
rect 340322 218832 340328 218844
rect 340380 218832 340386 218884
rect 344986 218872 345014 218980
rect 357066 218968 357072 219020
rect 357124 219008 357130 219020
rect 369118 219008 369124 219020
rect 357124 218980 369124 219008
rect 357124 218968 357130 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 370314 218968 370320 219020
rect 370372 219008 370378 219020
rect 380066 219008 380072 219020
rect 370372 218980 380072 219008
rect 370372 218968 370378 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 380250 218968 380256 219020
rect 380308 219008 380314 219020
rect 388622 219008 388628 219020
rect 380308 218980 388628 219008
rect 380308 218968 380314 218980
rect 388622 218968 388628 218980
rect 388680 218968 388686 219020
rect 552474 218968 552480 219020
rect 552532 219008 552538 219020
rect 552532 218980 569448 219008
rect 552532 218968 552538 218980
rect 345658 218872 345664 218884
rect 344986 218844 345664 218872
rect 345658 218832 345664 218844
rect 345716 218832 345722 218884
rect 347038 218832 347044 218884
rect 347096 218872 347102 218884
rect 363506 218872 363512 218884
rect 347096 218844 363512 218872
rect 347096 218832 347102 218844
rect 363506 218832 363512 218844
rect 363564 218832 363570 218884
rect 368658 218832 368664 218884
rect 368716 218872 368722 218884
rect 378778 218872 378784 218884
rect 368716 218844 378784 218872
rect 368716 218832 368722 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383562 218872 383568 218884
rect 382792 218844 383568 218872
rect 382792 218832 382798 218844
rect 383562 218832 383568 218844
rect 383620 218832 383626 218884
rect 386874 218832 386880 218884
rect 386932 218872 386938 218884
rect 398098 218872 398104 218884
rect 386932 218844 398104 218872
rect 386932 218832 386938 218844
rect 398098 218832 398104 218844
rect 398156 218832 398162 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 544930 218832 544936 218884
rect 544988 218872 544994 218884
rect 555970 218872 555976 218884
rect 544988 218844 555976 218872
rect 544988 218832 544994 218844
rect 555970 218832 555976 218844
rect 556028 218832 556034 218884
rect 569218 218872 569224 218884
rect 556172 218844 569224 218872
rect 291654 218696 291660 218748
rect 291712 218736 291718 218748
rect 324590 218736 324596 218748
rect 291712 218708 324596 218736
rect 291712 218696 291718 218708
rect 324590 218696 324596 218708
rect 324648 218696 324654 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 371786 218736 371792 218748
rect 353812 218708 371792 218736
rect 353812 218696 353818 218708
rect 371786 218696 371792 218708
rect 371844 218696 371850 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 540606 218696 540612 218748
rect 540664 218736 540670 218748
rect 540664 218708 543136 218736
rect 540664 218696 540670 218708
rect 282288 218572 296714 218600
rect 288986 218464 288992 218476
rect 282196 218436 288992 218464
rect 288986 218424 288992 218436
rect 289044 218424 289050 218476
rect 296686 218464 296714 218572
rect 300486 218560 300492 218612
rect 300544 218600 300550 218612
rect 310974 218600 310980 218612
rect 300544 218572 310980 218600
rect 300544 218560 300550 218572
rect 310974 218560 310980 218572
rect 311032 218560 311038 218612
rect 311158 218560 311164 218612
rect 311216 218600 311222 218612
rect 316678 218600 316684 218612
rect 311216 218572 316684 218600
rect 311216 218560 311222 218572
rect 316678 218560 316684 218572
rect 316736 218560 316742 218612
rect 320634 218560 320640 218612
rect 320692 218600 320698 218612
rect 330478 218600 330484 218612
rect 320692 218572 330484 218600
rect 320692 218560 320698 218572
rect 330478 218560 330484 218572
rect 330536 218560 330542 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 537478 218560 537484 218612
rect 537536 218600 537542 218612
rect 543108 218600 543136 218708
rect 547506 218696 547512 218748
rect 547564 218736 547570 218748
rect 556172 218736 556200 218844
rect 569218 218832 569224 218844
rect 569276 218832 569282 218884
rect 569420 218872 569448 218980
rect 569586 218968 569592 219020
rect 569644 219008 569650 219020
rect 601878 219008 601884 219020
rect 569644 218980 601884 219008
rect 569644 218968 569650 218980
rect 601878 218968 601884 218980
rect 601936 218968 601942 219020
rect 676030 218968 676036 219020
rect 676088 219008 676094 219020
rect 676858 219008 676864 219020
rect 676088 218980 676864 219008
rect 676088 218968 676094 218980
rect 676858 218968 676864 218980
rect 676916 218968 676922 219020
rect 572438 218872 572444 218884
rect 569420 218844 572444 218872
rect 572438 218832 572444 218844
rect 572496 218832 572502 218884
rect 572622 218832 572628 218884
rect 572680 218872 572686 218884
rect 575014 218872 575020 218884
rect 572680 218844 575020 218872
rect 572680 218832 572686 218844
rect 575014 218832 575020 218844
rect 575072 218832 575078 218884
rect 582374 218832 582380 218884
rect 582432 218872 582438 218884
rect 597922 218872 597928 218884
rect 582432 218844 597928 218872
rect 582432 218832 582438 218844
rect 597922 218832 597928 218844
rect 597980 218832 597986 218884
rect 547564 218708 556200 218736
rect 547564 218696 547570 218708
rect 558178 218696 558184 218748
rect 558236 218736 558242 218748
rect 571702 218736 571708 218748
rect 558236 218708 571708 218736
rect 558236 218696 558242 218708
rect 571702 218696 571708 218708
rect 571760 218696 571766 218748
rect 571978 218696 571984 218748
rect 572036 218736 572042 218748
rect 575474 218736 575480 218748
rect 572036 218708 575480 218736
rect 572036 218696 572042 218708
rect 575474 218696 575480 218708
rect 575532 218696 575538 218748
rect 552474 218600 552480 218612
rect 537536 218572 543044 218600
rect 543108 218572 552480 218600
rect 537536 218560 537542 218572
rect 304258 218464 304264 218476
rect 296686 218436 304264 218464
rect 304258 218424 304264 218436
rect 304316 218424 304322 218476
rect 512730 218424 512736 218476
rect 512788 218464 512794 218476
rect 540606 218464 540612 218476
rect 512788 218436 540612 218464
rect 512788 218424 512794 218436
rect 540606 218424 540612 218436
rect 540664 218424 540670 218476
rect 543016 218464 543044 218572
rect 552474 218560 552480 218572
rect 552532 218560 552538 218612
rect 555970 218560 555976 218612
rect 556028 218600 556034 218612
rect 598842 218600 598848 218612
rect 556028 218572 598848 218600
rect 556028 218560 556034 218572
rect 598842 218560 598848 218572
rect 598900 218560 598906 218612
rect 568390 218464 568396 218476
rect 543016 218436 568396 218464
rect 568390 218424 568396 218436
rect 568448 218424 568454 218476
rect 568574 218424 568580 218476
rect 568632 218464 568638 218476
rect 569770 218464 569776 218476
rect 568632 218436 569776 218464
rect 568632 218424 568638 218436
rect 569770 218424 569776 218436
rect 569828 218424 569834 218476
rect 571334 218424 571340 218476
rect 571392 218464 571398 218476
rect 572254 218464 572260 218476
rect 571392 218436 572260 218464
rect 571392 218424 571398 218436
rect 572254 218424 572260 218436
rect 572312 218424 572318 218476
rect 572438 218424 572444 218476
rect 572496 218464 572502 218476
rect 604454 218464 604460 218476
rect 572496 218436 604460 218464
rect 572496 218424 572502 218436
rect 604454 218424 604460 218436
rect 604512 218424 604518 218476
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 117958 218288 117964 218340
rect 118016 218328 118022 218340
rect 123478 218328 123484 218340
rect 118016 218300 123484 218328
rect 118016 218288 118022 218300
rect 123478 218288 123484 218300
rect 123536 218288 123542 218340
rect 131850 218288 131856 218340
rect 131908 218328 131914 218340
rect 132402 218328 132408 218340
rect 131908 218300 132408 218328
rect 131908 218288 131914 218300
rect 132402 218288 132408 218300
rect 132460 218288 132466 218340
rect 136818 218288 136824 218340
rect 136876 218328 136882 218340
rect 139486 218328 139492 218340
rect 136876 218300 139492 218328
rect 136876 218288 136882 218300
rect 139486 218288 139492 218300
rect 139544 218288 139550 218340
rect 140130 218288 140136 218340
rect 140188 218328 140194 218340
rect 181162 218328 181168 218340
rect 140188 218300 181168 218328
rect 140188 218288 140194 218300
rect 181162 218288 181168 218300
rect 181220 218288 181226 218340
rect 181530 218288 181536 218340
rect 181588 218328 181594 218340
rect 181990 218328 181996 218340
rect 181588 218300 181996 218328
rect 181588 218288 181594 218300
rect 181990 218288 181996 218300
rect 182048 218288 182054 218340
rect 184014 218288 184020 218340
rect 184072 218328 184078 218340
rect 184934 218328 184940 218340
rect 184072 218300 184940 218328
rect 184072 218288 184078 218300
rect 184934 218288 184940 218300
rect 184992 218288 184998 218340
rect 185670 218288 185676 218340
rect 185728 218328 185734 218340
rect 186130 218328 186136 218340
rect 185728 218300 186136 218328
rect 185728 218288 185734 218300
rect 186130 218288 186136 218300
rect 186188 218288 186194 218340
rect 196434 218288 196440 218340
rect 196492 218328 196498 218340
rect 210142 218328 210148 218340
rect 196492 218300 210148 218328
rect 196492 218288 196498 218300
rect 210142 218288 210148 218300
rect 210200 218288 210206 218340
rect 210326 218288 210332 218340
rect 210384 218328 210390 218340
rect 213178 218328 213184 218340
rect 210384 218300 213184 218328
rect 210384 218288 210390 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 222930 218288 222936 218340
rect 222988 218328 222994 218340
rect 231026 218328 231032 218340
rect 222988 218300 231032 218328
rect 222988 218288 222994 218300
rect 231026 218288 231032 218300
rect 231084 218288 231090 218340
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 270770 218328 270776 218340
rect 232924 218300 270776 218328
rect 232924 218288 232930 218300
rect 270770 218288 270776 218300
rect 270828 218288 270834 218340
rect 340506 218288 340512 218340
rect 340564 218328 340570 218340
rect 352558 218328 352564 218340
rect 340564 218300 352564 218328
rect 340564 218288 340570 218300
rect 352558 218288 352564 218300
rect 352616 218288 352622 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429378 218328 429384 218340
rect 426676 218300 429384 218328
rect 426676 218288 426682 218300
rect 429378 218288 429384 218300
rect 429436 218288 429442 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 503162 218288 503168 218340
rect 503220 218328 503226 218340
rect 614482 218328 614488 218340
rect 503220 218300 614488 218328
rect 503220 218288 503226 218300
rect 614482 218288 614488 218300
rect 614540 218288 614546 218340
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61654 218192 61660 218204
rect 57480 218164 61660 218192
rect 57480 218152 57486 218164
rect 61654 218152 61660 218164
rect 61712 218152 61718 218204
rect 67266 218152 67272 218204
rect 67324 218192 67330 218204
rect 68278 218192 68284 218204
rect 67324 218164 68284 218192
rect 67324 218152 67330 218164
rect 68278 218152 68284 218164
rect 68336 218152 68342 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 123570 218152 123576 218204
rect 123628 218192 123634 218204
rect 165982 218192 165988 218204
rect 123628 218164 165988 218192
rect 123628 218152 123634 218164
rect 165982 218152 165988 218164
rect 166040 218152 166046 218204
rect 171410 218192 171416 218204
rect 166966 218164 171416 218192
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62022 218056 62028 218068
rect 61528 218028 62028 218056
rect 61528 218016 61534 218028
rect 62022 218016 62028 218028
rect 62080 218016 62086 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 66438 218016 66444 218068
rect 66496 218056 66502 218068
rect 67542 218056 67548 218068
rect 66496 218028 67548 218056
rect 66496 218016 66502 218028
rect 67542 218016 67548 218028
rect 67600 218016 67606 218068
rect 68094 218016 68100 218068
rect 68152 218056 68158 218068
rect 68738 218056 68744 218068
rect 68152 218028 68744 218056
rect 68152 218016 68158 218028
rect 68738 218016 68744 218028
rect 68796 218016 68802 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 90450 218016 90456 218068
rect 90508 218056 90514 218068
rect 91738 218056 91744 218068
rect 90508 218028 91744 218056
rect 90508 218016 90514 218028
rect 91738 218016 91744 218028
rect 91796 218016 91802 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93762 218056 93768 218068
rect 92992 218028 93768 218056
rect 92992 218016 92998 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 117774 218016 117780 218068
rect 117832 218056 117838 218068
rect 118694 218056 118700 218068
rect 117832 218028 118700 218056
rect 117832 218016 117838 218028
rect 118694 218016 118700 218028
rect 118752 218016 118758 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 126054 218016 126060 218068
rect 126112 218056 126118 218068
rect 126698 218056 126704 218068
rect 126112 218028 126704 218056
rect 126112 218016 126118 218028
rect 126698 218016 126704 218028
rect 126756 218016 126762 218068
rect 127710 218016 127716 218068
rect 127768 218056 127774 218068
rect 128262 218056 128268 218068
rect 127768 218028 128268 218056
rect 127768 218016 127774 218028
rect 128262 218016 128268 218028
rect 128320 218016 128326 218068
rect 128538 218016 128544 218068
rect 128596 218056 128602 218068
rect 129366 218056 129372 218068
rect 128596 218028 129372 218056
rect 128596 218016 128602 218028
rect 129366 218016 129372 218028
rect 129424 218016 129430 218068
rect 130194 218016 130200 218068
rect 130252 218056 130258 218068
rect 132494 218056 132500 218068
rect 130252 218028 132500 218056
rect 130252 218016 130258 218028
rect 132494 218016 132500 218028
rect 132552 218016 132558 218068
rect 132678 218016 132684 218068
rect 132736 218056 132742 218068
rect 133506 218056 133512 218068
rect 132736 218028 133512 218056
rect 132736 218016 132742 218028
rect 133506 218016 133512 218028
rect 133564 218016 133570 218068
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 136542 218056 136548 218068
rect 136048 218028 136548 218056
rect 136048 218016 136054 218028
rect 136542 218016 136548 218028
rect 136600 218016 136606 218068
rect 138474 218016 138480 218068
rect 138532 218056 138538 218068
rect 139118 218056 139124 218068
rect 138532 218028 139124 218056
rect 138532 218016 138538 218028
rect 139118 218016 139124 218028
rect 139176 218016 139182 218068
rect 139486 218016 139492 218068
rect 139544 218056 139550 218068
rect 166966 218056 166994 218164
rect 171410 218152 171416 218164
rect 171468 218152 171474 218204
rect 173250 218152 173256 218204
rect 173308 218192 173314 218204
rect 173308 218164 179552 218192
rect 173308 218152 173314 218164
rect 139544 218028 166994 218056
rect 139544 218016 139550 218028
rect 170766 218016 170772 218068
rect 170824 218056 170830 218068
rect 176470 218056 176476 218068
rect 170824 218028 176476 218056
rect 170824 218016 170830 218028
rect 176470 218016 176476 218028
rect 176528 218016 176534 218068
rect 178218 218016 178224 218068
rect 178276 218056 178282 218068
rect 179322 218056 179328 218068
rect 178276 218028 179328 218056
rect 178276 218016 178282 218028
rect 179322 218016 179328 218028
rect 179380 218016 179386 218068
rect 179524 218056 179552 218164
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 225598 218192 225604 218204
rect 179932 218164 225604 218192
rect 179932 218152 179938 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 241974 218152 241980 218204
rect 242032 218192 242038 218204
rect 242894 218192 242900 218204
rect 242032 218164 242900 218192
rect 242032 218152 242038 218164
rect 242894 218152 242900 218164
rect 242952 218152 242958 218204
rect 243538 218152 243544 218204
rect 243596 218192 243602 218204
rect 249058 218192 249064 218204
rect 243596 218164 249064 218192
rect 243596 218152 243602 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 297450 218152 297456 218204
rect 297508 218192 297514 218204
rect 302878 218192 302884 218204
rect 297508 218164 302884 218192
rect 297508 218152 297514 218164
rect 302878 218152 302884 218164
rect 302936 218152 302942 218204
rect 333054 218152 333060 218204
rect 333112 218192 333118 218204
rect 333882 218192 333888 218204
rect 333112 218164 333888 218192
rect 333112 218152 333118 218164
rect 333882 218152 333888 218164
rect 333940 218152 333946 218204
rect 335538 218152 335544 218204
rect 335596 218192 335602 218204
rect 338666 218192 338672 218204
rect 335596 218164 338672 218192
rect 335596 218152 335602 218164
rect 338666 218152 338672 218164
rect 338724 218152 338730 218204
rect 358722 218152 358728 218204
rect 358780 218192 358786 218204
rect 359458 218192 359464 218204
rect 358780 218164 359464 218192
rect 358780 218152 358786 218164
rect 359458 218152 359464 218164
rect 359516 218152 359522 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 400950 218152 400956 218204
rect 401008 218192 401014 218204
rect 402238 218192 402244 218204
rect 401008 218164 402244 218192
rect 401008 218152 401014 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 428458 218192 428464 218204
rect 425848 218164 428464 218192
rect 425848 218152 425854 218164
rect 428458 218152 428464 218164
rect 428516 218152 428522 218204
rect 429102 218152 429108 218204
rect 429160 218192 429166 218204
rect 430574 218192 430580 218204
rect 429160 218164 430580 218192
rect 429160 218152 429166 218164
rect 430574 218152 430580 218164
rect 430632 218152 430638 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 434714 218192 434720 218204
rect 433300 218164 434720 218192
rect 433300 218152 433306 218164
rect 434714 218152 434720 218164
rect 434772 218152 434778 218204
rect 435726 218152 435732 218204
rect 435784 218192 435790 218204
rect 436646 218192 436652 218204
rect 435784 218164 436652 218192
rect 435784 218152 435790 218164
rect 436646 218152 436652 218164
rect 436704 218152 436710 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 500034 218152 500040 218204
rect 500092 218192 500098 218204
rect 609882 218192 609888 218204
rect 500092 218164 609888 218192
rect 500092 218152 500098 218164
rect 609882 218152 609888 218164
rect 609940 218152 609946 218204
rect 210326 218056 210332 218068
rect 179524 218028 210332 218056
rect 210326 218016 210332 218028
rect 210384 218016 210390 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216122 218056 216128 218068
rect 215536 218028 216128 218056
rect 215536 218016 215542 218028
rect 216122 218016 216128 218028
rect 216180 218016 216186 218068
rect 218790 218016 218796 218068
rect 218848 218056 218854 218068
rect 219342 218056 219348 218068
rect 218848 218028 219348 218056
rect 218848 218016 218854 218028
rect 219342 218016 219348 218028
rect 219400 218016 219406 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 227070 218016 227076 218068
rect 227128 218056 227134 218068
rect 227530 218056 227536 218068
rect 227128 218028 227536 218056
rect 227128 218016 227134 218028
rect 227530 218016 227536 218028
rect 227588 218016 227594 218068
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 230474 218056 230480 218068
rect 229612 218028 230480 218056
rect 229612 218016 229618 218028
rect 230474 218016 230480 218028
rect 230532 218016 230538 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 245286 218056 245292 218068
rect 244516 218028 245292 218056
rect 244516 218016 244522 218028
rect 245286 218016 245292 218028
rect 245344 218016 245350 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248322 218056 248328 218068
rect 247828 218028 248328 218056
rect 247828 218016 247834 218028
rect 248322 218016 248328 218028
rect 248380 218016 248386 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249242 218056 249248 218068
rect 248656 218028 249248 218056
rect 248656 218016 248662 218028
rect 249242 218016 249248 218028
rect 249300 218016 249306 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257890 218056 257896 218068
rect 256936 218028 257896 218056
rect 256936 218016 256942 218028
rect 257890 218016 257896 218028
rect 257948 218016 257954 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259362 218056 259368 218068
rect 258592 218028 259368 218056
rect 258592 218016 258598 218028
rect 259362 218016 259368 218028
rect 259420 218016 259426 218068
rect 260190 218016 260196 218068
rect 260248 218056 260254 218068
rect 260742 218056 260748 218068
rect 260248 218028 260748 218056
rect 260248 218016 260254 218028
rect 260742 218016 260748 218028
rect 260800 218016 260806 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270218 218056 270224 218068
rect 269356 218028 270224 218056
rect 269356 218016 269362 218028
rect 270218 218016 270224 218028
rect 270276 218016 270282 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282730 218056 282736 218068
rect 281776 218028 282736 218056
rect 281776 218016 281782 218028
rect 282730 218016 282736 218028
rect 282788 218016 282794 218068
rect 283374 218016 283380 218068
rect 283432 218056 283438 218068
rect 284294 218056 284300 218068
rect 283432 218028 284300 218056
rect 283432 218016 283438 218028
rect 284294 218016 284300 218028
rect 284352 218016 284358 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288066 218056 288072 218068
rect 287572 218028 288072 218056
rect 287572 218016 287578 218028
rect 288066 218016 288072 218028
rect 288124 218016 288130 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289722 218056 289728 218068
rect 289228 218028 289728 218056
rect 289228 218016 289234 218028
rect 289722 218016 289728 218028
rect 289780 218016 289786 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299382 218056 299388 218068
rect 298336 218028 299388 218056
rect 298336 218016 298342 218028
rect 299382 218016 299388 218028
rect 299440 218016 299446 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310330 218056 310336 218068
rect 309928 218028 310336 218056
rect 309928 218016 309934 218028
rect 310330 218016 310336 218028
rect 310388 218016 310394 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315482 218056 315488 218068
rect 314896 218028 315488 218056
rect 314896 218016 314902 218028
rect 315482 218016 315488 218028
rect 315540 218016 315546 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 320082 218056 320088 218068
rect 319036 218028 320088 218056
rect 319036 218016 319042 218028
rect 320082 218016 320088 218028
rect 320140 218016 320146 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 323946 218056 323952 218068
rect 323176 218028 323952 218056
rect 323176 218016 323182 218028
rect 323946 218016 323952 218028
rect 324004 218016 324010 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325510 218056 325516 218068
rect 324832 218028 325516 218056
rect 324832 218016 324838 218028
rect 325510 218016 325516 218028
rect 325568 218016 325574 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 332226 218016 332232 218068
rect 332284 218056 332290 218068
rect 333422 218056 333428 218068
rect 332284 218028 333428 218056
rect 332284 218016 332290 218028
rect 333422 218016 333428 218028
rect 333480 218016 333486 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 337194 218016 337200 218068
rect 337252 218056 337258 218068
rect 337746 218056 337752 218068
rect 337252 218028 337752 218056
rect 337252 218016 337258 218028
rect 337746 218016 337752 218028
rect 337804 218016 337810 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347222 218056 347228 218068
rect 345532 218028 347228 218056
rect 345532 218016 345538 218028
rect 347222 218016 347228 218028
rect 347280 218016 347286 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 352098 218016 352104 218068
rect 352156 218056 352162 218068
rect 353294 218056 353300 218068
rect 352156 218028 353300 218056
rect 352156 218016 352162 218028
rect 353294 218016 353300 218028
rect 353352 218016 353358 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357250 218056 357256 218068
rect 356296 218028 357256 218056
rect 356296 218016 356302 218028
rect 357250 218016 357256 218028
rect 357308 218016 357314 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 358538 218056 358544 218068
rect 357952 218028 358544 218056
rect 357952 218016 357958 218028
rect 358538 218016 358544 218028
rect 358596 218016 358602 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373534 218056 373540 218068
rect 372856 218028 373540 218056
rect 372856 218016 372862 218028
rect 373534 218016 373540 218028
rect 373592 218016 373598 218068
rect 374454 218016 374460 218068
rect 374512 218056 374518 218068
rect 375006 218056 375012 218068
rect 374512 218028 375012 218056
rect 374512 218016 374518 218028
rect 375006 218016 375012 218028
rect 375064 218016 375070 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386046 218056 386052 218068
rect 385276 218028 386052 218056
rect 385276 218016 385282 218028
rect 386046 218016 386052 218028
rect 386104 218016 386110 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390462 218056 390468 218068
rect 389416 218028 390468 218056
rect 389416 218016 389422 218028
rect 390462 218016 390468 218028
rect 390520 218016 390526 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 401318 218056 401324 218068
rect 397696 218028 401324 218056
rect 397696 218016 397702 218028
rect 401318 218016 401324 218028
rect 401376 218016 401382 218068
rect 401778 218016 401784 218068
rect 401836 218056 401842 218068
rect 402790 218056 402796 218068
rect 401836 218028 402796 218056
rect 401836 218016 401842 218028
rect 402790 218016 402796 218028
rect 402848 218016 402854 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 428274 218016 428280 218068
rect 428332 218056 428338 218068
rect 429562 218056 429568 218068
rect 428332 218028 429568 218056
rect 428332 218016 428338 218028
rect 429562 218016 429568 218028
rect 429620 218016 429626 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434898 218016 434904 218068
rect 434956 218056 434962 218068
rect 436278 218056 436284 218068
rect 434956 218028 436284 218056
rect 434956 218016 434962 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437750 218056 437756 218068
rect 436612 218028 437756 218056
rect 436612 218016 436618 218028
rect 437750 218016 437756 218028
rect 437808 218016 437814 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 471422 218016 471428 218068
rect 471480 218056 471486 218068
rect 472894 218056 472900 218068
rect 471480 218028 472900 218056
rect 471480 218016 471486 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 492030 218016 492036 218068
rect 492088 218056 492094 218068
rect 505646 218056 505652 218068
rect 492088 218028 505652 218056
rect 492088 218016 492094 218028
rect 505646 218016 505652 218028
rect 505704 218016 505710 218068
rect 507670 218016 507676 218068
rect 507728 218056 507734 218068
rect 615678 218056 615684 218068
rect 507728 218028 615684 218056
rect 507728 218016 507734 218028
rect 615678 218016 615684 218028
rect 615736 218016 615742 218068
rect 646590 218016 646596 218068
rect 646648 218056 646654 218068
rect 653398 218056 653404 218068
rect 646648 218028 653404 218056
rect 646648 218016 646654 218028
rect 653398 218016 653404 218028
rect 653456 218016 653462 218068
rect 131022 217812 131028 217864
rect 131080 217852 131086 217864
rect 197722 217852 197728 217864
rect 131080 217824 197728 217852
rect 131080 217812 131086 217824
rect 197722 217812 197728 217824
rect 197780 217812 197786 217864
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 535454 217812 535460 217864
rect 535512 217852 535518 217864
rect 536650 217852 536656 217864
rect 535512 217824 536656 217852
rect 535512 217812 535518 217824
rect 536650 217812 536656 217824
rect 536708 217812 536714 217864
rect 536834 217812 536840 217864
rect 536892 217852 536898 217864
rect 536892 217824 603120 217852
rect 536892 217812 536898 217824
rect 116946 217676 116952 217728
rect 117004 217716 117010 217728
rect 189258 217716 189264 217728
rect 117004 217688 189264 217716
rect 117004 217676 117010 217688
rect 189258 217676 189264 217688
rect 189316 217676 189322 217728
rect 525978 217676 525984 217728
rect 526036 217716 526042 217728
rect 526530 217716 526536 217728
rect 526036 217688 526536 217716
rect 526036 217676 526042 217688
rect 526530 217676 526536 217688
rect 526588 217676 526594 217728
rect 533430 217676 533436 217728
rect 533488 217716 533494 217728
rect 602890 217716 602896 217728
rect 533488 217688 602896 217716
rect 533488 217676 533494 217688
rect 602890 217676 602896 217688
rect 602948 217676 602954 217728
rect 603092 217716 603120 217824
rect 603258 217812 603264 217864
rect 603316 217852 603322 217864
rect 613378 217852 613384 217864
rect 603316 217824 613384 217852
rect 603316 217812 603322 217824
rect 613378 217812 613384 217824
rect 613436 217812 613442 217864
rect 603442 217716 603448 217728
rect 603092 217688 603448 217716
rect 603442 217676 603448 217688
rect 603500 217676 603506 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 616874 217716 616880 217728
rect 604512 217688 616880 217716
rect 604512 217676 604518 217688
rect 616874 217676 616880 217688
rect 616932 217676 616938 217728
rect 103698 217540 103704 217592
rect 103756 217580 103762 217592
rect 178402 217580 178408 217592
rect 103756 217552 178408 217580
rect 103756 217540 103762 217552
rect 178402 217540 178408 217552
rect 178460 217540 178466 217592
rect 530578 217540 530584 217592
rect 530636 217580 530642 217592
rect 530946 217580 530952 217592
rect 530636 217552 530952 217580
rect 530636 217540 530642 217552
rect 530946 217540 530952 217552
rect 531004 217580 531010 217592
rect 536834 217580 536840 217592
rect 531004 217552 536840 217580
rect 531004 217540 531010 217552
rect 536834 217540 536840 217552
rect 536892 217540 536898 217592
rect 538214 217540 538220 217592
rect 538272 217580 538278 217592
rect 539134 217580 539140 217592
rect 538272 217552 539140 217580
rect 538272 217540 538278 217552
rect 539134 217540 539140 217552
rect 539192 217540 539198 217592
rect 545758 217540 545764 217592
rect 545816 217580 545822 217592
rect 606754 217580 606760 217592
rect 545816 217552 606760 217580
rect 545816 217540 545822 217552
rect 606754 217540 606760 217552
rect 606812 217540 606818 217592
rect 675846 217540 675852 217592
rect 675904 217580 675910 217592
rect 676582 217580 676588 217592
rect 675904 217552 676588 217580
rect 675904 217540 675910 217552
rect 676582 217540 676588 217552
rect 676640 217540 676646 217592
rect 93762 217404 93768 217456
rect 93820 217444 93826 217456
rect 171226 217444 171232 217456
rect 93820 217416 171232 217444
rect 93820 217404 93826 217416
rect 171226 217404 171232 217416
rect 171284 217404 171290 217456
rect 526530 217404 526536 217456
rect 526588 217444 526594 217456
rect 526588 217416 601602 217444
rect 526588 217404 526594 217416
rect 170306 217308 170312 217320
rect 93826 217280 170312 217308
rect 92060 217200 92066 217252
rect 92118 217240 92124 217252
rect 93826 217240 93854 217280
rect 170306 217268 170312 217280
rect 170364 217268 170370 217320
rect 535822 217268 535828 217320
rect 535880 217308 535886 217320
rect 598658 217308 598664 217320
rect 535880 217280 598664 217308
rect 535880 217268 535886 217280
rect 598658 217268 598664 217280
rect 598716 217268 598722 217320
rect 598842 217268 598848 217320
rect 598900 217308 598906 217320
rect 601326 217308 601332 217320
rect 598900 217280 601332 217308
rect 598900 217268 598906 217280
rect 601326 217268 601332 217280
rect 601384 217268 601390 217320
rect 601574 217308 601602 217416
rect 601878 217404 601884 217456
rect 601936 217444 601942 217456
rect 628282 217444 628288 217456
rect 601936 217416 628288 217444
rect 601936 217404 601942 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 602338 217308 602344 217320
rect 601574 217280 602344 217308
rect 602338 217268 602344 217280
rect 602396 217268 602402 217320
rect 602890 217268 602896 217320
rect 602948 217308 602954 217320
rect 603994 217308 604000 217320
rect 602948 217280 604000 217308
rect 602948 217268 602954 217280
rect 603994 217268 604000 217280
rect 604052 217268 604058 217320
rect 642174 217268 642180 217320
rect 642232 217308 642238 217320
rect 658918 217308 658924 217320
rect 642232 217280 658924 217308
rect 642232 217268 642238 217280
rect 658918 217268 658924 217280
rect 658976 217268 658982 217320
rect 92118 217212 93854 217240
rect 92118 217200 92124 217212
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 448606 217200 448612 217252
rect 448664 217240 448670 217252
rect 449756 217240 449762 217252
rect 448664 217212 449762 217240
rect 448664 217200 448670 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 489914 217200 489920 217252
rect 489972 217240 489978 217252
rect 491156 217240 491162 217252
rect 489972 217212 491162 217240
rect 489972 217200 489978 217212
rect 491156 217200 491162 217212
rect 491214 217200 491220 217252
rect 498286 217200 498292 217252
rect 498344 217240 498350 217252
rect 499436 217240 499442 217252
rect 498344 217212 499442 217240
rect 498344 217200 498350 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 502978 217200 502984 217252
rect 503036 217240 503042 217252
rect 503576 217240 503582 217252
rect 503036 217212 503582 217240
rect 503036 217200 503042 217212
rect 503576 217200 503582 217212
rect 503634 217200 503640 217252
rect 511028 217132 511034 217184
rect 511086 217172 511092 217184
rect 561858 217172 561864 217184
rect 511086 217144 561864 217172
rect 511086 217132 511092 217144
rect 561858 217132 561864 217144
rect 561916 217132 561922 217184
rect 562870 217132 562876 217184
rect 562928 217132 562934 217184
rect 565078 217132 565084 217184
rect 565136 217172 565142 217184
rect 599026 217172 599032 217184
rect 565136 217144 599032 217172
rect 565136 217132 565142 217144
rect 599026 217132 599032 217144
rect 599084 217132 599090 217184
rect 600774 217132 600780 217184
rect 600832 217172 600838 217184
rect 604546 217172 604552 217184
rect 600832 217144 604552 217172
rect 600832 217132 600838 217144
rect 604546 217132 604552 217144
rect 604604 217132 604610 217184
rect 503576 217064 503582 217116
rect 503634 217104 503640 217116
rect 562502 217104 562508 217116
rect 503634 217076 505094 217104
rect 503634 217064 503640 217076
rect 505066 217036 505094 217076
rect 562060 217076 562508 217104
rect 562060 217036 562088 217076
rect 562502 217064 562508 217076
rect 562560 217064 562566 217116
rect 505066 217008 562088 217036
rect 562888 217036 562916 217132
rect 608962 217036 608968 217048
rect 562888 217008 608968 217036
rect 608962 216996 608968 217008
rect 609020 216996 609026 217048
rect 609882 216996 609888 217048
rect 609940 217036 609946 217048
rect 614114 217036 614120 217048
rect 609940 217008 614120 217036
rect 609940 216996 609946 217008
rect 614114 216996 614120 217008
rect 614172 216996 614178 217048
rect 574094 216860 574100 216912
rect 574152 216900 574158 216912
rect 597554 216900 597560 216912
rect 574152 216872 597560 216900
rect 574152 216860 574158 216872
rect 597554 216860 597560 216872
rect 597612 216860 597618 216912
rect 598658 216860 598664 216912
rect 598716 216900 598722 216912
rect 600774 216900 600780 216912
rect 598716 216872 600780 216900
rect 598716 216860 598722 216872
rect 600774 216860 600780 216872
rect 600832 216860 600838 216912
rect 612274 216900 612280 216912
rect 600976 216872 612280 216900
rect 594794 216724 594800 216776
rect 594852 216764 594858 216776
rect 600976 216764 601004 216872
rect 612274 216860 612280 216872
rect 612332 216860 612338 216912
rect 594852 216736 601004 216764
rect 594852 216724 594858 216736
rect 601326 216724 601332 216776
rect 601384 216764 601390 216776
rect 623866 216764 623872 216776
rect 601384 216736 623872 216764
rect 601384 216724 601390 216736
rect 623866 216724 623872 216736
rect 623924 216724 623930 216776
rect 648246 216588 648252 216640
rect 648304 216628 648310 216640
rect 656158 216628 656164 216640
rect 648304 216600 656164 216628
rect 648304 216588 648310 216600
rect 656158 216588 656164 216600
rect 656216 216588 656222 216640
rect 675938 215500 675944 215552
rect 675996 215540 676002 215552
rect 677042 215540 677048 215552
rect 675996 215512 677048 215540
rect 675996 215500 676002 215512
rect 677042 215500 677048 215512
rect 677100 215500 677106 215552
rect 663150 215296 663156 215348
rect 663208 215336 663214 215348
rect 663702 215336 663708 215348
rect 663208 215308 663708 215336
rect 663208 215296 663214 215308
rect 663702 215296 663708 215308
rect 663760 215296 663766 215348
rect 575474 214820 575480 214872
rect 575532 214860 575538 214872
rect 622302 214860 622308 214872
rect 575532 214832 622308 214860
rect 575532 214820 575538 214832
rect 622302 214820 622308 214832
rect 622360 214820 622366 214872
rect 575014 214684 575020 214736
rect 575072 214724 575078 214736
rect 616690 214724 616696 214736
rect 575072 214696 616696 214724
rect 575072 214684 575078 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 617058 214684 617064 214736
rect 617116 214724 617122 214736
rect 617794 214724 617800 214736
rect 617116 214696 617800 214724
rect 617116 214684 617122 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 619818 214684 619824 214736
rect 619876 214724 619882 214736
rect 620554 214724 620560 214736
rect 619876 214696 620560 214724
rect 619876 214684 619882 214696
rect 620554 214684 620560 214696
rect 620612 214684 620618 214736
rect 621014 214684 621020 214736
rect 621072 214724 621078 214736
rect 621658 214724 621664 214736
rect 621072 214696 621664 214724
rect 621072 214684 621078 214696
rect 621658 214684 621664 214696
rect 621716 214684 621722 214736
rect 622486 214684 622492 214736
rect 622544 214724 622550 214736
rect 623314 214724 623320 214736
rect 622544 214696 623320 214724
rect 622544 214684 622550 214696
rect 623314 214684 623320 214696
rect 623372 214684 623378 214736
rect 625246 214684 625252 214736
rect 625304 214724 625310 214736
rect 626074 214724 626080 214736
rect 625304 214696 626080 214724
rect 625304 214684 625310 214696
rect 626074 214684 626080 214696
rect 626132 214684 626138 214736
rect 630030 214684 630036 214736
rect 630088 214724 630094 214736
rect 632882 214724 632888 214736
rect 630088 214696 632888 214724
rect 630088 214684 630094 214696
rect 632882 214684 632888 214696
rect 632940 214684 632946 214736
rect 644566 214684 644572 214736
rect 644624 214724 644630 214736
rect 654778 214724 654784 214736
rect 644624 214696 654784 214724
rect 644624 214684 644630 214696
rect 654778 214684 654784 214696
rect 654836 214684 654842 214736
rect 574646 214548 574652 214600
rect 574704 214588 574710 214600
rect 625614 214588 625620 214600
rect 574704 214560 625620 214588
rect 574704 214548 574710 214560
rect 625614 214548 625620 214560
rect 625672 214548 625678 214600
rect 654870 214548 654876 214600
rect 654928 214588 654934 214600
rect 664438 214588 664444 214600
rect 654928 214560 664444 214588
rect 654928 214548 654934 214560
rect 664438 214548 664444 214560
rect 664496 214548 664502 214600
rect 605926 214412 605932 214464
rect 605984 214452 605990 214464
rect 606294 214452 606300 214464
rect 605984 214424 606300 214452
rect 605984 214412 605990 214424
rect 606294 214412 606300 214424
rect 606352 214412 606358 214464
rect 607306 214412 607312 214464
rect 607364 214452 607370 214464
rect 607858 214452 607864 214464
rect 607364 214424 607864 214452
rect 607364 214412 607370 214424
rect 607858 214412 607864 214424
rect 607916 214412 607922 214464
rect 616690 214412 616696 214464
rect 616748 214452 616754 214464
rect 624418 214452 624424 214464
rect 616748 214424 624424 214452
rect 616748 214412 616754 214424
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 626350 214412 626356 214464
rect 626408 214452 626414 214464
rect 628834 214452 628840 214464
rect 626408 214424 628840 214452
rect 626408 214412 626414 214424
rect 628834 214412 628840 214424
rect 628892 214412 628898 214464
rect 664806 214344 664812 214396
rect 664864 214384 664870 214396
rect 665818 214384 665824 214396
rect 664864 214356 665824 214384
rect 664864 214344 664870 214356
rect 665818 214344 665824 214356
rect 665876 214344 665882 214396
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 41690 213976 41696 213988
rect 35860 213948 41696 213976
rect 35860 213936 35866 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 627454 213936 627460 213988
rect 627512 213976 627518 213988
rect 629386 213976 629392 213988
rect 627512 213948 629392 213976
rect 627512 213936 627518 213948
rect 629386 213936 629392 213948
rect 629444 213936 629450 213988
rect 649902 213868 649908 213920
rect 649960 213908 649966 213920
rect 652018 213908 652024 213920
rect 649960 213880 652024 213908
rect 649960 213868 649966 213880
rect 652018 213868 652024 213880
rect 652076 213868 652082 213920
rect 659562 213664 659568 213716
rect 659620 213704 659626 213716
rect 665542 213704 665548 213716
rect 659620 213676 665548 213704
rect 659620 213664 659626 213676
rect 665542 213664 665548 213676
rect 665600 213664 665606 213716
rect 647142 213596 647148 213648
rect 647200 213636 647206 213648
rect 649718 213636 649724 213648
rect 647200 213608 649724 213636
rect 647200 213596 647206 213608
rect 649718 213596 649724 213608
rect 649776 213596 649782 213648
rect 574094 213460 574100 213512
rect 574152 213500 574158 213512
rect 594794 213500 594800 213512
rect 574152 213472 594800 213500
rect 574152 213460 574158 213472
rect 594794 213460 594800 213472
rect 594852 213460 594858 213512
rect 574370 213324 574376 213376
rect 574428 213364 574434 213376
rect 612826 213364 612832 213376
rect 574428 213336 612832 213364
rect 574428 213324 574434 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 651098 213324 651104 213376
rect 651156 213364 651162 213376
rect 657538 213364 657544 213376
rect 651156 213336 657544 213364
rect 651156 213324 651162 213336
rect 657538 213324 657544 213336
rect 657596 213324 657602 213376
rect 574830 213188 574836 213240
rect 574888 213228 574894 213240
rect 616138 213228 616144 213240
rect 574888 213200 616144 213228
rect 574888 213188 574894 213200
rect 616138 213188 616144 213200
rect 616196 213188 616202 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 650638 213228 650644 213240
rect 643888 213200 650644 213228
rect 643888 213188 643894 213200
rect 650638 213188 650644 213200
rect 650696 213188 650702 213240
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 658182 212712 658188 212764
rect 658240 212752 658246 212764
rect 659102 212752 659108 212764
rect 658240 212724 659108 212752
rect 658240 212712 658246 212724
rect 659102 212712 659108 212724
rect 659160 212712 659166 212764
rect 664254 212712 664260 212764
rect 664312 212752 664318 212764
rect 665082 212752 665088 212764
rect 664312 212724 665088 212752
rect 664312 212712 664318 212724
rect 665082 212712 665088 212724
rect 665140 212712 665146 212764
rect 632698 212508 632704 212560
rect 632756 212548 632762 212560
rect 634354 212548 634360 212560
rect 632756 212520 634360 212548
rect 632756 212508 632762 212520
rect 634354 212508 634360 212520
rect 634412 212508 634418 212560
rect 630674 212372 630680 212424
rect 630732 212412 630738 212424
rect 631594 212412 631600 212424
rect 630732 212384 631600 212412
rect 630732 212372 630738 212384
rect 631594 212372 631600 212384
rect 631652 212372 631658 212424
rect 35802 211556 35808 211608
rect 35860 211596 35866 211608
rect 39574 211596 39580 211608
rect 35860 211568 39580 211596
rect 35860 211556 35866 211568
rect 39574 211556 39580 211568
rect 39632 211556 39638 211608
rect 35618 211284 35624 211336
rect 35676 211324 35682 211336
rect 41690 211324 41696 211336
rect 35676 211296 41696 211324
rect 35676 211284 35682 211296
rect 41690 211284 41696 211296
rect 41748 211284 41754 211336
rect 35434 211148 35440 211200
rect 35492 211188 35498 211200
rect 41322 211188 41328 211200
rect 35492 211160 41328 211188
rect 35492 211148 35498 211160
rect 41322 211148 41328 211160
rect 41380 211148 41386 211200
rect 578326 211148 578332 211200
rect 578384 211188 578390 211200
rect 580902 211188 580908 211200
rect 578384 211160 580908 211188
rect 578384 211148 578390 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 680354 211148 680360 211200
rect 680412 211188 680418 211200
rect 683114 211188 683120 211200
rect 680412 211160 683120 211188
rect 680412 211148 680418 211160
rect 683114 211148 683120 211160
rect 683172 211148 683178 211200
rect 600314 211012 600320 211064
rect 600372 211052 600378 211064
rect 600682 211052 600688 211064
rect 600372 211024 600688 211052
rect 600372 211012 600378 211024
rect 600682 211012 600688 211024
rect 600740 211012 600746 211064
rect 633434 211012 633440 211064
rect 633492 211052 633498 211064
rect 633802 211052 633808 211064
rect 633492 211024 633808 211052
rect 633492 211012 633498 211024
rect 633802 211012 633808 211024
rect 633860 211012 633866 211064
rect 635550 210128 635556 210180
rect 635608 210168 635614 210180
rect 636562 210168 636568 210180
rect 635608 210140 636568 210168
rect 635608 210128 635614 210140
rect 636562 210128 636568 210140
rect 636620 210128 636626 210180
rect 35802 209788 35808 209840
rect 35860 209828 35866 209840
rect 40310 209828 40316 209840
rect 35860 209800 40316 209828
rect 35860 209788 35866 209800
rect 40310 209788 40316 209800
rect 40368 209788 40374 209840
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 35802 208496 35808 208548
rect 35860 208536 35866 208548
rect 40678 208536 40684 208548
rect 35860 208508 40684 208536
rect 35860 208496 35866 208508
rect 40678 208496 40684 208508
rect 40736 208496 40742 208548
rect 35618 208360 35624 208412
rect 35676 208400 35682 208412
rect 40034 208400 40040 208412
rect 35676 208372 40040 208400
rect 35676 208360 35682 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207136 35808 207188
rect 35860 207176 35866 207188
rect 41138 207176 41144 207188
rect 35860 207148 41144 207176
rect 35860 207136 35866 207148
rect 41138 207136 41144 207148
rect 41196 207136 41202 207188
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 35802 205776 35808 205828
rect 35860 205816 35866 205828
rect 40678 205816 40684 205828
rect 35860 205788 40684 205816
rect 35860 205776 35866 205788
rect 40678 205776 40684 205788
rect 40736 205776 40742 205828
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204620 35808 204672
rect 35860 204660 35866 204672
rect 35860 204620 35894 204660
rect 35866 204592 35894 204620
rect 35866 204564 41414 204592
rect 41386 204524 41414 204564
rect 41690 204524 41696 204536
rect 41386 204496 41696 204524
rect 41690 204484 41696 204496
rect 41748 204484 41754 204536
rect 35802 204280 35808 204332
rect 35860 204320 35866 204332
rect 41690 204320 41696 204332
rect 35860 204292 41696 204320
rect 35860 204280 35866 204292
rect 41690 204280 41696 204292
rect 41748 204280 41754 204332
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 672902 192992 672908 193044
rect 672960 193032 672966 193044
rect 673362 193032 673368 193044
rect 672960 193004 673368 193032
rect 672960 192992 672966 193004
rect 673362 192992 673368 193004
rect 673420 192992 673426 193044
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 668210 165180 668216 165232
rect 668268 165220 668274 165232
rect 669590 165220 669596 165232
rect 668268 165192 669596 165220
rect 668268 165180 668274 165192
rect 669590 165180 669596 165192
rect 669648 165180 669654 165232
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 668210 163276 668216 163328
rect 668268 163316 668274 163328
rect 669774 163316 669780 163328
rect 668268 163288 669780 163316
rect 668268 163276 668274 163288
rect 669774 163276 669780 163288
rect 669832 163276 669838 163328
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 675846 162800 675852 162852
rect 675904 162840 675910 162852
rect 678238 162840 678244 162852
rect 675904 162812 678244 162840
rect 675904 162800 675910 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 668210 160012 668216 160064
rect 668268 160052 668274 160064
rect 670326 160052 670332 160064
rect 668268 160024 670332 160052
rect 668268 160012 668274 160024
rect 670326 160012 670332 160024
rect 670384 160012 670390 160064
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 668302 155116 668308 155168
rect 668360 155156 668366 155168
rect 670786 155156 670792 155168
rect 668360 155128 670792 155156
rect 668360 155116 668366 155128
rect 670786 155116 670792 155128
rect 670844 155116 670850 155168
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 668210 148724 668216 148776
rect 668268 148764 668274 148776
rect 670142 148764 670148 148776
rect 668268 148736 670148 148764
rect 668268 148724 668274 148736
rect 670142 148724 670148 148736
rect 670200 148724 670206 148776
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585778 143556 585784 143608
rect 585836 143596 585842 143608
rect 589458 143596 589464 143608
rect 585836 143568 589464 143596
rect 585836 143556 585842 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 668210 136212 668216 136264
rect 668268 136252 668274 136264
rect 669958 136252 669964 136264
rect 668268 136224 669964 136252
rect 668268 136212 668274 136224
rect 669958 136212 669964 136224
rect 670016 136212 670022 136264
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 585962 132472 585968 132524
rect 586020 132512 586026 132524
rect 589458 132512 589464 132524
rect 586020 132484 589464 132512
rect 586020 132472 586026 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585778 131152 585784 131164
rect 578936 131124 585784 131152
rect 578936 131112 578942 131124
rect 585778 131112 585784 131124
rect 585836 131112 585842 131164
rect 583386 129140 583392 129192
rect 583444 129180 583450 129192
rect 590378 129180 590384 129192
rect 583444 129152 590384 129180
rect 583444 129140 583450 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 668578 129140 668584 129192
rect 668636 129180 668642 129192
rect 670786 129180 670792 129192
rect 668636 129152 670792 129180
rect 668636 129140 668642 129152
rect 670786 129140 670792 129152
rect 670844 129140 670850 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 587802 126964 587808 127016
rect 587860 127004 587866 127016
rect 589458 127004 589464 127016
rect 587860 126976 589464 127004
rect 587860 126964 587866 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 579062 124856 579068 124908
rect 579120 124896 579126 124908
rect 587802 124896 587808 124908
rect 579120 124868 587808 124896
rect 579120 124856 579126 124868
rect 587802 124856 587808 124868
rect 587860 124856 587866 124908
rect 578694 124108 578700 124160
rect 578752 124148 578758 124160
rect 583018 124148 583024 124160
rect 578752 124120 583024 124148
rect 578752 124108 578758 124120
rect 583018 124108 583024 124120
rect 583076 124108 583082 124160
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589550 122856 589556 122868
rect 584456 122828 589556 122856
rect 584456 122816 584462 122828
rect 589550 122816 589556 122828
rect 589608 122816 589614 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 589918 122040 589924 122052
rect 580684 122012 589924 122040
rect 580684 122000 580690 122012
rect 589918 122000 589924 122012
rect 589976 122000 589982 122052
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589550 121496 589556 121508
rect 587400 121468 589556 121496
rect 587400 121456 587406 121468
rect 589550 121456 589556 121468
rect 589608 121456 589614 121508
rect 583202 120708 583208 120760
rect 583260 120748 583266 120760
rect 589366 120748 589372 120760
rect 583260 120720 589372 120748
rect 583260 120708 583266 120720
rect 589366 120708 589372 120720
rect 589424 120708 589430 120760
rect 578510 118532 578516 118584
rect 578568 118572 578574 118584
rect 580258 118572 580264 118584
rect 578568 118544 580264 118572
rect 578568 118532 578574 118544
rect 580258 118532 580264 118544
rect 580316 118532 580322 118584
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 682378 117280 682384 117292
rect 675904 117252 682384 117280
rect 675904 117240 675910 117252
rect 682378 117240 682384 117252
rect 682436 117240 682442 117292
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583386 116940 583392 116952
rect 579580 116912 583392 116940
rect 579580 116900 579586 116912
rect 583386 116900 583392 116912
rect 583444 116900 583450 116952
rect 585778 115948 585784 116000
rect 585836 115988 585842 116000
rect 589458 115988 589464 116000
rect 585836 115960 589464 115988
rect 585836 115948 585842 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 584582 115200 584588 115252
rect 584640 115240 584646 115252
rect 589642 115240 589648 115252
rect 584640 115212 589648 115240
rect 584640 115200 584646 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585962 112860 585968 112872
rect 579580 112832 585968 112860
rect 579580 112820 579586 112832
rect 585962 112820 585968 112832
rect 586020 112820 586026 112872
rect 586146 112412 586152 112464
rect 586204 112452 586210 112464
rect 590102 112452 590108 112464
rect 586204 112424 590108 112452
rect 586204 112412 586210 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110236 579344 110288
rect 579396 110276 579402 110288
rect 581822 110276 581828 110288
rect 579396 110248 581828 110276
rect 579396 110236 579402 110248
rect 581822 110236 581828 110248
rect 581880 110236 581886 110288
rect 580442 109080 580448 109132
rect 580500 109120 580506 109132
rect 589458 109120 589464 109132
rect 580500 109092 589464 109120
rect 580500 109080 580506 109092
rect 589458 109080 589464 109092
rect 589516 109080 589522 109132
rect 578326 108944 578332 108996
rect 578384 108984 578390 108996
rect 580626 108984 580632 108996
rect 578384 108956 580632 108984
rect 578384 108944 578390 108956
rect 580626 108944 580632 108956
rect 580684 108944 580690 108996
rect 667934 108808 667940 108860
rect 667992 108848 667998 108860
rect 669958 108848 669964 108860
rect 667992 108820 669964 108848
rect 667992 108808 667998 108820
rect 669958 108808 669964 108820
rect 670016 108808 670022 108860
rect 582282 107652 582288 107704
rect 582340 107692 582346 107704
rect 589458 107692 589464 107704
rect 582340 107664 589464 107692
rect 582340 107652 582346 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 580258 106292 580264 106344
rect 580316 106332 580322 106344
rect 589458 106332 589464 106344
rect 580316 106304 589464 106332
rect 580316 106292 580322 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 579338 105612 579344 105664
rect 579396 105652 579402 105664
rect 582282 105652 582288 105664
rect 579396 105624 582288 105652
rect 579396 105612 579402 105624
rect 582282 105612 582288 105624
rect 582340 105612 582346 105664
rect 587158 104864 587164 104916
rect 587216 104904 587222 104916
rect 589826 104904 589832 104916
rect 587216 104876 589832 104904
rect 587216 104864 587222 104876
rect 589826 104864 589832 104876
rect 589884 104864 589890 104916
rect 668210 104796 668216 104848
rect 668268 104836 668274 104848
rect 670786 104836 670792 104848
rect 668268 104808 670792 104836
rect 668268 104796 668274 104808
rect 670786 104796 670792 104808
rect 670844 104796 670850 104848
rect 578510 103368 578516 103420
rect 578568 103408 578574 103420
rect 588722 103408 588728 103420
rect 578568 103380 588728 103408
rect 578568 103368 578574 103380
rect 588722 103368 588728 103380
rect 588780 103368 588786 103420
rect 579154 102076 579160 102128
rect 579212 102116 579218 102128
rect 584398 102116 584404 102128
rect 579212 102088 584404 102116
rect 579212 102076 579218 102088
rect 584398 102076 584404 102088
rect 584456 102076 584462 102128
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 578602 99968 578608 100020
rect 578660 100008 578666 100020
rect 587342 100008 587348 100020
rect 578660 99980 587348 100008
rect 578660 99968 578666 99980
rect 587342 99968 587348 99980
rect 587400 99968 587406 100020
rect 592678 99968 592684 100020
rect 592736 100008 592742 100020
rect 667934 100008 667940 100020
rect 592736 99980 667940 100008
rect 592736 99968 592742 99980
rect 667934 99968 667940 99980
rect 667992 99968 667998 100020
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 579522 99220 579528 99272
rect 579580 99260 579586 99272
rect 583202 99260 583208 99272
rect 579580 99232 583208 99260
rect 579580 99220 579586 99232
rect 583202 99220 583208 99232
rect 583260 99220 583266 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 624602 99016 624608 99068
rect 624660 99056 624666 99068
rect 634998 99056 635004 99068
rect 624660 99028 635004 99056
rect 624660 99016 624666 99028
rect 634998 99016 635004 99028
rect 635056 99016 635062 99068
rect 625062 98880 625068 98932
rect 625120 98920 625126 98932
rect 636286 98920 636292 98932
rect 625120 98892 636292 98920
rect 625120 98880 625126 98892
rect 636286 98880 636292 98892
rect 636344 98880 636350 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98608 647148 98660
rect 647200 98648 647206 98660
rect 661954 98648 661960 98660
rect 647200 98620 661960 98648
rect 647200 98608 647206 98620
rect 661954 98608 661960 98620
rect 662012 98608 662018 98660
rect 630490 98540 630496 98592
rect 630548 98580 630554 98592
rect 646590 98580 646596 98592
rect 630548 98552 646596 98580
rect 630548 98540 630554 98552
rect 646590 98540 646596 98552
rect 646648 98540 646654 98592
rect 629754 98268 629760 98320
rect 629812 98308 629818 98320
rect 645302 98308 645308 98320
rect 629812 98280 645308 98308
rect 629812 98268 629818 98280
rect 645302 98268 645308 98280
rect 645360 98268 645366 98320
rect 633618 98132 633624 98184
rect 633676 98172 633682 98184
rect 640702 98172 640708 98184
rect 633676 98144 640708 98172
rect 633676 98132 633682 98144
rect 640702 98132 640708 98144
rect 640760 98132 640766 98184
rect 631980 98076 632100 98104
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 628282 97928 628288 97980
rect 628340 97968 628346 97980
rect 631980 97968 632008 98076
rect 632072 98036 632100 98076
rect 642174 98036 642180 98048
rect 632072 98008 642180 98036
rect 642174 97996 642180 98008
rect 642232 97996 642238 98048
rect 628340 97940 632008 97968
rect 628340 97928 628346 97940
rect 659930 97928 659936 97980
rect 659988 97968 659994 97980
rect 665358 97968 665364 97980
rect 659988 97940 665364 97968
rect 659988 97928 659994 97940
rect 665358 97928 665364 97940
rect 665416 97928 665422 97980
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 647510 97832 647516 97844
rect 632756 97804 647516 97832
rect 632756 97792 632762 97804
rect 647510 97792 647516 97804
rect 647568 97792 647574 97844
rect 653950 97792 653956 97844
rect 654008 97832 654014 97844
rect 655054 97832 655060 97844
rect 654008 97804 655060 97832
rect 654008 97792 654014 97804
rect 655054 97792 655060 97804
rect 655112 97792 655118 97844
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 662506 97832 662512 97844
rect 655480 97804 662512 97832
rect 655480 97792 655486 97804
rect 662506 97792 662512 97804
rect 662564 97792 662570 97844
rect 631226 97656 631232 97708
rect 631284 97696 631290 97708
rect 647326 97696 647332 97708
rect 631284 97668 647332 97696
rect 631284 97656 631290 97668
rect 647326 97656 647332 97668
rect 647384 97656 647390 97708
rect 650362 97656 650368 97708
rect 650420 97696 650426 97708
rect 658274 97696 658280 97708
rect 650420 97668 658280 97696
rect 650420 97656 650426 97668
rect 658274 97656 658280 97668
rect 658332 97656 658338 97708
rect 659838 97696 659844 97708
rect 658844 97668 659844 97696
rect 627546 97520 627552 97572
rect 627604 97560 627610 97572
rect 633618 97560 633624 97572
rect 627604 97532 633624 97560
rect 627604 97520 627610 97532
rect 633618 97520 633624 97532
rect 633676 97520 633682 97572
rect 633802 97520 633808 97572
rect 633860 97560 633866 97572
rect 639230 97560 639236 97572
rect 633860 97532 639236 97560
rect 633860 97520 633866 97532
rect 639230 97520 639236 97532
rect 639288 97520 639294 97572
rect 643002 97520 643008 97572
rect 643060 97560 643066 97572
rect 658844 97560 658872 97668
rect 659838 97656 659844 97668
rect 659896 97656 659902 97708
rect 659562 97560 659568 97572
rect 643060 97532 658872 97560
rect 659028 97532 659568 97560
rect 643060 97520 643066 97532
rect 605466 97384 605472 97436
rect 605524 97424 605530 97436
rect 611906 97424 611912 97436
rect 605524 97396 611912 97424
rect 605524 97384 605530 97396
rect 611906 97384 611912 97396
rect 611964 97384 611970 97436
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 620278 97424 620284 97436
rect 612700 97396 620284 97424
rect 612700 97384 612706 97396
rect 620278 97384 620284 97396
rect 620336 97384 620342 97436
rect 623130 97384 623136 97436
rect 623188 97424 623194 97436
rect 632054 97424 632060 97436
rect 623188 97396 632060 97424
rect 623188 97384 623194 97396
rect 632054 97384 632060 97396
rect 632112 97384 632118 97436
rect 633250 97384 633256 97436
rect 633308 97424 633314 97436
rect 650546 97424 650552 97436
rect 633308 97396 650552 97424
rect 633308 97384 633314 97396
rect 650546 97384 650552 97396
rect 650604 97384 650610 97436
rect 651834 97384 651840 97436
rect 651892 97424 651898 97436
rect 659028 97424 659056 97532
rect 659562 97520 659568 97532
rect 659620 97520 659626 97572
rect 651892 97396 659056 97424
rect 651892 97384 651898 97396
rect 659194 97384 659200 97436
rect 659252 97424 659258 97436
rect 664346 97424 664352 97436
rect 659252 97396 664352 97424
rect 659252 97384 659258 97396
rect 664346 97384 664352 97396
rect 664404 97384 664410 97436
rect 592126 97248 592132 97300
rect 592184 97288 592190 97300
rect 598934 97288 598940 97300
rect 592184 97260 598940 97288
rect 592184 97248 592190 97260
rect 598934 97248 598940 97260
rect 598992 97248 598998 97300
rect 621658 97248 621664 97300
rect 621716 97288 621722 97300
rect 629294 97288 629300 97300
rect 621716 97260 629300 97288
rect 621716 97248 621722 97260
rect 629294 97248 629300 97260
rect 629352 97248 629358 97300
rect 631870 97248 631876 97300
rect 631928 97288 631934 97300
rect 648614 97288 648620 97300
rect 631928 97260 648620 97288
rect 631928 97248 631934 97260
rect 648614 97248 648620 97260
rect 648672 97248 648678 97300
rect 656802 97180 656808 97232
rect 656860 97220 656866 97232
rect 661402 97220 661408 97232
rect 656860 97192 661408 97220
rect 656860 97180 656866 97192
rect 661402 97180 661408 97192
rect 661460 97180 661466 97232
rect 620094 97112 620100 97164
rect 620152 97152 620158 97164
rect 626350 97152 626356 97164
rect 620152 97124 626356 97152
rect 620152 97112 620158 97124
rect 626350 97112 626356 97124
rect 626408 97112 626414 97164
rect 626810 97112 626816 97164
rect 626868 97152 626874 97164
rect 633802 97152 633808 97164
rect 626868 97124 633808 97152
rect 626868 97112 626874 97124
rect 633802 97112 633808 97124
rect 633860 97112 633866 97164
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 649074 97152 649080 97164
rect 634228 97124 649080 97152
rect 634228 97112 634234 97124
rect 649074 97112 649080 97124
rect 649132 97112 649138 97164
rect 658090 97044 658096 97096
rect 658148 97084 658154 97096
rect 663058 97084 663064 97096
rect 658148 97056 663064 97084
rect 658148 97044 658154 97056
rect 663058 97044 663064 97056
rect 663116 97044 663122 97096
rect 634722 96976 634728 97028
rect 634780 97016 634786 97028
rect 647050 97016 647056 97028
rect 634780 96988 647056 97016
rect 634780 96976 634786 96988
rect 647050 96976 647056 96988
rect 647108 96976 647114 97028
rect 596174 96908 596180 96960
rect 596232 96948 596238 96960
rect 596726 96948 596732 96960
rect 596232 96920 596732 96948
rect 596232 96908 596238 96920
rect 596726 96908 596732 96920
rect 596784 96908 596790 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 656710 96908 656716 96960
rect 656768 96948 656774 96960
rect 660114 96948 660120 96960
rect 656768 96920 660120 96948
rect 656768 96908 656774 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 626074 96840 626080 96892
rect 626132 96880 626138 96892
rect 637758 96880 637764 96892
rect 626132 96852 637764 96880
rect 626132 96840 626138 96852
rect 637758 96840 637764 96852
rect 637816 96840 637822 96892
rect 644290 96772 644296 96824
rect 644348 96812 644354 96824
rect 658826 96812 658832 96824
rect 644348 96784 658832 96812
rect 644348 96772 644354 96784
rect 658826 96772 658832 96784
rect 658884 96772 658890 96824
rect 609146 96704 609152 96756
rect 609204 96744 609210 96756
rect 609698 96744 609704 96756
rect 609204 96716 609704 96744
rect 609204 96704 609210 96716
rect 609698 96704 609704 96716
rect 609756 96704 609762 96756
rect 640058 96568 640064 96620
rect 640116 96608 640122 96620
rect 645118 96608 645124 96620
rect 640116 96580 645124 96608
rect 640116 96568 640122 96580
rect 645118 96568 645124 96580
rect 645176 96568 645182 96620
rect 646406 96568 646412 96620
rect 646464 96608 646470 96620
rect 652018 96608 652024 96620
rect 646464 96580 652024 96608
rect 646464 96568 646470 96580
rect 652018 96568 652024 96580
rect 652076 96568 652082 96620
rect 653306 96568 653312 96620
rect 653364 96608 653370 96620
rect 665174 96608 665180 96620
rect 653364 96580 665180 96608
rect 653364 96568 653370 96580
rect 665174 96568 665180 96580
rect 665232 96568 665238 96620
rect 638586 96432 638592 96484
rect 638644 96472 638650 96484
rect 641346 96472 641352 96484
rect 638644 96444 641352 96472
rect 638644 96432 638650 96444
rect 641346 96432 641352 96444
rect 641404 96432 641410 96484
rect 641530 96432 641536 96484
rect 641588 96472 641594 96484
rect 648062 96472 648068 96484
rect 641588 96444 648068 96472
rect 641588 96432 641594 96444
rect 648062 96432 648068 96444
rect 648120 96432 648126 96484
rect 648890 96432 648896 96484
rect 648948 96472 648954 96484
rect 664530 96472 664536 96484
rect 648948 96444 664536 96472
rect 648948 96432 648954 96444
rect 664530 96432 664536 96444
rect 664588 96432 664594 96484
rect 648264 96376 648568 96404
rect 637574 96296 637580 96348
rect 637632 96336 637638 96348
rect 648264 96336 648292 96376
rect 637632 96308 648292 96336
rect 648540 96336 648568 96376
rect 660666 96336 660672 96348
rect 648540 96308 660672 96336
rect 637632 96296 637638 96308
rect 660666 96296 660672 96308
rect 660724 96296 660730 96348
rect 644934 96160 644940 96212
rect 644992 96200 644998 96212
rect 647878 96200 647884 96212
rect 644992 96172 647884 96200
rect 644992 96160 644998 96172
rect 647878 96160 647884 96172
rect 647936 96160 647942 96212
rect 649258 96160 649264 96212
rect 649316 96200 649322 96212
rect 663978 96200 663984 96212
rect 649316 96172 663984 96200
rect 649316 96160 649322 96172
rect 663978 96160 663984 96172
rect 664036 96160 664042 96212
rect 591298 96024 591304 96076
rect 591356 96064 591362 96076
rect 602614 96064 602620 96076
rect 591356 96036 602620 96064
rect 591356 96024 591362 96036
rect 602614 96024 602620 96036
rect 602672 96024 602678 96076
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 621658 96064 621664 96076
rect 610676 96036 621664 96064
rect 610676 96024 610682 96036
rect 621658 96024 621664 96036
rect 621716 96024 621722 96076
rect 640518 96024 640524 96076
rect 640576 96064 640582 96076
rect 645578 96064 645584 96076
rect 640576 96036 645584 96064
rect 640576 96024 640582 96036
rect 645578 96024 645584 96036
rect 645636 96024 645642 96076
rect 645762 96024 645768 96076
rect 645820 96064 645826 96076
rect 648062 96064 648068 96076
rect 645820 96036 648068 96064
rect 645820 96024 645826 96036
rect 648062 96024 648068 96036
rect 648120 96024 648126 96076
rect 648798 96024 648804 96076
rect 648856 96064 648862 96076
rect 664162 96064 664168 96076
rect 648856 96036 664168 96064
rect 648856 96024 648862 96036
rect 664162 96024 664168 96036
rect 664220 96024 664226 96076
rect 594058 95888 594064 95940
rect 594116 95928 594122 95940
rect 668026 95928 668032 95940
rect 594116 95900 668032 95928
rect 594116 95888 594122 95900
rect 668026 95888 668032 95900
rect 668084 95888 668090 95940
rect 639046 95752 639052 95804
rect 639104 95792 639110 95804
rect 648798 95792 648804 95804
rect 639104 95764 648804 95792
rect 639104 95752 639110 95764
rect 648798 95752 648804 95764
rect 648856 95752 648862 95804
rect 652570 95752 652576 95804
rect 652628 95792 652634 95804
rect 663794 95792 663800 95804
rect 652628 95764 663800 95792
rect 652628 95752 652634 95764
rect 663794 95752 663800 95764
rect 663852 95752 663858 95804
rect 645118 95616 645124 95668
rect 645176 95656 645182 95668
rect 652202 95656 652208 95668
rect 645176 95628 652208 95656
rect 645176 95616 645182 95628
rect 652202 95616 652208 95628
rect 652260 95616 652266 95668
rect 656158 95520 656164 95532
rect 654106 95492 656164 95520
rect 641346 95412 641352 95464
rect 641404 95412 641410 95464
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 647878 95452 647884 95464
rect 643520 95424 647884 95452
rect 643520 95412 643526 95424
rect 647878 95412 647884 95424
rect 647936 95412 647942 95464
rect 641364 95316 641392 95412
rect 648062 95344 648068 95396
rect 648120 95384 648126 95396
rect 654106 95384 654134 95492
rect 656158 95480 656164 95492
rect 656216 95480 656222 95532
rect 648120 95356 654134 95384
rect 648120 95344 648126 95356
rect 647694 95316 647700 95328
rect 641364 95288 647700 95316
rect 647694 95276 647700 95288
rect 647752 95276 647758 95328
rect 578326 95140 578332 95192
rect 578384 95180 578390 95192
rect 584582 95180 584588 95192
rect 578384 95152 584588 95180
rect 578384 95140 578390 95152
rect 584582 95140 584588 95152
rect 584640 95140 584646 95192
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 625430 95180 625436 95192
rect 620980 95152 625436 95180
rect 620980 95140 620986 95152
rect 625430 95140 625436 95152
rect 625488 95140 625494 95192
rect 647050 95140 647056 95192
rect 647108 95180 647114 95192
rect 650270 95180 650276 95192
rect 647108 95152 650276 95180
rect 647108 95140 647114 95152
rect 650270 95140 650276 95152
rect 650328 95140 650334 95192
rect 590930 94936 590936 94988
rect 590988 94976 590994 94988
rect 592126 94976 592132 94988
rect 590988 94948 592132 94976
rect 590988 94936 590994 94948
rect 592126 94936 592132 94948
rect 592184 94936 592190 94988
rect 616506 94936 616512 94988
rect 616564 94976 616570 94988
rect 624970 94976 624976 94988
rect 616564 94948 624976 94976
rect 616564 94936 616570 94948
rect 624970 94936 624976 94948
rect 625028 94936 625034 94988
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 620922 94500 620928 94512
rect 607732 94472 620928 94500
rect 607732 94460 607738 94472
rect 620922 94460 620928 94472
rect 620980 94460 620986 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626166 93820 626172 93832
rect 619600 93792 626172 93820
rect 619600 93780 619606 93792
rect 626166 93780 626172 93792
rect 626224 93780 626230 93832
rect 647510 93712 647516 93764
rect 647568 93752 647574 93764
rect 648246 93752 648252 93764
rect 647568 93724 648252 93752
rect 647568 93712 647574 93724
rect 648246 93712 648252 93724
rect 648304 93712 648310 93764
rect 651282 93576 651288 93628
rect 651340 93616 651346 93628
rect 654686 93616 654692 93628
rect 651340 93588 654692 93616
rect 651340 93576 651346 93588
rect 654686 93576 654692 93588
rect 654744 93576 654750 93628
rect 579246 93372 579252 93424
rect 579304 93412 579310 93424
rect 586146 93412 586152 93424
rect 579304 93384 586152 93412
rect 579304 93372 579310 93384
rect 586146 93372 586152 93384
rect 586204 93372 586210 93424
rect 609698 93100 609704 93152
rect 609756 93140 609762 93152
rect 618622 93140 618628 93152
rect 609756 93112 618628 93140
rect 609756 93100 609762 93112
rect 618622 93100 618628 93112
rect 618680 93100 618686 93152
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647694 92420 647700 92472
rect 647752 92460 647758 92472
rect 655422 92460 655428 92472
rect 647752 92432 655428 92460
rect 647752 92420 647758 92432
rect 655422 92420 655428 92432
rect 655480 92420 655486 92472
rect 577498 91740 577504 91792
rect 577556 91780 577562 91792
rect 590930 91780 590936 91792
rect 577556 91752 590936 91780
rect 577556 91740 577562 91752
rect 590930 91740 590936 91752
rect 590988 91740 590994 91792
rect 606938 91740 606944 91792
rect 606996 91780 607002 91792
rect 622394 91780 622400 91792
rect 606996 91752 622400 91780
rect 606996 91740 607002 91752
rect 622394 91740 622400 91752
rect 622452 91740 622458 91792
rect 578694 91400 578700 91452
rect 578752 91440 578758 91452
rect 585778 91440 585784 91452
rect 578752 91412 585784 91440
rect 578752 91400 578758 91412
rect 585778 91400 585784 91412
rect 585836 91400 585842 91452
rect 618162 91128 618168 91180
rect 618220 91168 618226 91180
rect 618220 91140 618392 91168
rect 618220 91128 618226 91140
rect 611262 90992 611268 91044
rect 611320 91032 611326 91044
rect 618162 91032 618168 91044
rect 611320 91004 618168 91032
rect 611320 90992 611326 91004
rect 618162 90992 618168 91004
rect 618220 90992 618226 91044
rect 618364 91032 618392 91140
rect 626442 91032 626448 91044
rect 618364 91004 626448 91032
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 648798 90788 648804 90840
rect 648856 90828 648862 90840
rect 655422 90828 655428 90840
rect 648856 90800 655428 90828
rect 648856 90788 648862 90800
rect 655422 90788 655428 90800
rect 655480 90788 655486 90840
rect 620922 89632 620928 89684
rect 620980 89672 620986 89684
rect 625430 89672 625436 89684
rect 620980 89644 625436 89672
rect 620980 89632 620986 89644
rect 625430 89632 625436 89644
rect 625488 89632 625494 89684
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664346 88788 664352 88800
rect 662380 88760 664352 88788
rect 662380 88748 662386 88760
rect 664346 88748 664352 88760
rect 664404 88748 664410 88800
rect 656158 88612 656164 88664
rect 656216 88652 656222 88664
rect 657446 88652 657452 88664
rect 656216 88624 657452 88652
rect 656216 88612 656222 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 579246 88272 579252 88324
rect 579304 88312 579310 88324
rect 589918 88312 589924 88324
rect 579304 88284 589924 88312
rect 579304 88272 579310 88284
rect 589918 88272 589924 88284
rect 589976 88272 589982 88324
rect 618162 88272 618168 88324
rect 618220 88312 618226 88324
rect 625614 88312 625620 88324
rect 618220 88284 625620 88312
rect 618220 88272 618226 88284
rect 625614 88272 625620 88284
rect 625672 88272 625678 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 622394 88136 622400 88188
rect 622452 88176 622458 88188
rect 626442 88176 626448 88188
rect 622452 88148 626448 88176
rect 622452 88136 622458 88148
rect 626442 88136 626448 88148
rect 626500 88136 626506 88188
rect 648430 86980 648436 87032
rect 648488 87020 648494 87032
rect 662506 87020 662512 87032
rect 648488 86992 662512 87020
rect 648488 86980 648494 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 652202 86708 652208 86760
rect 652260 86748 652266 86760
rect 660114 86748 660120 86760
rect 652260 86720 660120 86748
rect 652260 86708 652266 86720
rect 660114 86708 660120 86720
rect 660172 86708 660178 86760
rect 647878 86572 647884 86624
rect 647936 86612 647942 86624
rect 661402 86612 661408 86624
rect 647936 86584 661408 86612
rect 647936 86572 647942 86584
rect 661402 86572 661408 86584
rect 661460 86572 661466 86624
rect 652018 86436 652024 86488
rect 652076 86476 652082 86488
rect 657170 86476 657176 86488
rect 652076 86448 657176 86476
rect 652076 86436 652082 86448
rect 657170 86436 657176 86448
rect 657228 86436 657234 86488
rect 621658 86300 621664 86352
rect 621716 86340 621722 86352
rect 626442 86340 626448 86352
rect 621716 86312 626448 86340
rect 621716 86300 621722 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 656342 86300 656348 86352
rect 656400 86340 656406 86352
rect 660666 86340 660672 86352
rect 656400 86312 660672 86340
rect 656400 86300 656406 86312
rect 660666 86300 660672 86312
rect 660724 86300 660730 86352
rect 618622 85484 618628 85536
rect 618680 85524 618686 85536
rect 626442 85524 626448 85536
rect 618680 85496 626448 85524
rect 618680 85484 618686 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 609882 85348 609888 85400
rect 609940 85388 609946 85400
rect 609940 85360 625154 85388
rect 609940 85348 609946 85360
rect 625126 85320 625154 85360
rect 625338 85320 625344 85332
rect 625126 85292 625344 85320
rect 625338 85280 625344 85292
rect 625396 85280 625402 85332
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625798 84164 625804 84176
rect 608560 84136 625804 84164
rect 608560 84124 608566 84136
rect 625798 84124 625804 84136
rect 625856 84124 625862 84176
rect 579246 83988 579252 84040
rect 579304 84028 579310 84040
rect 581638 84028 581644 84040
rect 579304 84000 581644 84028
rect 579304 83988 579310 84000
rect 581638 83988 581644 84000
rect 581696 83988 581702 84040
rect 578694 82764 578700 82816
rect 578752 82804 578758 82816
rect 583018 82804 583024 82816
rect 578752 82776 583024 82804
rect 578752 82764 578758 82776
rect 583018 82764 583024 82776
rect 583076 82764 583082 82816
rect 579062 82084 579068 82136
rect 579120 82124 579126 82136
rect 587158 82124 587164 82136
rect 579120 82096 587164 82124
rect 579120 82084 579126 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 81064 628748 81116
rect 628800 81104 628806 81116
rect 642450 81104 642456 81116
rect 628800 81076 642456 81104
rect 628800 81064 628806 81076
rect 642450 81064 642456 81076
rect 642508 81064 642514 81116
rect 615402 80928 615408 80980
rect 615460 80968 615466 80980
rect 646130 80968 646136 80980
rect 615460 80940 646136 80968
rect 615460 80928 615466 80940
rect 646130 80928 646136 80940
rect 646188 80928 646194 80980
rect 613838 80792 613844 80844
rect 613896 80832 613902 80844
rect 647326 80832 647332 80844
rect 613896 80804 647332 80832
rect 613896 80792 613902 80804
rect 647326 80792 647332 80804
rect 647384 80792 647390 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 614022 79432 614028 79484
rect 614080 79472 614086 79484
rect 645946 79472 645952 79484
rect 614080 79444 645952 79472
rect 614080 79432 614086 79444
rect 645946 79432 645952 79444
rect 646004 79432 646010 79484
rect 583018 79296 583024 79348
rect 583076 79336 583082 79348
rect 600498 79336 600504 79348
rect 583076 79308 600504 79336
rect 583076 79296 583082 79308
rect 600498 79296 600504 79308
rect 600556 79296 600562 79348
rect 612642 79296 612648 79348
rect 612700 79336 612706 79348
rect 648614 79336 648620 79348
rect 612700 79308 648620 79336
rect 612700 79296 612706 79308
rect 648614 79296 648620 79308
rect 648672 79296 648678 79348
rect 578510 78412 578516 78464
rect 578568 78452 578574 78464
rect 580258 78452 580264 78464
rect 578568 78424 580264 78452
rect 578568 78412 578574 78424
rect 580258 78412 580264 78424
rect 580316 78412 580322 78464
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77664 628472 77716
rect 628524 77704 628530 77716
rect 632790 77704 632796 77716
rect 628524 77676 632796 77704
rect 628524 77664 628530 77676
rect 632790 77664 632796 77676
rect 632848 77664 632854 77716
rect 624418 77392 624424 77444
rect 624476 77432 624482 77444
rect 628466 77432 628472 77444
rect 624476 77404 628472 77432
rect 624476 77392 624482 77404
rect 628466 77392 628472 77404
rect 628524 77392 628530 77444
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 620278 76780 620284 76832
rect 620336 76820 620342 76832
rect 648982 76820 648988 76832
rect 620336 76792 648988 76820
rect 620336 76780 620342 76792
rect 648982 76780 648988 76792
rect 649040 76780 649046 76832
rect 611998 76644 612004 76696
rect 612056 76684 612062 76696
rect 662414 76684 662420 76696
rect 612056 76656 662420 76684
rect 612056 76644 612062 76656
rect 662414 76644 662420 76656
rect 662472 76644 662478 76696
rect 587158 76508 587164 76560
rect 587216 76548 587222 76560
rect 668210 76548 668216 76560
rect 587216 76520 668216 76548
rect 587216 76508 587222 76520
rect 668210 76508 668216 76520
rect 668268 76508 668274 76560
rect 616782 75420 616788 75472
rect 616840 75460 616846 75472
rect 646498 75460 646504 75472
rect 616840 75432 646504 75460
rect 616840 75420 616846 75432
rect 646498 75420 646504 75432
rect 646556 75420 646562 75472
rect 607122 75284 607128 75336
rect 607180 75324 607186 75336
rect 646314 75324 646320 75336
rect 607180 75296 646320 75324
rect 607180 75284 607186 75296
rect 646314 75284 646320 75296
rect 646372 75284 646378 75336
rect 578878 75148 578884 75200
rect 578936 75188 578942 75200
rect 666554 75188 666560 75200
rect 578936 75160 666560 75188
rect 578936 75148 578942 75160
rect 666554 75148 666560 75160
rect 666612 75148 666618 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 588538 73148 588544 73160
rect 579580 73120 588544 73148
rect 579580 73108 579586 73120
rect 588538 73108 588544 73120
rect 588596 73108 588602 73160
rect 578510 71544 578516 71596
rect 578568 71584 578574 71596
rect 584398 71584 584404 71596
rect 578568 71556 584404 71584
rect 578568 71544 578574 71556
rect 584398 71544 584404 71556
rect 584456 71544 584462 71596
rect 579522 66852 579528 66904
rect 579580 66892 579586 66904
rect 625982 66892 625988 66904
rect 579580 66864 625988 66892
rect 579580 66852 579586 66864
rect 625982 66852 625988 66864
rect 626040 66852 626046 66904
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 592678 64852 592684 64864
rect 579580 64824 592684 64852
rect 579580 64812 579586 64824
rect 592678 64812 592684 64824
rect 592736 64812 592742 64864
rect 579522 62024 579528 62076
rect 579580 62064 579586 62076
rect 587158 62064 587164 62076
rect 579580 62036 587164 62064
rect 579580 62024 579586 62036
rect 587158 62024 587164 62036
rect 587216 62024 587222 62076
rect 578326 59984 578332 60036
rect 578384 60024 578390 60036
rect 624418 60024 624424 60036
rect 578384 59996 624424 60024
rect 578384 59984 578390 59996
rect 624418 59984 624424 59996
rect 624476 59984 624482 60036
rect 577682 58760 577688 58812
rect 577740 58800 577746 58812
rect 604454 58800 604460 58812
rect 577740 58772 604460 58800
rect 577740 58760 577746 58772
rect 604454 58760 604460 58772
rect 604512 58760 604518 58812
rect 576118 58624 576124 58676
rect 576176 58664 576182 58676
rect 603074 58664 603080 58676
rect 576176 58636 603080 58664
rect 576176 58624 576182 58636
rect 603074 58624 603080 58636
rect 603132 58624 603138 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 594058 57916 594064 57928
rect 579580 57888 594064 57916
rect 579580 57876 579586 57888
rect 594058 57876 594064 57888
rect 594116 57876 594122 57928
rect 577314 57196 577320 57248
rect 577372 57236 577378 57248
rect 600314 57236 600320 57248
rect 577372 57208 600320 57236
rect 577372 57196 577378 57208
rect 600314 57196 600320 57208
rect 600372 57196 600378 57248
rect 574278 55972 574284 56024
rect 574336 56012 574342 56024
rect 598934 56012 598940 56024
rect 574336 55984 598940 56012
rect 574336 55972 574342 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 577130 55836 577136 55888
rect 577188 55876 577194 55888
rect 601878 55876 601884 55888
rect 577188 55848 601884 55876
rect 577188 55836 577194 55848
rect 601878 55836 601884 55848
rect 601936 55836 601942 55888
rect 577314 55604 577320 55616
rect 564452 55576 577320 55604
rect 466426 55508 483014 55536
rect 466426 55332 466454 55508
rect 464080 55304 466454 55332
rect 470704 55372 478184 55400
rect 460768 54080 460934 54108
rect 460382 53592 460388 53644
rect 460440 53632 460446 53644
rect 460768 53632 460796 54080
rect 460440 53604 460796 53632
rect 460906 53632 460934 54080
rect 461946 53632 461952 53644
rect 460906 53604 461952 53632
rect 460440 53592 460446 53604
rect 461946 53592 461952 53604
rect 462004 53592 462010 53644
rect 462222 53592 462228 53644
rect 462280 53632 462286 53644
rect 464080 53632 464108 55304
rect 470704 55196 470732 55372
rect 464724 55168 470732 55196
rect 470796 55236 478092 55264
rect 464724 53904 464752 55168
rect 470796 54992 470824 55236
rect 478064 55060 478092 55236
rect 478156 55196 478184 55372
rect 482986 55332 483014 55508
rect 564452 55332 564480 55576
rect 577314 55564 577320 55576
rect 577372 55564 577378 55616
rect 482986 55304 564480 55332
rect 569236 55440 579614 55468
rect 569236 55196 569264 55440
rect 478156 55168 569264 55196
rect 569328 55304 574968 55332
rect 569328 55060 569356 55304
rect 465138 54964 470824 54992
rect 473096 55032 475792 55060
rect 478064 55032 569356 55060
rect 574940 55060 574968 55304
rect 579586 55196 579614 55440
rect 596450 55196 596456 55208
rect 579586 55168 596456 55196
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 596174 55060 596180 55072
rect 574940 55032 596180 55060
rect 464724 53876 464936 53904
rect 464908 53644 464936 53876
rect 465138 53644 465166 54964
rect 473096 54924 473124 55032
rect 475764 54992 475792 55032
rect 596174 55020 596180 55032
rect 596232 55020 596238 55072
rect 475764 54964 476344 54992
rect 472820 54896 473124 54924
rect 476316 54924 476344 54964
rect 597646 54924 597652 54936
rect 476316 54896 597652 54924
rect 472820 54856 472848 54896
rect 597646 54884 597652 54896
rect 597704 54884 597710 54936
rect 465552 54828 472848 54856
rect 465552 53644 465580 54828
rect 597922 54788 597928 54800
rect 473326 54760 597928 54788
rect 473326 54720 473354 54760
rect 597922 54748 597928 54760
rect 597980 54748 597986 54800
rect 465736 54692 473354 54720
rect 465736 53644 465764 54692
rect 580442 54652 580448 54664
rect 475672 54624 580448 54652
rect 475672 54584 475700 54624
rect 580442 54612 580448 54624
rect 580500 54612 580506 54664
rect 473280 54556 475700 54584
rect 473280 54312 473308 54556
rect 625798 54516 625804 54528
rect 475764 54488 565676 54516
rect 475764 54380 475792 54488
rect 565648 54448 565676 54488
rect 574296 54488 625804 54516
rect 574296 54448 574324 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 565648 54420 574324 54448
rect 583018 54380 583024 54392
rect 469968 54284 473308 54312
rect 473924 54352 475792 54380
rect 476316 54352 565032 54380
rect 469968 53644 469996 54284
rect 473924 54176 473952 54352
rect 472820 54148 473952 54176
rect 472820 53644 472848 54148
rect 476316 54108 476344 54352
rect 476086 54080 476344 54108
rect 476592 54216 564756 54244
rect 476086 54040 476114 54080
rect 473924 54012 476114 54040
rect 473004 53808 473354 53836
rect 462280 53604 464108 53632
rect 462280 53592 462286 53604
rect 464890 53592 464896 53644
rect 464948 53592 464954 53644
rect 465074 53592 465080 53644
rect 465132 53604 465166 53644
rect 465132 53592 465138 53604
rect 465534 53592 465540 53644
rect 465592 53592 465598 53644
rect 465718 53592 465724 53644
rect 465776 53592 465782 53644
rect 469950 53592 469956 53644
rect 470008 53592 470014 53644
rect 472802 53592 472808 53644
rect 472860 53592 472866 53644
rect 459462 53456 459468 53508
rect 459520 53496 459526 53508
rect 473004 53496 473032 53808
rect 459520 53468 473032 53496
rect 473326 53496 473354 53808
rect 473924 53644 473952 54012
rect 476592 53836 476620 54216
rect 564728 54176 564756 54216
rect 565004 54176 565032 54352
rect 579586 54352 583024 54380
rect 579586 54312 579614 54352
rect 583018 54340 583024 54352
rect 583076 54340 583082 54392
rect 565464 54284 579614 54312
rect 565464 54176 565492 54284
rect 577498 54176 577504 54188
rect 564728 54148 564940 54176
rect 565004 54148 565492 54176
rect 574066 54148 577504 54176
rect 476086 53808 476620 53836
rect 476684 54080 564664 54108
rect 473906 53592 473912 53644
rect 473964 53592 473970 53644
rect 476086 53496 476114 53808
rect 476684 53644 476712 54080
rect 478156 53944 564434 53972
rect 478156 53644 478184 53944
rect 564406 53904 564434 53944
rect 564406 53876 564572 53904
rect 482986 53808 563054 53836
rect 476666 53592 476672 53644
rect 476724 53592 476730 53644
rect 478138 53592 478144 53644
rect 478196 53592 478202 53644
rect 473326 53468 476114 53496
rect 459520 53456 459526 53468
rect 50522 53320 50528 53372
rect 50580 53360 50586 53372
rect 130378 53360 130384 53372
rect 50580 53332 130384 53360
rect 50580 53320 50586 53332
rect 130378 53320 130384 53332
rect 130436 53320 130442 53372
rect 461302 53320 461308 53372
rect 461360 53360 461366 53372
rect 482986 53360 483014 53808
rect 461360 53332 483014 53360
rect 461360 53320 461366 53332
rect 563026 53292 563054 53808
rect 564544 53644 564572 53876
rect 564636 53768 564664 54080
rect 564912 54040 564940 54148
rect 574066 54108 574094 54148
rect 577498 54136 577504 54148
rect 577556 54136 577562 54188
rect 569052 54080 574094 54108
rect 569052 54040 569080 54080
rect 564912 54012 569080 54040
rect 574738 53932 574744 53984
rect 574796 53972 574802 53984
rect 623038 53972 623044 53984
rect 574796 53944 623044 53972
rect 574796 53932 574802 53944
rect 623038 53932 623044 53944
rect 623096 53932 623102 53984
rect 564636 53740 572714 53768
rect 564526 53592 564532 53644
rect 564584 53592 564590 53644
rect 572686 53496 572714 53740
rect 577130 53496 577136 53508
rect 572686 53468 577136 53496
rect 577130 53456 577136 53468
rect 577188 53456 577194 53508
rect 574278 53292 574284 53304
rect 563026 53264 574284 53292
rect 574278 53252 574284 53264
rect 574336 53252 574342 53304
rect 48958 53184 48964 53236
rect 49016 53224 49022 53236
rect 129182 53224 129188 53236
rect 49016 53196 129188 53224
rect 49016 53184 49022 53196
rect 129182 53184 129188 53196
rect 129240 53184 129246 53236
rect 464522 53184 464528 53236
rect 464580 53224 464586 53236
rect 465534 53224 465540 53236
rect 464580 53196 465540 53224
rect 464580 53184 464586 53196
rect 465534 53184 465540 53196
rect 465592 53184 465598 53236
rect 465902 53184 465908 53236
rect 465960 53224 465966 53236
rect 478138 53224 478144 53236
rect 465960 53196 478144 53224
rect 465960 53184 465966 53196
rect 478138 53184 478144 53196
rect 478196 53184 478202 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 47578 53048 47584 53100
rect 47636 53088 47642 53100
rect 128998 53088 129004 53100
rect 47636 53060 129004 53088
rect 47636 53048 47642 53060
rect 128998 53048 129004 53060
rect 129056 53048 129062 53100
rect 476666 53088 476672 53100
rect 462286 53060 476672 53088
rect 459600 52776 459606 52828
rect 459658 52816 459664 52828
rect 462286 52816 462314 53060
rect 476666 53048 476672 53060
rect 476724 53048 476730 53100
rect 463602 52912 463608 52964
rect 463660 52952 463666 52964
rect 465718 52952 465724 52964
rect 463660 52924 465724 52952
rect 463660 52912 463666 52924
rect 465718 52912 465724 52924
rect 465776 52912 465782 52964
rect 459658 52788 462314 52816
rect 459658 52776 459664 52788
rect 463740 52776 463746 52828
rect 463798 52816 463804 52828
rect 465074 52816 465080 52828
rect 463798 52788 465080 52816
rect 463798 52776 463804 52788
rect 465074 52776 465080 52788
rect 465132 52776 465138 52828
rect 465442 52776 465448 52828
rect 465500 52816 465506 52828
rect 469950 52816 469956 52828
rect 465500 52788 469956 52816
rect 465500 52776 465506 52788
rect 469950 52776 469956 52788
rect 470008 52776 470014 52828
rect 50338 51824 50344 51876
rect 50396 51864 50402 51876
rect 129366 51864 129372 51876
rect 50396 51836 129372 51864
rect 50396 51824 50402 51836
rect 129366 51824 129372 51836
rect 129424 51824 129430 51876
rect 46198 51688 46204 51740
rect 46256 51728 46262 51740
rect 130562 51728 130568 51740
rect 46256 51700 130568 51728
rect 46256 51688 46262 51700
rect 130562 51688 130568 51700
rect 130620 51688 130626 51740
rect 145374 51688 145380 51740
rect 145432 51728 145438 51740
rect 306006 51728 306012 51740
rect 145432 51700 306012 51728
rect 145432 51688 145438 51700
rect 306006 51688 306012 51700
rect 306064 51688 306070 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 49142 50328 49148 50380
rect 49200 50368 49206 50380
rect 131022 50368 131028 50380
rect 49200 50340 131028 50368
rect 49200 50328 49206 50340
rect 131022 50328 131028 50340
rect 131080 50328 131086 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 129642 49144 129648 49156
rect 51776 49116 129648 49144
rect 51776 49104 51782 49116
rect 129642 49104 129648 49116
rect 129700 49104 129706 49156
rect 45462 48968 45468 49020
rect 45520 49008 45526 49020
rect 128998 49008 129004 49020
rect 45520 48980 129004 49008
rect 45520 48968 45526 48980
rect 128998 48968 129004 48980
rect 129056 48968 129062 49020
rect 625982 46452 625988 46504
rect 626040 46492 626046 46504
rect 661770 46492 661776 46504
rect 626040 46464 661776 46492
rect 626040 46452 626046 46464
rect 661770 46452 661776 46464
rect 661828 46452 661834 46504
rect 128998 46044 129004 46096
rect 129056 46084 129062 46096
rect 132402 46084 132408 46096
rect 129056 46056 132408 46084
rect 129056 46044 129062 46056
rect 132402 46044 132408 46056
rect 132460 46044 132466 46096
rect 130562 45908 130568 45960
rect 130620 45948 130626 45960
rect 132586 45948 132592 45960
rect 130620 45920 132592 45948
rect 130620 45908 130626 45920
rect 132586 45908 132592 45920
rect 132644 45908 132650 45960
rect 129642 45364 129648 45416
rect 129700 45404 129706 45416
rect 129700 45376 131206 45404
rect 129700 45364 129706 45376
rect 131178 45336 131206 45376
rect 131178 45308 131298 45336
rect 43806 45160 43812 45212
rect 43864 45200 43870 45212
rect 131114 45200 131120 45212
rect 43864 45172 131120 45200
rect 43864 45160 43870 45172
rect 131114 45160 131120 45172
rect 131172 45160 131178 45212
rect 131270 45090 131298 45308
rect 131390 45296 131396 45348
rect 131448 45336 131454 45348
rect 132954 45336 132960 45348
rect 131448 45308 132960 45336
rect 131448 45296 131454 45308
rect 132954 45296 132960 45308
rect 133012 45296 133018 45348
rect 131390 45160 131396 45212
rect 131448 45200 131454 45212
rect 133138 45200 133144 45212
rect 131448 45172 133144 45200
rect 131448 45160 131454 45172
rect 133138 45160 133144 45172
rect 133196 45160 133202 45212
rect 129366 45024 129372 45076
rect 129424 45064 129430 45076
rect 129424 45036 131068 45064
rect 129424 45024 129430 45036
rect 131040 45020 131068 45036
rect 131040 44992 131330 45020
rect 126422 44888 126428 44940
rect 126480 44928 126486 44940
rect 126480 44900 131620 44928
rect 126480 44888 126486 44900
rect 131684 44824 131790 44852
rect 129182 44752 129188 44804
rect 129240 44792 129246 44804
rect 131684 44792 131712 44824
rect 129240 44764 131712 44792
rect 129240 44752 129246 44764
rect 131868 44740 131974 44768
rect 131868 44600 131896 44740
rect 132144 44656 132172 44670
rect 131776 44588 131896 44600
rect 125566 44572 131896 44588
rect 132052 44628 132172 44656
rect 125566 44560 131804 44572
rect 43622 44276 43628 44328
rect 43680 44316 43686 44328
rect 125566 44316 125594 44560
rect 128814 44344 128820 44396
rect 128872 44384 128878 44396
rect 132052 44384 132080 44628
rect 132420 44464 132448 44586
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 132604 44416 132632 44502
rect 128872 44356 132080 44384
rect 132586 44364 132592 44416
rect 132644 44364 132650 44416
rect 128872 44344 128878 44356
rect 43680 44288 125594 44316
rect 43680 44276 43686 44288
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 126422 44180 126428 44192
rect 43496 44152 126428 44180
rect 43496 44140 43502 44152
rect 126422 44140 126428 44152
rect 126480 44140 126486 44192
rect 132742 44180 132770 44390
rect 132954 44252 132960 44304
rect 133012 44252 133018 44304
rect 131776 44152 132770 44180
rect 130378 44004 130384 44056
rect 130436 44044 130442 44056
rect 131776 44044 131804 44152
rect 133138 44140 133144 44192
rect 133196 44140 133202 44192
rect 130436 44016 131804 44044
rect 130436 44004 130442 44016
rect 440234 43800 440240 43852
rect 440292 43840 440298 43852
rect 441062 43840 441068 43852
rect 440292 43812 441068 43840
rect 440292 43800 440298 43812
rect 441062 43800 441068 43812
rect 441120 43800 441126 43852
rect 410886 42848 410892 42900
rect 410944 42888 410950 42900
rect 415578 42888 415584 42900
rect 410944 42860 415584 42888
rect 410944 42848 410950 42860
rect 415578 42848 415584 42860
rect 415636 42848 415642 42900
rect 187326 42780 187332 42832
rect 187384 42820 187390 42832
rect 255866 42820 255872 42832
rect 187384 42792 255872 42820
rect 187384 42780 187390 42792
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 310422 42712 310428 42764
rect 310480 42752 310486 42764
rect 364518 42752 364524 42764
rect 310480 42724 364524 42752
rect 310480 42712 310486 42724
rect 364518 42712 364524 42724
rect 364576 42712 364582 42764
rect 431218 42752 431224 42764
rect 364720 42724 431224 42752
rect 361758 42440 361764 42492
rect 361816 42480 361822 42492
rect 364720 42480 364748 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 453574 42712 453580 42764
rect 453632 42752 453638 42764
rect 464338 42752 464344 42764
rect 453632 42724 464344 42752
rect 453632 42712 453638 42724
rect 464338 42712 464344 42724
rect 464396 42712 464402 42764
rect 364886 42576 364892 42628
rect 364944 42616 364950 42628
rect 427078 42616 427084 42628
rect 364944 42588 427084 42616
rect 364944 42576 364950 42588
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 441246 42576 441252 42628
rect 441304 42616 441310 42628
rect 446398 42616 446404 42628
rect 441304 42588 446404 42616
rect 441304 42576 441310 42588
rect 446398 42576 446404 42588
rect 446456 42576 446462 42628
rect 454678 42576 454684 42628
rect 454736 42616 454742 42628
rect 462958 42616 462964 42628
rect 454736 42588 462964 42616
rect 454736 42576 454742 42588
rect 462958 42576 462964 42588
rect 463016 42576 463022 42628
rect 410886 42480 410892 42492
rect 361816 42452 364748 42480
rect 373966 42452 410892 42480
rect 361816 42440 361822 42452
rect 364518 42304 364524 42356
rect 364576 42344 364582 42356
rect 373966 42344 373994 42452
rect 410886 42440 410892 42452
rect 410944 42440 410950 42492
rect 429102 42480 429108 42492
rect 422266 42452 429108 42480
rect 364576 42316 373994 42344
rect 364576 42304 364582 42316
rect 415578 42304 415584 42356
rect 415636 42344 415642 42356
rect 422266 42344 422294 42452
rect 429102 42440 429108 42452
rect 429160 42440 429166 42492
rect 454494 42440 454500 42492
rect 454552 42480 454558 42492
rect 463694 42480 463700 42492
rect 454552 42452 463700 42480
rect 454552 42440 454558 42452
rect 463694 42440 463700 42452
rect 463752 42440 463758 42492
rect 415636 42316 422294 42344
rect 415636 42304 415642 42316
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 427078 41964 427084 42016
rect 427136 42004 427142 42016
rect 427136 41976 427814 42004
rect 427136 41964 427142 41976
rect 427786 41868 427814 41976
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 446398 41964 446404 42016
rect 446456 42004 446462 42016
rect 454494 42004 454500 42016
rect 446456 41976 454500 42004
rect 446456 41964 446462 41976
rect 454494 41964 454500 41976
rect 454552 41964 454558 42016
rect 441246 41868 441252 41880
rect 427786 41840 441252 41868
rect 441246 41828 441252 41840
rect 441304 41828 441310 41880
rect 454678 41868 454684 41880
rect 441586 41840 454684 41868
rect 429102 41692 429108 41744
rect 429160 41732 429166 41744
rect 441586 41732 441614 41840
rect 454678 41828 454684 41840
rect 454736 41828 454742 41880
rect 429160 41704 441614 41732
rect 429160 41692 429166 41704
rect 449158 41692 449164 41744
rect 449216 41732 449222 41744
rect 453574 41732 453580 41744
rect 449216 41704 453580 41732
rect 449216 41692 449222 41704
rect 453574 41692 453580 41704
rect 453632 41692 453638 41744
<< via1 >>
rect 652024 896996 652076 897048
rect 676036 897064 676088 897116
rect 654784 895772 654836 895824
rect 675852 895772 675904 895824
rect 672724 895636 672776 895688
rect 676036 895636 676088 895688
rect 671988 894412 672040 894464
rect 676036 894412 676088 894464
rect 671436 894276 671488 894328
rect 675852 894276 675904 894328
rect 672356 892984 672408 893036
rect 675852 892984 675904 893036
rect 673368 892848 673420 892900
rect 676036 892848 676088 892900
rect 676220 891488 676272 891540
rect 676864 891488 676916 891540
rect 676036 889992 676088 890044
rect 677048 889992 677100 890044
rect 674380 888904 674432 888956
rect 676036 888904 676088 888956
rect 674840 888700 674892 888752
rect 675668 888700 675720 888752
rect 674656 888496 674708 888548
rect 676036 888496 676088 888548
rect 674196 888088 674248 888140
rect 676036 888088 676088 888140
rect 671804 886864 671856 886916
rect 675484 886864 675536 886916
rect 673184 885640 673236 885692
rect 676036 885640 676088 885692
rect 675208 881084 675260 881136
rect 683304 881084 683356 881136
rect 653404 880472 653456 880524
rect 675576 880472 675628 880524
rect 675944 880132 675996 880184
rect 679624 880132 679676 880184
rect 675760 879316 675812 879368
rect 677048 879316 677100 879368
rect 674932 879112 674984 879164
rect 678244 879112 678296 879164
rect 675392 878976 675444 879028
rect 676864 878976 676916 879028
rect 675760 878364 675812 878416
rect 675484 877208 675536 877260
rect 674196 873604 674248 873656
rect 675116 873604 675168 873656
rect 674840 872380 674892 872432
rect 675300 872380 675352 872432
rect 674656 869796 674708 869848
rect 675208 869796 675260 869848
rect 674380 869592 674432 869644
rect 674840 869592 674892 869644
rect 657544 869388 657596 869440
rect 675024 869388 675076 869440
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 654140 868028 654192 868080
rect 674748 868028 674800 868080
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35808 817096 35860 817148
rect 46204 817096 46256 817148
rect 35624 816960 35676 817012
rect 61384 816960 61436 817012
rect 35808 815736 35860 815788
rect 44272 815736 44324 815788
rect 35440 815600 35492 815652
rect 44824 815600 44876 815652
rect 35624 814376 35676 814428
rect 44548 814376 44600 814428
rect 35808 814240 35860 814292
rect 45100 814240 45152 814292
rect 41328 812812 41380 812864
rect 43352 812812 43404 812864
rect 40960 810704 41012 810756
rect 42524 810704 42576 810756
rect 41144 807440 41196 807492
rect 43168 807440 43220 807492
rect 40960 807304 41012 807356
rect 45284 807304 45336 807356
rect 31760 806624 31812 806676
rect 35624 806624 35676 806676
rect 44824 806556 44876 806608
rect 62764 806556 62816 806608
rect 44916 806420 44968 806472
rect 45284 806420 45336 806472
rect 41328 805944 41380 805996
rect 43812 805944 43864 805996
rect 35624 802612 35676 802664
rect 42340 802612 42392 802664
rect 33048 802408 33100 802460
rect 42156 802408 42208 802460
rect 33784 801252 33836 801304
rect 39856 801252 39908 801304
rect 31024 801048 31076 801100
rect 40684 801048 40736 801100
rect 43536 799076 43588 799128
rect 53104 799076 53156 799128
rect 42892 797648 42944 797700
rect 57244 797648 57296 797700
rect 42248 796288 42300 796340
rect 42892 796288 42944 796340
rect 43536 794996 43588 795048
rect 44916 794996 44968 795048
rect 42248 794792 42300 794844
rect 43076 794792 43128 794844
rect 42340 793772 42392 793824
rect 43444 793772 43496 793824
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 671620 789352 671672 789404
rect 675116 789352 675168 789404
rect 57244 789148 57296 789200
rect 62120 789148 62172 789200
rect 42708 786632 42760 786684
rect 62120 786632 62172 786684
rect 46204 785136 46256 785188
rect 62120 785136 62172 785188
rect 673000 783844 673052 783896
rect 675116 783844 675168 783896
rect 673736 782620 673788 782672
rect 675116 782620 675168 782672
rect 669228 782484 669280 782536
rect 675300 782484 675352 782536
rect 655520 781192 655572 781244
rect 675024 781192 675076 781244
rect 673920 779968 673972 780020
rect 675116 779968 675168 780020
rect 673552 778540 673604 778592
rect 675300 778540 675352 778592
rect 655060 778336 655112 778388
rect 675116 778336 675168 778388
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 674288 776976 674340 777028
rect 675300 776976 675352 777028
rect 674656 775684 674708 775736
rect 675116 775684 675168 775736
rect 651472 775548 651524 775600
rect 669964 775548 670016 775600
rect 672172 775548 672224 775600
rect 675024 775548 675076 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 669780 774256 669832 774308
rect 675116 774256 675168 774308
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 60004 774188 60056 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655060 773780 655112 773832
rect 35808 773304 35860 773356
rect 41696 773304 41748 773356
rect 35808 773100 35860 773152
rect 41052 773100 41104 773152
rect 35624 772964 35676 773016
rect 41512 772964 41564 773016
rect 35440 772828 35492 772880
rect 41328 772828 41380 772880
rect 42064 772828 42116 772880
rect 61384 772828 61436 772880
rect 35532 771808 35584 771860
rect 39764 771808 39816 771860
rect 42064 771604 42116 771656
rect 45100 771604 45152 771656
rect 35808 771536 35860 771588
rect 41696 771536 41748 771588
rect 35348 771400 35400 771452
rect 41696 771400 41748 771452
rect 42064 771400 42116 771452
rect 44548 771400 44600 771452
rect 35808 770448 35860 770500
rect 40316 770448 40368 770500
rect 35624 770176 35676 770228
rect 41696 770244 41748 770296
rect 42064 770244 42116 770296
rect 43260 770244 43312 770296
rect 35808 770040 35860 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44272 770040 44324 770092
rect 35808 768952 35860 769004
rect 39580 768952 39632 769004
rect 35532 768816 35584 768868
rect 40684 768816 40736 768868
rect 35348 768680 35400 768732
rect 41696 768680 41748 768732
rect 35808 767524 35860 767576
rect 35808 767320 35860 767372
rect 36544 767320 36596 767372
rect 41696 767252 41748 767304
rect 35808 766096 35860 766148
rect 41236 766096 41288 766148
rect 35808 764804 35860 764856
rect 40868 764804 40920 764856
rect 35808 764532 35860 764584
rect 41512 764532 41564 764584
rect 35808 763308 35860 763360
rect 39304 763308 39356 763360
rect 35624 763172 35676 763224
rect 41512 763240 41564 763292
rect 35808 761880 35860 761932
rect 38936 761880 38988 761932
rect 33048 760996 33100 761048
rect 41512 760996 41564 761048
rect 35164 759636 35216 759688
rect 40040 759636 40092 759688
rect 39304 757732 39356 757784
rect 41604 757732 41656 757784
rect 44732 755488 44784 755540
rect 62764 755488 62816 755540
rect 43444 754876 43496 754928
rect 45284 754876 45336 754928
rect 42248 754264 42300 754316
rect 44732 754264 44784 754316
rect 42248 753856 42300 753908
rect 42984 753856 43036 753908
rect 43628 753652 43680 753704
rect 45100 753652 45152 753704
rect 61384 746988 61436 747040
rect 62396 746988 62448 747040
rect 45100 746512 45152 746564
rect 62120 746512 62172 746564
rect 670792 745220 670844 745272
rect 675024 745220 675076 745272
rect 42708 743996 42760 744048
rect 62120 743860 62172 743912
rect 671252 743792 671304 743844
rect 675116 743792 675168 743844
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 60004 742364 60056 742416
rect 62120 742364 62172 742416
rect 670148 739100 670200 739152
rect 675392 739100 675444 739152
rect 674196 738624 674248 738676
rect 675392 738624 675444 738676
rect 668400 736924 668452 736976
rect 675300 736924 675352 736976
rect 652024 736176 652076 736228
rect 653404 736176 653456 736228
rect 657544 735564 657596 735616
rect 667480 735564 667532 735616
rect 667480 734816 667532 734868
rect 675208 734816 675260 734868
rect 673644 734272 673696 734324
rect 675300 734272 675352 734324
rect 654784 734136 654836 734188
rect 670976 734136 671028 734188
rect 675300 733592 675352 733644
rect 651472 733388 651524 733440
rect 668584 733388 668636 733440
rect 675300 733252 675352 733304
rect 651472 732776 651524 732828
rect 661684 732776 661736 732828
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 651472 731280 651524 731332
rect 671252 731280 671304 731332
rect 672540 730464 672592 730516
rect 675208 730464 675260 730516
rect 43444 730328 43496 730380
rect 61384 730328 61436 730380
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 667848 729920 667900 729972
rect 675208 729920 675260 729972
rect 42248 729308 42300 729360
rect 62764 729308 62816 729360
rect 41328 729036 41380 729088
rect 41696 729036 41748 729088
rect 42064 728628 42116 728680
rect 43076 728628 43128 728680
rect 670332 728628 670384 728680
rect 675300 728628 675352 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 673184 728288 673236 728340
rect 671804 728084 671856 728136
rect 674656 727880 674708 727932
rect 683304 727880 683356 727932
rect 672816 727812 672868 727864
rect 673460 727812 673512 727864
rect 675116 727744 675168 727796
rect 677324 727744 677376 727796
rect 675024 727608 675076 727660
rect 40868 727404 40920 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 44548 727404 44600 727456
rect 674840 727404 674892 727456
rect 41328 727268 41380 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 45008 727268 45060 727320
rect 674656 727268 674708 727320
rect 675024 727268 675076 727320
rect 674380 726588 674432 726640
rect 683488 726588 683540 726640
rect 41328 726180 41380 726232
rect 41696 726180 41748 726232
rect 41144 725908 41196 725960
rect 41604 725908 41656 725960
rect 672816 723120 672868 723172
rect 673552 723120 673604 723172
rect 673736 722168 673788 722220
rect 673736 722032 673788 722084
rect 673920 721964 673972 722016
rect 673920 721760 673972 721812
rect 675760 721692 675812 721744
rect 675944 721692 675996 721744
rect 675760 721216 675812 721268
rect 675944 721216 675996 721268
rect 675760 720808 675812 720860
rect 675944 720808 675996 720860
rect 673920 720536 673972 720588
rect 675760 720468 675812 720520
rect 675944 720468 675996 720520
rect 673920 720400 673972 720452
rect 43076 719720 43128 719772
rect 42892 719516 42944 719568
rect 42708 719380 42760 719432
rect 43076 719380 43128 719432
rect 674288 716456 674340 716508
rect 676036 716456 676088 716508
rect 653404 716252 653456 716304
rect 674012 716252 674064 716304
rect 35164 715776 35216 715828
rect 41696 715776 41748 715828
rect 669964 715708 670016 715760
rect 674012 715708 674064 715760
rect 33784 715640 33836 715692
rect 40408 715640 40460 715692
rect 32956 715504 33008 715556
rect 40592 715504 40644 715556
rect 671436 715300 671488 715352
rect 674012 715300 674064 715352
rect 671068 714960 671120 715012
rect 674012 714960 674064 715012
rect 674288 714892 674340 714944
rect 676036 714892 676088 714944
rect 660304 714824 660356 714876
rect 674012 714824 674064 714876
rect 671988 714484 672040 714536
rect 674012 714484 674064 714536
rect 672356 713668 672408 713720
rect 674012 713668 674064 713720
rect 671344 713192 671396 713244
rect 674012 713192 674064 713244
rect 671160 712376 671212 712428
rect 674012 712376 674064 712428
rect 42892 712104 42944 712156
rect 50344 712104 50396 712156
rect 676220 712036 676272 712088
rect 677324 712036 677376 712088
rect 672172 709996 672224 710048
rect 674012 709996 674064 710048
rect 42248 709724 42300 709776
rect 44640 709724 44692 709776
rect 671620 709588 671672 709640
rect 674012 709588 674064 709640
rect 674288 709520 674340 709572
rect 676036 709520 676088 709572
rect 669228 709316 669280 709368
rect 674012 709316 674064 709368
rect 42248 707956 42300 708008
rect 44640 707956 44692 708008
rect 674288 707956 674340 708008
rect 675852 707956 675904 708008
rect 674472 707548 674524 707600
rect 676036 707548 676088 707600
rect 674656 707140 674708 707192
rect 676036 707140 676088 707192
rect 42248 705508 42300 705560
rect 43628 705508 43680 705560
rect 669780 705372 669832 705424
rect 674012 705372 674064 705424
rect 674288 705304 674340 705356
rect 683120 705304 683172 705356
rect 50344 705100 50396 705152
rect 62120 705100 62172 705152
rect 669228 703808 669280 703860
rect 674012 703808 674064 703860
rect 674288 703808 674340 703860
rect 676036 703808 676088 703860
rect 44456 703740 44508 703792
rect 62120 703740 62172 703792
rect 673460 701428 673512 701480
rect 673920 701428 673972 701480
rect 666468 701224 666520 701276
rect 674012 701224 674064 701276
rect 674288 701224 674340 701276
rect 675116 701224 675168 701276
rect 42708 701020 42760 701072
rect 62212 701020 62264 701072
rect 654784 701020 654836 701072
rect 674012 701020 674064 701072
rect 674288 701020 674340 701072
rect 675392 701020 675444 701072
rect 42892 700408 42944 700460
rect 43076 700340 43128 700392
rect 43076 700204 43128 700256
rect 42892 700068 42944 700120
rect 46204 698164 46256 698216
rect 62120 698164 62172 698216
rect 666284 696940 666336 696992
rect 673736 696940 673788 696992
rect 674472 693472 674524 693524
rect 675392 693472 675444 693524
rect 674288 692996 674340 693048
rect 675116 692996 675168 693048
rect 656440 690072 656492 690124
rect 673736 690072 673788 690124
rect 652760 688780 652812 688832
rect 673736 688780 673788 688832
rect 651472 688644 651524 688696
rect 657544 688644 657596 688696
rect 42708 687284 42760 687336
rect 61384 687216 61436 687268
rect 651472 687216 651524 687268
rect 669964 687216 670016 687268
rect 651472 687012 651524 687064
rect 654784 687012 654836 687064
rect 43444 686468 43496 686520
rect 62764 686468 62816 686520
rect 651656 686468 651708 686520
rect 667204 686468 667256 686520
rect 41328 686264 41380 686316
rect 41696 686264 41748 686316
rect 42064 686264 42116 686316
rect 43076 686264 43128 686316
rect 41144 686060 41196 686112
rect 41696 686060 41748 686112
rect 42064 686060 42116 686112
rect 45192 686060 45244 686112
rect 40868 685856 40920 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45192 685856 45244 685908
rect 668768 685856 668820 685908
rect 672172 685856 672224 685908
rect 651472 685516 651524 685568
rect 656440 685516 656492 685568
rect 41052 684700 41104 684752
rect 41696 684700 41748 684752
rect 41328 683408 41380 683460
rect 41696 683408 41748 683460
rect 42064 683408 42116 683460
rect 42708 683408 42760 683460
rect 41144 683272 41196 683324
rect 41696 683272 41748 683324
rect 42064 683272 42116 683324
rect 44272 683272 44324 683324
rect 40776 683136 40828 683188
rect 41696 683136 41748 683188
rect 42064 683136 42116 683188
rect 45008 683136 45060 683188
rect 674564 682388 674616 682440
rect 683212 682388 683264 682440
rect 41328 681980 41380 682032
rect 41696 681980 41748 682032
rect 42064 681980 42116 682032
rect 42524 681980 42576 682032
rect 40960 679124 41012 679176
rect 41328 679124 41380 679176
rect 41144 678988 41196 679040
rect 41696 678988 41748 679040
rect 42064 678988 42116 679040
rect 45008 678988 45060 679040
rect 40960 677696 41012 677748
rect 41604 677696 41656 677748
rect 35164 672868 35216 672920
rect 38844 672868 38896 672920
rect 33784 672732 33836 672784
rect 37924 672732 37976 672784
rect 42432 671508 42484 671560
rect 42708 671100 42760 671152
rect 668584 671100 668636 671152
rect 673920 671100 673972 671152
rect 661684 670692 661736 670744
rect 673552 670692 673604 670744
rect 670976 670080 671028 670132
rect 673920 670080 673972 670132
rect 658924 669468 658976 669520
rect 673552 669468 673604 669520
rect 45376 669332 45428 669384
rect 53104 669332 53156 669384
rect 669596 669332 669648 669384
rect 673920 669332 673972 669384
rect 671344 668516 671396 668568
rect 673920 668516 673972 668568
rect 671528 668176 671580 668228
rect 673552 668176 673604 668228
rect 45744 667904 45796 667956
rect 57244 667904 57296 667956
rect 671344 667904 671396 667956
rect 673920 667904 673972 667956
rect 42248 667428 42300 667480
rect 45376 667428 45428 667480
rect 671160 666884 671212 666936
rect 673920 666884 673972 666936
rect 669412 666544 669464 666596
rect 673552 666544 673604 666596
rect 670884 666000 670936 666052
rect 673920 666000 673972 666052
rect 42340 665796 42392 665848
rect 45744 665796 45796 665848
rect 42248 665388 42300 665440
rect 43996 665388 44048 665440
rect 672540 665388 672592 665440
rect 673552 665388 673604 665440
rect 668952 665184 669004 665236
rect 673920 665184 673972 665236
rect 670332 664436 670384 664488
rect 673920 664436 673972 664488
rect 670148 663960 670200 664012
rect 673920 663960 673972 664012
rect 674932 663960 674984 664012
rect 676220 663960 676272 664012
rect 42432 663552 42484 663604
rect 42432 663076 42484 663128
rect 668400 661920 668452 661972
rect 673920 661920 673972 661972
rect 670516 661580 670568 661632
rect 673920 661580 673972 661632
rect 667388 661104 667440 661156
rect 673920 661104 673972 661156
rect 53104 660900 53156 660952
rect 62120 660900 62172 660952
rect 42156 660492 42208 660544
rect 43628 660492 43680 660544
rect 667848 660152 667900 660204
rect 673920 660152 673972 660204
rect 674564 659812 674616 659864
rect 683120 659812 683172 659864
rect 672172 659676 672224 659728
rect 673920 659676 673972 659728
rect 57244 659540 57296 659592
rect 62120 659540 62172 659592
rect 42524 657228 42576 657280
rect 62120 657500 62172 657552
rect 653404 655528 653456 655580
rect 673920 655528 673972 655580
rect 44824 655460 44876 655512
rect 62120 655460 62172 655512
rect 667572 647232 667624 647284
rect 674012 647232 674064 647284
rect 655520 645872 655572 645924
rect 670976 645872 671028 645924
rect 35808 644444 35860 644496
rect 41696 644444 41748 644496
rect 42064 644444 42116 644496
rect 60004 644444 60056 644496
rect 674932 643560 674984 643612
rect 35808 643492 35860 643544
rect 40500 643492 40552 643544
rect 675116 643492 675168 643544
rect 674932 643424 674984 643476
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 45192 643288 45244 643340
rect 674748 643288 674800 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 61384 643084 61436 643136
rect 655336 643084 655388 643136
rect 674012 643084 674064 643136
rect 674564 642744 674616 642796
rect 675300 642744 675352 642796
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62764 642336 62816 642388
rect 651472 642336 651524 642388
rect 658924 642336 658976 642388
rect 35624 641996 35676 642048
rect 39580 641996 39632 642048
rect 35808 641724 35860 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 44640 641724 44692 641776
rect 35808 640704 35860 640756
rect 39948 640704 40000 640756
rect 35348 640432 35400 640484
rect 41696 640500 41748 640552
rect 42064 640500 42116 640552
rect 44640 640500 44692 640552
rect 35532 640296 35584 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 44272 640296 44324 640348
rect 651472 640296 651524 640348
rect 668584 640296 668636 640348
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 35808 639140 35860 639192
rect 37924 639072 37976 639124
rect 35808 638936 35860 638988
rect 41696 638868 41748 638920
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 35808 637576 35860 637628
rect 36544 637576 36596 637628
rect 35624 636828 35676 636880
rect 39120 636828 39172 636880
rect 674288 636828 674340 636880
rect 683304 636828 683356 636880
rect 35532 636488 35584 636540
rect 39764 636488 39816 636540
rect 35808 636216 35860 636268
rect 39948 636216 40000 636268
rect 669596 635604 669648 635656
rect 670240 635604 670292 635656
rect 35808 634924 35860 634976
rect 41420 634924 41472 634976
rect 35808 633700 35860 633752
rect 39120 633700 39172 633752
rect 35808 633428 35860 633480
rect 40408 633428 40460 633480
rect 669412 633088 669464 633140
rect 671160 633088 671212 633140
rect 669504 631320 669556 631372
rect 669872 631320 669924 631372
rect 36544 630708 36596 630760
rect 41512 630708 41564 630760
rect 32036 629892 32088 629944
rect 37740 629892 37792 629944
rect 42064 629484 42116 629536
rect 42708 629484 42760 629536
rect 674288 627852 674340 627904
rect 675392 627852 675444 627904
rect 670056 625948 670108 626000
rect 673552 625948 673604 626000
rect 45744 625812 45796 625864
rect 62948 625812 63000 625864
rect 667204 625676 667256 625728
rect 674012 625676 674064 625728
rect 674932 625676 674984 625728
rect 676496 625676 676548 625728
rect 657544 625132 657596 625184
rect 674012 625132 674064 625184
rect 670148 624656 670200 624708
rect 674012 624656 674064 624708
rect 42340 624452 42392 624504
rect 44364 624452 44416 624504
rect 671528 624316 671580 624368
rect 674012 624316 674064 624368
rect 671620 623840 671672 623892
rect 674012 623840 674064 623892
rect 671344 623500 671396 623552
rect 674012 623500 674064 623552
rect 669964 623024 670016 623076
rect 674012 623024 674064 623076
rect 669504 622888 669556 622940
rect 669504 622752 669556 622804
rect 670332 622208 670384 622260
rect 674012 622208 674064 622260
rect 668216 621732 668268 621784
rect 674012 621732 674064 621784
rect 666468 621052 666520 621104
rect 674012 621052 674064 621104
rect 674380 620848 674432 620900
rect 675392 620848 675444 620900
rect 668768 620236 668820 620288
rect 674012 620236 674064 620288
rect 42248 619624 42300 619676
rect 44180 619624 44232 619676
rect 666284 619624 666336 619676
rect 673644 619624 673696 619676
rect 672356 619012 672408 619064
rect 674012 619012 674064 619064
rect 42156 617244 42208 617296
rect 42708 617244 42760 617296
rect 668032 616904 668084 616956
rect 674012 616904 674064 616956
rect 44364 616768 44416 616820
rect 62120 616768 62172 616820
rect 670700 616564 670752 616616
rect 674012 616564 674064 616616
rect 669780 615476 669832 615528
rect 674012 615476 674064 615528
rect 675116 615476 675168 615528
rect 683120 615476 683172 615528
rect 670700 614864 670752 614916
rect 674012 614864 674064 614916
rect 43076 614252 43128 614304
rect 44456 614252 44508 614304
rect 42616 614116 42668 614168
rect 62120 614116 62172 614168
rect 43904 612688 43956 612740
rect 60004 612620 60056 612672
rect 62120 612620 62172 612672
rect 44088 612348 44140 612400
rect 43766 612144 43818 612196
rect 44088 612008 44140 612060
rect 43996 611736 44048 611788
rect 44272 611600 44324 611652
rect 44088 611532 44140 611584
rect 44211 611328 44263 611380
rect 44318 611124 44370 611176
rect 44824 611192 44876 611244
rect 653404 611328 653456 611380
rect 674012 611328 674064 611380
rect 674840 604528 674892 604580
rect 675300 604528 675352 604580
rect 35808 601672 35860 601724
rect 36544 601672 36596 601724
rect 657544 600312 657596 600364
rect 673828 600312 673880 600364
rect 654784 598952 654836 599004
rect 673828 599428 673880 599480
rect 651472 597524 651524 597576
rect 667204 597524 667256 597576
rect 42892 597388 42944 597440
rect 42892 596980 42944 597032
rect 651472 596164 651524 596216
rect 660304 596164 660356 596216
rect 39948 595756 40000 595808
rect 41696 595756 41748 595808
rect 651656 595416 651708 595468
rect 653404 595416 653456 595468
rect 675024 595212 675076 595264
rect 675208 595008 675260 595060
rect 651472 594872 651524 594924
rect 656164 594872 656216 594924
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 38568 594260 38620 594312
rect 41604 594260 41656 594312
rect 36544 593036 36596 593088
rect 41696 593036 41748 593088
rect 651472 593036 651524 593088
rect 654784 593036 654836 593088
rect 675484 591404 675536 591456
rect 683212 591404 683264 591456
rect 674380 591268 674432 591320
rect 683396 591268 683448 591320
rect 35624 587256 35676 587308
rect 39580 587256 39632 587308
rect 33048 587120 33100 587172
rect 41420 587120 41472 587172
rect 33784 585896 33836 585948
rect 40224 585896 40276 585948
rect 31024 585760 31076 585812
rect 39948 585760 40000 585812
rect 42156 585760 42208 585812
rect 42708 585760 42760 585812
rect 652024 581000 652076 581052
rect 674012 581000 674064 581052
rect 670148 580388 670200 580440
rect 674012 580388 674064 580440
rect 668584 580252 668636 580304
rect 674012 580252 674064 580304
rect 674288 580252 674340 580304
rect 676404 580252 676456 580304
rect 674288 580116 674340 580168
rect 676220 580116 676272 580168
rect 658924 579640 658976 579692
rect 674012 579640 674064 579692
rect 669780 579232 669832 579284
rect 674012 579232 674064 579284
rect 674288 579232 674340 579284
rect 676220 579232 676272 579284
rect 671620 579028 671672 579080
rect 674012 579028 674064 579080
rect 674288 578416 674340 578468
rect 676220 578416 676272 578468
rect 671528 578280 671580 578332
rect 674012 578280 674064 578332
rect 42248 578212 42300 578264
rect 42708 578212 42760 578264
rect 669964 578076 670016 578128
rect 674012 578076 674064 578128
rect 674288 578076 674340 578128
rect 676220 578076 676272 578128
rect 674840 577872 674892 577924
rect 675484 577872 675536 577924
rect 670332 577804 670384 577856
rect 674012 577804 674064 577856
rect 674288 577736 674340 577788
rect 675852 577736 675904 577788
rect 674288 577600 674340 577652
rect 676220 577600 676272 577652
rect 670240 577464 670292 577516
rect 674012 577464 674064 577516
rect 671160 576920 671212 576972
rect 674012 576920 674064 576972
rect 674288 575968 674340 576020
rect 676220 575968 676272 576020
rect 668400 575492 668452 575544
rect 674012 575492 674064 575544
rect 44640 575424 44692 575476
rect 62120 575424 62172 575476
rect 670976 574540 671028 574592
rect 674012 574540 674064 574592
rect 671988 574268 672040 574320
rect 674012 574268 674064 574320
rect 674288 574132 674340 574184
rect 676220 574132 676272 574184
rect 667572 574064 667624 574116
rect 674012 574064 674064 574116
rect 45560 573996 45612 574048
rect 62120 573996 62172 574048
rect 42156 573452 42208 573504
rect 42616 573452 42668 573504
rect 669504 573044 669556 573096
rect 674012 573044 674064 573096
rect 674288 572908 674340 572960
rect 676220 572908 676272 572960
rect 667756 572704 667808 572756
rect 674012 572704 674064 572756
rect 674288 571888 674340 571940
rect 676220 571888 676272 571940
rect 670424 571412 670476 571464
rect 674012 571412 674064 571464
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 674288 570052 674340 570104
rect 676220 570052 676272 570104
rect 671988 569916 672040 569968
rect 674012 569916 674064 569968
rect 674288 569236 674340 569288
rect 676220 569236 676272 569288
rect 670056 568556 670108 568608
rect 674012 568556 674064 568608
rect 653404 565836 653456 565888
rect 673828 565836 673880 565888
rect 674472 559308 674524 559360
rect 675116 559308 675168 559360
rect 674288 558220 674340 558272
rect 675392 558220 675444 558272
rect 674656 557540 674708 557592
rect 675116 557540 675168 557592
rect 657820 554752 657872 554804
rect 673828 554752 673880 554804
rect 674472 554684 674524 554736
rect 675116 554684 675168 554736
rect 655152 553392 655204 553444
rect 673828 553664 673880 553716
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 651472 552032 651524 552084
rect 658924 552032 658976 552084
rect 40040 550944 40092 550996
rect 41696 550944 41748 550996
rect 651472 550604 651524 550656
rect 669596 550604 669648 550656
rect 651380 550332 651432 550384
rect 653404 550332 653456 550384
rect 675024 549992 675076 550044
rect 675300 549788 675352 549840
rect 651472 549040 651524 549092
rect 657820 549040 657872 549092
rect 651472 548836 651524 548888
rect 655152 548836 655204 548888
rect 31760 547408 31812 547460
rect 41604 547408 41656 547460
rect 675484 547136 675536 547188
rect 684316 547136 684368 547188
rect 675116 546864 675168 546916
rect 675116 546660 675168 546712
rect 674840 546456 674892 546508
rect 681004 546456 681056 546508
rect 675668 545708 675720 545760
rect 683304 545708 683356 545760
rect 34428 544348 34480 544400
rect 37832 544348 37884 544400
rect 42984 538160 43036 538212
rect 42800 537888 42852 537940
rect 667204 535644 667256 535696
rect 674012 535644 674064 535696
rect 660304 535440 660356 535492
rect 674012 535440 674064 535492
rect 669780 534964 669832 535016
rect 672724 534964 672776 535016
rect 656164 534216 656216 534268
rect 674012 534216 674064 534268
rect 670792 534080 670844 534132
rect 674012 534080 674064 534132
rect 670240 532924 670292 532976
rect 674012 532924 674064 532976
rect 42432 532720 42484 532772
rect 43168 532720 43220 532772
rect 671620 532720 671672 532772
rect 674012 532720 674064 532772
rect 671160 531700 671212 531752
rect 674012 531700 674064 531752
rect 671160 531292 671212 531344
rect 674012 531292 674064 531344
rect 44732 531224 44784 531276
rect 62120 531224 62172 531276
rect 60004 531088 60056 531140
rect 62304 531088 62356 531140
rect 667020 530476 667072 530528
rect 674012 530476 674064 530528
rect 671804 530204 671856 530256
rect 674012 530204 674064 530256
rect 42156 530068 42208 530120
rect 42984 530068 43036 530120
rect 669044 530000 669096 530052
rect 674012 529864 674064 529916
rect 671344 528708 671396 528760
rect 674012 528708 674064 528760
rect 45100 528572 45152 528624
rect 62120 528572 62172 528624
rect 668860 528572 668912 528624
rect 674012 528572 674064 528624
rect 42064 527756 42116 527808
rect 42616 527756 42668 527808
rect 672540 527348 672592 527400
rect 674012 527348 674064 527400
rect 672356 527144 672408 527196
rect 673644 527144 673696 527196
rect 681004 525716 681056 525768
rect 683120 525716 683172 525768
rect 676864 518916 676916 518968
rect 683304 518916 683356 518968
rect 677876 518780 677928 518832
rect 675484 518644 675536 518696
rect 675668 503820 675720 503872
rect 678244 503820 678296 503872
rect 674288 494708 674340 494760
rect 683212 494708 683264 494760
rect 669596 491852 669648 491904
rect 674012 491852 674064 491904
rect 674288 491784 674340 491836
rect 675852 491784 675904 491836
rect 674288 491648 674340 491700
rect 676036 491648 676088 491700
rect 665824 491444 665876 491496
rect 674012 491444 674064 491496
rect 658924 491308 658976 491360
rect 673828 491308 673880 491360
rect 670792 490900 670844 490952
rect 674012 490900 674064 490952
rect 671620 489268 671672 489320
rect 673920 489268 673972 489320
rect 671160 488452 671212 488504
rect 673920 488452 673972 488504
rect 675208 488452 675260 488504
rect 676036 488452 676088 488504
rect 668676 485800 668728 485852
rect 673920 485800 673972 485852
rect 670976 485596 671028 485648
rect 674012 485596 674064 485648
rect 667756 484372 667808 484424
rect 674012 484372 674064 484424
rect 670424 483964 670476 484016
rect 674012 483964 674064 484016
rect 674932 480428 674984 480480
rect 683120 480428 683172 480480
rect 675300 475192 675352 475244
rect 680360 475192 680412 475244
rect 669228 456560 669280 456612
rect 673368 455948 673420 456000
rect 672172 455812 672224 455864
rect 667388 455608 667440 455660
rect 670608 455472 670660 455524
rect 673276 455336 673328 455388
rect 672080 455064 672132 455116
rect 673388 455200 673440 455252
rect 674288 454996 674340 455048
rect 675484 454996 675536 455048
rect 673046 454792 673098 454844
rect 672908 454656 672960 454708
rect 672816 454384 672868 454436
rect 674288 454724 674340 454776
rect 676864 454724 676916 454776
rect 674288 454452 674340 454504
rect 675668 454452 675720 454504
rect 672448 453908 672500 453960
rect 35808 429156 35860 429208
rect 41696 429156 41748 429208
rect 41328 425076 41380 425128
rect 41696 425076 41748 425128
rect 40960 424260 41012 424312
rect 41512 424260 41564 424312
rect 32036 416168 32088 416220
rect 41696 416168 41748 416220
rect 53840 404268 53892 404320
rect 62120 404268 62172 404320
rect 674564 403248 674616 403300
rect 676220 403248 676272 403300
rect 45284 402908 45336 402960
rect 62120 402908 62172 402960
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 60004 400052 60056 400104
rect 62120 400052 62172 400104
rect 674840 398828 674892 398880
rect 676036 398828 676088 398880
rect 675024 396176 675076 396228
rect 676220 396176 676272 396228
rect 674380 396040 674432 396092
rect 676036 396040 676088 396092
rect 674656 395088 674708 395140
rect 676220 395088 676272 395140
rect 675208 389104 675260 389156
rect 679624 389104 679676 389156
rect 675208 386316 675260 386368
rect 675484 385976 675536 386028
rect 674840 384752 674892 384804
rect 675484 384752 675536 384804
rect 41328 382236 41380 382288
rect 41696 382236 41748 382288
rect 674380 382168 674432 382220
rect 675116 382168 675168 382220
rect 674380 378088 674432 378140
rect 675116 378088 675168 378140
rect 40224 378020 40276 378072
rect 41696 378020 41748 378072
rect 42064 377952 42116 378004
rect 42708 377952 42760 378004
rect 651472 373940 651524 373992
rect 657544 373940 657596 373992
rect 35164 371832 35216 371884
rect 41696 371832 41748 371884
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 42248 365236 42300 365288
rect 42248 364896 42300 364948
rect 42248 364284 42300 364336
rect 42708 364148 42760 364200
rect 46572 361496 46624 361548
rect 62120 361496 62172 361548
rect 45376 360136 45428 360188
rect 62120 360136 62172 360188
rect 44640 359592 44692 359644
rect 45376 359592 45428 359644
rect 44824 359456 44876 359508
rect 45468 359456 45520 359508
rect 51724 357416 51776 357468
rect 62120 357416 62172 357468
rect 44640 354696 44692 354748
rect 44824 354696 44876 354748
rect 44732 354424 44784 354476
rect 44855 354424 44907 354476
rect 45836 353880 45888 353932
rect 45836 353676 45888 353728
rect 45303 353472 45355 353524
rect 45422 353200 45474 353252
rect 676036 347420 676088 347472
rect 676496 347420 676548 347472
rect 35808 344564 35860 344616
rect 39856 344564 39908 344616
rect 35624 343612 35676 343664
rect 40040 343612 40092 343664
rect 35808 342184 35860 342236
rect 40224 342184 40276 342236
rect 45468 342184 45520 342236
rect 63132 342184 63184 342236
rect 35808 341504 35860 341556
rect 40224 341504 40276 341556
rect 35808 341028 35860 341080
rect 40132 341028 40184 341080
rect 35532 339600 35584 339652
rect 37096 339600 37148 339652
rect 35808 339464 35860 339516
rect 38844 339464 38896 339516
rect 674840 339328 674892 339380
rect 675484 339328 675536 339380
rect 674380 336540 674432 336592
rect 675392 336540 675444 336592
rect 35808 335316 35860 335368
rect 39856 335316 39908 335368
rect 35808 334092 35860 334144
rect 40316 334092 40368 334144
rect 651380 328244 651432 328296
rect 654784 328244 654836 328296
rect 651380 325592 651432 325644
rect 653404 325592 653456 325644
rect 53840 317364 53892 317416
rect 62120 317364 62172 317416
rect 53104 315936 53156 315988
rect 62120 315936 62172 315988
rect 59912 314712 59964 314764
rect 62120 314712 62172 314764
rect 676220 307776 676272 307828
rect 676864 307776 676916 307828
rect 675852 304512 675904 304564
rect 676220 304512 676272 304564
rect 651380 303492 651432 303544
rect 653404 303492 653456 303544
rect 651472 300772 651524 300824
rect 664444 300772 664496 300824
rect 35624 298732 35676 298784
rect 41604 298732 41656 298784
rect 35808 298256 35860 298308
rect 41604 298256 41656 298308
rect 651472 298120 651524 298172
rect 662420 298120 662472 298172
rect 676128 298052 676180 298104
rect 676864 298052 676916 298104
rect 675944 297644 675996 297696
rect 677600 297644 677652 297696
rect 675852 297168 675904 297220
rect 679624 297168 679676 297220
rect 651472 297032 651524 297084
rect 656164 297032 656216 297084
rect 652668 295944 652720 295996
rect 665824 295944 665876 295996
rect 35808 295604 35860 295656
rect 40684 295604 40736 295656
rect 35440 295468 35492 295520
rect 40040 295468 40092 295520
rect 58624 295400 58676 295452
rect 62120 295400 62172 295452
rect 35624 295332 35676 295384
rect 41604 295332 41656 295384
rect 35808 294244 35860 294296
rect 41696 294244 41748 294296
rect 57244 294040 57296 294092
rect 62120 294040 62172 294092
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 35808 292884 35860 292936
rect 41328 292816 41380 292868
rect 35808 292544 35860 292596
rect 39212 292544 39264 292596
rect 54484 292544 54536 292596
rect 62304 292544 62356 292596
rect 651472 292544 651524 292596
rect 663064 292544 663116 292596
rect 46204 292408 46256 292460
rect 62120 292408 62172 292460
rect 40040 291320 40092 291372
rect 41696 291320 41748 291372
rect 42064 291184 42116 291236
rect 42616 291184 42668 291236
rect 53104 291116 53156 291168
rect 62120 291116 62172 291168
rect 35808 289892 35860 289944
rect 41696 289892 41748 289944
rect 42064 289824 42116 289876
rect 43352 289824 43404 289876
rect 651472 289824 651524 289876
rect 660304 289824 660356 289876
rect 35624 289076 35676 289128
rect 41696 289076 41748 289128
rect 55864 288464 55916 288516
rect 62120 288464 62172 288516
rect 651472 288396 651524 288448
rect 661684 288396 661736 288448
rect 651472 287036 651524 287088
rect 672448 287036 672500 287088
rect 674380 286968 674432 287020
rect 675116 286968 675168 287020
rect 33784 286288 33836 286340
rect 41696 286288 41748 286340
rect 46204 285676 46256 285728
rect 62120 285676 62172 285728
rect 651472 285676 651524 285728
rect 672080 285676 672132 285728
rect 60004 284384 60056 284436
rect 62120 284384 62172 284436
rect 651472 284316 651524 284368
rect 672632 284316 672684 284368
rect 651472 282888 651524 282940
rect 667204 282888 667256 282940
rect 42248 281732 42300 281784
rect 42616 281732 42668 281784
rect 47768 280304 47820 280356
rect 62120 280304 62172 280356
rect 651472 280168 651524 280220
rect 667388 280168 667440 280220
rect 42248 280100 42300 280152
rect 42984 280100 43036 280152
rect 482836 277312 482888 277364
rect 557540 277312 557592 277364
rect 485688 277176 485740 277228
rect 562324 277176 562376 277228
rect 495072 277040 495124 277092
rect 576492 277040 576544 277092
rect 511632 276904 511684 276956
rect 600136 276904 600188 276956
rect 42248 276768 42300 276820
rect 42616 276768 42668 276820
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 518716 276632 518768 276684
rect 609612 276632 609664 276684
rect 478512 276496 478564 276548
rect 551652 276496 551704 276548
rect 477040 276360 477092 276412
rect 550456 276360 550508 276412
rect 471612 276224 471664 276276
rect 543372 276224 543424 276276
rect 107200 275952 107252 276004
rect 162124 275952 162176 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 454408 275952 454460 276004
rect 100116 275816 100168 275868
rect 161388 275816 161440 275868
rect 161572 275816 161624 275868
rect 161756 275816 161808 275868
rect 167000 275816 167052 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 217140 275816 217192 275868
rect 224040 275816 224092 275868
rect 232504 275816 232556 275868
rect 239864 275816 239916 275868
rect 284576 275816 284628 275868
rect 290096 275816 290148 275868
rect 445024 275816 445076 275868
rect 457444 275952 457496 276004
rect 509056 275952 509108 276004
rect 517152 275952 517204 276004
rect 608416 275952 608468 276004
rect 93032 275680 93084 275732
rect 155960 275680 156012 275732
rect 163136 275680 163188 275732
rect 164056 275680 164108 275732
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 156880 275544 156932 275596
rect 171048 275680 171100 275732
rect 211068 275680 211120 275732
rect 224224 275680 224276 275732
rect 232780 275680 232832 275732
rect 236092 275680 236144 275732
rect 253388 275680 253440 275732
rect 435640 275680 435692 275732
rect 454408 275680 454460 275732
rect 475384 275816 475436 275868
rect 479524 275816 479576 275868
rect 523316 275816 523368 275868
rect 524144 275816 524196 275868
rect 615500 275816 615552 275868
rect 498476 275680 498528 275732
rect 507860 275680 507912 275732
rect 545764 275680 545816 275732
rect 277492 275612 277544 275664
rect 284300 275612 284352 275664
rect 81256 275408 81308 275460
rect 145564 275408 145616 275460
rect 160468 275408 160520 275460
rect 161848 275408 161900 275460
rect 206376 275544 206428 275596
rect 221924 275544 221976 275596
rect 239404 275544 239456 275596
rect 243176 275544 243228 275596
rect 255320 275544 255372 275596
rect 257344 275544 257396 275596
rect 262864 275544 262916 275596
rect 286876 275544 286928 275596
rect 291844 275544 291896 275596
rect 430212 275544 430264 275596
rect 484308 275544 484360 275596
rect 501604 275544 501656 275596
rect 512644 275544 512696 275596
rect 515404 275544 515456 275596
rect 526812 275544 526864 275596
rect 528192 275544 528244 275596
rect 622584 275544 622636 275596
rect 198740 275408 198792 275460
rect 214840 275408 214892 275460
rect 236644 275408 236696 275460
rect 239588 275408 239640 275460
rect 251916 275408 251968 275460
rect 263232 275408 263284 275460
rect 273260 275408 273312 275460
rect 285680 275408 285732 275460
rect 291200 275408 291252 275460
rect 291660 275408 291712 275460
rect 295432 275408 295484 275460
rect 386052 275408 386104 275460
rect 420460 275408 420512 275460
rect 423404 275408 423456 275460
rect 473360 275408 473412 275460
rect 475384 275408 475436 275460
rect 485044 275408 485096 275460
rect 485228 275408 485280 275460
rect 537484 275408 537536 275460
rect 297548 275340 297600 275392
rect 299572 275340 299624 275392
rect 299940 275340 299992 275392
rect 301136 275340 301188 275392
rect 71780 275272 71832 275324
rect 141056 275272 141108 275324
rect 146208 275272 146260 275324
rect 189080 275272 189132 275324
rect 218336 275272 218388 275324
rect 243084 275272 243136 275324
rect 256148 275272 256200 275324
rect 268660 275272 268712 275324
rect 273904 275272 273956 275324
rect 282920 275272 282972 275324
rect 361212 275272 361264 275324
rect 385040 275272 385092 275324
rect 416412 275272 416464 275324
rect 462964 275272 463016 275324
rect 463148 275272 463200 275324
rect 530400 275272 530452 275324
rect 532332 275272 532384 275324
rect 537300 275272 537352 275324
rect 537576 275272 537628 275324
rect 636752 275408 636804 275460
rect 537944 275272 537996 275324
rect 540980 275272 541032 275324
rect 543004 275272 543056 275324
rect 629668 275272 629720 275324
rect 290464 275204 290516 275256
rect 294144 275204 294196 275256
rect 298744 275204 298796 275256
rect 300032 275204 300084 275256
rect 139124 275136 139176 275188
rect 146944 275136 146996 275188
rect 149796 275136 149848 275188
rect 191748 275136 191800 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 485044 275136 485096 275188
rect 491392 275136 491444 275188
rect 493324 275136 493376 275188
rect 269212 275068 269264 275120
rect 274916 275068 274968 275120
rect 110788 275000 110840 275052
rect 149704 275000 149756 275052
rect 153384 275000 153436 275052
rect 154488 275000 154540 275052
rect 132040 274864 132092 274916
rect 161664 275000 161716 275052
rect 161848 275000 161900 275052
rect 175924 275000 175976 275052
rect 190000 275000 190052 275052
rect 218704 275000 218756 275052
rect 288072 275000 288124 275052
rect 292672 275000 292724 275052
rect 420644 275000 420696 275052
rect 470140 275000 470192 275052
rect 476120 275000 476172 275052
rect 485228 275000 485280 275052
rect 492404 275000 492456 275052
rect 494888 275000 494940 275052
rect 497464 275136 497516 275188
rect 505560 275136 505612 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 501972 275000 502024 275052
rect 503444 275000 503496 275052
rect 587072 275000 587124 275052
rect 293960 274932 294012 274984
rect 296812 274932 296864 274984
rect 167552 274864 167604 274916
rect 169024 274864 169076 274916
rect 289268 274864 289320 274916
rect 293408 274864 293460 274916
rect 413468 274864 413520 274916
rect 459468 274864 459520 274916
rect 473360 274864 473412 274916
rect 544568 274864 544620 274916
rect 103704 274728 103756 274780
rect 104808 274728 104860 274780
rect 74172 274660 74224 274712
rect 76748 274660 76800 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 96620 274524 96672 274576
rect 117688 274592 117740 274644
rect 117872 274592 117924 274644
rect 174636 274796 174688 274848
rect 182732 274796 182784 274848
rect 295156 274796 295208 274848
rect 297456 274796 297508 274848
rect 136824 274728 136876 274780
rect 137652 274728 137704 274780
rect 143908 274728 143960 274780
rect 144368 274728 144420 274780
rect 146944 274728 146996 274780
rect 174452 274728 174504 274780
rect 469864 274728 469916 274780
rect 516232 274728 516284 274780
rect 526444 274728 526496 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 537944 274728 537996 274780
rect 538128 274728 538180 274780
rect 543004 274728 543056 274780
rect 543188 274728 543240 274780
rect 643836 274728 643888 274780
rect 253848 274660 253900 274712
rect 258356 274660 258408 274712
rect 268016 274660 268068 274712
rect 272432 274660 272484 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 292856 274660 292908 274712
rect 295800 274660 295852 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 350724 274660 350776 274712
rect 353116 274660 353168 274712
rect 174176 274592 174228 274644
rect 182916 274592 182968 274644
rect 214564 274592 214616 274644
rect 382924 274592 382976 274644
rect 392124 274592 392176 274644
rect 404176 274592 404228 274644
rect 446496 274592 446548 274644
rect 450544 274592 450596 274644
rect 480720 274592 480772 274644
rect 488356 274592 488408 274644
rect 567016 274592 567068 274644
rect 67088 274320 67140 274372
rect 95884 274456 95936 274508
rect 105176 274456 105228 274508
rect 163320 274456 163372 274508
rect 168748 274456 168800 274508
rect 208492 274456 208544 274508
rect 227812 274456 227864 274508
rect 248880 274456 248932 274508
rect 358084 274456 358136 274508
rect 369584 274456 369636 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 166356 274320 166408 274372
rect 207296 274320 207348 274372
rect 207756 274320 207808 274372
rect 233884 274320 233936 274372
rect 249064 274320 249116 274372
rect 265256 274320 265308 274372
rect 333796 274320 333848 274372
rect 345940 274320 345992 274372
rect 347044 274320 347096 274372
rect 359004 274320 359056 274372
rect 369308 274320 369360 274372
rect 395620 274456 395672 274508
rect 409236 274456 409288 274508
rect 453580 274456 453632 274508
rect 453764 274456 453816 274508
rect 486608 274456 486660 274508
rect 536748 274456 536800 274508
rect 634360 274456 634412 274508
rect 373264 274320 373316 274372
rect 400312 274320 400364 274372
rect 413836 274320 413888 274372
rect 460664 274320 460716 274372
rect 465724 274320 465776 274372
rect 487804 274320 487856 274372
rect 508596 274320 508648 274372
rect 595076 274320 595128 274372
rect 595444 274320 595496 274372
rect 640340 274320 640392 274372
rect 282184 274252 282236 274304
rect 287704 274252 287756 274304
rect 89444 274184 89496 274236
rect 152004 274184 152056 274236
rect 155684 274184 155736 274236
rect 200120 274184 200172 274236
rect 205364 274184 205416 274236
rect 234712 274184 234764 274236
rect 237288 274184 237340 274236
rect 256976 274184 257028 274236
rect 325332 274184 325384 274236
rect 332968 274184 333020 274236
rect 343456 274184 343508 274236
rect 360200 274184 360252 274236
rect 364984 274184 365036 274236
rect 374368 274184 374420 274236
rect 379336 274184 379388 274236
rect 410984 274184 411036 274236
rect 416596 274184 416648 274236
rect 464160 274184 464212 274236
rect 474372 274184 474424 274236
rect 507860 274184 507912 274236
rect 511816 274184 511868 274236
rect 598940 274184 598992 274236
rect 77668 274048 77720 274100
rect 65892 273912 65944 273964
rect 136824 273912 136876 273964
rect 145104 274048 145156 274100
rect 192392 274048 192444 274100
rect 198280 274048 198332 274100
rect 229192 274048 229244 274100
rect 234896 274048 234948 274100
rect 145104 273912 145156 273964
rect 147404 273912 147456 273964
rect 193404 273912 193456 273964
rect 195888 273912 195940 273964
rect 227904 273912 227956 273964
rect 229008 273912 229060 273964
rect 250444 273912 250496 273964
rect 255320 274048 255372 274100
rect 261024 274048 261076 274100
rect 261208 274048 261260 274100
rect 273536 274048 273588 274100
rect 275100 274048 275152 274100
rect 283472 274048 283524 274100
rect 332324 274048 332376 274100
rect 343640 274048 343692 274100
rect 350356 274048 350408 274100
rect 368480 274048 368532 274100
rect 369124 274048 369176 274100
rect 387340 274048 387392 274100
rect 394332 274048 394384 274100
rect 432236 274048 432288 274100
rect 432604 274048 432656 274100
rect 485504 274048 485556 274100
rect 491208 274048 491260 274100
rect 569960 274048 570012 274100
rect 571984 274048 572036 274100
rect 583576 274048 583628 274100
rect 255412 273912 255464 273964
rect 258540 273912 258592 273964
rect 272064 273912 272116 273964
rect 272708 273912 272760 273964
rect 281816 273912 281868 273964
rect 324044 273912 324096 273964
rect 331772 273912 331824 273964
rect 331956 273912 332008 273964
rect 341248 273912 341300 273964
rect 342076 273912 342128 273964
rect 357808 273912 357860 273964
rect 360108 273912 360160 273964
rect 382648 273912 382700 273964
rect 387432 273912 387484 273964
rect 421656 273912 421708 273964
rect 421840 273912 421892 273964
rect 471244 273912 471296 273964
rect 475752 273912 475804 273964
rect 547512 273912 547564 273964
rect 547696 273912 547748 273964
rect 639144 273912 639196 273964
rect 113456 273776 113508 273828
rect 169944 273776 169996 273828
rect 175924 273776 175976 273828
rect 204260 273776 204312 273828
rect 206560 273776 206612 273828
rect 235448 273776 235500 273828
rect 400128 273776 400180 273828
rect 439320 273776 439372 273828
rect 442264 273776 442316 273828
rect 481916 273776 481968 273828
rect 487068 273776 487120 273828
rect 123760 273640 123812 273692
rect 177488 273640 177540 273692
rect 392584 273640 392636 273692
rect 409788 273640 409840 273692
rect 440884 273640 440936 273692
rect 474832 273640 474884 273692
rect 484308 273640 484360 273692
rect 552664 273640 552716 273692
rect 552848 273640 552900 273692
rect 562232 273640 562284 273692
rect 562600 273776 562652 273828
rect 571984 273776 572036 273828
rect 563428 273640 563480 273692
rect 563704 273640 563756 273692
rect 597744 273776 597796 273828
rect 134432 273504 134484 273556
rect 185124 273504 185176 273556
rect 446404 273504 446456 273556
rect 475936 273504 475988 273556
rect 481364 273504 481416 273556
rect 556344 273504 556396 273556
rect 556804 273504 556856 273556
rect 590660 273504 590712 273556
rect 135628 273368 135680 273420
rect 146944 273368 146996 273420
rect 460020 273368 460072 273420
rect 465724 273368 465776 273420
rect 467564 273368 467616 273420
rect 476120 273368 476172 273420
rect 478696 273368 478748 273420
rect 552480 273368 552532 273420
rect 552664 273368 552716 273420
rect 559932 273368 559984 273420
rect 374644 273300 374696 273352
rect 377864 273300 377916 273352
rect 453304 273300 453356 273352
rect 453764 273300 453816 273352
rect 318708 273232 318760 273284
rect 324688 273232 324740 273284
rect 327540 273232 327592 273284
rect 329472 273232 329524 273284
rect 114376 273164 114428 273216
rect 171600 273164 171652 273216
rect 184112 273164 184164 273216
rect 218888 273164 218940 273216
rect 366364 273164 366416 273216
rect 383844 273164 383896 273216
rect 401508 273164 401560 273216
rect 442908 273164 442960 273216
rect 452292 273164 452344 273216
rect 515036 273164 515088 273216
rect 515220 273164 515272 273216
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 278596 273096 278648 273148
rect 285864 273096 285916 273148
rect 101312 273028 101364 273080
rect 160192 273028 160244 273080
rect 172244 273028 172296 273080
rect 210608 273028 210660 273080
rect 224040 273028 224092 273080
rect 243268 273028 243320 273080
rect 329472 273028 329524 273080
rect 338856 273028 338908 273080
rect 349804 273028 349856 273080
rect 366088 273028 366140 273080
rect 377404 273028 377456 273080
rect 399208 273028 399260 273080
rect 408224 273028 408276 273080
rect 450820 273028 450872 273080
rect 451188 273028 451240 273080
rect 513840 273028 513892 273080
rect 526812 273028 526864 273080
rect 621388 273028 621440 273080
rect 99012 272892 99064 272944
rect 160376 272892 160428 272944
rect 162768 272892 162820 272944
rect 204720 272892 204772 272944
rect 219532 272892 219584 272944
rect 244464 272892 244516 272944
rect 251456 272892 251508 272944
rect 267004 272892 267056 272944
rect 335268 272892 335320 272944
rect 346860 272892 346912 272944
rect 362776 272892 362828 272944
rect 385868 272892 385920 272944
rect 406844 272892 406896 272944
rect 449992 272892 450044 272944
rect 455236 272892 455288 272944
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 158076 272756 158128 272808
rect 200672 272756 200724 272808
rect 208860 272756 208912 272808
rect 237380 272756 237432 272808
rect 252652 272756 252704 272808
rect 72976 272620 73028 272672
rect 142160 272620 142212 272672
rect 152188 272620 152240 272672
rect 197544 272620 197596 272672
rect 199476 272620 199528 272672
rect 230572 272620 230624 272672
rect 233700 272620 233752 272672
rect 253940 272620 253992 272672
rect 69388 272484 69440 272536
rect 139400 272484 139452 272536
rect 141516 272484 141568 272536
rect 120264 272348 120316 272400
rect 175280 272348 175332 272400
rect 189080 272484 189132 272536
rect 194048 272484 194100 272536
rect 194692 272484 194744 272536
rect 227168 272484 227220 272536
rect 238484 272484 238536 272536
rect 258080 272484 258132 272536
rect 271512 272756 271564 272808
rect 280344 272756 280396 272808
rect 336372 272756 336424 272808
rect 349528 272756 349580 272808
rect 352564 272756 352616 272808
rect 370780 272756 370832 272808
rect 375196 272756 375248 272808
rect 403900 272756 403952 272808
rect 412272 272756 412324 272808
rect 457076 272756 457128 272808
rect 458088 272892 458140 272944
rect 463332 272892 463384 272944
rect 518532 272892 518584 272944
rect 529848 272892 529900 272944
rect 624976 272892 625028 272944
rect 463884 272756 463936 272808
rect 522120 272756 522172 272808
rect 522764 272756 522816 272808
rect 524144 272756 524196 272808
rect 532516 272756 532568 272808
rect 628472 272756 628524 272808
rect 266820 272620 266872 272672
rect 277584 272620 277636 272672
rect 280988 272620 281040 272672
rect 286324 272620 286376 272672
rect 322756 272620 322808 272672
rect 330576 272620 330628 272672
rect 338028 272620 338080 272672
rect 351920 272620 351972 272672
rect 354496 272620 354548 272672
rect 375564 272620 375616 272672
rect 382004 272620 382056 272672
rect 414572 272620 414624 272672
rect 419172 272620 419224 272672
rect 467380 272620 467432 272672
rect 467748 272620 467800 272672
rect 470416 272620 470468 272672
rect 470600 272620 470652 272672
rect 536288 272620 536340 272672
rect 536564 272620 536616 272672
rect 635556 272620 635608 272672
rect 267924 272484 267976 272536
rect 325516 272484 325568 272536
rect 334164 272484 334216 272536
rect 344652 272484 344704 272536
rect 361396 272484 361448 272536
rect 363788 272484 363840 272536
rect 388536 272484 388588 272536
rect 397276 272484 397328 272536
rect 435824 272484 435876 272536
rect 438768 272484 438820 272536
rect 489874 272484 489926 272536
rect 490012 272484 490064 272536
rect 529204 272484 529256 272536
rect 533712 272484 533764 272536
rect 632060 272484 632112 272536
rect 189172 272348 189224 272400
rect 193588 272348 193640 272400
rect 224224 272348 224276 272400
rect 264428 272348 264480 272400
rect 276020 272348 276072 272400
rect 388996 272348 389048 272400
rect 425152 272348 425204 272400
rect 449716 272348 449768 272400
rect 511448 272348 511500 272400
rect 512644 272348 512696 272400
rect 515220 272348 515272 272400
rect 517336 272348 517388 272400
rect 607220 272348 607272 272400
rect 119068 272212 119120 272264
rect 173256 272212 173308 272264
rect 174452 272212 174504 272264
rect 189356 272212 189408 272264
rect 446956 272212 447008 272264
rect 508044 272212 508096 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 130844 272076 130896 272128
rect 182456 272076 182508 272128
rect 426348 272076 426400 272128
rect 470554 272076 470606 272128
rect 470784 272076 470836 272128
rect 489874 272076 489926 272128
rect 490012 272076 490064 272128
rect 558736 272076 558788 272128
rect 191472 271940 191524 271992
rect 108396 271804 108448 271856
rect 165896 271804 165948 271856
rect 188804 271804 188856 271856
rect 192576 271804 192628 271856
rect 447784 271940 447836 271992
rect 506756 271940 506808 271992
rect 507124 271940 507176 271992
rect 569408 271940 569460 271992
rect 268660 271872 268712 271924
rect 270500 271872 270552 271924
rect 225052 271804 225104 271856
rect 225420 271804 225472 271856
rect 228364 271804 228416 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 376576 271804 376628 271856
rect 407488 271804 407540 271856
rect 407764 271804 407816 271856
rect 437020 271804 437072 271856
rect 437204 271804 437256 271856
rect 493692 271804 493744 271856
rect 496544 271804 496596 271856
rect 578516 271804 578568 271856
rect 578884 271804 578936 271856
rect 611912 271804 611964 271856
rect 106096 271668 106148 271720
rect 164976 271668 165028 271720
rect 175740 271668 175792 271720
rect 213000 271668 213052 271720
rect 239864 271668 239916 271720
rect 254124 271668 254176 271720
rect 353944 271668 353996 271720
rect 372804 271668 372856 271720
rect 384948 271668 385000 271720
rect 418068 271668 418120 271720
rect 420184 271668 420236 271720
rect 431132 271668 431184 271720
rect 434628 271668 434680 271720
rect 485228 271668 485280 271720
rect 485412 271668 485464 271720
rect 490012 271668 490064 271720
rect 501972 271668 502024 271720
rect 585968 271668 586020 271720
rect 94228 271532 94280 271584
rect 156144 271532 156196 271584
rect 170128 271532 170180 271584
rect 209780 271532 209832 271584
rect 223120 271532 223172 271584
rect 247224 271532 247276 271584
rect 357164 271532 357216 271584
rect 379060 271532 379112 271584
rect 387616 271532 387668 271584
rect 422852 271532 422904 271584
rect 439964 271532 440016 271584
rect 497280 271532 497332 271584
rect 499304 271532 499356 271584
rect 582380 271532 582432 271584
rect 585784 271532 585836 271584
rect 626080 271532 626132 271584
rect 87144 271396 87196 271448
rect 152188 271396 152240 271448
rect 159272 271396 159324 271448
rect 202328 271396 202380 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 250260 271396 250312 271448
rect 75368 271260 75420 271312
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 142712 271260 142764 271312
rect 144184 271260 144236 271312
rect 154304 271260 154356 271312
rect 198096 271260 198148 271312
rect 212264 271260 212316 271312
rect 239312 271260 239364 271312
rect 244648 271260 244700 271312
rect 262220 271260 262272 271312
rect 265624 271396 265676 271448
rect 276848 271396 276900 271448
rect 329656 271396 329708 271448
rect 340052 271396 340104 271448
rect 340604 271396 340656 271448
rect 355140 271396 355192 271448
rect 358728 271396 358780 271448
rect 381452 271396 381504 271448
rect 393964 271396 394016 271448
rect 429936 271396 429988 271448
rect 442908 271396 442960 271448
rect 500868 271396 500920 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 266452 271260 266504 271312
rect 276664 271260 276716 271312
rect 284484 271260 284536 271312
rect 326436 271260 326488 271312
rect 335084 271260 335136 271312
rect 339408 271260 339460 271312
rect 354220 271260 354272 271312
rect 365444 271260 365496 271312
rect 390928 271260 390980 271312
rect 391848 271260 391900 271312
rect 428740 271260 428792 271312
rect 445668 271260 445720 271312
rect 504364 271260 504416 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 612004 271260 612056 271312
rect 618628 271260 618680 271312
rect 618904 271260 618956 271312
rect 633256 271260 633308 271312
rect 142712 271124 142764 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 197084 271124 197136 271176
rect 229284 271124 229336 271176
rect 230204 271124 230256 271176
rect 251732 271124 251784 271176
rect 254952 271124 255004 271176
rect 269304 271124 269356 271176
rect 270316 271124 270368 271176
rect 280528 271124 280580 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 347596 271124 347648 271176
rect 364524 271124 364576 271176
rect 366916 271124 366968 271176
rect 393320 271124 393372 271176
rect 402612 271124 402664 271176
rect 444104 271124 444156 271176
rect 459468 271124 459520 271176
rect 523868 271124 523920 271176
rect 524052 271124 524104 271176
rect 617800 271124 617852 271176
rect 625804 271124 625856 271176
rect 645032 271124 645084 271176
rect 116676 270988 116728 271040
rect 172520 270988 172572 271040
rect 192760 270988 192812 271040
rect 225512 270988 225564 271040
rect 381544 270988 381596 271040
rect 411812 270988 411864 271040
rect 414480 270988 414532 271040
rect 438124 270988 438176 271040
rect 438308 270988 438360 271040
rect 124956 270852 125008 270904
rect 178684 270852 178736 270904
rect 417424 270852 417476 270904
rect 427544 270852 427596 270904
rect 430396 270852 430448 270904
rect 483112 270852 483164 270904
rect 485228 270988 485280 271040
rect 490196 270988 490248 271040
rect 495256 270988 495308 271040
rect 575296 270988 575348 271040
rect 492404 270852 492456 270904
rect 492588 270852 492640 270904
rect 571708 270852 571760 270904
rect 571984 270852 572036 270904
rect 604828 270852 604880 270904
rect 127348 270716 127400 270768
rect 179880 270716 179932 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 427452 270716 427504 270768
rect 479156 270716 479208 270768
rect 486884 270716 486936 270768
rect 564624 270716 564676 270768
rect 137928 270580 137980 270632
rect 187700 270580 187752 270632
rect 422944 270580 422996 270632
rect 445300 270580 445352 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 129464 270444 129516 270496
rect 181168 270444 181220 270496
rect 191748 270444 191800 270496
rect 196900 270444 196952 270496
rect 201776 270444 201828 270496
rect 232228 270444 232280 270496
rect 395620 270444 395672 270496
rect 433616 270444 433668 270496
rect 453580 270444 453632 270496
rect 516784 270444 516836 270496
rect 517520 270444 517572 270496
rect 579620 270444 579672 270496
rect 581644 270444 581696 270496
rect 620284 270444 620336 270496
rect 88340 270308 88392 270360
rect 121460 270308 121512 270360
rect 122472 270308 122524 270360
rect 176200 270308 176252 270360
rect 180708 270308 180760 270360
rect 215300 270308 215352 270360
rect 232780 270308 232832 270360
rect 247868 270308 247920 270360
rect 262864 270308 262916 270360
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 179328 270172 179380 270224
rect 214104 270172 214156 270224
rect 226616 270172 226668 270224
rect 249892 270172 249944 270224
rect 259736 270172 259788 270224
rect 367468 270308 367520 270360
rect 393504 270308 393556 270360
rect 400864 270308 400916 270360
rect 441620 270308 441672 270360
rect 456064 270308 456116 270360
rect 520280 270308 520332 270360
rect 85488 270036 85540 270088
rect 149428 270036 149480 270088
rect 173716 270036 173768 270088
rect 212632 270036 212684 270088
rect 216496 270036 216548 270088
rect 242440 270036 242492 270088
rect 248328 270036 248380 270088
rect 264796 270036 264848 270088
rect 70584 269900 70636 269952
rect 79968 269900 80020 269952
rect 80152 269900 80204 269952
rect 146392 269900 146444 269952
rect 165436 269900 165488 269952
rect 206008 269900 206060 269952
rect 210056 269900 210108 269952
rect 238300 269900 238352 269952
rect 241980 269900 242032 269952
rect 260380 269900 260432 269952
rect 271420 270172 271472 270224
rect 345112 270172 345164 270224
rect 361580 270172 361632 270224
rect 364156 270172 364208 270224
rect 389180 270172 389232 270224
rect 390100 270172 390152 270224
rect 405740 270172 405792 270224
rect 409696 270172 409748 270224
rect 454040 270172 454092 270224
rect 458548 270172 458600 270224
rect 524420 270308 524472 270360
rect 525616 270308 525668 270360
rect 523132 270172 523184 270224
rect 533160 270172 533212 270224
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 619640 270172 619692 270224
rect 327724 270036 327776 270088
rect 336740 270036 336792 270088
rect 345940 270036 345992 270088
rect 362960 270036 363012 270088
rect 369952 270036 370004 270088
rect 396080 270036 396132 270088
rect 399944 270036 399996 270088
rect 412640 270036 412692 270088
rect 414664 270036 414716 270088
rect 460940 270036 460992 270088
rect 461400 270036 461452 270088
rect 527180 270036 527232 270088
rect 528376 270036 528428 270088
rect 623964 270172 624016 270224
rect 620284 270036 620336 270088
rect 630680 270036 630732 270088
rect 273076 269900 273128 269952
rect 335084 269900 335136 269952
rect 347780 269900 347832 269952
rect 351736 269900 351788 269952
rect 371240 269900 371292 269952
rect 372436 269900 372488 269952
rect 400496 269900 400548 269952
rect 401876 269900 401928 269952
rect 416780 269900 416832 269952
rect 417148 269900 417200 269952
rect 465080 269900 465132 269952
rect 468484 269900 468536 269952
rect 76748 269764 76800 269816
rect 143908 269764 143960 269816
rect 144368 269764 144420 269816
rect 190828 269764 190880 269816
rect 202972 269764 203024 269816
rect 233332 269764 233384 269816
rect 241428 269764 241480 269816
rect 259828 269764 259880 269816
rect 261944 269764 261996 269816
rect 274732 269764 274784 269816
rect 280068 269764 280120 269816
rect 287152 269764 287204 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336832 269764 336884 269816
rect 350540 269764 350592 269816
rect 355048 269764 355100 269816
rect 376944 269764 376996 269816
rect 377680 269764 377732 269816
rect 408500 269764 408552 269816
rect 412456 269764 412508 269816
rect 458272 269764 458324 269816
rect 463516 269764 463568 269816
rect 531320 269764 531372 269816
rect 531964 269900 532016 269952
rect 533528 269900 533580 269952
rect 533988 269900 534040 269952
rect 537760 269900 537812 269952
rect 537944 269900 537996 269952
rect 538496 269764 538548 269816
rect 538680 269764 538732 269816
rect 542820 269764 542872 269816
rect 543188 269900 543240 269952
rect 640524 269900 640576 269952
rect 637580 269764 637632 269816
rect 126888 269628 126940 269680
rect 178316 269628 178368 269680
rect 200488 269628 200540 269680
rect 226892 269628 226944 269680
rect 384764 269628 384816 269680
rect 418252 269628 418304 269680
rect 422116 269628 422168 269680
rect 471980 269628 472032 269680
rect 472624 269628 472676 269680
rect 473360 269628 473412 269680
rect 78864 269492 78916 269544
rect 130384 269492 130436 269544
rect 133788 269492 133840 269544
rect 183652 269492 183704 269544
rect 186412 269492 186464 269544
rect 204076 269492 204128 269544
rect 392032 269492 392084 269544
rect 401692 269492 401744 269544
rect 404544 269492 404596 269544
rect 423680 269492 423732 269544
rect 432236 269492 432288 269544
rect 466460 269492 466512 269544
rect 530400 269628 530452 269680
rect 530584 269628 530636 269680
rect 531964 269628 532016 269680
rect 533160 269628 533212 269680
rect 616144 269628 616196 269680
rect 140688 269356 140740 269408
rect 188620 269356 188672 269408
rect 429108 269356 429160 269408
rect 455420 269356 455472 269408
rect 466000 269356 466052 269408
rect 509056 269492 509108 269544
rect 596180 269492 596232 269544
rect 474648 269356 474700 269408
rect 538128 269356 538180 269408
rect 538312 269356 538364 269408
rect 581644 269356 581696 269408
rect 121644 269220 121696 269272
rect 167828 269220 167880 269272
rect 272432 269220 272484 269272
rect 278872 269220 278924 269272
rect 423956 269220 424008 269272
rect 448520 269220 448572 269272
rect 470968 269220 471020 269272
rect 540612 269220 540664 269272
rect 540796 269220 540848 269272
rect 543188 269220 543240 269272
rect 543372 269152 543424 269204
rect 546500 269152 546552 269204
rect 274916 269084 274968 269136
rect 279700 269084 279752 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 42156 269016 42208 269068
rect 43168 269016 43220 269068
rect 84108 269016 84160 269068
rect 137468 269016 137520 269068
rect 137652 269016 137704 269068
rect 186136 269016 186188 269068
rect 379704 269016 379756 269068
rect 404360 269016 404412 269068
rect 436192 269016 436244 269068
rect 491760 269016 491812 269068
rect 498292 269016 498344 269068
rect 581000 269016 581052 269068
rect 273260 268948 273312 269000
rect 275560 268948 275612 269000
rect 111984 268880 112036 268932
rect 168748 268880 168800 268932
rect 382372 268880 382424 268932
rect 415400 268880 415452 268932
rect 433708 268880 433760 268932
rect 488540 268880 488592 268932
rect 500776 268880 500828 268932
rect 583760 268880 583812 268932
rect 115848 268744 115900 268796
rect 110236 268608 110288 268660
rect 102508 268472 102560 268524
rect 162952 268472 163004 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 211344 268744 211396 268796
rect 223488 268744 223540 268796
rect 389824 268744 389876 268796
rect 425336 268744 425388 268796
rect 441160 268744 441212 268796
rect 499580 268744 499632 268796
rect 505744 268744 505796 268796
rect 590844 268744 590896 268796
rect 167000 268608 167052 268660
rect 184480 268608 184532 268660
rect 187332 268608 187384 268660
rect 219440 268608 219492 268660
rect 245568 268608 245620 268660
rect 263140 268608 263192 268660
rect 396172 268608 396224 268660
rect 433340 268608 433392 268660
rect 443644 268608 443696 268660
rect 502340 268608 502392 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 171232 268472 171284 268524
rect 176936 268472 176988 268524
rect 215116 268472 215168 268524
rect 220452 268472 220504 268524
rect 245752 268472 245804 268524
rect 338488 268472 338540 268524
rect 350724 268472 350776 268524
rect 359832 268472 359884 268524
rect 379520 268472 379572 268524
rect 403256 268472 403308 268524
rect 440240 268472 440292 268524
rect 448612 268472 448664 268524
rect 509240 268472 509292 268524
rect 513196 268472 513248 268524
rect 601700 268472 601752 268524
rect 167644 268336 167696 268388
rect 168012 268336 168064 268388
rect 203524 268336 203576 268388
rect 203892 268336 203944 268388
rect 230756 268336 230808 268388
rect 231676 268336 231728 268388
rect 253204 268336 253256 268388
rect 258356 268336 258408 268388
rect 268936 268336 268988 268388
rect 348424 268336 348476 268388
rect 367100 268336 367152 268388
rect 372160 268336 372212 268388
rect 397460 268336 397512 268388
rect 408040 268336 408092 268388
rect 451372 268336 451424 268388
rect 464344 268336 464396 268388
rect 532700 268336 532752 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 128544 268200 128596 268252
rect 150440 268200 150492 268252
rect 151728 268200 151780 268252
rect 196072 268200 196124 268252
rect 419632 268200 419684 268252
rect 467932 268200 467984 268252
rect 493600 268200 493652 268252
rect 574100 268200 574152 268252
rect 163136 268064 163188 268116
rect 168012 268064 168064 268116
rect 412640 268064 412692 268116
rect 447140 268064 447192 268116
rect 495808 268064 495860 268116
rect 576860 268064 576912 268116
rect 198740 267792 198792 267844
rect 201868 267792 201920 267844
rect 117688 267656 117740 267708
rect 159640 267656 159692 267708
rect 167828 267656 167880 267708
rect 177028 267656 177080 267708
rect 181996 267656 182048 267708
rect 95884 267520 95936 267572
rect 138112 267520 138164 267572
rect 150440 267520 150492 267572
rect 181996 267520 182048 267572
rect 182732 267656 182784 267708
rect 214288 267656 214340 267708
rect 378232 267656 378284 267708
rect 392584 267656 392636 267708
rect 398104 267656 398156 267708
rect 414480 267656 414532 267708
rect 423772 267656 423824 267708
rect 440884 267656 440936 267708
rect 450268 267656 450320 267708
rect 501604 267656 501656 267708
rect 514852 267656 514904 267708
rect 571984 267656 572036 267708
rect 219256 267520 219308 267572
rect 340972 267520 341024 267572
rect 355324 267520 355376 267572
rect 362500 267520 362552 267572
rect 369124 267520 369176 267572
rect 370780 267520 370832 267572
rect 377404 267520 377456 267572
rect 380716 267520 380768 267572
rect 399944 267520 399996 267572
rect 410524 267520 410576 267572
rect 429108 267520 429160 267572
rect 445300 267520 445352 267572
rect 497464 267520 497516 267572
rect 504824 267520 504876 267572
rect 517520 267520 517572 267572
rect 529664 267520 529716 267572
rect 585784 267520 585836 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 146944 267384 146996 267436
rect 186964 267384 187016 267436
rect 236644 267384 236696 267436
rect 241612 267384 241664 267436
rect 315304 267384 315356 267436
rect 319168 267384 319220 267436
rect 350080 267384 350132 267436
rect 358084 267384 358136 267436
rect 371608 267384 371660 267436
rect 373264 267384 373316 267436
rect 383200 267384 383252 267436
rect 401876 267384 401928 267436
rect 405556 267384 405608 267436
rect 423956 267384 424008 267436
rect 432052 267384 432104 267436
rect 453304 267384 453356 267436
rect 460204 267384 460256 267436
rect 515404 267384 515456 267436
rect 519820 267384 519872 267436
rect 578884 267384 578936 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 169024 267248 169076 267300
rect 209320 267248 209372 267300
rect 218704 267248 218756 267300
rect 223028 267248 223080 267300
rect 223488 267248 223540 267300
rect 239128 267248 239180 267300
rect 353392 267248 353444 267300
rect 364984 267248 365036 267300
rect 373264 267248 373316 267300
rect 392032 267248 392084 267300
rect 403072 267248 403124 267300
rect 422944 267248 422996 267300
rect 424600 267248 424652 267300
rect 446404 267248 446456 267300
rect 448152 267248 448204 267300
rect 457444 267248 457496 267300
rect 470140 267248 470192 267300
rect 534724 267248 534776 267300
rect 543004 267248 543056 267300
rect 625804 267248 625856 267300
rect 79968 267112 80020 267164
rect 140596 267112 140648 267164
rect 144184 267112 144236 267164
rect 191932 267112 191984 267164
rect 192576 267112 192628 267164
rect 223948 267112 224000 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 317788 267112 317840 267164
rect 322940 267112 322992 267164
rect 365812 267112 365864 267164
rect 382924 267112 382976 267164
rect 390652 267112 390704 267164
rect 417424 267112 417476 267164
rect 417976 267112 418028 267164
rect 432236 267112 432288 267164
rect 432880 267112 432932 267164
rect 460020 267112 460072 267164
rect 465172 267112 465224 267164
rect 526444 267112 526496 267164
rect 534724 267112 534776 267164
rect 618904 267112 618956 267164
rect 90364 266976 90416 267028
rect 151360 266976 151412 267028
rect 154488 266976 154540 267028
rect 199384 266976 199436 267028
rect 218888 266976 218940 267028
rect 220084 266976 220136 267028
rect 228364 266976 228416 267028
rect 121460 266840 121512 266892
rect 144920 266840 144972 266892
rect 145380 266840 145432 266892
rect 150532 266840 150584 266892
rect 204076 266840 204128 266892
rect 220912 266840 220964 266892
rect 314476 266976 314528 267028
rect 318984 266976 319036 267028
rect 355876 266976 355928 267028
rect 374644 266976 374696 267028
rect 375748 266976 375800 267028
rect 390100 266976 390152 267028
rect 393136 266976 393188 267028
rect 420184 266976 420236 267028
rect 431224 266976 431276 267028
rect 432604 266976 432656 267028
rect 249064 266840 249116 266892
rect 286324 266840 286376 266892
rect 287980 266840 288032 266892
rect 313648 266840 313700 266892
rect 317420 266840 317472 266892
rect 321928 266840 321980 266892
rect 327540 266840 327592 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 392308 266840 392360 266892
rect 393964 266840 394016 266892
rect 427912 266840 427964 266892
rect 450544 266976 450596 267028
rect 455052 266976 455104 267028
rect 512644 266976 512696 267028
rect 524788 266976 524840 267028
rect 612004 266976 612056 267028
rect 442724 266840 442776 266892
rect 493324 266840 493376 266892
rect 497464 266840 497516 266892
rect 517704 266840 517756 266892
rect 518992 266840 519044 266892
rect 520096 266840 520148 266892
rect 527272 266840 527324 266892
rect 528192 266840 528244 266892
rect 528928 266840 528980 266892
rect 529848 266840 529900 266892
rect 531412 266840 531464 266892
rect 532516 266840 532568 266892
rect 533068 266840 533120 266892
rect 533988 266840 534040 266892
rect 535552 266840 535604 266892
rect 536748 266840 536800 266892
rect 539692 266840 539744 266892
rect 595444 266840 595496 266892
rect 130384 266704 130436 266756
rect 147220 266704 147272 266756
rect 149704 266704 149756 266756
rect 169576 266704 169628 266756
rect 230756 266704 230808 266756
rect 234160 266704 234212 266756
rect 252008 266704 252060 266756
rect 259000 266704 259052 266756
rect 359648 266704 359700 266756
rect 366364 266704 366416 266756
rect 388168 266704 388220 266756
rect 214564 266636 214616 266688
rect 218428 266636 218480 266688
rect 308680 266636 308732 266688
rect 310612 266636 310664 266688
rect 312360 266636 312412 266688
rect 314660 266636 314712 266688
rect 316960 266636 317012 266688
rect 321560 266636 321612 266688
rect 342628 266636 342680 266688
rect 347044 266636 347096 266688
rect 137468 266568 137520 266620
rect 145380 266568 145432 266620
rect 145564 266568 145616 266620
rect 148048 266568 148100 266620
rect 226892 266568 226944 266620
rect 231676 266568 231728 266620
rect 397092 266704 397144 266756
rect 407764 266704 407816 266756
rect 428740 266704 428792 266756
rect 442264 266704 442316 266756
rect 457720 266704 457772 266756
rect 479524 266704 479576 266756
rect 490012 266704 490064 266756
rect 507124 266704 507176 266756
rect 509884 266704 509936 266756
rect 563704 266704 563756 266756
rect 404544 266568 404596 266620
rect 404728 266568 404780 266620
rect 412640 266568 412692 266620
rect 440332 266568 440384 266620
rect 445024 266568 445076 266620
rect 452752 266568 452804 266620
rect 469864 266568 469916 266620
rect 499948 266568 500000 266620
rect 214104 266500 214156 266552
rect 215944 266500 215996 266552
rect 248880 266500 248932 266552
rect 250720 266500 250772 266552
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312820 266500 312872 266552
rect 316040 266500 316092 266552
rect 316408 266500 316460 266552
rect 320180 266500 320232 266552
rect 347412 266500 347464 266552
rect 349804 266500 349856 266552
rect 350908 266500 350960 266552
rect 352564 266500 352616 266552
rect 357532 266500 357584 266552
rect 359832 266500 359884 266552
rect 369124 266500 369176 266552
rect 369952 266500 370004 266552
rect 374920 266500 374972 266552
rect 379704 266500 379756 266552
rect 482560 266500 482612 266552
rect 485044 266500 485096 266552
rect 144920 266432 144972 266484
rect 153844 266432 153896 266484
rect 491668 266432 491720 266484
rect 492588 266432 492640 266484
rect 494152 266432 494204 266484
rect 495256 266432 495308 266484
rect 502432 266432 502484 266484
rect 503444 266432 503496 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 510712 266568 510764 266620
rect 511816 266568 511868 266620
rect 516508 266568 516560 266620
rect 517336 266568 517388 266620
rect 517520 266568 517572 266620
rect 556804 266568 556856 266620
rect 549904 266432 549956 266484
rect 162124 266364 162176 266416
rect 167092 266364 167144 266416
rect 178684 266364 178736 266416
rect 179512 266364 179564 266416
rect 215300 266364 215352 266416
rect 217600 266364 217652 266416
rect 219440 266364 219492 266416
rect 222568 266364 222620 266416
rect 224224 266364 224276 266416
rect 226708 266364 226760 266416
rect 233884 266364 233936 266416
rect 236644 266364 236696 266416
rect 239588 266364 239640 266416
rect 246580 266364 246632 266416
rect 250444 266364 250496 266416
rect 251548 266364 251600 266416
rect 253388 266364 253440 266416
rect 256516 266364 256568 266416
rect 287704 266364 287756 266416
rect 288808 266364 288860 266416
rect 300952 266364 301004 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310980 266364 311032 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329472 266364 329524 266416
rect 330208 266364 330260 266416
rect 331956 266364 332008 266416
rect 334348 266364 334400 266416
rect 335268 266364 335320 266416
rect 346768 266364 346820 266416
rect 347596 266364 347648 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 352564 266364 352616 266416
rect 353944 266364 353996 266416
rect 359188 266364 359240 266416
rect 360108 266364 360160 266416
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 368296 266364 368348 266416
rect 369308 266364 369360 266416
rect 369952 266364 370004 266416
rect 372160 266364 372212 266416
rect 374092 266364 374144 266416
rect 375196 266364 375248 266416
rect 379888 266364 379940 266416
rect 381544 266364 381596 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387432 266364 387484 266416
rect 394792 266364 394844 266416
rect 396172 266364 396224 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 400128 266228 400180 266280
rect 403256 266364 403308 266416
rect 407212 266364 407264 266416
rect 408224 266364 408276 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 446128 266364 446180 266416
rect 447784 266364 447836 266416
rect 454408 266364 454460 266416
rect 455236 266364 455288 266416
rect 456892 266364 456944 266416
rect 458088 266364 458140 266416
rect 466828 266364 466880 266416
rect 467748 266364 467800 266416
rect 473452 266364 473504 266416
rect 474372 266364 474424 266416
rect 477592 266364 477644 266416
rect 478512 266364 478564 266416
rect 481732 266364 481784 266416
rect 482836 266364 482888 266416
rect 483388 266364 483440 266416
rect 484308 266364 484360 266416
rect 485872 266364 485924 266416
rect 487068 266364 487120 266416
rect 484216 266228 484268 266280
rect 560484 266296 560536 266348
rect 487528 266160 487580 266212
rect 565820 266160 565872 266212
rect 492496 266024 492548 266076
rect 572720 266024 572772 266076
rect 674472 265956 674524 266008
rect 675484 265956 675536 266008
rect 512368 265888 512420 265940
rect 600320 265888 600372 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 152004 265616 152056 265668
rect 152740 265616 152792 265668
rect 155960 265616 156012 265668
rect 156788 265616 156840 265668
rect 160192 265616 160244 265668
rect 161020 265616 161072 265668
rect 189172 265616 189224 265668
rect 189908 265616 189960 265668
rect 229100 265616 229152 265668
rect 229652 265616 229704 265668
rect 243084 265616 243136 265668
rect 243820 265616 243872 265668
rect 253940 265616 253992 265668
rect 254492 265616 254544 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 520648 265616 520700 265668
rect 612740 265616 612792 265668
rect 480076 265480 480128 265532
rect 554780 265480 554832 265532
rect 479248 265344 479300 265396
rect 553400 265344 553452 265396
rect 475108 265208 475160 265260
rect 547880 265208 547932 265260
rect 469312 265072 469364 265124
rect 539968 265072 540020 265124
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 675852 259564 675904 259616
rect 676220 259564 676272 259616
rect 554320 259428 554372 259480
rect 560944 259428 560996 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 563704 256708 563756 256760
rect 553492 255552 553544 255604
rect 555424 255552 555476 255604
rect 35808 255348 35860 255400
rect 39764 255348 39816 255400
rect 675852 254668 675904 254720
rect 683028 254668 683080 254720
rect 35808 254056 35860 254108
rect 39212 254056 39264 254108
rect 675852 253852 675904 253904
rect 681004 253852 681056 253904
rect 35808 252696 35860 252748
rect 41420 252696 41472 252748
rect 35624 252560 35676 252612
rect 40316 252560 40368 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 35808 251336 35860 251388
rect 41696 251336 41748 251388
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 35808 249908 35860 249960
rect 39672 249908 39724 249960
rect 35808 248616 35860 248668
rect 41512 248616 41564 248668
rect 674840 248072 674892 248124
rect 675300 247936 675352 247988
rect 35808 247188 35860 247240
rect 41696 247188 41748 247240
rect 35624 247052 35676 247104
rect 39856 247052 39908 247104
rect 558184 246304 558236 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 554504 244264 554556 244316
rect 573364 244264 573416 244316
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 674840 239912 674892 239964
rect 675208 239912 675260 239964
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 668768 237396 668820 237448
rect 671620 237396 671672 237448
rect 672172 236784 672224 236836
rect 671620 236580 671672 236632
rect 672954 236648 673006 236700
rect 671804 236376 671856 236428
rect 673184 236240 673236 236292
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 670148 235900 670200 235952
rect 672172 235900 672224 235952
rect 670976 235764 671028 235816
rect 673276 235900 673328 235952
rect 673000 235696 673052 235748
rect 673092 235492 673144 235544
rect 669596 235288 669648 235340
rect 668216 234880 668268 234932
rect 661684 234608 661736 234660
rect 673644 234744 673696 234796
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 668400 234472 668452 234524
rect 671160 234336 671212 234388
rect 671160 234200 671212 234252
rect 674196 234200 674248 234252
rect 675116 234064 675168 234116
rect 675852 233928 675904 233980
rect 683396 233996 683448 234048
rect 652208 233860 652260 233912
rect 672172 233860 672224 233912
rect 675852 233724 675904 233776
rect 678244 233724 678296 233776
rect 672264 233248 672316 233300
rect 673092 233248 673144 233300
rect 670332 233044 670384 233096
rect 673000 233044 673052 233096
rect 669412 232908 669464 232960
rect 674196 232908 674248 232960
rect 639604 232500 639656 232552
rect 654784 232500 654836 232552
rect 660304 232500 660356 232552
rect 675852 232500 675904 232552
rect 683212 232500 683264 232552
rect 670792 232432 670844 232484
rect 665456 231616 665508 231668
rect 674932 231616 674984 231668
rect 146208 231548 146260 231600
rect 150532 231548 150584 231600
rect 155500 231548 155552 231600
rect 156972 231548 157024 231600
rect 663064 231480 663116 231532
rect 670792 231480 670844 231532
rect 675852 231480 675904 231532
rect 683580 231480 683632 231532
rect 146760 231412 146812 231464
rect 147220 231412 147272 231464
rect 156604 231412 156656 231464
rect 163688 231412 163740 231464
rect 662328 231344 662380 231396
rect 675116 231344 675168 231396
rect 137928 231276 137980 231328
rect 152464 231276 152516 231328
rect 155776 231276 155828 231328
rect 161756 231276 161808 231328
rect 91744 231140 91796 231192
rect 168840 231140 168892 231192
rect 664996 231140 665048 231192
rect 596824 231072 596876 231124
rect 633624 231072 633676 231124
rect 636844 231072 636896 231124
rect 650644 231072 650696 231124
rect 128268 231004 128320 231056
rect 195888 231004 195940 231056
rect 675116 231004 675168 231056
rect 97908 230868 97960 230920
rect 173992 230868 174044 230920
rect 674956 230800 675008 230852
rect 110328 230732 110380 230784
rect 184296 230732 184348 230784
rect 118608 230596 118660 230648
rect 188160 230596 188212 230648
rect 195060 230596 195112 230648
rect 196900 230596 196952 230648
rect 672172 230596 672224 230648
rect 439320 230528 439372 230580
rect 152464 230460 152516 230512
rect 203616 230460 203668 230512
rect 42432 230392 42484 230444
rect 43168 230392 43220 230444
rect 130384 230392 130436 230444
rect 142436 230392 142488 230444
rect 142620 230392 142672 230444
rect 146208 230392 146260 230444
rect 147634 230392 147686 230444
rect 149520 230392 149572 230444
rect 206284 230392 206336 230444
rect 256424 230392 256476 230444
rect 287060 230392 287112 230444
rect 307944 230392 307996 230444
rect 308404 230392 308456 230444
rect 334992 230392 335044 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 444472 230392 444524 230444
rect 447600 230392 447652 230444
rect 526904 230392 526956 230444
rect 536104 230392 536156 230444
rect 673460 230392 673512 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 487620 230324 487672 230376
rect 488448 230324 488500 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 511448 230324 511500 230376
rect 517520 230324 517572 230376
rect 133788 230256 133840 230308
rect 202328 230256 202380 230308
rect 210424 230256 210476 230308
rect 261576 230256 261628 230308
rect 275652 230256 275704 230308
rect 313096 230256 313148 230308
rect 436100 230256 436152 230308
rect 436836 230256 436888 230308
rect 528836 230256 528888 230308
rect 539600 230256 539652 230308
rect 388444 230188 388496 230240
rect 391664 230188 391716 230240
rect 443828 230188 443880 230240
rect 444656 230188 444708 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 453488 230188 453540 230240
rect 455788 230188 455840 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 674380 230188 674432 230240
rect 95240 230120 95292 230172
rect 157294 230120 157346 230172
rect 157432 230120 157484 230172
rect 161112 230120 161164 230172
rect 176752 230120 176804 230172
rect 235816 230120 235868 230172
rect 264244 230120 264296 230172
rect 302792 230120 302844 230172
rect 312636 230120 312688 230172
rect 340144 230120 340196 230172
rect 521108 230120 521160 230172
rect 529204 230120 529256 230172
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 126888 229984 126940 230036
rect 195060 229984 195112 230036
rect 195428 229984 195480 230036
rect 214748 229984 214800 230036
rect 220084 229984 220136 230036
rect 230664 229984 230716 230036
rect 242532 229984 242584 230036
rect 287336 229984 287388 230036
rect 302884 229984 302936 230036
rect 329840 229984 329892 230036
rect 334256 229984 334308 230036
rect 355600 229984 355652 230036
rect 355784 229984 355836 230036
rect 371056 229984 371108 230036
rect 457352 229984 457404 230036
rect 463884 229984 463936 230036
rect 476672 229984 476724 230036
rect 481640 229984 481692 230036
rect 517244 229984 517296 230036
rect 526444 229984 526496 230036
rect 534632 229984 534684 230036
rect 549260 229984 549312 230036
rect 674196 229984 674248 230036
rect 86224 229848 86276 229900
rect 156788 229848 156840 229900
rect 68284 229712 68336 229764
rect 142620 229712 142672 229764
rect 147772 229712 147824 229764
rect 158536 229848 158588 229900
rect 163964 229848 164016 229900
rect 225512 229848 225564 229900
rect 230480 229848 230532 229900
rect 277032 229848 277084 229900
rect 282552 229848 282604 229900
rect 318248 229848 318300 229900
rect 324228 229848 324280 229900
rect 350448 229848 350500 229900
rect 366732 229848 366784 229900
rect 383936 229848 383988 229900
rect 449624 229848 449676 229900
rect 450544 229848 450596 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 479248 229848 479300 229900
rect 488080 229848 488132 229900
rect 492128 229848 492180 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 476028 229780 476080 229832
rect 478604 229780 478656 229832
rect 82084 229576 82136 229628
rect 147128 229508 147180 229560
rect 171048 229712 171100 229764
rect 220084 229712 220136 229764
rect 148140 229576 148192 229628
rect 155960 229576 156012 229628
rect 157340 229576 157392 229628
rect 102140 229440 102192 229492
rect 144000 229440 144052 229492
rect 144184 229440 144236 229492
rect 146944 229440 146996 229492
rect 111064 229304 111116 229356
rect 147588 229304 147640 229356
rect 147772 229304 147824 229356
rect 210056 229440 210108 229492
rect 214748 229576 214800 229628
rect 246120 229712 246172 229764
rect 256516 229712 256568 229764
rect 297640 229712 297692 229764
rect 318064 229712 318116 229764
rect 220360 229440 220412 229492
rect 220636 229440 220688 229492
rect 266728 229576 266780 229628
rect 276296 229576 276348 229628
rect 292488 229576 292540 229628
rect 296996 229576 297048 229628
rect 323400 229576 323452 229628
rect 345020 229712 345072 229764
rect 360752 229712 360804 229764
rect 361212 229712 361264 229764
rect 378784 229712 378836 229764
rect 391204 229712 391256 229764
rect 398748 229712 398800 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 410892 229712 410944 229764
rect 417424 229712 417476 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 469588 229712 469640 229764
rect 481824 229712 481876 229764
rect 489920 229712 489972 229764
rect 490196 229712 490248 229764
rect 493600 229712 493652 229764
rect 495992 229848 496044 229900
rect 507124 229848 507176 229900
rect 510804 229848 510856 229900
rect 511908 229848 511960 229900
rect 515312 229848 515364 229900
rect 525708 229848 525760 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 674452 229916 674504 229968
rect 505192 229712 505244 229764
rect 507584 229712 507636 229764
rect 516784 229712 516836 229764
rect 523040 229712 523092 229764
rect 534816 229712 534868 229764
rect 538496 229712 538548 229764
rect 566464 229712 566516 229764
rect 476764 229644 476816 229696
rect 345296 229576 345348 229628
rect 509516 229576 509568 229628
rect 515404 229576 515456 229628
rect 530124 229576 530176 229628
rect 531136 229576 531188 229628
rect 384304 229508 384356 229560
rect 389088 229508 389140 229560
rect 448980 229508 449032 229560
rect 451372 229508 451424 229560
rect 231124 229440 231176 229492
rect 271880 229440 271932 229492
rect 530768 229440 530820 229492
rect 538312 229576 538364 229628
rect 674334 229712 674386 229764
rect 446404 229372 446456 229424
rect 448796 229372 448848 229424
rect 450912 229372 450964 229424
rect 453028 229372 453080 229424
rect 673184 229372 673236 229424
rect 151176 229304 151228 229356
rect 123484 229168 123536 229220
rect 153384 229168 153436 229220
rect 153844 229304 153896 229356
rect 156604 229304 156656 229356
rect 159364 229304 159416 229356
rect 215208 229304 215260 229356
rect 246488 229304 246540 229356
rect 282184 229304 282236 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 472164 229304 472216 229356
rect 472992 229304 473044 229356
rect 488264 229304 488316 229356
rect 490380 229304 490432 229356
rect 450268 229236 450320 229288
rect 451832 229236 451884 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 505652 229236 505704 229288
rect 510620 229236 510672 229288
rect 513380 229236 513432 229288
rect 519360 229236 519412 229288
rect 155776 229168 155828 229220
rect 157616 229168 157668 229220
rect 166264 229168 166316 229220
rect 167368 229168 167420 229220
rect 174268 229168 174320 229220
rect 184664 229168 184716 229220
rect 240968 229168 241020 229220
rect 100668 229032 100720 229084
rect 106188 229032 106240 229084
rect 142988 229032 143040 229084
rect 143448 229032 143500 229084
rect 146208 229032 146260 229084
rect 146392 229032 146444 229084
rect 156880 229032 156932 229084
rect 157524 229032 157576 229084
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 519176 229100 519228 229152
rect 202880 229032 202932 229084
rect 204720 229032 204772 229084
rect 212356 229032 212408 229084
rect 213920 229032 213972 229084
rect 214564 229032 214616 229084
rect 214748 229032 214800 229084
rect 257068 229032 257120 229084
rect 257896 229032 257948 229084
rect 296352 229032 296404 229084
rect 302148 229032 302200 229084
rect 331128 229032 331180 229084
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 660948 229100 661000 229152
rect 665456 229100 665508 229152
rect 673368 229100 673420 229152
rect 167000 228896 167052 228948
rect 167368 228896 167420 228948
rect 169484 228896 169536 228948
rect 179696 228896 179748 228948
rect 180064 228896 180116 228948
rect 219900 228896 219952 228948
rect 93768 228760 93820 228812
rect 166816 228760 166868 228812
rect 166954 228760 167006 228812
rect 174820 228760 174872 228812
rect 218152 228760 218204 228812
rect 246764 228896 246816 228948
rect 257712 228896 257764 228948
rect 299572 228896 299624 228948
rect 300676 228896 300728 228948
rect 330484 228896 330536 228948
rect 502432 228896 502484 228948
rect 521016 228896 521068 228948
rect 542452 228896 542504 228948
rect 67548 228624 67600 228676
rect 61660 228488 61712 228540
rect 142620 228488 142672 228540
rect 57244 228352 57296 228404
rect 141148 228352 141200 228404
rect 142988 228624 143040 228676
rect 152464 228624 152516 228676
rect 153108 228624 153160 228676
rect 142988 228488 143040 228540
rect 145932 228488 145984 228540
rect 146116 228488 146168 228540
rect 210700 228488 210752 228540
rect 212356 228624 212408 228676
rect 238576 228760 238628 228812
rect 282828 228760 282880 228812
rect 296628 228760 296680 228812
rect 329196 228760 329248 228812
rect 336464 228760 336516 228812
rect 358820 228760 358872 228812
rect 359924 228760 359976 228812
rect 376852 228760 376904 228812
rect 478880 228760 478932 228812
rect 490196 228760 490248 228812
rect 518532 228760 518584 228812
rect 541624 228760 541676 228812
rect 215852 228488 215904 228540
rect 216220 228488 216272 228540
rect 264796 228624 264848 228676
rect 285496 228624 285548 228676
rect 318892 228624 318944 228676
rect 326896 228624 326948 228676
rect 351092 228624 351144 228676
rect 354588 228624 354640 228676
rect 372344 228624 372396 228676
rect 377772 228624 377824 228676
rect 390376 228624 390428 228676
rect 498568 228624 498620 228676
rect 515772 228624 515824 228676
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 554964 228624 555016 228676
rect 220176 228488 220228 228540
rect 260288 228488 260340 228540
rect 268936 228488 268988 228540
rect 306012 228488 306064 228540
rect 313924 228488 313976 228540
rect 320824 228488 320876 228540
rect 325516 228488 325568 228540
rect 349160 228488 349212 228540
rect 350448 228488 350500 228540
rect 369124 228488 369176 228540
rect 373448 228488 373500 228540
rect 387156 228488 387208 228540
rect 390468 228488 390520 228540
rect 400036 228488 400088 228540
rect 148876 228352 148928 228404
rect 152464 228352 152516 228404
rect 166816 228352 166868 228404
rect 166954 228352 167006 228404
rect 214564 228352 214616 228404
rect 218152 228352 218204 228404
rect 231308 228352 231360 228404
rect 233884 228352 233936 228404
rect 273812 228352 273864 228404
rect 274272 228352 274324 228404
rect 312452 228352 312504 228404
rect 320088 228352 320140 228404
rect 346860 228352 346912 228404
rect 347044 228352 347096 228404
rect 365904 228352 365956 228404
rect 371148 228352 371200 228404
rect 385224 228352 385276 228404
rect 386236 228352 386288 228404
rect 397460 228352 397512 228404
rect 112812 228216 112864 228268
rect 184940 228216 184992 228268
rect 189724 228216 189776 228268
rect 239036 228216 239088 228268
rect 254952 228216 255004 228268
rect 295708 228216 295760 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485688 228488 485740 228540
rect 498292 228488 498344 228540
rect 499856 228488 499908 228540
rect 517704 228488 517756 228540
rect 527548 228488 527600 228540
rect 553216 228488 553268 228540
rect 555424 228488 555476 228540
rect 571340 228488 571392 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484584 228352 484636 228404
rect 485044 228352 485096 228404
rect 498568 228352 498620 228404
rect 507124 228352 507176 228404
rect 512092 228352 512144 228404
rect 532976 228352 533028 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 663524 228352 663576 228404
rect 672172 228352 672224 228404
rect 512736 228216 512788 228268
rect 539416 228216 539468 228268
rect 540888 228216 540940 228268
rect 119988 228080 120040 228132
rect 190092 228080 190144 228132
rect 192944 228080 192996 228132
rect 204720 228080 204772 228132
rect 214564 228080 214616 228132
rect 126704 227944 126756 227996
rect 195152 227944 195204 227996
rect 205456 227944 205508 227996
rect 214748 227944 214800 227996
rect 217508 228080 217560 228132
rect 219440 228080 219492 228132
rect 219900 228080 219952 228132
rect 225788 228080 225840 228132
rect 225972 228080 226024 228132
rect 272524 228080 272576 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 221004 227944 221056 227996
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 200396 227808 200448 227860
rect 203524 227808 203576 227860
rect 42432 227672 42484 227724
rect 42984 227672 43036 227724
rect 64788 227672 64840 227724
rect 111064 227672 111116 227724
rect 117228 227672 117280 227724
rect 187516 227672 187568 227724
rect 187700 227672 187752 227724
rect 110144 227536 110196 227588
rect 182364 227536 182416 227588
rect 185400 227536 185452 227588
rect 192668 227536 192720 227588
rect 200028 227672 200080 227724
rect 204904 227672 204956 227724
rect 210976 227808 211028 227860
rect 220084 227808 220136 227860
rect 251272 227944 251324 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 217784 227672 217836 227724
rect 219440 227672 219492 227724
rect 224592 227740 224644 227792
rect 220452 227672 220504 227724
rect 223580 227672 223632 227724
rect 233884 227808 233936 227860
rect 239312 227808 239364 227860
rect 243544 227808 243596 227860
rect 246304 227808 246356 227860
rect 248696 227808 248748 227860
rect 249064 227808 249116 227860
rect 253848 227808 253900 227860
rect 331036 227740 331088 227792
rect 334256 227740 334308 227792
rect 351092 227740 351144 227792
rect 353024 227740 353076 227792
rect 371792 227740 371844 227792
rect 373632 227740 373684 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 489920 227740 489972 227792
rect 494520 227740 494572 227792
rect 660488 227740 660540 227792
rect 665272 227740 665324 227792
rect 669044 227740 669096 227792
rect 672908 227740 672960 227792
rect 226708 227672 226760 227724
rect 268016 227672 268068 227724
rect 293776 227672 293828 227724
rect 325332 227672 325384 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 214748 227536 214800 227588
rect 214932 227536 214984 227588
rect 262220 227536 262272 227588
rect 264796 227536 264848 227588
rect 304724 227536 304776 227588
rect 315488 227536 315540 227588
rect 341432 227536 341484 227588
rect 525708 227536 525760 227588
rect 537484 227536 537536 227588
rect 60648 227400 60700 227452
rect 102140 227400 102192 227452
rect 103428 227400 103480 227452
rect 171232 227400 171284 227452
rect 172152 227400 172204 227452
rect 177212 227400 177264 227452
rect 181352 227400 181404 227452
rect 96436 227264 96488 227316
rect 89628 227128 89680 227180
rect 156880 227128 156932 227180
rect 169484 227264 169536 227316
rect 160192 227128 160244 227180
rect 185584 227264 185636 227316
rect 186136 227400 186188 227452
rect 187700 227400 187752 227452
rect 189908 227400 189960 227452
rect 204720 227400 204772 227452
rect 204904 227400 204956 227452
rect 251916 227400 251968 227452
rect 259368 227400 259420 227452
rect 298284 227400 298336 227452
rect 306196 227400 306248 227452
rect 336924 227400 336976 227452
rect 337752 227400 337804 227452
rect 345020 227400 345072 227452
rect 352564 227400 352616 227452
rect 363236 227400 363288 227452
rect 494704 227400 494756 227452
rect 511080 227400 511132 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 536104 227400 536156 227452
rect 552480 227400 552532 227452
rect 219440 227264 219492 227316
rect 219808 227264 219860 227316
rect 241612 227264 241664 227316
rect 249248 227264 249300 227316
rect 290556 227264 290608 227316
rect 291016 227264 291068 227316
rect 322112 227264 322164 227316
rect 340696 227264 340748 227316
rect 361396 227264 361448 227316
rect 363604 227264 363656 227316
rect 368480 227264 368532 227316
rect 382096 227264 382148 227316
rect 392952 227264 393004 227316
rect 171600 227128 171652 227180
rect 56508 226992 56560 227044
rect 142160 226992 142212 227044
rect 143264 226992 143316 227044
rect 204076 226992 204128 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 214104 226992 214156 227044
rect 220268 227128 220320 227180
rect 233700 227128 233752 227180
rect 235816 227128 235868 227180
rect 280252 227128 280304 227180
rect 281356 227128 281408 227180
rect 317604 227128 317656 227180
rect 322204 227128 322256 227180
rect 332416 227128 332468 227180
rect 333888 227128 333940 227180
rect 356244 227128 356296 227180
rect 357256 227128 357308 227180
rect 374276 227128 374328 227180
rect 376668 227128 376720 227180
rect 389732 227128 389784 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 510620 227264 510672 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 551560 227264 551612 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 490380 227128 490432 227180
rect 503168 227128 503220 227180
rect 505008 227128 505060 227180
rect 523040 227128 523092 227180
rect 523684 227128 523736 227180
rect 548156 227128 548208 227180
rect 556804 227128 556856 227180
rect 570604 227128 570656 227180
rect 668584 227128 668636 227180
rect 673552 227128 673604 227180
rect 129556 226720 129608 226772
rect 197452 226720 197504 226772
rect 204720 226720 204772 226772
rect 214748 226856 214800 226908
rect 219808 226856 219860 226908
rect 228732 226992 228784 227044
rect 228916 226992 228968 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 310336 226992 310388 227044
rect 338212 226992 338264 227044
rect 338672 226992 338724 227044
rect 360108 226992 360160 227044
rect 362776 226992 362828 227044
rect 379060 226992 379112 227044
rect 391756 226992 391808 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 506296 226992 506348 227044
rect 526628 226992 526680 227044
rect 533344 226992 533396 227044
rect 560760 226992 560812 227044
rect 652024 226992 652076 227044
rect 673552 226992 673604 227044
rect 426440 226924 426492 226976
rect 426992 226924 427044 226976
rect 220268 226856 220320 226908
rect 214104 226720 214156 226772
rect 218428 226720 218480 226772
rect 219348 226720 219400 226772
rect 267372 226856 267424 226908
rect 378784 226788 378836 226840
rect 385868 226788 385920 226840
rect 225604 226720 225656 226772
rect 238392 226720 238444 226772
rect 241152 226720 241204 226772
rect 286692 226720 286744 226772
rect 136548 226584 136600 226636
rect 203156 226584 203208 226636
rect 204076 226584 204128 226636
rect 208124 226584 208176 226636
rect 212172 226584 212224 226636
rect 214932 226584 214984 226636
rect 220452 226584 220504 226636
rect 226708 226584 226760 226636
rect 670792 226516 670844 226568
rect 106924 226448 106976 226500
rect 146576 226448 146628 226500
rect 150072 226448 150124 226500
rect 213276 226448 213328 226500
rect 216404 226448 216456 226500
rect 220636 226448 220688 226500
rect 221832 226448 221884 226500
rect 228916 226448 228968 226500
rect 369124 226448 369176 226500
rect 376208 226448 376260 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 673000 226516 673052 226568
rect 386052 226380 386104 226432
rect 391204 226380 391256 226432
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 488080 226312 488132 226364
rect 490012 226312 490064 226364
rect 672156 226312 672208 226364
rect 122564 226244 122616 226296
rect 193956 226244 194008 226296
rect 194140 226244 194192 226296
rect 204904 226244 204956 226296
rect 205088 226244 205140 226296
rect 255136 226244 255188 226296
rect 260656 226244 260708 226296
rect 298928 226244 298980 226296
rect 308220 226244 308272 226296
rect 336280 226244 336332 226296
rect 388628 226244 388680 226296
rect 394240 226244 394292 226296
rect 72424 226108 72476 226160
rect 141148 226108 141200 226160
rect 141516 226108 141568 226160
rect 145012 226108 145064 226160
rect 145196 226108 145248 226160
rect 146760 226108 146812 226160
rect 148968 226108 149020 226160
rect 213460 226108 213512 226160
rect 213644 226108 213696 226160
rect 220084 226108 220136 226160
rect 222016 226108 222068 226160
rect 269948 226108 270000 226160
rect 270224 226108 270276 226160
rect 287060 226108 287112 226160
rect 288072 226108 288124 226160
rect 322756 226108 322808 226160
rect 526444 226108 526496 226160
rect 539968 226244 540020 226296
rect 563704 226244 563756 226296
rect 568120 226244 568172 226296
rect 83464 225972 83516 226024
rect 163044 225972 163096 226024
rect 196348 225972 196400 226024
rect 236460 225972 236512 226024
rect 252468 225972 252520 226024
rect 293132 225972 293184 226024
rect 299388 225972 299440 226024
rect 328552 225972 328604 226024
rect 335176 225972 335228 226024
rect 356888 225972 356940 226024
rect 361212 225972 361264 226024
rect 377496 225972 377548 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538496 226108 538548 226160
rect 670792 226040 670844 226092
rect 538312 225972 538364 226024
rect 556160 225972 556212 226024
rect 76564 225836 76616 225888
rect 157892 225836 157944 225888
rect 169668 225836 169720 225888
rect 171600 225836 171652 225888
rect 171784 225836 171836 225888
rect 204536 225836 204588 225888
rect 204904 225836 204956 225888
rect 213644 225836 213696 225888
rect 220084 225836 220136 225888
rect 244188 225836 244240 225888
rect 261852 225836 261904 225888
rect 300860 225836 300912 225888
rect 312912 225836 312964 225888
rect 341708 225836 341760 225888
rect 341984 225836 342036 225888
rect 365260 225836 365312 225888
rect 375012 225836 375064 225888
rect 387800 225836 387852 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 501144 225836 501196 225888
rect 519176 225836 519228 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 672264 225836 672316 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 66168 225700 66220 225752
rect 149796 225700 149848 225752
rect 151268 225700 151320 225752
rect 58992 225564 59044 225616
rect 141516 225564 141568 225616
rect 141792 225564 141844 225616
rect 203156 225564 203208 225616
rect 203892 225700 203944 225752
rect 204720 225700 204772 225752
rect 204904 225700 204956 225752
rect 248880 225700 248932 225752
rect 251088 225700 251140 225752
rect 294420 225700 294472 225752
rect 296444 225700 296496 225752
rect 327908 225700 327960 225752
rect 329748 225700 329800 225752
rect 353668 225700 353720 225752
rect 365352 225700 365404 225752
rect 383292 225700 383344 225752
rect 387708 225700 387760 225752
rect 397828 225700 397880 225752
rect 481180 225700 481232 225752
rect 492680 225700 492732 225752
rect 493600 225700 493652 225752
rect 505376 225700 505428 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563060 225700 563112 225752
rect 217140 225564 217192 225616
rect 220084 225564 220136 225616
rect 266084 225564 266136 225616
rect 267004 225564 267056 225616
rect 274456 225564 274508 225616
rect 278412 225564 278464 225616
rect 313280 225564 313332 225616
rect 327724 225564 327776 225616
rect 352380 225564 352432 225616
rect 352932 225564 352984 225616
rect 371608 225564 371660 225616
rect 382924 225564 382976 225616
rect 396172 225564 396224 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488724 225564 488776 225616
rect 489368 225564 489420 225616
rect 502984 225564 503036 225616
rect 510160 225564 510212 225616
rect 530584 225564 530636 225616
rect 531412 225564 531464 225616
rect 558184 225564 558236 225616
rect 672264 225496 672316 225548
rect 125232 225428 125284 225480
rect 196164 225428 196216 225480
rect 198004 225428 198056 225480
rect 204904 225428 204956 225480
rect 209596 225428 209648 225480
rect 259644 225428 259696 225480
rect 297364 225428 297416 225480
rect 310520 225428 310572 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 129372 225292 129424 225344
rect 199108 225292 199160 225344
rect 203156 225292 203208 225344
rect 209412 225292 209464 225344
rect 62028 225156 62080 225208
rect 130384 225156 130436 225208
rect 135076 225156 135128 225208
rect 204260 225156 204312 225208
rect 204536 225156 204588 225208
rect 222936 225292 222988 225344
rect 242900 225292 242952 225344
rect 285036 225292 285088 225344
rect 672156 225292 672208 225344
rect 671252 225224 671304 225276
rect 215208 225156 215260 225208
rect 220084 225156 220136 225208
rect 132408 225020 132460 225072
rect 201684 225020 201736 225072
rect 202604 225020 202656 225072
rect 254492 225020 254544 225072
rect 554964 225020 555016 225072
rect 559104 225020 559156 225072
rect 666468 225020 666520 225072
rect 355232 224952 355284 225004
rect 358176 224952 358228 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 96252 224884 96304 224936
rect 172980 224884 173032 224936
rect 177488 224884 177540 224936
rect 199752 224884 199804 224936
rect 199936 224884 199988 224936
rect 248052 224884 248104 224936
rect 266268 224884 266320 224936
rect 303436 224884 303488 224936
rect 304264 224884 304316 224936
rect 315304 224884 315356 224936
rect 319812 224884 319864 224936
rect 345940 224884 345992 224936
rect 460572 224884 460624 224936
rect 463148 224884 463200 224936
rect 519360 224884 519412 224936
rect 535000 224884 535052 224936
rect 621020 224884 621072 224936
rect 350264 224816 350316 224868
rect 355784 224816 355836 224868
rect 670792 224816 670844 224868
rect 89444 224748 89496 224800
rect 168196 224748 168248 224800
rect 79968 224612 80020 224664
rect 160468 224612 160520 224664
rect 165160 224612 165212 224664
rect 171968 224748 172020 224800
rect 172152 224748 172204 224800
rect 178960 224748 179012 224800
rect 179328 224748 179380 224800
rect 237748 224748 237800 224800
rect 248328 224748 248380 224800
rect 291844 224748 291896 224800
rect 294880 224748 294932 224800
rect 325976 224748 326028 224800
rect 331864 224748 331916 224800
rect 337568 224748 337620 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526352 224748 526404 224800
rect 529940 224748 529992 224800
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 224868 224612 224920 224664
rect 227536 224612 227588 224664
rect 272340 224612 272392 224664
rect 272524 224612 272576 224664
rect 309876 224612 309928 224664
rect 311532 224612 311584 224664
rect 338856 224612 338908 224664
rect 346308 224612 346360 224664
rect 366548 224612 366600 224664
rect 494060 224612 494112 224664
rect 510160 224612 510212 224664
rect 520464 224612 520516 224664
rect 544108 224612 544160 224664
rect 548340 224748 548392 224800
rect 550824 224748 550876 224800
rect 549076 224612 549128 224664
rect 549260 224612 549312 224664
rect 555792 224748 555844 224800
rect 556160 224748 556212 224800
rect 557356 224748 557408 224800
rect 558828 224748 558880 224800
rect 559104 224748 559156 224800
rect 562692 224748 562744 224800
rect 571524 224748 571576 224800
rect 557816 224612 557868 224664
rect 562140 224612 562192 224664
rect 610992 224748 611044 224800
rect 610624 224612 610676 224664
rect 617064 224612 617116 224664
rect 73712 224340 73764 224392
rect 155316 224340 155368 224392
rect 156696 224340 156748 224392
rect 157340 224340 157392 224392
rect 161664 224340 161716 224392
rect 171600 224476 171652 224528
rect 178500 224476 178552 224528
rect 178960 224476 179012 224528
rect 232596 224476 232648 224528
rect 233148 224476 233200 224528
rect 272340 224476 272392 224528
rect 165988 224340 166040 224392
rect 171784 224340 171836 224392
rect 171968 224340 172020 224392
rect 227076 224340 227128 224392
rect 228732 224340 228784 224392
rect 275100 224476 275152 224528
rect 286324 224476 286376 224528
rect 289912 224476 289964 224528
rect 290832 224476 290884 224528
rect 324044 224476 324096 224528
rect 342168 224476 342220 224528
rect 362040 224476 362092 224528
rect 366732 224476 366784 224528
rect 381636 224476 381688 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506020 224476 506072 224528
rect 535276 224476 535328 224528
rect 562140 224476 562192 224528
rect 562324 224476 562376 224528
rect 610808 224476 610860 224528
rect 671712 224476 671764 224528
rect 670608 224408 670660 224460
rect 275100 224340 275152 224392
rect 311164 224340 311216 224392
rect 322848 224340 322900 224392
rect 349804 224340 349856 224392
rect 359464 224340 359516 224392
rect 378140 224340 378192 224392
rect 379244 224340 379296 224392
rect 393596 224340 393648 224392
rect 394516 224340 394568 224392
rect 404544 224340 404596 224392
rect 480536 224340 480588 224392
rect 492864 224340 492916 224392
rect 499212 224340 499264 224392
rect 516600 224340 516652 224392
rect 525524 224340 525576 224392
rect 548340 224340 548392 224392
rect 548524 224340 548576 224392
rect 558184 224340 558236 224392
rect 558828 224340 558880 224392
rect 626540 224340 626592 224392
rect 68928 224204 68980 224256
rect 152740 224204 152792 224256
rect 155776 224204 155828 224256
rect 160192 224204 160244 224256
rect 168288 224204 168340 224256
rect 230020 224204 230072 224256
rect 231676 224204 231728 224256
rect 102048 224068 102100 224120
rect 171600 224068 171652 224120
rect 171784 224068 171836 224120
rect 194600 224068 194652 224120
rect 194784 224068 194836 224120
rect 250628 224068 250680 224120
rect 272340 224204 272392 224256
rect 277676 224204 277728 224256
rect 289728 224204 289780 224256
rect 296996 224204 297048 224256
rect 299112 224204 299164 224256
rect 331404 224204 331456 224256
rect 339408 224204 339460 224256
rect 362316 224204 362368 224256
rect 372528 224204 372580 224256
rect 387432 224204 387484 224256
rect 390192 224204 390244 224256
rect 401968 224204 402020 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 427912 224204 427964 224256
rect 428740 224204 428792 224256
rect 451372 224204 451424 224256
rect 452200 224204 452252 224256
rect 470232 224204 470284 224256
rect 480352 224204 480404 224256
rect 483756 224204 483808 224256
rect 496912 224204 496964 224256
rect 278964 224068 279016 224120
rect 504364 224068 504416 224120
rect 523500 224204 523552 224256
rect 524420 224204 524472 224256
rect 525064 224204 525116 224256
rect 619640 224204 619692 224256
rect 651288 224204 651340 224256
rect 666468 224204 666520 224256
rect 668032 224204 668084 224256
rect 620192 224136 620244 224188
rect 625436 224136 625488 224188
rect 667848 224068 667900 224120
rect 279424 224000 279476 224052
rect 284760 224000 284812 224052
rect 517704 224000 517756 224052
rect 610624 224000 610676 224052
rect 610992 224000 611044 224052
rect 106004 223932 106056 223984
rect 181076 223932 181128 223984
rect 191564 223932 191616 223984
rect 199844 223932 199896 223984
rect 201408 223932 201460 223984
rect 255780 223932 255832 223984
rect 515956 223864 516008 223916
rect 538496 223864 538548 223916
rect 539508 223864 539560 223916
rect 542452 223864 542504 223916
rect 548524 223864 548576 223916
rect 549260 223864 549312 223916
rect 549904 223864 549956 223916
rect 557816 223864 557868 223916
rect 558184 223864 558236 223916
rect 610624 223864 610676 223916
rect 610808 223864 610860 223916
rect 620192 223864 620244 223916
rect 625252 223864 625304 223916
rect 108672 223796 108724 223848
rect 183652 223796 183704 223848
rect 184388 223796 184440 223848
rect 207480 223796 207532 223848
rect 207664 223796 207716 223848
rect 228088 223796 228140 223848
rect 245476 223796 245528 223848
rect 287612 223796 287664 223848
rect 505192 223728 505244 223780
rect 507676 223728 507728 223780
rect 539968 223728 540020 223780
rect 622676 223728 622728 223780
rect 115296 223660 115348 223712
rect 188804 223660 188856 223712
rect 505376 223592 505428 223644
rect 99288 223524 99340 223576
rect 175740 223524 175792 223576
rect 183192 223524 183244 223576
rect 184664 223524 184716 223576
rect 187332 223524 187384 223576
rect 242256 223524 242308 223576
rect 249432 223524 249484 223576
rect 276296 223524 276348 223576
rect 278596 223524 278648 223576
rect 315028 223524 315080 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 610624 223592 610676 223644
rect 622492 223592 622544 223644
rect 614948 223456 615000 223508
rect 81348 223388 81400 223440
rect 157248 223388 157300 223440
rect 157432 223388 157484 223440
rect 159824 223388 159876 223440
rect 162124 223388 162176 223440
rect 85304 223252 85356 223304
rect 162400 223252 162452 223304
rect 171784 223388 171836 223440
rect 181720 223388 181772 223440
rect 184848 223388 184900 223440
rect 239680 223388 239732 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 186872 223252 186924 223304
rect 188160 223252 188212 223304
rect 245108 223252 245160 223304
rect 250904 223252 250956 223304
rect 291200 223388 291252 223440
rect 316684 223388 316736 223440
rect 327264 223388 327316 223440
rect 517520 223388 517572 223440
rect 532516 223388 532568 223440
rect 534816 223388 534868 223440
rect 547512 223388 547564 223440
rect 297548 223320 297600 223372
rect 305368 223320 305420 223372
rect 288992 223252 289044 223304
rect 295064 223252 295116 223304
rect 307668 223252 307720 223304
rect 335636 223252 335688 223304
rect 337936 223252 337988 223304
rect 359188 223252 359240 223304
rect 493048 223252 493100 223304
rect 508504 223252 508556 223304
rect 514668 223252 514720 223304
rect 535460 223252 535512 223304
rect 68744 223116 68796 223168
rect 146576 223116 146628 223168
rect 146760 223116 146812 223168
rect 147634 223116 147686 223168
rect 147772 223116 147824 223168
rect 176292 223116 176344 223168
rect 181996 223116 182048 223168
rect 240324 223116 240376 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321468 223116 321520 223168
rect 323952 223116 324004 223168
rect 348516 223116 348568 223168
rect 358544 223116 358596 223168
rect 374644 223116 374696 223168
rect 483112 223116 483164 223168
rect 496084 223116 496136 223168
rect 503352 223116 503404 223168
rect 521752 223116 521804 223168
rect 529480 223116 529532 223168
rect 555700 223116 555752 223168
rect 557540 223116 557592 223168
rect 559932 223116 559984 223168
rect 562876 223116 562928 223168
rect 75828 222980 75880 223032
rect 154948 222980 155000 223032
rect 155132 222980 155184 223032
rect 71412 222844 71464 222896
rect 152096 222844 152148 222896
rect 152280 222844 152332 222896
rect 155500 222844 155552 222896
rect 157524 222980 157576 223032
rect 219072 222980 219124 223032
rect 245292 222980 245344 223032
rect 289268 222980 289320 223032
rect 291476 222980 291528 223032
rect 300216 222980 300268 223032
rect 315672 222980 315724 223032
rect 344652 222980 344704 223032
rect 349068 222980 349120 223032
rect 367192 222980 367244 223032
rect 368388 222980 368440 223032
rect 382648 222980 382700 223032
rect 383568 222980 383620 223032
rect 394884 222980 394936 223032
rect 486608 222980 486660 223032
rect 500040 222980 500092 223032
rect 508228 222980 508280 223032
rect 527180 222980 527232 223032
rect 532056 222980 532108 223032
rect 559012 222980 559064 223032
rect 171784 222844 171836 222896
rect 172888 222844 172940 222896
rect 212632 222844 212684 222896
rect 213184 222844 213236 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282736 222844 282788 222896
rect 316316 222844 316368 222896
rect 321468 222844 321520 222896
rect 346584 222844 346636 222896
rect 347228 222844 347280 222896
rect 367836 222844 367888 222896
rect 375196 222844 375248 222896
rect 391020 222844 391072 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 492036 222844 492088 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 543372 222844 543424 222896
rect 554044 222844 554096 222896
rect 632704 222844 632756 222896
rect 78588 222708 78640 222760
rect 98552 222708 98604 222760
rect 87972 222572 88024 222624
rect 164976 222708 165028 222760
rect 165620 222708 165672 222760
rect 192024 222708 192076 222760
rect 193956 222708 194008 222760
rect 247408 222708 247460 222760
rect 284208 222708 284260 222760
rect 316960 222708 317012 222760
rect 345664 222708 345716 222760
rect 347872 222708 347924 222760
rect 532516 222708 532568 222760
rect 533528 222708 533580 222760
rect 558184 222708 558236 222760
rect 98552 222436 98604 222488
rect 126520 222572 126572 222624
rect 118424 222436 118476 222488
rect 191380 222572 191432 222624
rect 197176 222572 197228 222624
rect 249984 222572 250036 222624
rect 482744 222572 482796 222624
rect 593972 222572 594024 222624
rect 670792 223592 670844 223644
rect 671022 223320 671074 223372
rect 670792 223116 670844 223168
rect 630680 222572 630732 222624
rect 126520 222300 126572 222352
rect 146760 222436 146812 222488
rect 139124 222300 139176 222352
rect 206836 222436 206888 222488
rect 207848 222436 207900 222488
rect 258356 222436 258408 222488
rect 500224 222436 500276 222488
rect 533344 222436 533396 222488
rect 533528 222436 533580 222488
rect 621204 222436 621256 222488
rect 490012 222368 490064 222420
rect 147128 222300 147180 222352
rect 211988 222300 212040 222352
rect 237012 222300 237064 222352
rect 280896 222300 280948 222352
rect 484584 222300 484636 222352
rect 670792 222368 670844 222420
rect 629852 222300 629904 222352
rect 500224 222164 500276 222216
rect 533344 222164 533396 222216
rect 558184 222164 558236 222216
rect 562876 222164 562928 222216
rect 627092 222164 627144 222216
rect 111984 222096 112036 222148
rect 185860 222096 185912 222148
rect 200396 222096 200448 222148
rect 252928 222096 252980 222148
rect 258080 222096 258132 222148
rect 263876 222096 263928 222148
rect 270040 222096 270092 222148
rect 306380 222096 306432 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353944 222096 353996 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 560944 222096 560996 222148
rect 562508 222096 562560 222148
rect 533160 222028 533212 222080
rect 538772 222028 538824 222080
rect 539508 222028 539560 222080
rect 543188 222028 543240 222080
rect 543372 222028 543424 222080
rect 546960 222028 547012 222080
rect 547144 222028 547196 222080
rect 547696 222028 547748 222080
rect 547880 222028 547932 222080
rect 91284 221960 91336 222012
rect 167184 221960 167236 222012
rect 167460 221960 167512 222012
rect 220636 221960 220688 222012
rect 220820 221960 220872 222012
rect 222200 221960 222252 222012
rect 232136 221960 232188 222012
rect 234712 221960 234764 222012
rect 261024 221960 261076 222012
rect 301688 221960 301740 222012
rect 313188 221960 313240 222012
rect 340420 221960 340472 222012
rect 516784 221960 516836 222012
rect 527548 221960 527600 222012
rect 598572 222028 598624 222080
rect 598756 221960 598808 222012
rect 603080 221960 603132 222012
rect 533988 221892 534040 221944
rect 94596 221824 94648 221876
rect 169852 221824 169904 221876
rect 97724 221688 97776 221740
rect 172704 221824 172756 221876
rect 174084 221824 174136 221876
rect 231952 221824 232004 221876
rect 233700 221824 233752 221876
rect 277952 221824 278004 221876
rect 280068 221824 280120 221876
rect 313740 221824 313792 221876
rect 318248 221824 318300 221876
rect 343824 221824 343876 221876
rect 353300 221824 353352 221876
rect 372712 221824 372764 221876
rect 171600 221688 171652 221740
rect 73896 221552 73948 221604
rect 82084 221552 82136 221604
rect 86316 221552 86368 221604
rect 164332 221552 164384 221604
rect 164516 221552 164568 221604
rect 171784 221552 171836 221604
rect 174912 221688 174964 221740
rect 185768 221688 185820 221740
rect 243084 221688 243136 221740
rect 182640 221552 182692 221604
rect 232136 221552 232188 221604
rect 263140 221688 263192 221740
rect 263508 221688 263560 221740
rect 301044 221688 301096 221740
rect 303252 221688 303304 221740
rect 332784 221688 332836 221740
rect 344652 221688 344704 221740
rect 364524 221688 364576 221740
rect 370964 221688 371016 221740
rect 380348 221824 380400 221876
rect 492496 221824 492548 221876
rect 506848 221824 506900 221876
rect 523500 221824 523552 221876
rect 533712 221824 533764 221876
rect 424968 221756 425020 221808
rect 429200 221756 429252 221808
rect 547880 221756 547932 221808
rect 553492 221756 553544 221808
rect 380072 221688 380124 221740
rect 386512 221688 386564 221740
rect 475844 221688 475896 221740
rect 486148 221688 486200 221740
rect 496268 221688 496320 221740
rect 513564 221688 513616 221740
rect 524236 221688 524288 221740
rect 547696 221688 547748 221740
rect 553860 221824 553912 221876
rect 598940 221824 598992 221876
rect 599124 221824 599176 221876
rect 606116 221824 606168 221876
rect 559380 221688 559432 221740
rect 559564 221688 559616 221740
rect 562692 221688 562744 221740
rect 562876 221688 562928 221740
rect 567016 221688 567068 221740
rect 567200 221688 567252 221740
rect 609428 221688 609480 221740
rect 59360 221416 59412 221468
rect 141332 221416 141384 221468
rect 147588 221416 147640 221468
rect 204904 221416 204956 221468
rect 205088 221416 205140 221468
rect 220820 221416 220872 221468
rect 221004 221416 221056 221468
rect 243728 221552 243780 221604
rect 283748 221552 283800 221604
rect 302424 221552 302476 221604
rect 334072 221552 334124 221604
rect 348792 221552 348844 221604
rect 370044 221552 370096 221604
rect 373724 221552 373776 221604
rect 384304 221552 384356 221604
rect 391020 221552 391072 221604
rect 400404 221552 400456 221604
rect 401324 221552 401376 221604
rect 405832 221552 405884 221604
rect 484768 221552 484820 221604
rect 498108 221552 498160 221604
rect 501328 221552 501380 221604
rect 520188 221552 520240 221604
rect 522672 221552 522724 221604
rect 234068 221416 234120 221468
rect 276112 221416 276164 221468
rect 284024 221416 284076 221468
rect 320364 221416 320416 221468
rect 333428 221416 333480 221468
rect 357532 221416 357584 221468
rect 369492 221416 369544 221468
rect 384120 221416 384172 221468
rect 384396 221416 384448 221468
rect 395160 221416 395212 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 533160 221416 533212 221468
rect 533528 221552 533580 221604
rect 598756 221552 598808 221604
rect 598940 221552 598992 221604
rect 605932 221552 605984 221604
rect 546592 221416 546644 221468
rect 546776 221416 546828 221468
rect 599124 221416 599176 221468
rect 599308 221348 599360 221400
rect 605012 221348 605064 221400
rect 104532 221280 104584 221332
rect 176476 221280 176528 221332
rect 111156 221144 111208 221196
rect 171600 221144 171652 221196
rect 171784 221144 171836 221196
rect 185860 221280 185912 221332
rect 234252 221280 234304 221332
rect 237840 221280 237892 221332
rect 243728 221280 243780 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 527180 221280 527232 221332
rect 528192 221280 528244 221332
rect 533528 221280 533580 221332
rect 177304 221144 177356 221196
rect 185308 221144 185360 221196
rect 533712 221212 533764 221264
rect 601700 221212 601752 221264
rect 124404 221008 124456 221060
rect 193312 221008 193364 221060
rect 204904 221144 204956 221196
rect 211160 221144 211212 221196
rect 211528 221144 211580 221196
rect 260840 221144 260892 221196
rect 521016 221076 521068 221128
rect 601148 221076 601200 221128
rect 205088 221008 205140 221060
rect 218060 221008 218112 221060
rect 221004 221008 221056 221060
rect 83004 220940 83056 220992
rect 151084 220872 151136 220924
rect 155040 220872 155092 220924
rect 219624 220872 219676 220924
rect 220636 220872 220688 220924
rect 226524 221008 226576 221060
rect 227904 221008 227956 221060
rect 234068 221008 234120 221060
rect 223488 220872 223540 220924
rect 268200 221008 268252 221060
rect 517520 220940 517572 220992
rect 518440 220940 518492 220992
rect 600320 220940 600372 220992
rect 253848 220872 253900 220924
rect 258632 220872 258684 220924
rect 80520 220804 80572 220856
rect 86132 220804 86184 220856
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 456708 220804 456760 220856
rect 462136 220804 462188 220856
rect 466092 220804 466144 220856
rect 471428 220804 471480 220856
rect 515772 220804 515824 220856
rect 600504 220804 600556 220856
rect 101220 220736 101272 220788
rect 166954 220736 167006 220788
rect 167184 220736 167236 220788
rect 176476 220736 176528 220788
rect 176614 220736 176666 220788
rect 180524 220736 180576 220788
rect 180708 220736 180760 220788
rect 236736 220736 236788 220788
rect 254400 220736 254452 220788
rect 296812 220736 296864 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 455328 220668 455380 220720
rect 458824 220668 458876 220720
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 511816 220668 511868 220720
rect 76380 220600 76432 220652
rect 149244 220600 149296 220652
rect 149428 220600 149480 220652
rect 166356 220600 166408 220652
rect 166540 220600 166592 220652
rect 221280 220600 221332 220652
rect 79692 220464 79744 220516
rect 158904 220464 158956 220516
rect 164148 220464 164200 220516
rect 166908 220464 166960 220516
rect 167092 220464 167144 220516
rect 223764 220600 223816 220652
rect 236184 220600 236236 220652
rect 246488 220600 246540 220652
rect 246948 220600 247000 220652
rect 288624 220600 288676 220652
rect 304908 220600 304960 220652
rect 333244 220600 333296 220652
rect 500408 220600 500460 220652
rect 511816 220532 511868 220584
rect 223764 220464 223816 220516
rect 270592 220464 270644 220516
rect 276756 220464 276808 220516
rect 311348 220464 311400 220516
rect 328092 220464 328144 220516
rect 351276 220464 351328 220516
rect 364524 220464 364576 220516
rect 379704 220464 379756 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 567016 220668 567068 220720
rect 567200 220668 567252 220720
rect 529020 220600 529072 220652
rect 544936 220600 544988 220652
rect 550824 220600 550876 220652
rect 531688 220464 531740 220516
rect 548340 220464 548392 220516
rect 551192 220464 551244 220516
rect 560760 220464 560812 220516
rect 562876 220464 562928 220516
rect 563244 220600 563296 220652
rect 566832 220600 566884 220652
rect 567384 220600 567436 220652
rect 611452 220600 611504 220652
rect 607312 220464 607364 220516
rect 64604 220328 64656 220380
rect 141976 220328 142028 220380
rect 69756 220192 69808 220244
rect 144644 220328 144696 220380
rect 144828 220328 144880 220380
rect 202420 220328 202472 220380
rect 202788 220328 202840 220380
rect 214564 220328 214616 220380
rect 142252 220192 142304 220244
rect 149428 220192 149480 220244
rect 150900 220192 150952 220244
rect 73068 220056 73120 220108
rect 153568 220056 153620 220108
rect 154212 220056 154264 220108
rect 211712 220056 211764 220108
rect 213828 220192 213880 220244
rect 262404 220328 262456 220380
rect 262680 220328 262732 220380
rect 264244 220328 264296 220380
rect 264612 220328 264664 220380
rect 269304 220328 269356 220380
rect 273444 220328 273496 220380
rect 309232 220328 309284 220380
rect 316500 220328 316552 220380
rect 217140 220192 217192 220244
rect 265164 220192 265216 220244
rect 267648 220192 267700 220244
rect 306840 220192 306892 220244
rect 308956 220192 309008 220244
rect 339684 220192 339736 220244
rect 340328 220328 340380 220380
rect 342444 220328 342496 220380
rect 342996 220328 343048 220380
rect 351276 220328 351328 220380
rect 369308 220328 369360 220380
rect 376944 220328 376996 220380
rect 388444 220328 388496 220380
rect 436284 220328 436336 220380
rect 437020 220328 437072 220380
rect 472992 220328 473044 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 509884 220328 509936 220380
rect 522580 220328 522632 220380
rect 528376 220328 528428 220380
rect 553952 220328 554004 220380
rect 558184 220328 558236 220380
rect 566464 220328 566516 220380
rect 567844 220328 567896 220380
rect 610532 220328 610584 220380
rect 566648 220260 566700 220312
rect 567154 220260 567206 220312
rect 342996 220192 343048 220244
rect 363328 220192 363380 220244
rect 363696 220192 363748 220244
rect 381084 220192 381136 220244
rect 388444 220192 388496 220244
rect 400956 220192 401008 220244
rect 429568 220192 429620 220244
rect 432052 220192 432104 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 473176 220192 473228 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495348 220192 495400 220244
rect 497464 220192 497516 220244
rect 515220 220192 515272 220244
rect 515404 220192 515456 220244
rect 530032 220192 530084 220244
rect 531136 220192 531188 220244
rect 552296 220192 552348 220244
rect 552664 220192 552716 220244
rect 576768 220192 576820 220244
rect 610072 220192 610124 220244
rect 576584 220124 576636 220176
rect 214288 220056 214340 220108
rect 214564 220056 214616 220108
rect 229284 220056 229336 220108
rect 230204 220056 230256 220108
rect 275284 220056 275336 220108
rect 292488 220056 292540 220108
rect 326160 220056 326212 220108
rect 328920 220056 328972 220108
rect 354772 220056 354824 220108
rect 355416 220056 355468 220108
rect 375564 220056 375616 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426716 220056 426768 220108
rect 431960 220056 432012 220108
rect 434812 220056 434864 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 489644 220056 489696 220108
rect 504364 220056 504416 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 558184 220056 558236 220108
rect 582472 220056 582524 220108
rect 633440 220056 633492 220108
rect 558368 219988 558420 220040
rect 576768 219988 576820 220040
rect 576952 219988 577004 220040
rect 581644 219988 581696 220040
rect 581828 219988 581880 220040
rect 582334 219988 582386 220040
rect 107844 219920 107896 219972
rect 127624 219920 127676 219972
rect 127808 219920 127860 219972
rect 185768 219920 185820 219972
rect 114468 219784 114520 219836
rect 185124 219784 185176 219836
rect 190092 219784 190144 219836
rect 190644 219920 190696 219972
rect 244464 219920 244516 219972
rect 253572 219920 253624 219972
rect 293316 219920 293368 219972
rect 527548 219852 527600 219904
rect 202788 219784 202840 219836
rect 121092 219648 121144 219700
rect 127624 219648 127676 219700
rect 140780 219648 140832 219700
rect 140964 219648 141016 219700
rect 127808 219512 127860 219564
rect 134340 219512 134392 219564
rect 200764 219512 200816 219564
rect 201132 219648 201184 219700
rect 252744 219784 252796 219836
rect 270776 219784 270828 219836
rect 279148 219784 279200 219836
rect 286692 219784 286744 219836
rect 319076 219784 319128 219836
rect 530032 219852 530084 219904
rect 552664 219852 552716 219904
rect 552848 219852 552900 219904
rect 598388 219852 598440 219904
rect 598572 219852 598624 219904
rect 558368 219716 558420 219768
rect 558552 219716 558604 219768
rect 608600 219716 608652 219768
rect 620008 219716 620060 219768
rect 203156 219648 203208 219700
rect 205824 219512 205876 219564
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 506020 219580 506072 219632
rect 576768 219580 576820 219632
rect 581644 219580 581696 219632
rect 582334 219580 582386 219632
rect 582472 219580 582524 219632
rect 598572 219580 598624 219632
rect 208584 219512 208636 219564
rect 211712 219512 211764 219564
rect 215944 219512 215996 219564
rect 366732 219512 366784 219564
rect 105820 219444 105872 219496
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 147128 219376 147180 219428
rect 148416 219376 148468 219428
rect 148968 219376 149020 219428
rect 149244 219376 149296 219428
rect 149980 219376 150032 219428
rect 152556 219376 152608 219428
rect 153108 219376 153160 219428
rect 159180 219376 159232 219428
rect 160008 219376 160060 219428
rect 163320 219376 163372 219428
rect 163964 219376 164016 219428
rect 63132 219104 63184 219156
rect 106924 219240 106976 219292
rect 113640 219240 113692 219292
rect 152372 219240 152424 219292
rect 153200 219240 153252 219292
rect 153844 219240 153896 219292
rect 160008 219240 160060 219292
rect 204536 219376 204588 219428
rect 209688 219376 209740 219428
rect 210424 219376 210476 219428
rect 213000 219376 213052 219428
rect 258080 219376 258132 219428
rect 272892 219376 272944 219428
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 297364 219376 297416 219428
rect 304080 219376 304132 219428
rect 308404 219376 308456 219428
rect 310980 219376 311032 219428
rect 322204 219376 322256 219428
rect 341340 219376 341392 219428
rect 342260 219376 342312 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 349620 219376 349672 219428
rect 350540 219376 350592 219428
rect 366180 219376 366232 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 501052 219444 501104 219496
rect 438216 219376 438268 219428
rect 438860 219376 438912 219428
rect 439872 219376 439924 219428
rect 440332 219376 440384 219428
rect 577136 219394 577188 219446
rect 591580 219444 591632 219496
rect 619824 219580 619876 219632
rect 553216 219308 553268 219360
rect 558552 219308 558604 219360
rect 572444 219308 572496 219360
rect 574652 219308 574704 219360
rect 582472 219308 582524 219360
rect 582656 219308 582708 219360
rect 598940 219444 598992 219496
rect 607496 219444 607548 219496
rect 673000 219376 673052 219428
rect 673460 219376 673512 219428
rect 591948 219308 592000 219360
rect 596824 219308 596876 219360
rect 169116 219240 169168 219292
rect 169668 219240 169720 219292
rect 171600 219240 171652 219292
rect 172152 219240 172204 219292
rect 172428 219240 172480 219292
rect 173348 219240 173400 219292
rect 182364 219240 182416 219292
rect 189724 219240 189776 219292
rect 192300 219240 192352 219292
rect 192944 219240 192996 219292
rect 193128 219240 193180 219292
rect 198188 219240 198240 219292
rect 198924 219240 198976 219292
rect 200028 219240 200080 219292
rect 202604 219240 202656 219292
rect 207664 219240 207716 219292
rect 211344 219240 211396 219292
rect 218060 219240 218112 219292
rect 239496 219240 239548 219292
rect 272708 219240 272760 219292
rect 279056 219240 279108 219292
rect 286324 219240 286376 219292
rect 291660 219240 291712 219292
rect 313924 219240 313976 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 561864 219240 561916 219292
rect 565084 219240 565136 219292
rect 568396 219240 568448 219292
rect 571984 219240 572036 219292
rect 70584 219104 70636 219156
rect 117964 219104 118016 219156
rect 132592 219104 132644 219156
rect 177488 219104 177540 219156
rect 179052 219104 179104 219156
rect 195888 219104 195940 219156
rect 199752 219104 199804 219156
rect 243544 219104 243596 219156
rect 272340 219104 272392 219156
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 77208 218968 77260 219020
rect 140044 218968 140096 219020
rect 50712 218832 50764 218884
rect 62764 218832 62816 218884
rect 83832 218832 83884 218884
rect 153200 218968 153252 219020
rect 153384 218968 153436 219020
rect 203524 218968 203576 219020
rect 206376 218968 206428 219020
rect 253848 218968 253900 219020
rect 259184 218968 259236 219020
rect 291476 218968 291528 219020
rect 142436 218832 142488 218884
rect 152188 218832 152240 218884
rect 152372 218832 152424 218884
rect 162124 218832 162176 218884
rect 162492 218832 162544 218884
rect 169760 218832 169812 218884
rect 169944 218832 169996 218884
rect 171048 218832 171100 218884
rect 59820 218696 59872 218748
rect 143724 218696 143776 218748
rect 146760 218696 146812 218748
rect 161940 218696 161992 218748
rect 165804 218696 165856 218748
rect 180064 218832 180116 218884
rect 175740 218696 175792 218748
rect 181168 218696 181220 218748
rect 184388 218696 184440 218748
rect 188988 218832 189040 218884
rect 194140 218832 194192 218884
rect 194324 218832 194376 218884
rect 239312 218832 239364 218884
rect 246120 218832 246172 218884
rect 279056 218832 279108 218884
rect 279240 218832 279292 218884
rect 189632 218696 189684 218748
rect 189816 218696 189868 218748
rect 195336 218696 195388 218748
rect 195612 218696 195664 218748
rect 198004 218696 198056 218748
rect 198188 218696 198240 218748
rect 246304 218696 246356 218748
rect 252744 218696 252796 218748
rect 100392 218560 100444 218612
rect 105820 218560 105872 218612
rect 107016 218560 107068 218612
rect 142436 218560 142488 218612
rect 142620 218560 142672 218612
rect 143264 218560 143316 218612
rect 144276 218560 144328 218612
rect 144828 218560 144880 218612
rect 145104 218560 145156 218612
rect 145932 218560 145984 218612
rect 120264 218424 120316 218476
rect 165620 218560 165672 218612
rect 166632 218560 166684 218612
rect 202604 218560 202656 218612
rect 203064 218560 203116 218612
rect 206192 218560 206244 218612
rect 208032 218560 208084 218612
rect 161940 218424 161992 218476
rect 169576 218424 169628 218476
rect 169760 218424 169812 218476
rect 181352 218424 181404 218476
rect 186504 218424 186556 218476
rect 194324 218424 194376 218476
rect 198096 218424 198148 218476
rect 200396 218424 200448 218476
rect 202236 218424 202288 218476
rect 202788 218424 202840 218476
rect 204720 218424 204772 218476
rect 207848 218424 207900 218476
rect 208860 218424 208912 218476
rect 209504 218424 209556 218476
rect 210148 218560 210200 218612
rect 217324 218560 217376 218612
rect 219624 218560 219676 218612
rect 264612 218560 264664 218612
rect 265992 218560 266044 218612
rect 272340 218560 272392 218612
rect 272708 218560 272760 218612
rect 279424 218560 279476 218612
rect 211528 218424 211580 218476
rect 217968 218424 218020 218476
rect 223488 218424 223540 218476
rect 225972 218424 226024 218476
rect 267004 218424 267056 218476
rect 285864 218832 285916 218884
rect 291660 218832 291712 218884
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 307392 219104 307444 219156
rect 331864 219104 331916 219156
rect 333704 219104 333756 219156
rect 355232 219172 355284 219224
rect 362040 219104 362092 219156
rect 370964 219104 371016 219156
rect 552664 219104 552716 219156
rect 558184 219104 558236 219156
rect 563060 219104 563112 219156
rect 563980 219104 564032 219156
rect 567292 219104 567344 219156
rect 626356 219104 626408 219156
rect 294144 218968 294196 219020
rect 311164 218968 311216 219020
rect 325332 218968 325384 219020
rect 327724 218968 327776 219020
rect 330484 218968 330536 219020
rect 297548 218832 297600 218884
rect 314016 218832 314068 218884
rect 340328 218832 340380 218884
rect 357072 218968 357124 219020
rect 369124 218968 369176 219020
rect 370320 218968 370372 219020
rect 380072 218968 380124 219020
rect 380256 218968 380308 219020
rect 388628 218968 388680 219020
rect 552480 218968 552532 219020
rect 345664 218832 345716 218884
rect 347044 218832 347096 218884
rect 363512 218832 363564 218884
rect 368664 218832 368716 218884
rect 378784 218832 378836 218884
rect 382740 218832 382792 218884
rect 383568 218832 383620 218884
rect 386880 218832 386932 218884
rect 398104 218832 398156 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 544936 218832 544988 218884
rect 555976 218832 556028 218884
rect 291660 218696 291712 218748
rect 324596 218696 324648 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 371792 218696 371844 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 540612 218696 540664 218748
rect 288992 218424 289044 218476
rect 300492 218560 300544 218612
rect 310980 218560 311032 218612
rect 311164 218560 311216 218612
rect 316684 218560 316736 218612
rect 320640 218560 320692 218612
rect 330484 218560 330536 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 537484 218560 537536 218612
rect 547512 218696 547564 218748
rect 569224 218832 569276 218884
rect 569592 218968 569644 219020
rect 601884 218968 601936 219020
rect 676036 218968 676088 219020
rect 676864 218968 676916 219020
rect 572444 218832 572496 218884
rect 572628 218832 572680 218884
rect 575020 218832 575072 218884
rect 582380 218832 582432 218884
rect 597928 218832 597980 218884
rect 558184 218696 558236 218748
rect 571708 218696 571760 218748
rect 571984 218696 572036 218748
rect 575480 218696 575532 218748
rect 304264 218424 304316 218476
rect 512736 218424 512788 218476
rect 540612 218424 540664 218476
rect 552480 218560 552532 218612
rect 555976 218560 556028 218612
rect 598848 218560 598900 218612
rect 568396 218424 568448 218476
rect 568580 218424 568632 218476
rect 569776 218424 569828 218476
rect 571340 218424 571392 218476
rect 572260 218424 572312 218476
rect 572444 218424 572496 218476
rect 604460 218424 604512 218476
rect 458180 218356 458232 218408
rect 117964 218288 118016 218340
rect 123484 218288 123536 218340
rect 131856 218288 131908 218340
rect 132408 218288 132460 218340
rect 136824 218288 136876 218340
rect 139492 218288 139544 218340
rect 140136 218288 140188 218340
rect 181168 218288 181220 218340
rect 181536 218288 181588 218340
rect 181996 218288 182048 218340
rect 184020 218288 184072 218340
rect 184940 218288 184992 218340
rect 185676 218288 185728 218340
rect 186136 218288 186188 218340
rect 196440 218288 196492 218340
rect 210148 218288 210200 218340
rect 210332 218288 210384 218340
rect 213184 218288 213236 218340
rect 222936 218288 222988 218340
rect 231032 218288 231084 218340
rect 232872 218288 232924 218340
rect 270776 218288 270828 218340
rect 340512 218288 340564 218340
rect 352564 218288 352616 218340
rect 426624 218288 426676 218340
rect 429384 218288 429436 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 503168 218288 503220 218340
rect 614488 218288 614540 218340
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61660 218152 61712 218204
rect 67272 218152 67324 218204
rect 68284 218152 68336 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 123576 218152 123628 218204
rect 165988 218152 166040 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62028 218016 62080 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 66444 218016 66496 218068
rect 67548 218016 67600 218068
rect 68100 218016 68152 218068
rect 68744 218016 68796 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 90456 218016 90508 218068
rect 91744 218016 91796 218068
rect 92940 218016 92992 218068
rect 93768 218016 93820 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 117780 218016 117832 218068
rect 118700 218016 118752 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 126060 218016 126112 218068
rect 126704 218016 126756 218068
rect 127716 218016 127768 218068
rect 128268 218016 128320 218068
rect 128544 218016 128596 218068
rect 129372 218016 129424 218068
rect 130200 218016 130252 218068
rect 132500 218016 132552 218068
rect 132684 218016 132736 218068
rect 133512 218016 133564 218068
rect 135996 218016 136048 218068
rect 136548 218016 136600 218068
rect 138480 218016 138532 218068
rect 139124 218016 139176 218068
rect 139492 218016 139544 218068
rect 171416 218152 171468 218204
rect 173256 218152 173308 218204
rect 170772 218016 170824 218068
rect 176476 218016 176528 218068
rect 178224 218016 178276 218068
rect 179328 218016 179380 218068
rect 179880 218152 179932 218204
rect 225604 218152 225656 218204
rect 241980 218152 242032 218204
rect 242900 218152 242952 218204
rect 243544 218152 243596 218204
rect 249064 218152 249116 218204
rect 297456 218152 297508 218204
rect 302884 218152 302936 218204
rect 333060 218152 333112 218204
rect 333888 218152 333940 218204
rect 335544 218152 335596 218204
rect 338672 218152 338724 218204
rect 358728 218152 358780 218204
rect 359464 218152 359516 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 400956 218152 401008 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 428464 218152 428516 218204
rect 429108 218152 429160 218204
rect 430580 218152 430632 218204
rect 433248 218152 433300 218204
rect 434720 218152 434772 218204
rect 435732 218152 435784 218204
rect 436652 218152 436704 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 500040 218152 500092 218204
rect 609888 218152 609940 218204
rect 210332 218016 210384 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216128 218016 216180 218068
rect 218796 218016 218848 218068
rect 219348 218016 219400 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 227076 218016 227128 218068
rect 227536 218016 227588 218068
rect 229560 218016 229612 218068
rect 230480 218016 230532 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 244464 218016 244516 218068
rect 245292 218016 245344 218068
rect 247776 218016 247828 218068
rect 248328 218016 248380 218068
rect 248604 218016 248656 218068
rect 249248 218016 249300 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257896 218016 257948 218068
rect 258540 218016 258592 218068
rect 259368 218016 259420 218068
rect 260196 218016 260248 218068
rect 260748 218016 260800 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270224 218016 270276 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282736 218016 282788 218068
rect 283380 218016 283432 218068
rect 284300 218016 284352 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288072 218016 288124 218068
rect 289176 218016 289228 218068
rect 289728 218016 289780 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 298284 218016 298336 218068
rect 299388 218016 299440 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 309876 218016 309928 218068
rect 310336 218016 310388 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 314844 218016 314896 218068
rect 315488 218016 315540 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 320088 218016 320140 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 323952 218016 324004 218068
rect 324780 218016 324832 218068
rect 325516 218016 325568 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 332232 218016 332284 218068
rect 333428 218016 333480 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 337200 218016 337252 218068
rect 337752 218016 337804 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347228 218016 347280 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 352104 218016 352156 218068
rect 353300 218016 353352 218068
rect 356244 218016 356296 218068
rect 357256 218016 357308 218068
rect 357900 218016 357952 218068
rect 358544 218016 358596 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373540 218016 373592 218068
rect 374460 218016 374512 218068
rect 375012 218016 375064 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 385224 218016 385276 218068
rect 386052 218016 386104 218068
rect 389364 218016 389416 218068
rect 390468 218016 390520 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 401324 218016 401376 218068
rect 401784 218016 401836 218068
rect 402796 218016 402848 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 428280 218016 428332 218068
rect 429568 218016 429620 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 434904 218016 434956 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437756 218016 437808 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 471428 218016 471480 218068
rect 472900 218016 472952 218068
rect 492036 218016 492088 218068
rect 505652 218016 505704 218068
rect 507676 218016 507728 218068
rect 615684 218016 615736 218068
rect 646596 218016 646648 218068
rect 653404 218016 653456 218068
rect 131028 217812 131080 217864
rect 197728 217812 197780 217864
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 535460 217812 535512 217864
rect 536656 217812 536708 217864
rect 536840 217812 536892 217864
rect 116952 217676 117004 217728
rect 189264 217676 189316 217728
rect 525984 217676 526036 217728
rect 526536 217676 526588 217728
rect 533436 217676 533488 217728
rect 602896 217676 602948 217728
rect 603264 217812 603316 217864
rect 613384 217812 613436 217864
rect 603448 217676 603500 217728
rect 604460 217676 604512 217728
rect 616880 217676 616932 217728
rect 103704 217540 103756 217592
rect 178408 217540 178460 217592
rect 530584 217540 530636 217592
rect 530952 217540 531004 217592
rect 536840 217540 536892 217592
rect 538220 217540 538272 217592
rect 539140 217540 539192 217592
rect 545764 217540 545816 217592
rect 606760 217540 606812 217592
rect 675852 217540 675904 217592
rect 676588 217540 676640 217592
rect 93768 217404 93820 217456
rect 171232 217404 171284 217456
rect 526536 217404 526588 217456
rect 92066 217200 92118 217252
rect 170312 217268 170364 217320
rect 535828 217268 535880 217320
rect 598664 217268 598716 217320
rect 598848 217268 598900 217320
rect 601332 217268 601384 217320
rect 601884 217404 601936 217456
rect 628288 217404 628340 217456
rect 602344 217268 602396 217320
rect 602896 217268 602948 217320
rect 604000 217268 604052 217320
rect 642180 217268 642232 217320
rect 658924 217268 658976 217320
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 448612 217200 448664 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 489920 217200 489972 217252
rect 491162 217200 491214 217252
rect 498292 217200 498344 217252
rect 499442 217200 499494 217252
rect 502984 217200 503036 217252
rect 503582 217200 503634 217252
rect 511034 217132 511086 217184
rect 561864 217132 561916 217184
rect 562876 217132 562928 217184
rect 565084 217132 565136 217184
rect 599032 217132 599084 217184
rect 600780 217132 600832 217184
rect 604552 217132 604604 217184
rect 503582 217064 503634 217116
rect 562508 217064 562560 217116
rect 608968 216996 609020 217048
rect 609888 216996 609940 217048
rect 614120 216996 614172 217048
rect 574100 216860 574152 216912
rect 597560 216860 597612 216912
rect 598664 216860 598716 216912
rect 600780 216860 600832 216912
rect 594800 216724 594852 216776
rect 612280 216860 612332 216912
rect 601332 216724 601384 216776
rect 623872 216724 623924 216776
rect 648252 216588 648304 216640
rect 656164 216588 656216 216640
rect 675944 215500 675996 215552
rect 677048 215500 677100 215552
rect 663156 215296 663208 215348
rect 663708 215296 663760 215348
rect 575480 214820 575532 214872
rect 622308 214820 622360 214872
rect 575020 214684 575072 214736
rect 616696 214684 616748 214736
rect 617064 214684 617116 214736
rect 617800 214684 617852 214736
rect 619824 214684 619876 214736
rect 620560 214684 620612 214736
rect 621020 214684 621072 214736
rect 621664 214684 621716 214736
rect 622492 214684 622544 214736
rect 623320 214684 623372 214736
rect 625252 214684 625304 214736
rect 626080 214684 626132 214736
rect 630036 214684 630088 214736
rect 632888 214684 632940 214736
rect 644572 214684 644624 214736
rect 654784 214684 654836 214736
rect 574652 214548 574704 214600
rect 625620 214548 625672 214600
rect 654876 214548 654928 214600
rect 664444 214548 664496 214600
rect 605932 214412 605984 214464
rect 606300 214412 606352 214464
rect 607312 214412 607364 214464
rect 607864 214412 607916 214464
rect 616696 214412 616748 214464
rect 624424 214412 624476 214464
rect 626356 214412 626408 214464
rect 628840 214412 628892 214464
rect 664812 214344 664864 214396
rect 665824 214344 665876 214396
rect 35808 213936 35860 213988
rect 41696 213936 41748 213988
rect 627460 213936 627512 213988
rect 629392 213936 629444 213988
rect 649908 213868 649960 213920
rect 652024 213868 652076 213920
rect 659568 213664 659620 213716
rect 665548 213664 665600 213716
rect 647148 213596 647200 213648
rect 649724 213596 649776 213648
rect 574100 213460 574152 213512
rect 594800 213460 594852 213512
rect 574376 213324 574428 213376
rect 612832 213324 612884 213376
rect 651104 213324 651156 213376
rect 657544 213324 657596 213376
rect 574836 213188 574888 213240
rect 616144 213188 616196 213240
rect 643836 213188 643888 213240
rect 650644 213188 650696 213240
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 658188 212712 658240 212764
rect 659108 212712 659160 212764
rect 664260 212712 664312 212764
rect 665088 212712 665140 212764
rect 632704 212508 632756 212560
rect 634360 212508 634412 212560
rect 630680 212372 630732 212424
rect 631600 212372 631652 212424
rect 35808 211556 35860 211608
rect 39580 211556 39632 211608
rect 35624 211284 35676 211336
rect 41696 211284 41748 211336
rect 35440 211148 35492 211200
rect 41328 211148 41380 211200
rect 578332 211148 578384 211200
rect 580908 211148 580960 211200
rect 680360 211148 680412 211200
rect 683120 211148 683172 211200
rect 600320 211012 600372 211064
rect 600688 211012 600740 211064
rect 633440 211012 633492 211064
rect 633808 211012 633860 211064
rect 635556 210128 635608 210180
rect 636568 210128 636620 210180
rect 35808 209788 35860 209840
rect 40316 209788 40368 209840
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 35808 208496 35860 208548
rect 40684 208496 40736 208548
rect 35624 208360 35676 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207136 35860 207188
rect 41144 207136 41196 207188
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 35808 205776 35860 205828
rect 40684 205776 40736 205828
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204620 35860 204672
rect 41696 204484 41748 204536
rect 35808 204280 35860 204332
rect 41696 204280 41748 204332
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 672908 192992 672960 193044
rect 673368 192992 673420 193044
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 668216 165180 668268 165232
rect 669596 165180 669648 165232
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 668216 163276 668268 163328
rect 669780 163276 669832 163328
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 675852 162800 675904 162852
rect 678244 162800 678296 162852
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 668216 160012 668268 160064
rect 670332 160012 670384 160064
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 668308 155116 668360 155168
rect 670792 155116 670844 155168
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 668216 148724 668268 148776
rect 670148 148724 670200 148776
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585784 143556 585836 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 668216 136212 668268 136264
rect 669964 136212 670016 136264
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 585968 132472 586020 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585784 131112 585836 131164
rect 583392 129140 583444 129192
rect 590384 129140 590436 129192
rect 668584 129140 668636 129192
rect 670792 129140 670844 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 587808 126964 587860 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 579068 124856 579120 124908
rect 587808 124856 587860 124908
rect 578700 124108 578752 124160
rect 583024 124108 583076 124160
rect 584404 122816 584456 122868
rect 589556 122816 589608 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 589924 122000 589976 122052
rect 587348 121456 587400 121508
rect 589556 121456 589608 121508
rect 583208 120708 583260 120760
rect 589372 120708 589424 120760
rect 578516 118532 578568 118584
rect 580264 118532 580316 118584
rect 675852 117240 675904 117292
rect 682384 117240 682436 117292
rect 579528 116900 579580 116952
rect 583392 116900 583444 116952
rect 585784 115948 585836 116000
rect 589464 115948 589516 116000
rect 584588 115200 584640 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 579528 112820 579580 112872
rect 585968 112820 586020 112872
rect 586152 112412 586204 112464
rect 590108 112412 590160 112464
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110236 579396 110288
rect 581828 110236 581880 110288
rect 580448 109080 580500 109132
rect 589464 109080 589516 109132
rect 578332 108944 578384 108996
rect 580632 108944 580684 108996
rect 667940 108808 667992 108860
rect 669964 108808 670016 108860
rect 582288 107652 582340 107704
rect 589464 107652 589516 107704
rect 580264 106292 580316 106344
rect 589464 106292 589516 106344
rect 579344 105612 579396 105664
rect 582288 105612 582340 105664
rect 587164 104864 587216 104916
rect 589832 104864 589884 104916
rect 668216 104796 668268 104848
rect 670792 104796 670844 104848
rect 578516 103368 578568 103420
rect 588728 103368 588780 103420
rect 579160 102076 579212 102128
rect 584404 102076 584456 102128
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 578608 99968 578660 100020
rect 587348 99968 587400 100020
rect 592684 99968 592736 100020
rect 667940 99968 667992 100020
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 579528 99220 579580 99272
rect 583208 99220 583260 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 624608 99016 624660 99068
rect 635004 99016 635056 99068
rect 625068 98880 625120 98932
rect 636292 98880 636344 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98608 647200 98660
rect 661960 98608 662012 98660
rect 630496 98540 630548 98592
rect 646596 98540 646648 98592
rect 629760 98268 629812 98320
rect 645308 98268 645360 98320
rect 633624 98132 633676 98184
rect 640708 98132 640760 98184
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 628288 97928 628340 97980
rect 642180 97996 642232 98048
rect 659936 97928 659988 97980
rect 665364 97928 665416 97980
rect 632704 97792 632756 97844
rect 647516 97792 647568 97844
rect 653956 97792 654008 97844
rect 655060 97792 655112 97844
rect 655428 97792 655480 97844
rect 662512 97792 662564 97844
rect 631232 97656 631284 97708
rect 647332 97656 647384 97708
rect 650368 97656 650420 97708
rect 658280 97656 658332 97708
rect 627552 97520 627604 97572
rect 633624 97520 633676 97572
rect 633808 97520 633860 97572
rect 639236 97520 639288 97572
rect 643008 97520 643060 97572
rect 659844 97656 659896 97708
rect 605472 97384 605524 97436
rect 611912 97384 611964 97436
rect 612648 97384 612700 97436
rect 620284 97384 620336 97436
rect 623136 97384 623188 97436
rect 632060 97384 632112 97436
rect 633256 97384 633308 97436
rect 650552 97384 650604 97436
rect 651840 97384 651892 97436
rect 659568 97520 659620 97572
rect 659200 97384 659252 97436
rect 664352 97384 664404 97436
rect 592132 97248 592184 97300
rect 598940 97248 598992 97300
rect 621664 97248 621716 97300
rect 629300 97248 629352 97300
rect 631876 97248 631928 97300
rect 648620 97248 648672 97300
rect 656808 97180 656860 97232
rect 661408 97180 661460 97232
rect 620100 97112 620152 97164
rect 626356 97112 626408 97164
rect 626816 97112 626868 97164
rect 633808 97112 633860 97164
rect 634176 97112 634228 97164
rect 649080 97112 649132 97164
rect 658096 97044 658148 97096
rect 663064 97044 663116 97096
rect 634728 96976 634780 97028
rect 647056 96976 647108 97028
rect 596180 96908 596232 96960
rect 596732 96908 596784 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 656716 96908 656768 96960
rect 660120 96908 660172 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 626080 96840 626132 96892
rect 637764 96840 637816 96892
rect 644296 96772 644348 96824
rect 658832 96772 658884 96824
rect 609152 96704 609204 96756
rect 609704 96704 609756 96756
rect 640064 96568 640116 96620
rect 645124 96568 645176 96620
rect 646412 96568 646464 96620
rect 652024 96568 652076 96620
rect 653312 96568 653364 96620
rect 665180 96568 665232 96620
rect 638592 96432 638644 96484
rect 641352 96432 641404 96484
rect 641536 96432 641588 96484
rect 648068 96432 648120 96484
rect 648896 96432 648948 96484
rect 664536 96432 664588 96484
rect 637580 96296 637632 96348
rect 660672 96296 660724 96348
rect 644940 96160 644992 96212
rect 647884 96160 647936 96212
rect 649264 96160 649316 96212
rect 663984 96160 664036 96212
rect 591304 96024 591356 96076
rect 602620 96024 602672 96076
rect 610624 96024 610676 96076
rect 621664 96024 621716 96076
rect 640524 96024 640576 96076
rect 645584 96024 645636 96076
rect 645768 96024 645820 96076
rect 648068 96024 648120 96076
rect 648804 96024 648856 96076
rect 664168 96024 664220 96076
rect 594064 95888 594116 95940
rect 668032 95888 668084 95940
rect 639052 95752 639104 95804
rect 648804 95752 648856 95804
rect 652576 95752 652628 95804
rect 663800 95752 663852 95804
rect 645124 95616 645176 95668
rect 652208 95616 652260 95668
rect 641352 95412 641404 95464
rect 643468 95412 643520 95464
rect 647884 95412 647936 95464
rect 648068 95344 648120 95396
rect 656164 95480 656216 95532
rect 647700 95276 647752 95328
rect 578332 95140 578384 95192
rect 584588 95140 584640 95192
rect 620928 95140 620980 95192
rect 625436 95140 625488 95192
rect 647056 95140 647108 95192
rect 650276 95140 650328 95192
rect 590936 94936 590988 94988
rect 592132 94936 592184 94988
rect 616512 94936 616564 94988
rect 624976 94936 625028 94988
rect 607680 94460 607732 94512
rect 620928 94460 620980 94512
rect 619548 93780 619600 93832
rect 626172 93780 626224 93832
rect 647516 93712 647568 93764
rect 648252 93712 648304 93764
rect 651288 93576 651340 93628
rect 654692 93576 654744 93628
rect 579252 93372 579304 93424
rect 586152 93372 586204 93424
rect 609704 93100 609756 93152
rect 618628 93100 618680 93152
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 647700 92420 647752 92472
rect 655428 92420 655480 92472
rect 577504 91740 577556 91792
rect 590936 91740 590988 91792
rect 606944 91740 606996 91792
rect 622400 91740 622452 91792
rect 578700 91400 578752 91452
rect 585784 91400 585836 91452
rect 618168 91128 618220 91180
rect 611268 90992 611320 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 648804 90788 648856 90840
rect 655428 90788 655480 90840
rect 620928 89632 620980 89684
rect 625436 89632 625488 89684
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 664352 88748 664404 88800
rect 656164 88612 656216 88664
rect 657452 88612 657504 88664
rect 579252 88272 579304 88324
rect 589924 88272 589976 88324
rect 618168 88272 618220 88324
rect 625620 88272 625672 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 622400 88136 622452 88188
rect 626448 88136 626500 88188
rect 648436 86980 648488 87032
rect 662512 86980 662564 87032
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 652208 86708 652260 86760
rect 660120 86708 660172 86760
rect 647884 86572 647936 86624
rect 661408 86572 661460 86624
rect 652024 86436 652076 86488
rect 657176 86436 657228 86488
rect 621664 86300 621716 86352
rect 626448 86300 626500 86352
rect 656348 86300 656400 86352
rect 660672 86300 660724 86352
rect 618628 85484 618680 85536
rect 626448 85484 626500 85536
rect 609888 85348 609940 85400
rect 625344 85280 625396 85332
rect 608508 84124 608560 84176
rect 625804 84124 625856 84176
rect 579252 83988 579304 84040
rect 581644 83988 581696 84040
rect 578700 82764 578752 82816
rect 583024 82764 583076 82816
rect 579068 82084 579120 82136
rect 587164 82084 587216 82136
rect 628748 81064 628800 81116
rect 642456 81064 642508 81116
rect 615408 80928 615460 80980
rect 646136 80928 646188 80980
rect 613844 80792 613896 80844
rect 647332 80792 647384 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 614028 79432 614080 79484
rect 645952 79432 646004 79484
rect 583024 79296 583076 79348
rect 600504 79296 600556 79348
rect 612648 79296 612700 79348
rect 648620 79296 648672 79348
rect 578516 78412 578568 78464
rect 580264 78412 580316 78464
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77664 628524 77716
rect 632796 77664 632848 77716
rect 624424 77392 624476 77444
rect 628472 77392 628524 77444
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 620284 76780 620336 76832
rect 648988 76780 649040 76832
rect 612004 76644 612056 76696
rect 662420 76644 662472 76696
rect 587164 76508 587216 76560
rect 668216 76508 668268 76560
rect 616788 75420 616840 75472
rect 646504 75420 646556 75472
rect 607128 75284 607180 75336
rect 646320 75284 646372 75336
rect 578884 75148 578936 75200
rect 666560 75148 666612 75200
rect 579528 73108 579580 73160
rect 588544 73108 588596 73160
rect 578516 71544 578568 71596
rect 584404 71544 584456 71596
rect 579528 66852 579580 66904
rect 625988 66852 626040 66904
rect 579528 64812 579580 64864
rect 592684 64812 592736 64864
rect 579528 62024 579580 62076
rect 587164 62024 587216 62076
rect 578332 59984 578384 60036
rect 624424 59984 624476 60036
rect 577688 58760 577740 58812
rect 604460 58760 604512 58812
rect 576124 58624 576176 58676
rect 603080 58624 603132 58676
rect 579528 57876 579580 57928
rect 594064 57876 594116 57928
rect 577320 57196 577372 57248
rect 600320 57196 600372 57248
rect 574284 55972 574336 56024
rect 598940 55972 598992 56024
rect 577136 55836 577188 55888
rect 601884 55836 601936 55888
rect 460388 53592 460440 53644
rect 461952 53592 462004 53644
rect 462228 53592 462280 53644
rect 577320 55564 577372 55616
rect 596456 55156 596508 55208
rect 596180 55020 596232 55072
rect 597652 54884 597704 54936
rect 597928 54748 597980 54800
rect 580448 54612 580500 54664
rect 625804 54476 625856 54528
rect 464896 53592 464948 53644
rect 465080 53592 465132 53644
rect 465540 53592 465592 53644
rect 465724 53592 465776 53644
rect 469956 53592 470008 53644
rect 472808 53592 472860 53644
rect 459468 53456 459520 53508
rect 583024 54340 583076 54392
rect 473912 53592 473964 53644
rect 476672 53592 476724 53644
rect 478144 53592 478196 53644
rect 50528 53320 50580 53372
rect 130384 53320 130436 53372
rect 461308 53320 461360 53372
rect 577504 54136 577556 54188
rect 574744 53932 574796 53984
rect 623044 53932 623096 53984
rect 564532 53592 564584 53644
rect 577136 53456 577188 53508
rect 574284 53252 574336 53304
rect 48964 53184 49016 53236
rect 129188 53184 129240 53236
rect 464528 53184 464580 53236
rect 465540 53184 465592 53236
rect 465908 53184 465960 53236
rect 478144 53184 478196 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 47584 53048 47636 53100
rect 129004 53048 129056 53100
rect 459606 52776 459658 52828
rect 476672 53048 476724 53100
rect 463608 52912 463660 52964
rect 465724 52912 465776 52964
rect 463746 52776 463798 52828
rect 465080 52776 465132 52828
rect 465448 52776 465500 52828
rect 469956 52776 470008 52828
rect 50344 51824 50396 51876
rect 129372 51824 129424 51876
rect 46204 51688 46256 51740
rect 130568 51688 130620 51740
rect 145380 51688 145432 51740
rect 306012 51688 306064 51740
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 49148 50328 49200 50380
rect 131028 50328 131080 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 51724 49104 51776 49156
rect 129648 49104 129700 49156
rect 45468 48968 45520 49020
rect 129004 48968 129056 49020
rect 625988 46452 626040 46504
rect 661776 46452 661828 46504
rect 129004 46044 129056 46096
rect 132408 46044 132460 46096
rect 130568 45908 130620 45960
rect 132592 45908 132644 45960
rect 129648 45364 129700 45416
rect 43812 45160 43864 45212
rect 131120 45160 131172 45212
rect 131396 45296 131448 45348
rect 132960 45296 133012 45348
rect 131396 45160 131448 45212
rect 133144 45160 133196 45212
rect 129372 45024 129424 45076
rect 126428 44888 126480 44940
rect 129188 44752 129240 44804
rect 43628 44276 43680 44328
rect 128820 44344 128872 44396
rect 132408 44412 132460 44464
rect 132592 44364 132644 44416
rect 43444 44140 43496 44192
rect 126428 44140 126480 44192
rect 132960 44252 133012 44304
rect 130384 44004 130436 44056
rect 133144 44140 133196 44192
rect 440240 43800 440292 43852
rect 441068 43800 441120 43852
rect 410892 42848 410944 42900
rect 415584 42848 415636 42900
rect 187332 42780 187384 42832
rect 255872 42780 255924 42832
rect 310428 42712 310480 42764
rect 364524 42712 364576 42764
rect 361764 42440 361816 42492
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 453580 42712 453632 42764
rect 464344 42712 464396 42764
rect 364892 42576 364944 42628
rect 427084 42576 427136 42628
rect 441252 42576 441304 42628
rect 446404 42576 446456 42628
rect 454684 42576 454736 42628
rect 462964 42576 463016 42628
rect 364524 42304 364576 42356
rect 410892 42440 410944 42492
rect 415584 42304 415636 42356
rect 429108 42440 429160 42492
rect 454500 42440 454552 42492
rect 463700 42440 463752 42492
rect 661408 42129 661460 42181
rect 427084 41964 427136 42016
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 446404 41964 446456 42016
rect 454500 41964 454552 42016
rect 441252 41828 441304 41880
rect 429108 41692 429160 41744
rect 454684 41828 454736 41880
rect 449164 41692 449216 41744
rect 453580 41692 453632 41744
<< metal2 >>
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 652024 897048 652076 897054
rect 652024 896990 652076 896996
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 652036 867649 652064 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 675864 895830 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 654784 895824 654836 895830
rect 654784 895766 654836 895772
rect 675852 895824 675904 895830
rect 675852 895766 675904 895772
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 652022 867640 652078 867649
rect 652022 867575 652078 867584
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895766
rect 676048 895694 676076 896271
rect 672724 895688 672776 895694
rect 672724 895630 672776 895636
rect 676036 895688 676088 895694
rect 676036 895630 676088 895636
rect 671988 894464 672040 894470
rect 671988 894406 672040 894412
rect 671436 894328 671488 894334
rect 671436 894270 671488 894276
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817018 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 46204 817148 46256 817154
rect 46204 817090 46256 817096
rect 35624 817012 35676 817018
rect 35624 816954 35676 816960
rect 35438 816912 35494 816921
rect 35438 816847 35494 816856
rect 35452 815658 35480 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35820 815794 35848 816031
rect 35808 815788 35860 815794
rect 35808 815730 35860 815736
rect 44272 815788 44324 815794
rect 44272 815730 44324 815736
rect 35440 815652 35492 815658
rect 35440 815594 35492 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814434 35664 815215
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 35806 814399 35862 814408
rect 35624 814370 35676 814376
rect 35820 814298 35848 814399
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 40958 812832 41014 812841
rect 41328 812806 41380 812812
rect 43352 812864 43404 812870
rect 43352 812806 43404 812812
rect 40958 812767 41014 812776
rect 39302 811608 39358 811617
rect 39302 811543 39358 811552
rect 33046 811200 33102 811209
rect 33046 811135 33102 811144
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 31036 801106 31064 809911
rect 31758 806712 31814 806721
rect 31758 806647 31760 806656
rect 31812 806647 31814 806656
rect 31760 806618 31812 806624
rect 33060 802466 33088 811135
rect 33782 809568 33838 809577
rect 33782 809503 33838 809512
rect 33048 802460 33100 802466
rect 33048 802402 33100 802408
rect 33796 801310 33824 809503
rect 35624 806676 35676 806682
rect 35624 806618 35676 806624
rect 35636 802670 35664 806618
rect 35624 802664 35676 802670
rect 35624 802606 35676 802612
rect 33784 801304 33836 801310
rect 33784 801246 33836 801252
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 39316 800601 39344 811543
rect 40972 810762 41000 812767
rect 41142 812424 41198 812433
rect 41142 812359 41198 812368
rect 40960 810756 41012 810762
rect 40960 810698 41012 810704
rect 41156 809282 41184 812359
rect 42154 810792 42210 810801
rect 42154 810727 42210 810736
rect 42524 810756 42576 810762
rect 41970 810384 42026 810393
rect 41970 810319 42026 810328
rect 41786 809296 41842 809305
rect 41156 809254 41786 809282
rect 41786 809231 41842 809240
rect 40682 809160 40738 809169
rect 40682 809095 40738 809104
rect 40696 801553 40724 809095
rect 41786 808752 41842 808761
rect 41786 808687 41842 808696
rect 40958 808344 41014 808353
rect 40958 808279 41014 808288
rect 40972 807362 41000 808279
rect 41142 807936 41198 807945
rect 41142 807871 41198 807880
rect 41156 807498 41184 807871
rect 41144 807492 41196 807498
rect 41144 807434 41196 807440
rect 40960 807356 41012 807362
rect 40960 807298 41012 807304
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806002 41368 806239
rect 41328 805996 41380 806002
rect 41328 805938 41380 805944
rect 41800 805225 41828 808687
rect 41984 805633 42012 810319
rect 41970 805624 42026 805633
rect 41970 805559 42026 805568
rect 41786 805216 41842 805225
rect 41786 805151 41842 805160
rect 42168 804953 42196 810727
rect 42524 810698 42576 810704
rect 42154 804944 42210 804953
rect 42154 804879 42210 804888
rect 42340 802664 42392 802670
rect 42392 802612 42472 802618
rect 42340 802606 42472 802612
rect 42352 802590 42472 802606
rect 42156 802460 42208 802466
rect 42156 802402 42208 802408
rect 40682 801544 40738 801553
rect 42168 801530 42196 802402
rect 42168 801502 42288 801530
rect 40682 801479 40738 801488
rect 39856 801304 39908 801310
rect 39854 801272 39856 801281
rect 39908 801272 39910 801281
rect 39854 801207 39910 801216
rect 40684 801100 40736 801106
rect 40684 801042 40736 801048
rect 40696 800873 40724 801042
rect 40682 800864 40738 800873
rect 40682 800799 40738 800808
rect 39302 800592 39358 800601
rect 39302 800527 39358 800536
rect 42260 799898 42288 801502
rect 42168 799870 42288 799898
rect 42168 799445 42196 799870
rect 42444 799490 42472 802590
rect 42352 799462 42472 799490
rect 42352 799459 42380 799462
rect 42260 799431 42380 799459
rect 42260 798266 42288 799431
rect 42536 799218 42564 810698
rect 42982 807528 43038 807537
rect 42982 807463 43038 807472
rect 43168 807492 43220 807498
rect 42996 801666 43024 807463
rect 43168 807434 43220 807440
rect 43180 804554 43208 807434
rect 43180 804526 43300 804554
rect 42996 801638 43208 801666
rect 42182 798238 42288 798266
rect 42352 799190 42564 799218
rect 42352 797994 42380 799190
rect 42260 797966 42380 797994
rect 42260 797619 42288 797966
rect 42892 797700 42944 797706
rect 42892 797642 42944 797648
rect 42182 797591 42288 797619
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 42706 796920 42762 796929
rect 42706 796855 42762 796864
rect 42248 796340 42300 796346
rect 42248 796282 42300 796288
rect 41786 796240 41842 796249
rect 41786 796175 41842 796184
rect 41800 795765 41828 796175
rect 42260 795138 42288 796282
rect 42182 795110 42288 795138
rect 42248 794844 42300 794850
rect 42248 794786 42300 794792
rect 42260 794594 42288 794786
rect 42182 794566 42288 794594
rect 42062 794472 42118 794481
rect 42062 794407 42118 794416
rect 42076 793900 42104 794407
rect 42340 793824 42392 793830
rect 42340 793766 42392 793772
rect 42352 793302 42380 793766
rect 42182 793274 42380 793302
rect 41786 793112 41842 793121
rect 41786 793047 41842 793056
rect 41800 792744 41828 793047
rect 41786 790664 41842 790673
rect 41786 790599 41842 790608
rect 41800 790228 41828 790599
rect 42338 790256 42394 790265
rect 42338 790191 42394 790200
rect 42062 789848 42118 789857
rect 42062 789783 42118 789792
rect 42076 789616 42104 789783
rect 41800 788769 41828 788936
rect 41786 788760 41842 788769
rect 41786 788695 41842 788704
rect 42352 788406 42380 790191
rect 42720 789857 42748 796855
rect 42904 796346 42932 797642
rect 42892 796340 42944 796346
rect 42892 796282 42944 796288
rect 43180 795410 43208 801638
rect 42904 795382 43208 795410
rect 42706 789848 42762 789857
rect 42706 789783 42762 789792
rect 42522 789440 42578 789449
rect 42522 789375 42578 789384
rect 42536 789290 42564 789375
rect 42182 788378 42380 788406
rect 42444 789262 42564 789290
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42260 786570 42288 788151
rect 42182 786542 42288 786570
rect 42444 785958 42472 789262
rect 42706 789168 42762 789177
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42536 789126 42706 789154
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 789126
rect 42706 789103 42762 789112
rect 42708 786684 42760 786690
rect 42708 786626 42760 786632
rect 42182 785250 42564 785278
rect 42720 784734 42748 786626
rect 42182 784706 42748 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 41050 774752 41106 774761
rect 41050 774687 41106 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 35438 773936 35494 773945
rect 35438 773871 35494 773880
rect 35452 772886 35480 773871
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 773362 35848 773463
rect 35808 773356 35860 773362
rect 35808 773298 35860 773304
rect 41064 773158 41092 774687
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 41326 773528 41382 773537
rect 41326 773463 41382 773472
rect 42062 773528 42118 773537
rect 42062 773463 42118 773472
rect 35808 773152 35860 773158
rect 35806 773120 35808 773129
rect 41052 773152 41104 773158
rect 35860 773120 35862 773129
rect 41052 773094 41104 773100
rect 35806 773055 35862 773064
rect 35624 773016 35676 773022
rect 35624 772958 35676 772964
rect 35440 772880 35492 772886
rect 35440 772822 35492 772828
rect 35636 772721 35664 772958
rect 41340 772886 41368 773463
rect 41696 773356 41748 773362
rect 41696 773298 41748 773304
rect 41708 773129 41736 773298
rect 41694 773120 41750 773129
rect 41694 773055 41750 773064
rect 41512 773016 41564 773022
rect 41512 772958 41564 772964
rect 41328 772880 41380 772886
rect 41328 772822 41380 772828
rect 41524 772834 41552 772958
rect 42076 772886 42104 773463
rect 42064 772880 42116 772886
rect 41786 772848 41842 772857
rect 41524 772806 41786 772834
rect 42064 772822 42116 772828
rect 41786 772783 41842 772792
rect 35622 772712 35678 772721
rect 35622 772647 35678 772656
rect 35346 772304 35402 772313
rect 35346 772239 35402 772248
rect 35360 771458 35388 772239
rect 35530 771896 35586 771905
rect 35530 771831 35532 771840
rect 35584 771831 35586 771840
rect 35806 771896 35862 771905
rect 35806 771831 35862 771840
rect 39764 771860 39816 771866
rect 35532 771802 35584 771808
rect 35820 771594 35848 771831
rect 39764 771802 39816 771808
rect 35808 771588 35860 771594
rect 35808 771530 35860 771536
rect 35348 771452 35400 771458
rect 35348 771394 35400 771400
rect 35806 771080 35862 771089
rect 35806 771015 35862 771024
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35636 770234 35664 770607
rect 35820 770506 35848 771015
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 35806 770264 35862 770273
rect 35624 770228 35676 770234
rect 35806 770199 35862 770208
rect 35624 770170 35676 770176
rect 35820 770098 35848 770199
rect 35808 770092 35860 770098
rect 35808 770034 35860 770040
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768738 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35544 768874 35572 768975
rect 35860 768975 35862 768984
rect 39580 769004 39632 769010
rect 35808 768946 35860 768952
rect 39580 768946 39632 768952
rect 35532 768868 35584 768874
rect 35532 768810 35584 768816
rect 35348 768732 35400 768738
rect 35348 768674 35400 768680
rect 39592 768641 39620 768946
rect 39578 768632 39634 768641
rect 39578 768567 39634 768576
rect 35806 768224 35862 768233
rect 35806 768159 35862 768168
rect 33046 767816 33102 767825
rect 33046 767751 33102 767760
rect 33060 761054 33088 767751
rect 35820 767582 35848 768159
rect 35808 767576 35860 767582
rect 35808 767518 35860 767524
rect 35806 767408 35862 767417
rect 35806 767343 35808 767352
rect 35860 767343 35862 767352
rect 36544 767372 36596 767378
rect 35808 767314 35860 767320
rect 36544 767314 36596 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 33048 761048 33100 761054
rect 33048 760990 33100 760996
rect 35176 759694 35204 766935
rect 35806 766184 35862 766193
rect 35806 766119 35808 766128
rect 35860 766119 35862 766128
rect 35808 766090 35860 766096
rect 35806 765776 35862 765785
rect 35806 765711 35862 765720
rect 35820 764862 35848 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35808 764584 35860 764590
rect 35806 764552 35808 764561
rect 35860 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763230 35664 764079
rect 35808 763360 35860 763366
rect 35806 763328 35808 763337
rect 35860 763328 35862 763337
rect 35806 763263 35862 763272
rect 35624 763224 35676 763230
rect 35624 763166 35676 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761938 35848 762855
rect 35808 761932 35860 761938
rect 35808 761874 35860 761880
rect 35164 759688 35216 759694
rect 35164 759630 35216 759636
rect 36556 759121 36584 767314
rect 39776 764153 39804 771802
rect 42064 771656 42116 771662
rect 41708 771604 42064 771610
rect 41708 771598 42116 771604
rect 41708 771594 42104 771598
rect 41696 771588 42104 771594
rect 41748 771582 42104 771588
rect 41696 771530 41748 771536
rect 41708 771458 42104 771474
rect 41696 771452 42116 771458
rect 41748 771446 42064 771452
rect 41696 771394 41748 771400
rect 42064 771394 42116 771400
rect 40316 770500 40368 770506
rect 40316 770442 40368 770448
rect 40328 770273 40356 770442
rect 41696 770296 41748 770302
rect 40314 770264 40370 770273
rect 42064 770296 42116 770302
rect 41748 770244 42064 770250
rect 41696 770238 42116 770244
rect 41708 770222 42104 770238
rect 40314 770199 40370 770208
rect 41708 770098 42104 770114
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 40684 768868 40736 768874
rect 40684 768810 40736 768816
rect 39762 764144 39818 764153
rect 39762 764079 39818 764088
rect 39304 763360 39356 763366
rect 39304 763302 39356 763308
rect 38936 761932 38988 761938
rect 38936 761874 38988 761880
rect 36542 759112 36598 759121
rect 36542 759047 36598 759056
rect 38948 757489 38976 761874
rect 39316 757790 39344 763302
rect 40040 759688 40092 759694
rect 40040 759630 40092 759636
rect 39304 757784 39356 757790
rect 40052 757761 40080 759630
rect 40696 757761 40724 768810
rect 41696 768732 41748 768738
rect 41696 768674 41748 768680
rect 41708 768618 41736 768674
rect 42706 768632 42762 768641
rect 41708 768590 41920 768618
rect 41696 767304 41748 767310
rect 41696 767246 41748 767252
rect 41236 766148 41288 766154
rect 41236 766090 41288 766096
rect 40868 764856 40920 764862
rect 40868 764798 40920 764804
rect 40880 763745 40908 764798
rect 41248 764561 41276 766090
rect 41510 764960 41566 764969
rect 41510 764895 41566 764904
rect 41524 764590 41552 764895
rect 41512 764584 41564 764590
rect 41234 764552 41290 764561
rect 41512 764526 41564 764532
rect 41234 764487 41290 764496
rect 40866 763736 40922 763745
rect 40866 763671 40922 763680
rect 41510 763328 41566 763337
rect 41510 763263 41512 763272
rect 41564 763263 41566 763272
rect 41512 763234 41564 763240
rect 41708 761161 41736 767246
rect 41694 761152 41750 761161
rect 41694 761087 41750 761096
rect 41512 761048 41564 761054
rect 41512 760990 41564 760996
rect 41524 758826 41552 760990
rect 41892 758985 41920 768590
rect 42706 768567 42762 768576
rect 42720 761274 42748 768567
rect 42720 761246 42840 761274
rect 42614 761152 42670 761161
rect 42614 761087 42670 761096
rect 41878 758976 41934 758985
rect 41878 758911 41934 758920
rect 42430 758976 42486 758985
rect 42430 758911 42486 758920
rect 41524 758798 42380 758826
rect 41604 757784 41656 757790
rect 39304 757726 39356 757732
rect 40038 757752 40094 757761
rect 40038 757687 40094 757696
rect 40682 757752 40738 757761
rect 41656 757732 41828 757738
rect 41604 757726 41828 757732
rect 41616 757710 41828 757726
rect 40682 757687 40738 757696
rect 38934 757480 38990 757489
rect 38934 757415 38990 757424
rect 41800 757081 41828 757710
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 42352 756650 42380 758798
rect 42168 756622 42380 756650
rect 42168 756226 42196 756622
rect 42444 756514 42472 758911
rect 42260 756486 42472 756514
rect 41878 755440 41934 755449
rect 41878 755375 41934 755384
rect 41892 755072 41920 755375
rect 42260 754406 42288 756486
rect 42628 756378 42656 761087
rect 42812 761002 42840 761246
rect 42352 756350 42656 756378
rect 42720 760974 42840 761002
rect 42352 755018 42380 756350
rect 42522 755168 42578 755177
rect 42522 755103 42578 755112
rect 42352 754990 42472 755018
rect 42182 754378 42288 754406
rect 42248 754316 42300 754322
rect 42248 754258 42300 754264
rect 42260 754066 42288 754258
rect 42076 754038 42288 754066
rect 42076 753780 42104 754038
rect 42248 753908 42300 753914
rect 42248 753850 42300 753856
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42168 751754 42196 751944
rect 42260 751890 42288 753850
rect 42260 751862 42380 751890
rect 42168 751726 42288 751754
rect 42062 751632 42118 751641
rect 42062 751567 42118 751576
rect 42076 751369 42104 751567
rect 42260 751210 42288 751726
rect 42076 751182 42288 751210
rect 42076 751097 42104 751182
rect 42062 751088 42118 751097
rect 42062 751023 42118 751032
rect 42352 750938 42380 751862
rect 42168 750910 42380 750938
rect 42168 750720 42196 750910
rect 41970 750408 42026 750417
rect 41970 750343 42026 750352
rect 41984 750108 42012 750343
rect 42444 750258 42472 754990
rect 42536 753494 42564 755103
rect 42536 753466 42656 753494
rect 42260 750230 42472 750258
rect 42260 749714 42288 750230
rect 42168 749686 42288 749714
rect 42168 749529 42196 749686
rect 42430 749592 42486 749601
rect 42430 749527 42486 749536
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 747062 42288 749391
rect 42182 747034 42288 747062
rect 42444 746594 42472 749527
rect 42076 746566 42472 746594
rect 42076 746401 42104 746566
rect 42628 746314 42656 753466
rect 42720 751958 42748 760974
rect 42904 756254 42932 795382
rect 43272 795274 43300 804526
rect 43088 795246 43300 795274
rect 43088 794850 43116 795246
rect 43364 794894 43392 812806
rect 43812 805996 43864 806002
rect 43812 805938 43864 805944
rect 43536 799128 43588 799134
rect 43536 799070 43588 799076
rect 43548 797337 43576 799070
rect 43534 797328 43590 797337
rect 43534 797263 43590 797272
rect 43536 795048 43588 795054
rect 43272 794866 43392 794894
rect 43456 794996 43536 795002
rect 43456 794990 43588 794996
rect 43456 794974 43576 794990
rect 43076 794844 43128 794850
rect 43076 794786 43128 794792
rect 43272 770302 43300 794866
rect 43456 793830 43484 794974
rect 43444 793824 43496 793830
rect 43444 793766 43496 793772
rect 43260 770296 43312 770302
rect 43260 770238 43312 770244
rect 43258 764144 43314 764153
rect 43258 764079 43314 764088
rect 43074 763736 43130 763745
rect 43074 763671 43130 763680
rect 43088 756254 43116 763671
rect 43272 763154 43300 764079
rect 42812 756226 42932 756254
rect 42996 756226 43116 756254
rect 43180 763126 43300 763154
rect 42812 753658 42840 756226
rect 42996 753914 43024 756226
rect 42984 753908 43036 753914
rect 42984 753850 43036 753856
rect 42812 753630 42932 753658
rect 42720 751930 42840 751958
rect 42812 751754 42840 751930
rect 42260 746286 42656 746314
rect 42720 751726 42840 751754
rect 42260 746042 42288 746286
rect 42720 746178 42748 751726
rect 42168 746014 42288 746042
rect 42352 746150 42748 746178
rect 42168 745756 42196 746014
rect 42352 745634 42380 746150
rect 42168 745606 42380 745634
rect 42168 745212 42196 745606
rect 42338 745376 42394 745385
rect 42338 745311 42394 745320
rect 42522 745376 42578 745385
rect 42522 745311 42578 745320
rect 42352 743390 42380 745311
rect 42536 745090 42564 745311
rect 42182 743362 42380 743390
rect 42444 745062 42564 745090
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42444 742710 42472 745062
rect 42706 744968 42762 744977
rect 42260 742682 42472 742710
rect 42536 744926 42706 744954
rect 42536 742098 42564 744926
rect 42706 744903 42762 744912
rect 42708 744048 42760 744054
rect 42708 743990 42760 743996
rect 42182 742070 42564 742098
rect 42720 741554 42748 743990
rect 42182 741526 42748 741554
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42246 730552 42302 730561
rect 42246 730487 42302 730496
rect 42260 729366 42288 730487
rect 42248 729360 42300 729366
rect 42248 729302 42300 729308
rect 41328 729088 41380 729094
rect 41328 729030 41380 729036
rect 41696 729088 41748 729094
rect 41696 729030 41748 729036
rect 41340 728691 41368 729030
rect 40866 728682 40922 728691
rect 40866 728617 40922 728626
rect 41326 728682 41382 728691
rect 41708 728668 41736 729030
rect 42064 728680 42116 728686
rect 41708 728640 42064 728668
rect 41326 728617 41382 728626
rect 42064 728622 42116 728628
rect 40880 727462 40908 728617
rect 40868 727456 40920 727462
rect 40868 727398 40920 727404
rect 41326 727458 41382 727467
rect 41326 727393 41382 727402
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727416 42064 727444
rect 41696 727398 41748 727404
rect 42064 727398 42116 727404
rect 41340 727326 41368 727393
rect 41328 727320 41380 727326
rect 41328 727262 41380 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727280 42064 727308
rect 41696 727262 41748 727268
rect 42064 727262 42116 727268
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 39302 726234 39358 726243
rect 39302 726169 39358 726178
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 31666 724432 31722 724441
rect 31666 724367 31722 724376
rect 31680 718321 31708 724367
rect 32954 724024 33010 724033
rect 32954 723959 33010 723968
rect 31666 718312 31722 718321
rect 31666 718247 31722 718256
rect 32968 715562 32996 723959
rect 33782 723208 33838 723217
rect 33782 723143 33838 723152
rect 33796 715698 33824 723143
rect 35176 715834 35204 724775
rect 39316 716145 39344 726169
rect 41156 725966 41184 726815
rect 41326 726234 41382 726243
rect 41326 726169 41382 726178
rect 41696 726232 41748 726238
rect 41748 726180 42196 726186
rect 41696 726174 42196 726180
rect 41708 726158 42196 726174
rect 41144 725960 41196 725966
rect 41144 725902 41196 725908
rect 41604 725960 41656 725966
rect 41604 725902 41656 725908
rect 41616 725778 41644 725902
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41142 725248 41198 725257
rect 41142 725183 41198 725192
rect 41156 720474 41184 725183
rect 41340 724514 41368 725591
rect 41340 724486 41552 724514
rect 41156 720446 41368 720474
rect 41142 720352 41198 720361
rect 41142 720287 41198 720296
rect 41156 717614 41184 720287
rect 41340 719273 41368 720446
rect 41326 719264 41382 719273
rect 41326 719199 41382 719208
rect 41156 717586 41276 717614
rect 39302 716136 39358 716145
rect 39302 716071 39358 716080
rect 35164 715828 35216 715834
rect 35164 715770 35216 715776
rect 40590 715728 40646 715737
rect 33784 715692 33836 715698
rect 33784 715634 33836 715640
rect 40408 715692 40460 715698
rect 40590 715663 40646 715672
rect 40408 715634 40460 715640
rect 32956 715556 33008 715562
rect 32956 715498 33008 715504
rect 40420 715465 40448 715634
rect 40604 715562 40632 715663
rect 40592 715556 40644 715562
rect 40592 715498 40644 715504
rect 40406 715456 40462 715465
rect 40406 715391 40462 715400
rect 41248 714241 41276 717586
rect 41524 714921 41552 724486
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41800 718593 41828 722327
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 42168 718434 42196 726158
rect 42904 724514 42932 753630
rect 43180 741074 43208 763126
rect 43442 757480 43498 757489
rect 43088 741046 43208 741074
rect 43272 757438 43442 757466
rect 43088 729337 43116 741046
rect 43074 729328 43130 729337
rect 43074 729263 43130 729272
rect 43076 728680 43128 728686
rect 43076 728622 43128 728628
rect 42720 724486 42932 724514
rect 42720 719438 42748 724486
rect 43088 719778 43116 728622
rect 43076 719772 43128 719778
rect 43076 719714 43128 719720
rect 42892 719568 42944 719574
rect 42892 719510 42944 719516
rect 42708 719432 42760 719438
rect 42708 719374 42760 719380
rect 42522 719264 42578 719273
rect 42522 719199 42578 719208
rect 41892 718406 42196 718434
rect 41696 715828 41748 715834
rect 41696 715770 41748 715776
rect 41510 714912 41566 714921
rect 41510 714847 41566 714856
rect 41708 714854 41736 715770
rect 41892 715034 41920 718406
rect 42246 715456 42302 715465
rect 42302 715414 42472 715442
rect 42246 715391 42302 715400
rect 41892 715006 42380 715034
rect 41708 714826 41828 714854
rect 41800 714762 41828 714826
rect 41800 714734 42288 714762
rect 41234 714232 41290 714241
rect 41234 714167 41290 714176
rect 42260 713062 42288 714734
rect 42182 713034 42288 713062
rect 41786 712192 41842 712201
rect 41786 712127 41842 712136
rect 41800 711824 41828 712127
rect 42352 711226 42380 715006
rect 42182 711198 42380 711226
rect 42062 710832 42118 710841
rect 42062 710767 42118 710776
rect 42076 710561 42104 710767
rect 42444 710002 42472 715414
rect 42260 709974 42472 710002
rect 42260 709866 42288 709974
rect 42076 709838 42288 709866
rect 42076 709376 42104 709838
rect 42248 709776 42300 709782
rect 42248 709718 42300 709724
rect 42076 708393 42104 708696
rect 42062 708384 42118 708393
rect 42062 708319 42118 708328
rect 42260 708234 42288 709718
rect 42536 709594 42564 719199
rect 42706 716000 42762 716009
rect 42706 715935 42762 715944
rect 42720 715850 42748 715935
rect 42168 708206 42288 708234
rect 42352 709566 42564 709594
rect 42628 715822 42748 715850
rect 42168 708152 42196 708206
rect 42352 708098 42380 709566
rect 42628 709390 42656 715822
rect 42904 715340 42932 719510
rect 43076 719432 43128 719438
rect 43128 719380 43208 719386
rect 43076 719374 43208 719380
rect 43088 719358 43208 719374
rect 42904 715312 43116 715340
rect 42798 714912 42854 714921
rect 42798 714854 42854 714856
rect 42444 709362 42656 709390
rect 42720 714847 42854 714854
rect 42720 714826 42840 714847
rect 42444 708710 42472 709362
rect 42720 708914 42748 714826
rect 42892 712156 42944 712162
rect 42892 712098 42944 712104
rect 42904 710841 42932 712098
rect 42890 710832 42946 710841
rect 42890 710767 42946 710776
rect 42720 708886 42932 708914
rect 42444 708682 42564 708710
rect 42352 708070 42472 708098
rect 42248 708008 42300 708014
rect 42248 707950 42300 707956
rect 42260 707554 42288 707950
rect 42182 707526 42288 707554
rect 41786 707160 41842 707169
rect 41786 707095 41842 707104
rect 41800 706860 41828 707095
rect 42444 706738 42472 708070
rect 42352 706710 42472 706738
rect 42352 706330 42380 706710
rect 42182 706302 42380 706330
rect 42248 705560 42300 705566
rect 42248 705502 42300 705508
rect 41786 704304 41842 704313
rect 41786 704239 41842 704248
rect 41800 703868 41828 704239
rect 42260 703610 42288 705502
rect 42168 703582 42288 703610
rect 42168 703188 42196 703582
rect 42536 702590 42564 708682
rect 42904 708506 42932 708886
rect 42168 702522 42196 702576
rect 42260 702562 42564 702590
rect 42628 708478 42932 708506
rect 42260 702522 42288 702562
rect 42168 702494 42288 702522
rect 42628 702386 42656 708478
rect 43088 705194 43116 715312
rect 42260 702358 42656 702386
rect 42904 705166 43116 705194
rect 42260 702250 42288 702358
rect 41984 702222 42288 702250
rect 41984 702032 42012 702222
rect 42706 702128 42762 702137
rect 42536 702086 42706 702114
rect 42246 701856 42302 701865
rect 42246 701791 42302 701800
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42260 699530 42288 701791
rect 42182 699502 42288 699530
rect 42536 698918 42564 702086
rect 42706 702063 42762 702072
rect 42708 701072 42760 701078
rect 42708 701014 42760 701020
rect 42168 698850 42196 698904
rect 42260 698890 42564 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42720 698339 42748 701014
rect 42904 700466 42932 705166
rect 43180 700482 43208 719358
rect 42892 700460 42944 700466
rect 42892 700402 42944 700408
rect 43088 700454 43208 700482
rect 43088 700398 43116 700454
rect 43076 700392 43128 700398
rect 43076 700334 43128 700340
rect 43076 700256 43128 700262
rect 43076 700198 43128 700204
rect 42892 700120 42944 700126
rect 42892 700062 42944 700068
rect 42182 698311 42748 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 42706 688120 42762 688129
rect 42706 688055 42762 688064
rect 42720 687342 42748 688055
rect 42708 687336 42760 687342
rect 42708 687278 42760 687284
rect 41142 686896 41198 686905
rect 41142 686831 41198 686840
rect 40866 686488 40922 686497
rect 40866 686423 40922 686432
rect 40880 685914 40908 686423
rect 41156 686118 41184 686831
rect 41328 686316 41380 686322
rect 41328 686258 41380 686264
rect 41696 686316 41748 686322
rect 42064 686316 42116 686322
rect 41748 686276 42064 686304
rect 41696 686258 41748 686264
rect 42064 686258 42116 686264
rect 41144 686112 41196 686118
rect 41144 686054 41196 686060
rect 41340 685919 41368 686258
rect 41696 686112 41748 686118
rect 42064 686112 42116 686118
rect 41748 686072 42064 686100
rect 41696 686054 41748 686060
rect 42064 686054 42116 686060
rect 40868 685908 40920 685914
rect 40868 685850 40920 685856
rect 41050 685910 41106 685919
rect 41050 685845 41106 685854
rect 41326 685910 41382 685919
rect 41326 685845 41382 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 41064 684758 41092 685845
rect 41052 684752 41104 684758
rect 40774 684686 40830 684695
rect 41052 684694 41104 684700
rect 41696 684752 41748 684758
rect 41696 684694 41748 684700
rect 40774 684621 40830 684630
rect 40788 683194 40816 684621
rect 41708 684321 41736 684694
rect 41694 684312 41750 684321
rect 41694 684247 41750 684256
rect 41142 684040 41198 684049
rect 41142 683975 41198 683984
rect 41156 683330 41184 683975
rect 41326 683462 41382 683471
rect 41326 683397 41382 683406
rect 41696 683460 41748 683466
rect 42064 683460 42116 683466
rect 41748 683420 42064 683448
rect 41696 683402 41748 683408
rect 42064 683402 42116 683408
rect 42708 683460 42760 683466
rect 42708 683402 42760 683408
rect 41144 683324 41196 683330
rect 41144 683266 41196 683272
rect 41696 683324 41748 683330
rect 42064 683324 42116 683330
rect 41748 683284 42064 683312
rect 41696 683266 41748 683272
rect 42064 683266 42116 683272
rect 41708 683194 42104 683210
rect 40776 683188 40828 683194
rect 40776 683130 40828 683136
rect 41696 683188 42116 683194
rect 41748 683182 42064 683188
rect 41696 683130 41748 683136
rect 42064 683130 42116 683136
rect 40958 682816 41014 682825
rect 40958 682751 41014 682760
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 32402 681184 32458 681193
rect 32402 681119 32458 681128
rect 32416 672761 32444 681119
rect 33782 680776 33838 680785
rect 33782 680711 33838 680720
rect 33796 672790 33824 680711
rect 35176 672926 35204 681935
rect 40972 679182 41000 682751
rect 41326 682408 41382 682417
rect 41326 682343 41382 682352
rect 41340 682038 41368 682343
rect 41328 682032 41380 682038
rect 41328 681974 41380 681980
rect 41696 682032 41748 682038
rect 42064 682032 42116 682038
rect 41748 681992 42064 682020
rect 41696 681974 41748 681980
rect 42064 681974 42116 681980
rect 42524 682032 42576 682038
rect 42524 681974 42576 681980
rect 42246 681592 42302 681601
rect 42246 681527 42302 681536
rect 41142 679960 41198 679969
rect 41142 679895 41198 679904
rect 40960 679176 41012 679182
rect 40960 679118 41012 679124
rect 41156 679046 41184 679895
rect 41328 679176 41380 679182
rect 41328 679118 41380 679124
rect 41144 679040 41196 679046
rect 41144 678982 41196 678988
rect 41340 678858 41368 679118
rect 41696 679040 41748 679046
rect 42064 679040 42116 679046
rect 41748 679000 42064 679028
rect 41696 678982 41748 678988
rect 42064 678982 42116 678988
rect 41786 678872 41842 678881
rect 41340 678830 41786 678858
rect 41786 678807 41842 678816
rect 41786 678328 41842 678337
rect 41616 678286 41786 678314
rect 40958 677750 41014 677759
rect 41616 677754 41644 678286
rect 41786 678263 41842 678272
rect 40958 677685 41014 677694
rect 41604 677748 41656 677754
rect 41604 677690 41656 677696
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 35164 672920 35216 672926
rect 35164 672862 35216 672868
rect 38844 672920 38896 672926
rect 38844 672862 38896 672868
rect 33784 672784 33836 672790
rect 32402 672752 32458 672761
rect 33784 672726 33836 672732
rect 37924 672784 37976 672790
rect 37924 672726 37976 672732
rect 32402 672687 32458 672696
rect 37936 671537 37964 672726
rect 37922 671528 37978 671537
rect 37922 671463 37978 671472
rect 38856 670993 38884 672862
rect 39960 672489 39988 677039
rect 39946 672480 40002 672489
rect 39946 672415 40002 672424
rect 38842 670984 38898 670993
rect 38842 670919 38898 670928
rect 42260 670290 42288 681527
rect 42536 674778 42564 681974
rect 42720 674834 42748 683402
rect 42904 674834 42932 700062
rect 43088 686322 43116 700198
rect 43076 686316 43128 686322
rect 43076 686258 43128 686264
rect 43074 677920 43130 677929
rect 43074 677855 43130 677864
rect 42444 674750 42564 674778
rect 42628 674806 42748 674834
rect 42812 674806 42932 674834
rect 42444 671566 42472 674750
rect 42432 671560 42484 671566
rect 42432 671502 42484 671508
rect 42628 671378 42656 674806
rect 42076 670262 42288 670290
rect 42352 671350 42656 671378
rect 42812 671378 42840 674806
rect 42812 671350 42932 671378
rect 42076 669868 42104 670262
rect 41786 669080 41842 669089
rect 41786 669015 41842 669024
rect 41800 668644 41828 669015
rect 42352 668046 42380 671350
rect 42708 671152 42760 671158
rect 42760 671100 42840 671106
rect 42708 671094 42840 671100
rect 42720 671078 42840 671094
rect 42522 670984 42578 670993
rect 42522 670919 42578 670928
rect 42168 667978 42196 668032
rect 42260 668018 42380 668046
rect 42260 667978 42288 668018
rect 42168 667950 42288 667978
rect 42536 667944 42564 670919
rect 42444 667916 42564 667944
rect 42248 667480 42300 667486
rect 42248 667422 42300 667428
rect 42260 667366 42288 667422
rect 42182 667338 42288 667366
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42444 666482 42472 667916
rect 42812 666482 42840 671078
rect 42444 666454 42656 666482
rect 42338 666360 42394 666369
rect 42394 666318 42564 666346
rect 42338 666295 42394 666304
rect 42340 665848 42392 665854
rect 42340 665790 42392 665796
rect 42352 665530 42380 665790
rect 42182 665502 42380 665530
rect 42248 665440 42300 665446
rect 42248 665382 42300 665388
rect 41786 665272 41842 665281
rect 41786 665207 41842 665216
rect 41800 664972 41828 665207
rect 42260 665174 42288 665382
rect 42260 665146 42472 665174
rect 42444 664339 42472 665146
rect 42182 664311 42472 664339
rect 41786 664184 41842 664193
rect 41786 664119 41842 664128
rect 41800 663680 41828 664119
rect 42536 663694 42564 666318
rect 42444 663666 42564 663694
rect 42444 663610 42472 663666
rect 42432 663604 42484 663610
rect 42432 663546 42484 663552
rect 42628 663354 42656 666454
rect 42444 663326 42656 663354
rect 42720 666454 42840 666482
rect 42444 663218 42472 663326
rect 42260 663190 42472 663218
rect 42260 663150 42288 663190
rect 42182 663122 42288 663150
rect 42432 663128 42484 663134
rect 42432 663070 42484 663076
rect 42154 662824 42210 662833
rect 42154 662759 42210 662768
rect 42168 662674 42196 662759
rect 42168 662646 42288 662674
rect 42260 661042 42288 662646
rect 42168 661014 42288 661042
rect 42168 660620 42196 661014
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42444 659371 42472 663070
rect 42182 659343 42472 659371
rect 42168 658838 42380 658866
rect 42168 658784 42196 658838
rect 42352 658798 42380 658838
rect 42720 658798 42748 666454
rect 42352 658770 42748 658798
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657280 42576 657286
rect 42524 657222 42576 657228
rect 42260 655642 42380 655670
rect 42536 655126 42564 657222
rect 42182 655098 42564 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 39578 644736 39634 644745
rect 39578 644671 39634 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35622 642696 35678 642705
rect 35622 642631 35678 642640
rect 35636 642054 35664 642631
rect 38580 642530 38608 644263
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 35806 642288 35862 642297
rect 35806 642223 35862 642232
rect 35624 642048 35676 642054
rect 35624 641990 35676 641996
rect 35820 641782 35848 642223
rect 39592 642054 39620 644671
rect 41696 644496 41748 644502
rect 42064 644496 42116 644502
rect 41748 644446 42064 644474
rect 41696 644438 41748 644444
rect 42064 644438 42116 644444
rect 40500 643544 40552 643550
rect 40498 643512 40500 643521
rect 40552 643512 40554 643521
rect 40498 643447 40554 643456
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 39580 642048 39632 642054
rect 39580 641990 39632 641996
rect 35808 641776 35860 641782
rect 35808 641718 35860 641724
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 35346 641472 35402 641481
rect 35346 641407 35402 641416
rect 35360 640490 35388 641407
rect 35530 641064 35586 641073
rect 35530 640999 35586 641008
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 35348 640484 35400 640490
rect 35348 640426 35400 640432
rect 35544 640354 35572 640999
rect 35820 640762 35848 640999
rect 35808 640756 35860 640762
rect 35808 640698 35860 640704
rect 39948 640756 40000 640762
rect 39948 640698 40000 640704
rect 35532 640348 35584 640354
rect 35532 640290 35584 640296
rect 39960 640257 39988 640698
rect 41696 640552 41748 640558
rect 42064 640552 42116 640558
rect 41748 640500 42064 640506
rect 41696 640494 42116 640500
rect 41708 640478 42104 640494
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 39946 640248 40002 640257
rect 39946 640183 40002 640192
rect 35806 639840 35862 639849
rect 35806 639775 35862 639784
rect 35820 639198 35848 639775
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 37924 639124 37976 639130
rect 37924 639066 37976 639072
rect 35806 639024 35862 639033
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 35808 638930 35860 638936
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 35162 637800 35218 637809
rect 35162 637735 35218 637744
rect 32034 636984 32090 636993
rect 32034 636919 32090 636928
rect 32048 629950 32076 636919
rect 32036 629944 32088 629950
rect 35176 629921 35204 637735
rect 35636 636886 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637634 35848 638143
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 36544 637628 36596 637634
rect 36544 637570 36596 637576
rect 35624 636880 35676 636886
rect 35624 636822 35676 636828
rect 35530 636576 35586 636585
rect 35530 636511 35532 636520
rect 35584 636511 35586 636520
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35532 636482 35584 636488
rect 35820 636274 35848 636511
rect 35808 636268 35860 636274
rect 35808 636210 35860 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634982 35848 635695
rect 35808 634976 35860 634982
rect 35808 634918 35860 634924
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633758 35848 634471
rect 35808 633752 35860 633758
rect 35808 633694 35860 633700
rect 35808 633480 35860 633486
rect 35808 633422 35860 633428
rect 35820 633321 35848 633422
rect 35806 633312 35862 633321
rect 35806 633247 35862 633256
rect 36556 630766 36584 637570
rect 36544 630760 36596 630766
rect 36544 630702 36596 630708
rect 37740 629944 37792 629950
rect 32036 629886 32088 629892
rect 35162 629912 35218 629921
rect 37740 629886 37792 629892
rect 35162 629847 35218 629856
rect 37752 629649 37780 629886
rect 37738 629640 37794 629649
rect 37738 629575 37794 629584
rect 37936 627745 37964 639066
rect 41696 638920 41748 638926
rect 41696 638862 41748 638868
rect 41708 637574 41736 638862
rect 41708 637546 42104 637574
rect 39120 636880 39172 636886
rect 39120 636822 39172 636828
rect 39132 636585 39160 636822
rect 39118 636576 39174 636585
rect 39118 636511 39174 636520
rect 39764 636540 39816 636546
rect 39764 636482 39816 636488
rect 39120 633752 39172 633758
rect 39120 633694 39172 633700
rect 39132 630465 39160 633694
rect 39776 632233 39804 636482
rect 39948 636268 40000 636274
rect 39948 636210 40000 636216
rect 39960 633729 39988 636210
rect 41420 634976 41472 634982
rect 41420 634918 41472 634924
rect 39946 633720 40002 633729
rect 39946 633655 40002 633664
rect 40408 633480 40460 633486
rect 40408 633422 40460 633428
rect 39762 632224 39818 632233
rect 39762 632159 39818 632168
rect 40420 630737 40448 633422
rect 41432 631417 41460 634918
rect 41878 633924 41934 633933
rect 41878 633859 41934 633868
rect 41418 631408 41474 631417
rect 41418 631343 41474 631352
rect 41512 630760 41564 630766
rect 40406 630728 40462 630737
rect 41512 630702 41564 630708
rect 40406 630663 40462 630672
rect 39118 630456 39174 630465
rect 39118 630391 39174 630400
rect 41524 628674 41552 630702
rect 41524 628646 41828 628674
rect 37922 627736 37978 627745
rect 37922 627671 37978 627680
rect 41800 627473 41828 628646
rect 41892 627586 41920 633859
rect 42076 629542 42104 637546
rect 42522 636576 42578 636585
rect 42522 636511 42578 636520
rect 42338 629640 42394 629649
rect 42338 629575 42394 629584
rect 42064 629536 42116 629542
rect 42064 629478 42116 629484
rect 42352 629252 42380 629575
rect 42536 629354 42564 636511
rect 42708 629536 42760 629542
rect 42708 629478 42760 629484
rect 42536 629326 42656 629354
rect 42352 629224 42564 629252
rect 42536 628946 42564 629224
rect 42444 628918 42564 628946
rect 42062 627736 42118 627745
rect 42118 627694 42380 627722
rect 42062 627671 42118 627680
rect 41892 627558 42288 627586
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 41786 627192 41842 627201
rect 41786 627127 41842 627136
rect 41800 626620 41828 627127
rect 42260 625478 42288 627558
rect 42182 625450 42288 625478
rect 42352 625274 42380 627694
rect 42260 625246 42380 625274
rect 42260 625138 42288 625246
rect 42168 625110 42288 625138
rect 42168 624784 42196 625110
rect 42444 624753 42472 628918
rect 42628 627914 42656 629326
rect 42536 627886 42656 627914
rect 42536 624866 42564 627886
rect 42720 625682 42748 629478
rect 42904 627914 42932 671350
rect 42812 627886 42932 627914
rect 42812 625954 42840 627886
rect 42812 625926 43024 625954
rect 42720 625654 42932 625682
rect 42536 624838 42656 624866
rect 42430 624744 42486 624753
rect 42430 624679 42486 624688
rect 42340 624504 42392 624510
rect 42062 624472 42118 624481
rect 42340 624446 42392 624452
rect 42062 624407 42118 624416
rect 42076 624172 42104 624407
rect 42062 623792 42118 623801
rect 42118 623750 42288 623778
rect 42062 623727 42118 623736
rect 42062 623384 42118 623393
rect 42062 623319 42118 623328
rect 42076 622948 42104 623319
rect 42076 622169 42104 622336
rect 42062 622160 42118 622169
rect 42062 622095 42118 622104
rect 42168 621738 42196 621792
rect 42260 621738 42288 623750
rect 42168 621710 42288 621738
rect 42352 621602 42380 624446
rect 42628 623778 42656 624838
rect 42168 621574 42380 621602
rect 42536 623750 42656 623778
rect 42168 621112 42196 621574
rect 42536 621126 42564 623750
rect 42444 621098 42564 621126
rect 41786 620800 41842 620809
rect 41786 620735 41842 620744
rect 41800 620500 41828 620735
rect 42076 620078 42288 620106
rect 42076 619956 42104 620078
rect 42260 619970 42288 620078
rect 42444 619970 42472 621098
rect 42904 621014 42932 625654
rect 42628 620986 42932 621014
rect 42628 620922 42656 620986
rect 42260 619942 42472 619970
rect 42536 620894 42656 620922
rect 42246 619848 42302 619857
rect 42302 619806 42472 619834
rect 42246 619783 42302 619792
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 617454 42288 619618
rect 42182 617426 42288 617454
rect 42156 617296 42208 617302
rect 42156 617238 42208 617244
rect 42168 616978 42196 617238
rect 42076 616950 42196 616978
rect 42076 616828 42104 616950
rect 42444 616570 42472 619806
rect 42536 616842 42564 620894
rect 42706 620800 42762 620809
rect 42706 620735 42762 620744
rect 42720 617302 42748 620735
rect 42996 618338 43024 625926
rect 42904 618310 43024 618338
rect 42708 617296 42760 617302
rect 42708 617238 42760 617244
rect 42536 616814 42748 616842
rect 42168 616542 42472 616570
rect 42168 616148 42196 616542
rect 42338 616312 42394 616321
rect 42338 616247 42394 616256
rect 42352 616162 42380 616247
rect 42260 616134 42380 616162
rect 42062 615768 42118 615777
rect 42062 615703 42118 615712
rect 42076 615604 42104 615703
rect 42260 613782 42288 616134
rect 42522 616040 42578 616049
rect 42182 613754 42288 613782
rect 42352 615998 42522 616026
rect 42352 613135 42380 615998
rect 42522 615975 42578 615984
rect 42720 615777 42748 616814
rect 42706 615768 42762 615777
rect 42706 615703 42762 615712
rect 42522 615496 42578 615505
rect 42522 615431 42578 615440
rect 42536 615346 42564 615431
rect 42182 613107 42380 613135
rect 42444 615318 42564 615346
rect 42444 612490 42472 615318
rect 42616 614168 42668 614174
rect 42616 614110 42668 614116
rect 42182 612462 42472 612490
rect 42628 611946 42656 614110
rect 42904 614009 42932 618310
rect 43088 614310 43116 677855
rect 43076 614304 43128 614310
rect 43076 614246 43128 614252
rect 42890 614000 42946 614009
rect 42890 613935 42946 613944
rect 43272 612241 43300 757438
rect 43442 757415 43498 757424
rect 43444 754928 43496 754934
rect 43444 754870 43496 754876
rect 43456 753001 43484 754870
rect 43628 753704 43680 753710
rect 43628 753646 43680 753652
rect 43442 752992 43498 753001
rect 43442 752927 43498 752936
rect 43640 751641 43668 753646
rect 43626 751632 43682 751641
rect 43626 751567 43682 751576
rect 43442 731368 43498 731377
rect 43442 731303 43498 731312
rect 43456 730386 43484 731303
rect 43444 730380 43496 730386
rect 43444 730322 43496 730328
rect 43626 723616 43682 723625
rect 43626 723551 43682 723560
rect 43640 705566 43668 723551
rect 43628 705560 43680 705566
rect 43628 705502 43680 705508
rect 43442 687304 43498 687313
rect 43442 687239 43498 687248
rect 43456 686526 43484 687239
rect 43444 686520 43496 686526
rect 43444 686462 43496 686468
rect 43626 680368 43682 680377
rect 43626 680303 43682 680312
rect 43442 676696 43498 676705
rect 43442 676631 43498 676640
rect 43258 612232 43314 612241
rect 43258 612167 43314 612176
rect 42182 611918 42656 611946
rect 43456 611402 43484 676631
rect 43640 669314 43668 680303
rect 43548 669286 43668 669314
rect 43548 665174 43576 669286
rect 43548 665146 43668 665174
rect 43640 660550 43668 665146
rect 43628 660544 43680 660550
rect 43628 660486 43680 660492
rect 43824 630674 43852 805938
rect 44284 774761 44312 815730
rect 44824 815652 44876 815658
rect 44824 815594 44876 815600
rect 44548 814428 44600 814434
rect 44548 814370 44600 814376
rect 44270 774752 44326 774761
rect 44270 774687 44326 774696
rect 44560 771458 44588 814370
rect 44836 806614 44864 815594
rect 45100 814292 45152 814298
rect 45100 814234 45152 814240
rect 44824 806608 44876 806614
rect 44824 806550 44876 806556
rect 44916 806472 44968 806478
rect 44916 806414 44968 806420
rect 44928 795054 44956 806414
rect 44916 795048 44968 795054
rect 44916 794990 44968 794996
rect 44914 772848 44970 772857
rect 44914 772783 44970 772792
rect 44548 771452 44600 771458
rect 44548 771394 44600 771400
rect 44546 770264 44602 770273
rect 44546 770199 44602 770208
rect 44272 770092 44324 770098
rect 44272 770034 44324 770040
rect 44284 736934 44312 770034
rect 44284 736906 44404 736934
rect 44178 728104 44234 728113
rect 44178 728039 44234 728048
rect 44192 724514 44220 728039
rect 44376 727705 44404 736906
rect 44362 727696 44418 727705
rect 44362 727631 44418 727640
rect 44560 727462 44588 770199
rect 44732 755540 44784 755546
rect 44732 755482 44784 755488
rect 44744 754322 44772 755482
rect 44732 754316 44784 754322
rect 44732 754258 44784 754264
rect 44928 730153 44956 772783
rect 45112 771662 45140 814234
rect 45284 807356 45336 807362
rect 45284 807298 45336 807304
rect 45296 806478 45324 807298
rect 45284 806472 45336 806478
rect 45284 806414 45336 806420
rect 46216 785194 46244 817090
rect 61384 817012 61436 817018
rect 61384 816954 61436 816960
rect 53104 799128 53156 799134
rect 53104 799070 53156 799076
rect 53116 790770 53144 799070
rect 57244 797700 57296 797706
rect 57244 797642 57296 797648
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 57256 789206 57284 797642
rect 57244 789200 57296 789206
rect 57244 789142 57296 789148
rect 61396 786185 61424 816954
rect 62764 806608 62816 806614
rect 62764 806550 62816 806556
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 62120 789200 62172 789206
rect 62118 789168 62120 789177
rect 62172 789168 62174 789177
rect 62118 789103 62174 789112
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62776 787137 62804 806550
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 62762 787128 62818 787137
rect 62762 787063 62818 787072
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 61382 786176 61438 786185
rect 61382 786111 61438 786120
rect 46204 785188 46256 785194
rect 46204 785130 46256 785136
rect 62120 785188 62172 785194
rect 62120 785130 62172 785136
rect 62132 784961 62160 785130
rect 62118 784952 62174 784961
rect 62118 784887 62174 784896
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775606 651512 776047
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 60004 774240 60056 774246
rect 60004 774182 60056 774188
rect 651470 774208 651526 774217
rect 46202 773120 46258 773129
rect 46202 773055 46258 773064
rect 45100 771656 45152 771662
rect 45100 771598 45152 771604
rect 45098 764960 45154 764969
rect 45098 764895 45154 764904
rect 45112 753710 45140 764895
rect 45282 764552 45338 764561
rect 45282 764487 45338 764496
rect 45296 754934 45324 764487
rect 45558 763328 45614 763337
rect 45558 763263 45614 763272
rect 45284 754928 45336 754934
rect 45284 754870 45336 754876
rect 45100 753704 45152 753710
rect 45100 753646 45152 753652
rect 45098 751088 45154 751097
rect 45098 751023 45154 751032
rect 45112 746570 45140 751023
rect 45100 746564 45152 746570
rect 45100 746506 45152 746512
rect 44914 730144 44970 730153
rect 44914 730079 44970 730088
rect 45190 729736 45246 729745
rect 45190 729671 45246 729680
rect 44548 727456 44600 727462
rect 44548 727398 44600 727404
rect 45008 727320 45060 727326
rect 45008 727262 45060 727268
rect 44192 724486 44312 724514
rect 44284 685273 44312 724486
rect 44454 722800 44510 722809
rect 44454 722735 44510 722744
rect 44468 708710 44496 722735
rect 44638 721576 44694 721585
rect 44638 721511 44694 721520
rect 44652 709782 44680 721511
rect 44640 709776 44692 709782
rect 44640 709718 44692 709724
rect 44468 708682 44680 708710
rect 44454 708384 44510 708393
rect 44454 708319 44510 708328
rect 44468 703798 44496 708319
rect 44652 708014 44680 708682
rect 44640 708008 44692 708014
rect 44640 707950 44692 707956
rect 44456 703792 44508 703798
rect 44456 703734 44508 703740
rect 44822 687712 44878 687721
rect 44822 687647 44878 687656
rect 44270 685264 44326 685273
rect 44270 685199 44326 685208
rect 44454 684312 44510 684321
rect 44454 684247 44510 684256
rect 44272 683324 44324 683330
rect 44272 683266 44324 683272
rect 43994 679552 44050 679561
rect 43994 679487 44050 679496
rect 44008 665446 44036 679487
rect 43996 665440 44048 665446
rect 43996 665382 44048 665388
rect 44284 640354 44312 683266
rect 44468 644745 44496 684247
rect 44638 683904 44694 683913
rect 44638 683839 44694 683848
rect 44454 644736 44510 644745
rect 44454 644671 44510 644680
rect 44652 641782 44680 683839
rect 44836 655518 44864 687647
rect 45020 683194 45048 727262
rect 45204 686118 45232 729671
rect 45192 686112 45244 686118
rect 45192 686054 45244 686060
rect 45192 685908 45244 685914
rect 45192 685850 45244 685856
rect 45008 683188 45060 683194
rect 45008 683130 45060 683136
rect 45008 679040 45060 679046
rect 45008 678982 45060 678988
rect 45020 666641 45048 678982
rect 45006 666632 45062 666641
rect 45006 666567 45062 666576
rect 44824 655512 44876 655518
rect 44824 655454 44876 655460
rect 45006 643512 45062 643521
rect 45006 643447 45062 643456
rect 44640 641776 44692 641782
rect 44640 641718 44692 641724
rect 44640 640552 44692 640558
rect 44640 640494 44692 640500
rect 44272 640348 44324 640354
rect 44272 640290 44324 640296
rect 44362 633720 44418 633729
rect 44362 633655 44418 633664
rect 43994 632224 44050 632233
rect 43994 632159 44050 632168
rect 43824 630646 43944 630674
rect 43718 630456 43774 630465
rect 43718 630391 43774 630400
rect 43732 612626 43760 630391
rect 43916 612746 43944 630646
rect 44008 627914 44036 632159
rect 44178 631408 44234 631417
rect 44178 631343 44234 631352
rect 44008 627886 44128 627914
rect 44100 623393 44128 627886
rect 44192 623778 44220 631343
rect 44376 624510 44404 633655
rect 44364 624504 44416 624510
rect 44364 624446 44416 624452
rect 44192 623750 44588 623778
rect 44086 623384 44142 623393
rect 44086 623319 44142 623328
rect 44560 623234 44588 623750
rect 44192 623206 44588 623234
rect 44192 619682 44220 623206
rect 44362 622160 44418 622169
rect 44362 622095 44418 622104
rect 44180 619676 44232 619682
rect 44180 619618 44232 619624
rect 44376 616826 44404 622095
rect 44364 616820 44416 616826
rect 44364 616762 44416 616768
rect 44456 614304 44508 614310
rect 44456 614246 44508 614252
rect 44086 614000 44142 614009
rect 44086 613935 44142 613944
rect 43904 612740 43956 612746
rect 43904 612682 43956 612688
rect 43732 612598 43944 612626
rect 43764 612232 43820 612241
rect 43764 612167 43766 612176
rect 43818 612167 43820 612176
rect 43766 612138 43818 612144
rect 43916 611946 43944 612598
rect 44100 612406 44128 613935
rect 44088 612400 44140 612406
rect 44088 612342 44140 612348
rect 44086 612096 44142 612105
rect 44086 612031 44088 612040
rect 44140 612031 44142 612040
rect 44088 612002 44140 612008
rect 43916 611918 44312 611946
rect 43994 611824 44050 611833
rect 43994 611759 43996 611768
rect 44048 611759 44050 611768
rect 43996 611730 44048 611736
rect 44284 611658 44312 611918
rect 44272 611652 44324 611658
rect 44272 611594 44324 611600
rect 44088 611584 44140 611590
rect 44086 611552 44088 611561
rect 44140 611552 44142 611561
rect 44086 611487 44142 611496
rect 43456 611386 44251 611402
rect 43456 611380 44263 611386
rect 43456 611374 44211 611380
rect 44211 611322 44263 611328
rect 44468 611266 44496 614246
rect 44330 611238 44496 611266
rect 44330 611182 44358 611238
rect 44318 611176 44370 611182
rect 44318 611118 44370 611124
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 35806 601760 35862 601769
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 36544 601724 36596 601730
rect 35808 601666 35860 601672
rect 36544 601666 36596 601672
rect 35622 595810 35678 595819
rect 35622 595745 35678 595754
rect 33046 595232 33102 595241
rect 33046 595167 33102 595176
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595167
rect 33782 593600 33838 593609
rect 33782 593535 33838 593544
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 33796 585954 33824 593535
rect 35636 587314 35664 595745
rect 36556 593094 36584 601666
rect 38566 601352 38622 601361
rect 38566 601287 38622 601296
rect 38580 594318 38608 601287
rect 39946 600944 40002 600953
rect 39946 600879 40002 600888
rect 39960 595814 39988 600879
rect 44652 598913 44680 640494
rect 44822 630728 44878 630737
rect 44822 630663 44878 630672
rect 44836 627914 44864 630663
rect 44836 627886 44956 627914
rect 44928 611354 44956 627886
rect 44836 611326 44956 611354
rect 44836 611250 44864 611326
rect 44824 611244 44876 611250
rect 44824 611186 44876 611192
rect 45020 600545 45048 643447
rect 45204 643346 45232 685850
rect 45376 669384 45428 669390
rect 45376 669326 45428 669332
rect 45388 667486 45416 669326
rect 45376 667480 45428 667486
rect 45376 667422 45428 667428
rect 45192 643340 45244 643346
rect 45192 643282 45244 643288
rect 45282 640248 45338 640257
rect 45282 640183 45338 640192
rect 45006 600536 45062 600545
rect 45006 600471 45062 600480
rect 45098 600128 45154 600137
rect 45098 600063 45154 600072
rect 44638 598904 44694 598913
rect 44638 598839 44694 598848
rect 44914 598496 44970 598505
rect 44914 598431 44970 598440
rect 42890 597680 42946 597689
rect 42890 597615 42946 597624
rect 42904 597446 42932 597615
rect 42892 597440 42944 597446
rect 42892 597382 42944 597388
rect 42892 597032 42944 597038
rect 42892 596974 42944 596980
rect 43074 597000 43130 597009
rect 42430 596864 42486 596873
rect 42430 596799 42486 596808
rect 41142 596456 41198 596465
rect 41142 596391 41198 596400
rect 39948 595808 40000 595814
rect 39948 595750 40000 595756
rect 39302 594824 39358 594833
rect 39302 594759 39358 594768
rect 38568 594312 38620 594318
rect 38568 594254 38620 594260
rect 36544 593088 36596 593094
rect 36544 593030 36596 593036
rect 35624 587308 35676 587314
rect 35624 587250 35676 587256
rect 33784 585948 33836 585954
rect 33784 585890 33836 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 39316 585177 39344 594759
rect 41156 591410 41184 596391
rect 41970 596048 42026 596057
rect 41970 595983 42026 595992
rect 41696 595808 41748 595814
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41694 595711 41750 595720
rect 41604 594312 41656 594318
rect 41786 594280 41842 594289
rect 41656 594260 41786 594266
rect 41604 594254 41786 594260
rect 41616 594238 41786 594254
rect 41786 594215 41842 594224
rect 41696 593088 41748 593094
rect 41696 593030 41748 593036
rect 41708 592929 41736 593030
rect 41694 592920 41750 592929
rect 41694 592855 41750 592864
rect 41156 591382 41552 591410
rect 41524 591274 41552 591382
rect 41694 591288 41750 591297
rect 41524 591246 41694 591274
rect 41694 591223 41750 591232
rect 41050 590744 41106 590753
rect 41050 590679 41106 590688
rect 39580 587308 39632 587314
rect 39580 587250 39632 587256
rect 39592 585857 39620 587250
rect 40224 585948 40276 585954
rect 40224 585890 40276 585896
rect 39578 585848 39634 585857
rect 39578 585783 39634 585792
rect 39948 585812 40000 585818
rect 39948 585754 40000 585760
rect 39302 585168 39358 585177
rect 39302 585103 39358 585112
rect 39960 584633 39988 585754
rect 40236 584905 40264 585890
rect 41064 585449 41092 590679
rect 41420 587172 41472 587178
rect 41420 587114 41472 587120
rect 41050 585440 41106 585449
rect 41050 585375 41106 585384
rect 40222 584896 40278 584905
rect 40222 584831 40278 584840
rect 39946 584624 40002 584633
rect 39946 584559 40002 584568
rect 41432 584474 41460 587114
rect 41984 586129 42012 595983
rect 41970 586120 42026 586129
rect 41970 586055 42026 586064
rect 42154 585848 42210 585857
rect 42154 585783 42156 585792
rect 42208 585783 42210 585792
rect 42156 585754 42208 585760
rect 42246 585440 42302 585449
rect 42246 585375 42302 585384
rect 42260 584882 42288 585375
rect 42444 585120 42472 596799
rect 42708 585812 42760 585818
rect 42708 585754 42760 585760
rect 42720 585698 42748 585754
rect 42720 585670 42840 585698
rect 42444 585092 42564 585120
rect 42260 584854 42472 584882
rect 41432 584446 41828 584474
rect 41800 584361 41828 584446
rect 41786 584352 41842 584361
rect 41786 584287 41842 584296
rect 41786 583944 41842 583953
rect 41786 583879 41842 583888
rect 41800 583440 41828 583879
rect 42444 582263 42472 584854
rect 42182 582235 42472 582263
rect 42536 581754 42564 585092
rect 42444 581726 42564 581754
rect 42444 581618 42472 581726
rect 42182 581590 42472 581618
rect 42614 581632 42670 581641
rect 42614 581567 42670 581576
rect 42338 581224 42394 581233
rect 42338 581159 42394 581168
rect 42076 580689 42104 580961
rect 42062 580680 42118 580689
rect 42062 580615 42118 580624
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42168 578921 42196 579121
rect 42154 578912 42210 578921
rect 42154 578847 42210 578856
rect 42352 578626 42380 581159
rect 42168 578598 42380 578626
rect 42168 578544 42196 578598
rect 42628 578354 42656 581567
rect 42812 579614 42840 585670
rect 42536 578326 42656 578354
rect 42720 579586 42840 579614
rect 42248 578264 42300 578270
rect 42248 578206 42300 578212
rect 42062 578096 42118 578105
rect 42062 578031 42118 578040
rect 42076 577932 42104 578031
rect 41786 577824 41842 577833
rect 41786 577759 41842 577768
rect 41800 577281 41828 577759
rect 42260 576858 42288 578206
rect 42168 576830 42288 576858
rect 42168 576708 42196 576830
rect 42246 575784 42302 575793
rect 42246 575719 42302 575728
rect 41786 574696 41842 574705
rect 41786 574631 41842 574640
rect 41800 574260 41828 574631
rect 42260 573866 42288 575719
rect 42168 573838 42288 573866
rect 42168 573580 42196 573838
rect 42536 573594 42564 578326
rect 42720 578270 42748 579586
rect 42708 578264 42760 578270
rect 42708 578206 42760 578212
rect 42536 573566 42656 573594
rect 42628 573510 42656 573566
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42616 573504 42668 573510
rect 42616 573446 42668 573452
rect 42168 572968 42196 573446
rect 42614 572792 42670 572801
rect 42614 572727 42670 572736
rect 41984 572257 42012 572424
rect 41970 572248 42026 572257
rect 41970 572183 42026 572192
rect 42062 571568 42118 571577
rect 42062 571503 42118 571512
rect 42076 571282 42104 571503
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42076 571254 42380 571282
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42352 569310 42380 571254
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 571367
rect 42628 570994 42656 572727
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 42904 567194 42932 596974
rect 43074 596935 43130 596944
rect 43088 582374 43116 596935
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 44178 591968 44234 591977
rect 44178 591903 44234 591912
rect 43350 591560 43406 591569
rect 43350 591495 43406 591504
rect 42812 567166 42932 567194
rect 42996 582346 43116 582374
rect 43364 582374 43392 591495
rect 43626 590336 43682 590345
rect 43626 590271 43682 590280
rect 43364 582346 43484 582374
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 42246 558104 42302 558113
rect 42246 558039 42302 558048
rect 40038 553408 40094 553417
rect 40038 553343 40094 553352
rect 40866 553408 40922 553417
rect 40922 553366 41092 553394
rect 40866 553343 40922 553352
rect 34426 551984 34482 551993
rect 34426 551919 34482 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 34440 544406 34468 551919
rect 40052 551002 40080 553343
rect 40040 550996 40092 551002
rect 40040 550938 40092 550944
rect 41064 550610 41092 553366
rect 42260 552673 42288 558039
rect 42812 554849 42840 567166
rect 42996 556481 43024 582346
rect 42982 556472 43038 556481
rect 42982 556407 43038 556416
rect 42798 554840 42854 554849
rect 42798 554775 42854 554784
rect 42246 552664 42302 552673
rect 42246 552599 42302 552608
rect 42982 552392 43038 552401
rect 42982 552327 43038 552336
rect 42798 551168 42854 551177
rect 42798 551103 42854 551112
rect 41696 550996 41748 551002
rect 41748 550956 42380 550984
rect 41696 550938 41748 550944
rect 41786 550624 41842 550633
rect 41064 550582 41786 550610
rect 41786 550559 41842 550568
rect 41878 550352 41934 550361
rect 41878 550287 41934 550296
rect 41604 547460 41656 547466
rect 41604 547402 41656 547408
rect 41616 545578 41644 547402
rect 41892 545737 41920 550287
rect 42062 549944 42118 549953
rect 42062 549879 42118 549888
rect 41878 545728 41934 545737
rect 41878 545663 41934 545672
rect 41616 545550 41828 545578
rect 34428 544400 34480 544406
rect 34428 544342 34480 544348
rect 37832 544400 37884 544406
rect 37832 544342 37884 544348
rect 37844 541385 37872 544342
rect 37830 541376 37886 541385
rect 37830 541311 37886 541320
rect 41800 541113 41828 545550
rect 42076 545465 42104 549879
rect 42062 545456 42118 545465
rect 42062 545391 42118 545400
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42352 540818 42380 550956
rect 42352 540790 42472 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 42246 540696 42302 540705
rect 42246 540631 42302 540640
rect 41800 540260 41828 540631
rect 42260 539050 42288 540631
rect 42444 540410 42472 540790
rect 42182 539022 42288 539050
rect 42352 540382 42472 540410
rect 42352 538438 42380 540382
rect 42522 539608 42578 539617
rect 42522 539543 42578 539552
rect 42168 538370 42196 538424
rect 42260 538410 42380 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42536 538234 42564 539543
rect 42352 538206 42564 538234
rect 42168 537798 42288 537826
rect 42168 537744 42196 537798
rect 42260 537758 42288 537798
rect 42352 537758 42380 538206
rect 42614 538112 42670 538121
rect 42812 538098 42840 551103
rect 42996 550634 43024 552327
rect 42904 550606 43024 550634
rect 42904 540974 42932 550606
rect 43074 549536 43130 549545
rect 43074 549471 43130 549480
rect 43088 540974 43116 549471
rect 42904 540946 43024 540974
rect 43088 540946 43208 540974
rect 42996 538218 43024 540946
rect 42984 538212 43036 538218
rect 42984 538154 43036 538160
rect 42812 538070 43024 538098
rect 42614 538047 42670 538056
rect 42260 537730 42380 537758
rect 42430 537432 42486 537441
rect 42430 537367 42486 537376
rect 41786 537024 41842 537033
rect 41786 536959 41842 536968
rect 41800 536588 41828 536959
rect 42246 536480 42302 536489
rect 42246 536415 42302 536424
rect 42076 535673 42104 535908
rect 42062 535664 42118 535673
rect 42062 535599 42118 535608
rect 42260 535514 42288 536415
rect 42168 535486 42288 535514
rect 42168 535364 42196 535486
rect 42444 534766 42472 537367
rect 42628 536874 42656 538047
rect 42800 537940 42852 537946
rect 42800 537882 42852 537888
rect 42812 537758 42840 537882
rect 42168 534698 42196 534752
rect 42260 534738 42472 534766
rect 42536 536846 42656 536874
rect 42720 537730 42840 537758
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42536 534290 42564 536846
rect 42444 534262 42564 534290
rect 42444 534086 42472 534262
rect 42182 534058 42472 534086
rect 42720 533610 42748 537730
rect 42536 533582 42748 533610
rect 42536 533542 42564 533582
rect 42182 533514 42564 533542
rect 42706 532808 42762 532817
rect 42432 532772 42484 532778
rect 42706 532743 42762 532752
rect 42432 532714 42484 532720
rect 42444 531059 42472 532714
rect 42182 531031 42472 531059
rect 42720 530890 42748 532743
rect 42444 530862 42748 530890
rect 42444 530414 42472 530862
rect 42614 530768 42670 530777
rect 42614 530703 42670 530712
rect 42168 530346 42196 530400
rect 42352 530386 42472 530414
rect 42352 530346 42380 530386
rect 42168 530318 42380 530346
rect 42156 530120 42208 530126
rect 42156 530062 42208 530068
rect 42168 529757 42196 530062
rect 42430 529544 42486 529553
rect 42430 529479 42486 529488
rect 41892 529009 41920 529205
rect 41878 529000 41934 529009
rect 41878 528935 41934 528944
rect 42246 529000 42302 529009
rect 42246 528935 42302 528944
rect 42064 527808 42116 527814
rect 42064 527750 42116 527756
rect 42076 527340 42104 527750
rect 42260 526742 42288 528935
rect 42182 526714 42288 526742
rect 42444 526091 42472 529479
rect 42628 527814 42656 530703
rect 42996 530126 43024 538070
rect 43180 532778 43208 540946
rect 43168 532772 43220 532778
rect 43168 532714 43220 532720
rect 42984 530120 43036 530126
rect 42984 530062 43036 530068
rect 42616 527808 42668 527814
rect 42616 527750 42668 527756
rect 42614 527232 42670 527241
rect 42614 527167 42670 527176
rect 42182 526063 42472 526091
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42628 525518 42656 527167
rect 42260 525490 42656 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41696 429208 41748 429214
rect 41696 429150 41748 429156
rect 41708 427122 41736 429150
rect 41970 427136 42026 427145
rect 41708 427094 41970 427122
rect 41970 427071 42026 427080
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 41142 425640 41198 425649
rect 41142 425575 41198 425584
rect 40958 425232 41014 425241
rect 40958 425167 41014 425176
rect 32034 424416 32090 424425
rect 32034 424351 32090 424360
rect 32048 416226 32076 424351
rect 40972 424318 41000 425167
rect 40960 424312 41012 424318
rect 40960 424254 41012 424260
rect 41156 418849 41184 425575
rect 41340 425134 41368 425983
rect 41328 425128 41380 425134
rect 41328 425070 41380 425076
rect 41696 425128 41748 425134
rect 41748 425076 42104 425082
rect 41696 425070 42104 425076
rect 41708 425054 42104 425070
rect 41512 424312 41564 424318
rect 41878 424280 41934 424289
rect 41564 424260 41878 424266
rect 41512 424254 41878 424260
rect 41524 424238 41878 424254
rect 41878 424215 41934 424224
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 42076 418154 42104 425054
rect 42798 423600 42854 423609
rect 42798 423535 42854 423544
rect 42522 419928 42578 419937
rect 42522 419863 42578 419872
rect 42076 418126 42380 418154
rect 32036 416220 32088 416226
rect 32036 416162 32088 416168
rect 41696 416220 41748 416226
rect 41696 416162 41748 416168
rect 41708 416106 41736 416162
rect 41708 416078 42288 416106
rect 42260 413114 42288 416078
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42352 411074 42380 418126
rect 42536 411913 42564 419863
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42380 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 41970 408096 42026 408105
rect 41970 408031 42026 408040
rect 41984 407796 42012 408031
rect 42168 407946 42196 408340
rect 42168 407918 42288 407946
rect 42260 407674 42288 407918
rect 42444 407833 42472 410162
rect 42430 407824 42486 407833
rect 42430 407759 42486 407768
rect 42260 407646 42472 407674
rect 42246 407552 42302 407561
rect 42246 407487 42302 407496
rect 42260 407130 42288 407487
rect 42182 407102 42288 407130
rect 42062 406736 42118 406745
rect 42062 406671 42118 406680
rect 42076 406504 42104 406671
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42444 405657 42472 407646
rect 42246 405648 42302 405657
rect 42246 405583 42302 405592
rect 42430 405648 42486 405657
rect 42430 405583 42486 405592
rect 42260 403458 42288 405583
rect 42182 403430 42288 403458
rect 42812 402974 42840 423535
rect 43258 420744 43314 420753
rect 43258 420679 43314 420688
rect 43074 419520 43130 419529
rect 43074 419455 43130 419464
rect 42536 402946 42840 402974
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42536 402166 42564 402946
rect 42182 402138 42564 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 42444 399135 42472 400143
rect 42182 399107 42472 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 42168 395729 42196 397936
rect 42154 395720 42210 395729
rect 42154 395655 42210 395664
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41142 387152 41198 387161
rect 41142 387087 41198 387096
rect 40774 385928 40830 385937
rect 40774 385863 40830 385872
rect 40788 381449 40816 385863
rect 41156 381857 41184 387087
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41340 385937 41368 386679
rect 41326 385928 41382 385937
rect 41326 385863 41382 385872
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382294 41368 382599
rect 41328 382288 41380 382294
rect 41328 382230 41380 382236
rect 41696 382288 41748 382294
rect 41696 382230 41748 382236
rect 40958 381848 41014 381857
rect 40958 381783 41014 381792
rect 41142 381848 41198 381857
rect 41142 381783 41198 381792
rect 40222 381440 40278 381449
rect 40222 381375 40278 381384
rect 40774 381440 40830 381449
rect 40774 381375 40830 381384
rect 35162 381032 35218 381041
rect 35162 380967 35218 380976
rect 33782 379808 33838 379817
rect 33782 379743 33838 379752
rect 33796 371929 33824 379743
rect 33782 371920 33838 371929
rect 35176 371890 35204 380967
rect 37922 380216 37978 380225
rect 37922 380151 37978 380160
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 374649 35848 376479
rect 35806 374640 35862 374649
rect 35806 374575 35862 374584
rect 37936 372745 37964 380151
rect 40236 378078 40264 381375
rect 40972 380882 41000 381783
rect 40972 380854 41368 380882
rect 41340 379794 41368 380854
rect 41510 379808 41566 379817
rect 41340 379766 41510 379794
rect 41510 379743 41566 379752
rect 41708 379514 41736 382230
rect 42890 379536 42946 379545
rect 41708 379486 42380 379514
rect 40224 378072 40276 378078
rect 40224 378014 40276 378020
rect 41696 378072 41748 378078
rect 41748 378020 42104 378026
rect 41696 378014 42104 378020
rect 41708 378010 42104 378014
rect 41708 378004 42116 378010
rect 41708 377998 42064 378004
rect 42064 377946 42116 377952
rect 37922 372736 37978 372745
rect 37922 372671 37978 372680
rect 33782 371855 33838 371864
rect 35164 371884 35216 371890
rect 35164 371826 35216 371832
rect 41696 371884 41748 371890
rect 41696 371826 41748 371832
rect 41708 371770 41736 371826
rect 41708 371742 42288 371770
rect 42260 369458 42288 371742
rect 42182 369430 42288 369458
rect 41786 368520 41842 368529
rect 41786 368455 41842 368464
rect 41800 368249 41828 368455
rect 42352 367622 42380 379486
rect 42890 379471 42946 379480
rect 42708 378004 42760 378010
rect 42708 377946 42760 377952
rect 42182 367594 42380 367622
rect 42182 366947 42288 366975
rect 42062 366208 42118 366217
rect 42062 366143 42118 366152
rect 42076 365772 42104 366143
rect 42260 365294 42288 366947
rect 42248 365288 42300 365294
rect 42248 365230 42300 365236
rect 42182 365107 42472 365135
rect 42248 364948 42300 364954
rect 42248 364890 42300 364896
rect 42062 364848 42118 364857
rect 42062 364783 42118 364792
rect 42076 364548 42104 364783
rect 42260 364342 42288 364890
rect 42248 364336 42300 364342
rect 42248 364278 42300 364284
rect 42246 364168 42302 364177
rect 42246 364103 42302 364112
rect 42260 363950 42288 364103
rect 42182 363922 42288 363950
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 42444 363066 42472 365107
rect 42720 364334 42748 377946
rect 42904 366217 42932 379471
rect 42890 366208 42946 366217
rect 42890 366143 42946 366152
rect 42260 363038 42472 363066
rect 42536 364306 42748 364334
rect 42260 362953 42288 363038
rect 42246 362944 42302 362953
rect 42246 362879 42302 362888
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 364306
rect 42708 364200 42760 364206
rect 42708 364142 42760 364148
rect 42720 363225 42748 364142
rect 42706 363216 42762 363225
rect 42706 363151 42762 363160
rect 42260 362698 42564 362726
rect 42430 361584 42486 361593
rect 42430 361519 42486 361528
rect 42444 360278 42472 361519
rect 42168 360210 42196 360264
rect 42260 360250 42472 360278
rect 42260 360210 42288 360250
rect 42168 360182 42288 360210
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 41800 359584 41828 360023
rect 41786 359272 41842 359281
rect 41786 359207 41842 359216
rect 41800 358972 41828 359207
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42168 356538 42196 356592
rect 42260 356578 42472 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 41786 356144 41842 356153
rect 41786 356079 41842 356088
rect 41800 355912 41828 356079
rect 42168 355042 42196 355300
rect 42168 355014 42288 355042
rect 42168 353297 42196 354725
rect 42260 353920 42288 355014
rect 42444 354385 42472 356578
rect 42430 354376 42486 354385
rect 42430 354311 42486 354320
rect 43088 353977 43116 419455
rect 43074 353968 43130 353977
rect 42260 353892 42380 353920
rect 43074 353903 43130 353912
rect 42154 353288 42210 353297
rect 42154 353223 42210 353232
rect 42352 353025 42380 353892
rect 43272 353705 43300 420679
rect 43456 354674 43484 582346
rect 43640 354929 43668 590271
rect 44192 581233 44220 591903
rect 44178 581224 44234 581233
rect 44178 581159 44234 581168
rect 44376 578105 44404 593127
rect 44638 580680 44694 580689
rect 44638 580615 44694 580624
rect 44362 578096 44418 578105
rect 44362 578031 44418 578040
rect 44652 575482 44680 580615
rect 44640 575476 44692 575482
rect 44640 575418 44692 575424
rect 44546 556880 44602 556889
rect 44546 556815 44602 556824
rect 44270 556064 44326 556073
rect 44270 555999 44326 556008
rect 43810 548312 43866 548321
rect 43810 548247 43866 548256
rect 43824 355201 43852 548247
rect 43994 547088 44050 547097
rect 43994 547023 44050 547032
rect 43810 355192 43866 355201
rect 43810 355127 43866 355136
rect 43626 354920 43682 354929
rect 43626 354855 43682 354864
rect 43456 354646 43760 354674
rect 43732 354634 43760 354646
rect 44008 354634 44036 547023
rect 44284 428913 44312 555999
rect 44560 429729 44588 556815
rect 44928 555665 44956 598431
rect 45112 558793 45140 600063
rect 45296 598097 45324 640183
rect 45572 612105 45600 763263
rect 46216 743782 46244 773055
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 60016 742422 60044 774182
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 61396 747046 61424 772822
rect 62764 755540 62816 755546
rect 62764 755482 62816 755488
rect 62776 747697 62804 755482
rect 62762 747688 62818 747697
rect 62762 747623 62818 747632
rect 61384 747040 61436 747046
rect 61384 746982 61436 746988
rect 62396 747040 62448 747046
rect 62396 746982 62448 746988
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 60004 742416 60056 742422
rect 62120 742416 62172 742422
rect 60004 742358 60056 742364
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 62408 741849 62436 746982
rect 62394 741840 62450 741849
rect 62394 741775 62450 741784
rect 652036 736234 652064 776999
rect 653416 775334 653444 790774
rect 669228 782536 669280 782542
rect 669228 782478 669280 782484
rect 655520 781244 655572 781250
rect 655520 781186 655572 781192
rect 655060 778388 655112 778394
rect 655060 778330 655112 778336
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655072 773838 655100 778330
rect 655532 774178 655560 781186
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655060 773832 655112 773838
rect 655060 773774 655112 773780
rect 652024 736228 652076 736234
rect 652024 736170 652076 736176
rect 653404 736228 653456 736234
rect 653404 736170 653456 736176
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 651470 733000 651526 733009
rect 651470 732935 651526 732944
rect 651484 732834 651512 732935
rect 651472 732828 651524 732834
rect 651472 732770 651524 732776
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651472 731332 651524 731338
rect 651472 731274 651524 731280
rect 651484 731105 651512 731274
rect 651470 731096 651526 731105
rect 651470 731031 651526 731040
rect 46202 730960 46258 730969
rect 46202 730895 46258 730904
rect 46216 698222 46244 730895
rect 61384 730380 61436 730386
rect 61384 730322 61436 730328
rect 47214 721168 47270 721177
rect 47214 721103 47270 721112
rect 47030 719944 47086 719953
rect 47030 719879 47086 719888
rect 46204 698216 46256 698222
rect 46204 698158 46256 698164
rect 45744 667956 45796 667962
rect 45744 667898 45796 667904
rect 45756 665854 45784 667898
rect 45744 665848 45796 665854
rect 45744 665790 45796 665796
rect 45744 625864 45796 625870
rect 45744 625806 45796 625812
rect 45756 624481 45784 625806
rect 45742 624472 45798 624481
rect 45742 624407 45798 624416
rect 45558 612096 45614 612105
rect 45558 612031 45614 612040
rect 47044 611833 47072 719879
rect 47030 611824 47086 611833
rect 47030 611759 47086 611768
rect 47228 611561 47256 721103
rect 50344 712156 50396 712162
rect 50344 712098 50396 712104
rect 50356 705158 50384 712098
rect 50344 705152 50396 705158
rect 50344 705094 50396 705100
rect 61396 699689 61424 730322
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 62764 729360 62816 729366
rect 62764 729302 62816 729308
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 62210 701312 62266 701321
rect 62210 701247 62266 701256
rect 62224 701078 62252 701247
rect 62212 701072 62264 701078
rect 62212 701014 62264 701020
rect 62776 700913 62804 729302
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 651524 728512 651526 728521
rect 651470 728447 651526 728456
rect 653416 716310 653444 736170
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 654796 728550 654824 734130
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 654784 728544 654836 728550
rect 654784 728486 654836 728492
rect 653404 716304 653456 716310
rect 653404 716246 653456 716252
rect 654784 701072 654836 701078
rect 654784 701014 654836 701020
rect 62762 700904 62818 700913
rect 62762 700839 62818 700848
rect 61382 699680 61438 699689
rect 61382 699615 61438 699624
rect 62120 698216 62172 698222
rect 62118 698184 62120 698193
rect 62172 698184 62174 698193
rect 62118 698119 62174 698128
rect 651470 689480 651526 689489
rect 651470 689415 651526 689424
rect 651484 688702 651512 689415
rect 652760 688832 652812 688838
rect 651654 688800 651710 688809
rect 652760 688774 652812 688780
rect 651654 688735 651710 688744
rect 651472 688696 651524 688702
rect 651472 688638 651524 688644
rect 651470 687440 651526 687449
rect 651470 687375 651526 687384
rect 651484 687274 651512 687375
rect 61384 687268 61436 687274
rect 61384 687210 61436 687216
rect 651472 687268 651524 687274
rect 651472 687210 651524 687216
rect 53104 669384 53156 669390
rect 53104 669326 53156 669332
rect 53116 660958 53144 669326
rect 57244 667956 57296 667962
rect 57244 667898 57296 667904
rect 53104 660952 53156 660958
rect 53104 660894 53156 660900
rect 57256 659598 57284 667898
rect 57244 659592 57296 659598
rect 57244 659534 57296 659540
rect 61396 656577 61424 687210
rect 651472 687064 651524 687070
rect 651472 687006 651524 687012
rect 651484 686769 651512 687006
rect 651470 686760 651526 686769
rect 651470 686695 651526 686704
rect 651668 686526 651696 688735
rect 62764 686520 62816 686526
rect 62764 686462 62816 686468
rect 651656 686520 651708 686526
rect 651656 686462 651708 686468
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 62120 659592 62172 659598
rect 62118 659560 62120 659569
rect 62172 659560 62174 659569
rect 62118 659495 62174 659504
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62776 657665 62804 686462
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687070 654824 701014
rect 656440 690124 656492 690130
rect 656440 690066 656492 690072
rect 654784 687064 654836 687070
rect 654784 687006 654836 687012
rect 656452 685574 656480 690066
rect 657544 688696 657596 688702
rect 657544 688638 657596 688644
rect 656440 685568 656492 685574
rect 656440 685510 656492 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 62762 657656 62818 657665
rect 62762 657591 62818 657600
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 61382 656568 61438 656577
rect 61382 656503 61438 656512
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 62120 655512 62172 655518
rect 62120 655454 62172 655460
rect 62132 655353 62160 655454
rect 62118 655344 62174 655353
rect 62118 655279 62174 655288
rect 60004 644496 60056 644502
rect 60004 644438 60056 644444
rect 60016 612678 60044 644438
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 61384 643136 61436 643142
rect 61384 643078 61436 643084
rect 61396 613873 61424 643078
rect 651484 642394 651512 643175
rect 62764 642388 62816 642394
rect 62764 642330 62816 642336
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 61382 613864 61438 613873
rect 61382 613799 61438 613808
rect 60004 612672 60056 612678
rect 62120 612672 62172 612678
rect 60004 612614 60056 612620
rect 62118 612640 62120 612649
rect 62172 612640 62174 612649
rect 62118 612575 62174 612584
rect 62776 612105 62804 642330
rect 652022 641880 652078 641889
rect 652022 641815 652078 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 62948 625864 63000 625870
rect 62948 625806 63000 625812
rect 62960 618089 62988 625806
rect 62946 618080 63002 618089
rect 62946 618015 63002 618024
rect 62762 612096 62818 612105
rect 62762 612031 62818 612040
rect 47214 611552 47270 611561
rect 47214 611487 47270 611496
rect 45282 598088 45338 598097
rect 45282 598023 45338 598032
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 62946 595776 63002 595785
rect 62946 595711 63002 595720
rect 62762 594144 62818 594153
rect 62762 594079 62818 594088
rect 45558 578912 45614 578921
rect 45558 578847 45614 578856
rect 45572 574054 45600 578847
rect 62120 575476 62172 575482
rect 62120 575418 62172 575424
rect 62132 574841 62160 575418
rect 62118 574832 62174 574841
rect 62118 574767 62174 574776
rect 45560 574048 45612 574054
rect 45560 573990 45612 573996
rect 62120 574048 62172 574054
rect 62120 573990 62172 573996
rect 62132 573617 62160 573990
rect 62118 573608 62174 573617
rect 62118 573543 62174 573552
rect 62776 568585 62804 594079
rect 62960 571169 62988 595711
rect 651470 595504 651526 595513
rect 651470 595439 651526 595448
rect 651656 595468 651708 595474
rect 651484 594930 651512 595439
rect 651656 595410 651708 595416
rect 651668 595241 651696 595410
rect 651654 595232 651710 595241
rect 651654 595167 651710 595176
rect 651472 594924 651524 594930
rect 651472 594866 651524 594872
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 651472 593088 651524 593094
rect 651472 593030 651524 593036
rect 63130 592920 63186 592929
rect 63130 592855 63186 592864
rect 62946 571160 63002 571169
rect 62946 571095 63002 571104
rect 63144 569945 63172 592855
rect 651484 592793 651512 593030
rect 651470 592784 651526 592793
rect 651470 592719 651526 592728
rect 652036 581058 652064 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 657556 625190 657584 688638
rect 658936 669526 658964 731410
rect 660316 714882 660344 777582
rect 668400 736976 668452 736982
rect 668400 736918 668452 736924
rect 667480 735616 667532 735622
rect 667480 735558 667532 735564
rect 667492 734874 667520 735558
rect 667480 734868 667532 734874
rect 667480 734810 667532 734816
rect 661684 732828 661736 732834
rect 661684 732770 661736 732776
rect 660304 714876 660356 714882
rect 660304 714818 660356 714824
rect 661696 670750 661724 732770
rect 667848 729972 667900 729978
rect 667848 729914 667900 729920
rect 666468 701276 666520 701282
rect 666468 701218 666520 701224
rect 666284 696992 666336 696998
rect 666284 696934 666336 696940
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 658924 669520 658976 669526
rect 658924 669462 658976 669468
rect 658924 642388 658976 642394
rect 658924 642330 658976 642336
rect 657544 625184 657596 625190
rect 657544 625126 657596 625132
rect 653404 611380 653456 611386
rect 653404 611322 653456 611328
rect 653416 595474 653444 611322
rect 657544 600364 657596 600370
rect 657544 600306 657596 600312
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 653404 595468 653456 595474
rect 653404 595410 653456 595416
rect 654796 593094 654824 598946
rect 656164 594924 656216 594930
rect 656164 594866 656216 594872
rect 654784 593088 654836 593094
rect 654784 593030 654836 593036
rect 652024 581052 652076 581058
rect 652024 580994 652076 581000
rect 63130 569936 63186 569945
rect 63130 569871 63186 569880
rect 62762 568576 62818 568585
rect 62762 568511 62818 568520
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 45098 558784 45154 558793
rect 45098 558719 45154 558728
rect 61382 557560 61438 557569
rect 61382 557495 61438 557504
rect 44914 555656 44970 555665
rect 44914 555591 44970 555600
rect 45650 555248 45706 555257
rect 45650 555183 45706 555192
rect 45190 551576 45246 551585
rect 45190 551511 45246 551520
rect 45006 549128 45062 549137
rect 45006 549063 45062 549072
rect 44730 548720 44786 548729
rect 44730 548655 44786 548664
rect 44744 536897 44772 548655
rect 45020 538121 45048 549063
rect 45006 538112 45062 538121
rect 45006 538047 45062 538056
rect 44730 536888 44786 536897
rect 44730 536823 44786 536832
rect 44730 535664 44786 535673
rect 44730 535599 44786 535608
rect 44744 531282 44772 535599
rect 44732 531276 44784 531282
rect 44732 531218 44784 531224
rect 45204 529009 45232 551511
rect 45374 550760 45430 550769
rect 45374 550695 45430 550704
rect 45388 532817 45416 550695
rect 45374 532808 45430 532817
rect 45374 532743 45430 532752
rect 45190 529000 45246 529009
rect 45190 528935 45246 528944
rect 45100 528624 45152 528630
rect 45100 528566 45152 528572
rect 45112 527241 45140 528566
rect 45098 527232 45154 527241
rect 45098 527167 45154 527176
rect 44546 429720 44602 429729
rect 44546 429655 44602 429664
rect 44638 429312 44694 429321
rect 44638 429247 44694 429256
rect 44270 428904 44326 428913
rect 44270 428839 44326 428848
rect 44270 428496 44326 428505
rect 44270 428431 44326 428440
rect 44284 385665 44312 428431
rect 44454 422376 44510 422385
rect 44454 422311 44510 422320
rect 44468 407561 44496 422311
rect 44454 407552 44510 407561
rect 44454 407487 44510 407496
rect 44652 386481 44680 429247
rect 45664 428097 45692 555183
rect 45834 554432 45890 554441
rect 45834 554367 45890 554376
rect 45650 428088 45706 428097
rect 45650 428023 45706 428032
rect 45650 427680 45706 427689
rect 45650 427615 45706 427624
rect 45664 427258 45692 427615
rect 45848 427417 45876 554367
rect 60002 539608 60058 539617
rect 60002 539543 60058 539552
rect 60016 531146 60044 539543
rect 60004 531140 60056 531146
rect 60004 531082 60056 531088
rect 61396 527105 61424 557495
rect 63406 556744 63462 556753
rect 63406 556679 63462 556688
rect 62946 552664 63002 552673
rect 62946 552599 63002 552608
rect 62120 531276 62172 531282
rect 62120 531218 62172 531224
rect 62132 530641 62160 531218
rect 62302 531176 62358 531185
rect 62302 531111 62304 531120
rect 62356 531111 62358 531120
rect 62304 531082 62356 531088
rect 62118 530632 62174 530641
rect 62118 530567 62174 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 61382 527096 61438 527105
rect 61382 527031 61438 527040
rect 62960 525745 62988 552599
rect 63420 528057 63448 556679
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 651470 552392 651526 552401
rect 651470 552327 651526 552336
rect 651484 552090 651512 552327
rect 651472 552084 651524 552090
rect 651472 552026 651524 552032
rect 651470 551168 651526 551177
rect 651470 551103 651526 551112
rect 651484 550662 651512 551103
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 653416 550390 653444 565830
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 651380 550384 651432 550390
rect 651378 550352 651380 550361
rect 653404 550384 653456 550390
rect 651432 550352 651434 550361
rect 653404 550326 653456 550332
rect 651378 550287 651434 550296
rect 651470 549128 651526 549137
rect 651470 549063 651472 549072
rect 651524 549063 651526 549072
rect 651472 549034 651524 549040
rect 655164 548894 655192 553386
rect 651472 548888 651524 548894
rect 651472 548830 651524 548836
rect 655152 548888 655204 548894
rect 655152 548830 655204 548836
rect 651484 548457 651512 548830
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 656176 534274 656204 594866
rect 657556 594726 657584 600306
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 658936 579698 658964 642330
rect 666296 619682 666324 696934
rect 666480 621110 666508 701218
rect 667204 686520 667256 686526
rect 667204 686462 667256 686468
rect 667216 625734 667244 686462
rect 667388 661156 667440 661162
rect 667388 661098 667440 661104
rect 667204 625728 667256 625734
rect 667204 625670 667256 625676
rect 666468 621104 666520 621110
rect 666468 621046 666520 621052
rect 666284 619676 666336 619682
rect 666284 619618 666336 619624
rect 667204 597576 667256 597582
rect 667204 597518 667256 597524
rect 660304 596216 660356 596222
rect 660304 596158 660356 596164
rect 658924 579692 658976 579698
rect 658924 579634 658976 579640
rect 657820 554804 657872 554810
rect 657820 554746 657872 554752
rect 657832 549098 657860 554746
rect 658924 552084 658976 552090
rect 658924 552026 658976 552032
rect 657820 549092 657872 549098
rect 657820 549034 657872 549040
rect 656164 534268 656216 534274
rect 656164 534210 656216 534216
rect 63406 528048 63462 528057
rect 63406 527983 63462 527992
rect 62946 525736 63002 525745
rect 62946 525671 63002 525680
rect 658936 491366 658964 552026
rect 660316 535498 660344 596158
rect 667018 595504 667074 595513
rect 667018 595439 667074 595448
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 660304 535492 660356 535498
rect 660304 535434 660356 535440
rect 665836 491502 665864 552638
rect 667032 530534 667060 595439
rect 667216 535702 667244 597518
rect 667204 535696 667256 535702
rect 667204 535638 667256 535644
rect 667020 530528 667072 530534
rect 667020 530470 667072 530476
rect 665824 491496 665876 491502
rect 665824 491438 665876 491444
rect 658924 491360 658976 491366
rect 658924 491302 658976 491308
rect 667400 455666 667428 661098
rect 667860 660210 667888 729914
rect 668030 689888 668086 689897
rect 668030 689823 668086 689832
rect 667848 660204 667900 660210
rect 667848 660146 667900 660152
rect 667754 649224 667810 649233
rect 667754 649159 667810 649168
rect 667572 647284 667624 647290
rect 667572 647226 667624 647232
rect 667584 574122 667612 647226
rect 667572 574116 667624 574122
rect 667572 574058 667624 574064
rect 667768 572762 667796 649159
rect 668044 616962 668072 689823
rect 668214 686488 668270 686497
rect 668214 686423 668270 686432
rect 668228 621790 668256 686423
rect 668412 661978 668440 736918
rect 668950 736128 669006 736137
rect 668950 736063 669006 736072
rect 668584 733440 668636 733446
rect 668584 733382 668636 733388
rect 668596 671158 668624 733382
rect 668768 685908 668820 685914
rect 668768 685850 668820 685856
rect 668584 671152 668636 671158
rect 668584 671094 668636 671100
rect 668400 661972 668452 661978
rect 668400 661914 668452 661920
rect 668398 640656 668454 640665
rect 668398 640591 668454 640600
rect 668216 621784 668268 621790
rect 668216 621726 668268 621732
rect 668032 616956 668084 616962
rect 668032 616898 668084 616904
rect 668412 575550 668440 640591
rect 668584 640348 668636 640354
rect 668584 640290 668636 640296
rect 668596 580310 668624 640290
rect 668780 620294 668808 685850
rect 668964 665242 668992 736063
rect 669240 709374 669268 782478
rect 669964 775600 670016 775606
rect 669964 775542 670016 775548
rect 669780 774308 669832 774314
rect 669780 774250 669832 774256
rect 669228 709368 669280 709374
rect 669228 709310 669280 709316
rect 669792 705430 669820 774250
rect 669976 715766 670004 775542
rect 670792 745272 670844 745278
rect 670792 745214 670844 745220
rect 670148 739152 670200 739158
rect 670148 739094 670200 739100
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 669780 705424 669832 705430
rect 669780 705366 669832 705372
rect 669228 703860 669280 703866
rect 669228 703802 669280 703808
rect 668952 665236 669004 665242
rect 668952 665178 669004 665184
rect 669240 627914 669268 703802
rect 669964 687268 670016 687274
rect 669964 687210 670016 687216
rect 669778 685808 669834 685817
rect 669778 685743 669834 685752
rect 669596 669384 669648 669390
rect 669596 669326 669648 669332
rect 669412 666596 669464 666602
rect 669412 666538 669464 666544
rect 669424 633146 669452 666538
rect 669608 635662 669636 669326
rect 669792 649994 669820 685743
rect 669976 654134 670004 687210
rect 670160 664018 670188 739094
rect 670514 733816 670570 733825
rect 670514 733751 670570 733760
rect 670332 728680 670384 728686
rect 670332 728622 670384 728628
rect 670344 717614 670372 728622
rect 670252 717586 670372 717614
rect 670252 673454 670280 717586
rect 670252 673426 670372 673454
rect 670344 664494 670372 673426
rect 670332 664488 670384 664494
rect 670332 664430 670384 664436
rect 670148 664012 670200 664018
rect 670148 663954 670200 663960
rect 670528 661638 670556 733751
rect 670804 727274 670832 745214
rect 671252 743844 671304 743850
rect 671252 743786 671304 743792
rect 670974 734224 671030 734233
rect 670974 734159 670976 734168
rect 671028 734159 671030 734168
rect 670976 734130 671028 734136
rect 671264 731338 671292 743786
rect 671252 731332 671304 731338
rect 671252 731274 671304 731280
rect 670804 727246 670924 727274
rect 670698 689208 670754 689217
rect 670698 689143 670754 689152
rect 670516 661632 670568 661638
rect 670516 661574 670568 661580
rect 669976 654106 670096 654134
rect 669700 649966 669820 649994
rect 669700 635712 669728 649966
rect 669870 641744 669926 641753
rect 669870 641679 669926 641688
rect 669884 640334 669912 641679
rect 669792 640306 669912 640334
rect 669792 636154 669820 640306
rect 669792 636126 670004 636154
rect 669700 635684 669912 635712
rect 669596 635656 669648 635662
rect 669596 635598 669648 635604
rect 669884 635338 669912 635684
rect 669700 635310 669912 635338
rect 669412 633140 669464 633146
rect 669412 633082 669464 633088
rect 669504 631372 669556 631378
rect 669504 631314 669556 631320
rect 669148 627886 669268 627914
rect 669148 623098 669176 627886
rect 669148 623070 669268 623098
rect 668768 620288 668820 620294
rect 668768 620230 668820 620236
rect 669042 608288 669098 608297
rect 669042 608223 669098 608232
rect 668858 593600 668914 593609
rect 668858 593535 668914 593544
rect 668584 580304 668636 580310
rect 668584 580246 668636 580252
rect 668400 575544 668452 575550
rect 668400 575486 668452 575492
rect 667756 572756 667808 572762
rect 667756 572698 667808 572704
rect 667754 561912 667810 561921
rect 667754 561847 667810 561856
rect 667768 484430 667796 561847
rect 668674 555248 668730 555257
rect 668674 555183 668730 555192
rect 668688 485858 668716 555183
rect 668872 528630 668900 593535
rect 669056 530058 669084 608223
rect 669044 530052 669096 530058
rect 669044 529994 669096 530000
rect 668860 528624 668912 528630
rect 668860 528566 668912 528572
rect 668676 485852 668728 485858
rect 668676 485794 668728 485800
rect 667756 484424 667808 484430
rect 667756 484366 667808 484372
rect 669240 456618 669268 623070
rect 669516 622946 669544 631314
rect 669700 627586 669728 635310
rect 669976 631394 670004 636126
rect 669884 631378 670004 631394
rect 669872 631372 670004 631378
rect 669924 631366 670004 631372
rect 669872 631314 669924 631320
rect 669700 627558 669912 627586
rect 669884 626534 669912 627558
rect 669792 626506 669912 626534
rect 669792 626362 669820 626506
rect 669700 626334 669820 626362
rect 669504 622940 669556 622946
rect 669504 622882 669556 622888
rect 669504 622804 669556 622810
rect 669504 622746 669556 622752
rect 669516 618254 669544 622746
rect 669700 618254 669728 626334
rect 670068 626006 670096 654106
rect 670514 647864 670570 647873
rect 670514 647799 670570 647808
rect 670240 635656 670292 635662
rect 670240 635598 670292 635604
rect 670056 626000 670108 626006
rect 670056 625942 670108 625948
rect 670252 625161 670280 635598
rect 670238 625152 670294 625161
rect 670238 625087 670294 625096
rect 670148 624708 670200 624714
rect 670148 624650 670200 624656
rect 669964 623076 670016 623082
rect 669964 623018 670016 623024
rect 669516 618226 669636 618254
rect 669700 618226 669820 618254
rect 669608 601694 669636 618226
rect 669792 615534 669820 618226
rect 669780 615528 669832 615534
rect 669780 615470 669832 615476
rect 669516 601666 669636 601694
rect 669516 573102 669544 601666
rect 669780 579284 669832 579290
rect 669780 579226 669832 579232
rect 669504 573096 669556 573102
rect 669504 573038 669556 573044
rect 669596 550656 669648 550662
rect 669596 550598 669648 550604
rect 669608 491910 669636 550598
rect 669792 535022 669820 579226
rect 669976 578134 670004 623018
rect 670160 580446 670188 624650
rect 670332 622260 670384 622266
rect 670332 622202 670384 622208
rect 670148 580440 670200 580446
rect 670148 580382 670200 580388
rect 669964 578128 670016 578134
rect 669964 578070 670016 578076
rect 670344 577862 670372 622202
rect 670332 577856 670384 577862
rect 670332 577798 670384 577804
rect 670240 577516 670292 577522
rect 670240 577458 670292 577464
rect 670056 568608 670108 568614
rect 670056 568550 670108 568556
rect 669780 535016 669832 535022
rect 669780 534958 669832 534964
rect 669596 491904 669648 491910
rect 669596 491846 669648 491852
rect 669228 456612 669280 456618
rect 669228 456554 669280 456560
rect 667388 455660 667440 455666
rect 667388 455602 667440 455608
rect 670068 455433 670096 568550
rect 670252 532982 670280 577458
rect 670528 572714 670556 647799
rect 670712 616622 670740 689143
rect 670896 683114 670924 727246
rect 671448 715358 671476 894270
rect 671804 886916 671856 886922
rect 671804 886858 671856 886864
rect 671620 789404 671672 789410
rect 671620 789346 671672 789352
rect 671436 715352 671488 715358
rect 671436 715294 671488 715300
rect 671068 715012 671120 715018
rect 671068 714954 671120 714960
rect 671080 712586 671108 714954
rect 671344 713244 671396 713250
rect 671344 713186 671396 713192
rect 670804 683086 670924 683114
rect 670988 712558 671108 712586
rect 670804 670018 670832 683086
rect 670988 670138 671016 712558
rect 671160 712428 671212 712434
rect 671160 712370 671212 712376
rect 670976 670132 671028 670138
rect 670976 670074 671028 670080
rect 670804 669990 670924 670018
rect 670896 666058 670924 669990
rect 671172 666942 671200 712370
rect 671356 668574 671384 713186
rect 671632 709646 671660 789346
rect 671816 728142 671844 886858
rect 671804 728136 671856 728142
rect 671804 728078 671856 728084
rect 672000 714542 672028 894406
rect 672356 893036 672408 893042
rect 672356 892978 672408 892984
rect 672172 775600 672224 775606
rect 672172 775542 672224 775548
rect 671988 714536 672040 714542
rect 671988 714478 672040 714484
rect 672184 710054 672212 775542
rect 672368 713726 672396 892978
rect 672736 866658 672764 895630
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894334 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 676048 894470 676076 894639
rect 676036 894464 676088 894470
rect 676036 894406 676088 894412
rect 675852 894328 675904 894334
rect 675852 894270 675904 894276
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 675864 893042 675892 893823
rect 676034 893072 676090 893081
rect 675852 893036 675904 893042
rect 676034 893007 676090 893016
rect 675852 892978 675904 892984
rect 676048 892906 676076 893007
rect 673368 892900 673420 892906
rect 673368 892842 673420 892848
rect 676036 892900 676088 892906
rect 676036 892842 676088 892848
rect 673184 885692 673236 885698
rect 673184 885634 673236 885640
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 673000 783896 673052 783902
rect 673000 783838 673052 783844
rect 672540 730516 672592 730522
rect 672540 730458 672592 730464
rect 672356 713720 672408 713726
rect 672356 713662 672408 713668
rect 672172 710048 672224 710054
rect 672172 709990 672224 709996
rect 671620 709640 671672 709646
rect 671620 709582 671672 709588
rect 672354 695464 672410 695473
rect 672354 695399 672410 695408
rect 671802 690432 671858 690441
rect 671802 690367 671858 690376
rect 671344 668568 671396 668574
rect 671344 668510 671396 668516
rect 671528 668228 671580 668234
rect 671528 668170 671580 668176
rect 671344 667956 671396 667962
rect 671344 667898 671396 667904
rect 671160 666936 671212 666942
rect 671160 666878 671212 666884
rect 670884 666052 670936 666058
rect 670884 665994 670936 666000
rect 670976 645924 671028 645930
rect 670976 645866 671028 645872
rect 670988 643521 671016 645866
rect 670974 643512 671030 643521
rect 670974 643447 671030 643456
rect 670974 638752 671030 638761
rect 670974 638687 671030 638696
rect 670700 616616 670752 616622
rect 670700 616558 670752 616564
rect 670700 614916 670752 614922
rect 670700 614858 670752 614864
rect 670712 614802 670740 614858
rect 670436 572686 670556 572714
rect 670620 614774 670740 614802
rect 670436 571470 670464 572686
rect 670424 571464 670476 571470
rect 670424 571406 670476 571412
rect 670422 552120 670478 552129
rect 670422 552055 670478 552064
rect 670240 532976 670292 532982
rect 670240 532918 670292 532924
rect 670436 484022 670464 552055
rect 670424 484016 670476 484022
rect 670424 483958 670476 483964
rect 670620 455530 670648 614774
rect 670988 574598 671016 638687
rect 671160 633140 671212 633146
rect 671160 633082 671212 633088
rect 671172 622713 671200 633082
rect 671356 623558 671384 667898
rect 671540 624374 671568 668170
rect 671528 624368 671580 624374
rect 671528 624310 671580 624316
rect 671620 623892 671672 623898
rect 671620 623834 671672 623840
rect 671344 623552 671396 623558
rect 671344 623494 671396 623500
rect 671158 622704 671214 622713
rect 671158 622639 671214 622648
rect 671342 607336 671398 607345
rect 671342 607271 671398 607280
rect 671160 576972 671212 576978
rect 671160 576914 671212 576920
rect 670976 574592 671028 574598
rect 670976 574534 671028 574540
rect 670974 548448 671030 548457
rect 670974 548383 671030 548392
rect 670792 534132 670844 534138
rect 670792 534074 670844 534080
rect 670804 490958 670832 534074
rect 670792 490952 670844 490958
rect 670792 490894 670844 490900
rect 670988 485654 671016 548383
rect 671172 531758 671200 576914
rect 671160 531752 671212 531758
rect 671160 531694 671212 531700
rect 671160 531344 671212 531350
rect 671160 531286 671212 531292
rect 671172 488510 671200 531286
rect 671356 528766 671384 607271
rect 671632 579086 671660 623834
rect 671816 620265 671844 690367
rect 672172 685908 672224 685914
rect 672172 685850 672224 685856
rect 672184 685409 672212 685850
rect 672170 685400 672226 685409
rect 672170 685335 672226 685344
rect 672172 659728 672224 659734
rect 672172 659670 672224 659676
rect 671986 652216 672042 652225
rect 671986 652151 672042 652160
rect 671802 620256 671858 620265
rect 671802 620191 671858 620200
rect 671802 600672 671858 600681
rect 671802 600607 671858 600616
rect 671620 579080 671672 579086
rect 671620 579022 671672 579028
rect 671528 578332 671580 578338
rect 671528 578274 671580 578280
rect 671540 534177 671568 578274
rect 671526 534168 671582 534177
rect 671526 534103 671582 534112
rect 671620 532772 671672 532778
rect 671620 532714 671672 532720
rect 671344 528760 671396 528766
rect 671344 528702 671396 528708
rect 671632 489326 671660 532714
rect 671816 530262 671844 600607
rect 672000 574326 672028 652151
rect 671988 574320 672040 574326
rect 671988 574262 672040 574268
rect 671988 569968 672040 569974
rect 671988 569910 672040 569916
rect 671804 530256 671856 530262
rect 671804 530198 671856 530204
rect 671620 489320 671672 489326
rect 671620 489262 671672 489268
rect 671160 488504 671212 488510
rect 671160 488446 671212 488452
rect 670976 485648 671028 485654
rect 670976 485590 671028 485596
rect 670608 455524 670660 455530
rect 670608 455466 670660 455472
rect 670054 455424 670110 455433
rect 670054 455359 670110 455368
rect 672000 455138 672028 569910
rect 672184 455870 672212 659670
rect 672368 619070 672396 695399
rect 672552 665446 672580 730458
rect 672816 727864 672868 727870
rect 672816 727806 672868 727812
rect 672828 723178 672856 727806
rect 672816 723172 672868 723178
rect 672816 723114 672868 723120
rect 673012 717614 673040 783838
rect 673196 728346 673224 885634
rect 673184 728340 673236 728346
rect 673184 728282 673236 728288
rect 673380 727954 673408 892842
rect 676034 892664 676090 892673
rect 676090 892622 676260 892650
rect 676034 892599 676090 892608
rect 676232 891546 676260 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676220 891540 676272 891546
rect 676220 891482 676272 891488
rect 676864 891540 676916 891546
rect 676864 891482 676916 891488
rect 675850 891440 675906 891449
rect 675850 891375 675906 891384
rect 675666 891032 675722 891041
rect 675666 890967 675722 890976
rect 674380 888956 674432 888962
rect 674380 888898 674432 888904
rect 674196 888140 674248 888146
rect 674196 888082 674248 888088
rect 674208 873662 674236 888082
rect 674196 873656 674248 873662
rect 674196 873598 674248 873604
rect 674392 869650 674420 888898
rect 675680 888758 675708 890967
rect 674840 888752 674892 888758
rect 674840 888694 674892 888700
rect 675668 888752 675720 888758
rect 675668 888694 675720 888700
rect 674656 888548 674708 888554
rect 674656 888490 674708 888496
rect 674668 869854 674696 888490
rect 674852 879322 674880 888694
rect 675482 886952 675538 886961
rect 675482 886887 675484 886896
rect 675536 886887 675538 886896
rect 675484 886858 675536 886864
rect 675864 881834 675892 891375
rect 676034 890624 676090 890633
rect 676090 890582 676260 890610
rect 676034 890559 676090 890568
rect 676034 890216 676090 890225
rect 676034 890151 676090 890160
rect 676048 890050 676076 890151
rect 676036 890044 676088 890050
rect 676036 889986 676088 889992
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 676034 888584 676090 888593
rect 676034 888519 676036 888528
rect 676088 888519 676090 888528
rect 676036 888490 676088 888496
rect 676034 888176 676090 888185
rect 676034 888111 676036 888120
rect 676088 888111 676090 888120
rect 676036 888082 676088 888088
rect 676034 887496 676090 887505
rect 676232 887482 676260 890582
rect 676090 887454 676260 887482
rect 676034 887431 676090 887440
rect 676678 887360 676734 887369
rect 676678 887295 676734 887304
rect 676034 885728 676090 885737
rect 676034 885663 676036 885672
rect 676088 885663 676090 885672
rect 676036 885634 676088 885640
rect 676692 882609 676720 887295
rect 676678 882600 676734 882609
rect 676678 882535 676734 882544
rect 674760 879294 674880 879322
rect 675036 881806 675892 881834
rect 675036 879322 675064 881806
rect 675208 881136 675260 881142
rect 675208 881078 675260 881084
rect 675036 879294 675156 879322
rect 674760 879050 674788 879294
rect 674932 879164 674984 879170
rect 674932 879106 674984 879112
rect 674760 879022 674880 879050
rect 674852 872438 674880 879022
rect 674944 874290 674972 879106
rect 675128 879016 675156 879294
rect 675036 878988 675156 879016
rect 675036 874426 675064 878988
rect 675220 876466 675248 881078
rect 675576 880524 675628 880530
rect 675576 880466 675628 880472
rect 675588 879186 675616 880466
rect 675944 880184 675996 880190
rect 675944 880126 675996 880132
rect 675760 879368 675812 879374
rect 675760 879310 675812 879316
rect 675588 879158 675708 879186
rect 675392 879028 675444 879034
rect 675392 878970 675444 878976
rect 675404 878234 675432 878970
rect 675680 878642 675708 879158
rect 675312 878206 675432 878234
rect 675588 878614 675708 878642
rect 675312 876738 675340 878206
rect 675588 878084 675616 878614
rect 675772 878422 675800 879310
rect 675956 878529 675984 880126
rect 676876 879034 676904 891482
rect 677048 890044 677100 890050
rect 677048 889986 677100 889992
rect 677060 879374 677088 889986
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 879368 677100 879374
rect 677048 879310 677100 879316
rect 678256 879170 678284 889743
rect 679636 880190 679664 891783
rect 683302 889400 683358 889409
rect 683302 889335 683358 889344
rect 683026 886136 683082 886145
rect 683026 886071 683082 886080
rect 683040 881929 683068 886071
rect 683026 881920 683082 881929
rect 683026 881855 683082 881864
rect 683316 881142 683344 889335
rect 683304 881136 683356 881142
rect 683304 881078 683356 881084
rect 679624 880184 679676 880190
rect 679624 880126 679676 880132
rect 678244 879164 678296 879170
rect 678244 879106 678296 879112
rect 676864 879028 676916 879034
rect 676864 878970 676916 878976
rect 675942 878520 675998 878529
rect 675942 878455 675998 878464
rect 675760 878416 675812 878422
rect 675760 878358 675812 878364
rect 675666 877840 675722 877849
rect 675666 877775 675722 877784
rect 675680 877540 675708 877775
rect 675484 877260 675536 877266
rect 675484 877202 675536 877208
rect 675496 876860 675524 877202
rect 675312 876710 675708 876738
rect 675482 876480 675538 876489
rect 675220 876438 675482 876466
rect 675482 876415 675538 876424
rect 675680 876248 675708 876710
rect 675036 874398 675340 874426
rect 675312 874290 675340 874398
rect 675404 874290 675432 874412
rect 674944 874262 675064 874290
rect 675312 874262 675432 874290
rect 675036 874177 675064 874262
rect 675022 874168 675078 874177
rect 675022 874103 675078 874112
rect 675482 874168 675538 874177
rect 675482 874103 675538 874112
rect 675496 873868 675524 874103
rect 675116 873656 675168 873662
rect 675116 873598 675168 873604
rect 675128 872590 675156 873598
rect 675574 873488 675630 873497
rect 675574 873423 675630 873432
rect 675588 873188 675616 873423
rect 675128 872562 675248 872590
rect 675220 872522 675248 872562
rect 675404 872522 675432 872576
rect 675220 872494 675432 872522
rect 674840 872432 674892 872438
rect 674840 872374 674892 872380
rect 675300 872432 675352 872438
rect 675300 872374 675352 872380
rect 675312 870074 675340 872374
rect 675312 870046 675418 870074
rect 674656 869848 674708 869854
rect 674656 869790 674708 869796
rect 675208 869848 675260 869854
rect 675208 869790 675260 869796
rect 675758 869816 675814 869825
rect 674380 869644 674432 869650
rect 674380 869586 674432 869592
rect 674840 869644 674892 869650
rect 674840 869586 674892 869592
rect 674852 869258 674880 869586
rect 675024 869440 675076 869446
rect 675024 869382 675076 869388
rect 674852 869230 674972 869258
rect 674748 868080 674800 868086
rect 674800 868028 674880 868034
rect 674748 868022 674880 868028
rect 674760 868006 674880 868022
rect 674852 866289 674880 868006
rect 674944 867354 674972 869230
rect 675036 867694 675064 869382
rect 675220 868889 675248 869790
rect 675758 869751 675814 869760
rect 675772 869516 675800 869751
rect 675220 868861 675418 868889
rect 675758 868728 675814 868737
rect 675758 868663 675814 868672
rect 675772 868224 675800 868663
rect 675036 867666 675418 867694
rect 674944 867326 675432 867354
rect 675114 867232 675170 867241
rect 675114 867167 675170 867176
rect 674838 866280 674894 866289
rect 674838 866215 674894 866224
rect 675128 866130 675156 867167
rect 675404 867035 675432 867326
rect 675390 866280 675446 866289
rect 675390 866215 675446 866224
rect 675128 866102 675340 866130
rect 675114 865736 675170 865745
rect 675114 865671 675170 865680
rect 675128 863342 675156 865671
rect 675312 864566 675340 866102
rect 675404 865844 675432 866215
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675312 864538 675418 864566
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675116 789404 675168 789410
rect 675116 789346 675168 789352
rect 675128 787693 675156 789346
rect 675404 788868 675432 790774
rect 675404 788089 675432 788324
rect 675390 788080 675446 788089
rect 675390 788015 675446 788024
rect 675128 787665 675418 787693
rect 675496 786729 675524 787032
rect 675482 786720 675538 786729
rect 675482 786655 675538 786664
rect 674852 785182 675418 785210
rect 673736 782672 673788 782678
rect 673736 782614 673788 782620
rect 673552 778592 673604 778598
rect 673552 778534 673604 778540
rect 673564 770054 673592 778534
rect 673564 770026 673684 770054
rect 673656 743834 673684 770026
rect 673104 727926 673408 727954
rect 673472 743806 673684 743834
rect 673748 743834 673776 782614
rect 673920 780020 673972 780026
rect 673920 779962 673972 779968
rect 673932 760394 673960 779962
rect 674288 777028 674340 777034
rect 674288 776970 674340 776976
rect 673840 760366 673960 760394
rect 673840 750734 673868 760366
rect 673840 750706 673960 750734
rect 673748 743806 673868 743834
rect 673104 723194 673132 727926
rect 673472 727870 673500 743806
rect 673644 734324 673696 734330
rect 673644 734266 673696 734272
rect 673656 734174 673684 734266
rect 673840 734174 673868 743806
rect 673564 734146 673684 734174
rect 673748 734146 673868 734174
rect 673564 732794 673592 734146
rect 673564 732766 673684 732794
rect 673460 727864 673512 727870
rect 673460 727806 673512 727812
rect 673656 723738 673684 732766
rect 673380 723710 673684 723738
rect 673104 723166 673316 723194
rect 673288 721698 673316 723166
rect 672920 717586 673040 717614
rect 673104 721670 673316 721698
rect 673380 721698 673408 723710
rect 673552 723172 673604 723178
rect 673472 723120 673552 723134
rect 673472 723114 673604 723120
rect 673472 723106 673592 723114
rect 673472 722378 673500 723106
rect 673472 722350 673592 722378
rect 673564 721970 673592 722350
rect 673748 722226 673776 734146
rect 673736 722220 673788 722226
rect 673736 722162 673788 722168
rect 673736 722084 673788 722090
rect 673736 722026 673788 722032
rect 673564 721942 673684 721970
rect 673380 721670 673500 721698
rect 672722 714096 672778 714105
rect 672722 714031 672778 714040
rect 672736 669497 672764 714031
rect 672920 709209 672948 717586
rect 673104 712881 673132 721670
rect 673274 721576 673330 721585
rect 673274 721511 673330 721520
rect 673288 714854 673316 721511
rect 673472 719522 673500 721670
rect 673472 719494 673592 719522
rect 673288 714826 673500 714854
rect 673090 712872 673146 712881
rect 673090 712807 673146 712816
rect 672906 709200 672962 709209
rect 672906 709135 672962 709144
rect 673274 706344 673330 706353
rect 673274 706279 673330 706288
rect 673288 698294 673316 706279
rect 673472 701486 673500 714826
rect 673564 705194 673592 719494
rect 673656 708914 673684 721942
rect 673748 712858 673776 722026
rect 673932 722022 673960 750706
rect 674300 746594 674328 776970
rect 674656 775736 674708 775742
rect 674656 775678 674708 775684
rect 674300 746566 674420 746594
rect 674196 738676 674248 738682
rect 674196 738618 674248 738624
rect 674208 727274 674236 738618
rect 674024 727246 674236 727274
rect 674024 722106 674052 727246
rect 674392 726646 674420 746566
rect 674668 727938 674696 775678
rect 674852 770054 674880 785182
rect 675128 784638 675418 784666
rect 675128 783902 675156 784638
rect 675116 783896 675168 783902
rect 675496 783873 675524 783972
rect 675116 783838 675168 783844
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675128 783346 675418 783374
rect 675128 782678 675156 783346
rect 675116 782672 675168 782678
rect 675116 782614 675168 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675024 781244 675076 781250
rect 675024 781186 675076 781192
rect 675036 781130 675064 781186
rect 674944 781102 675064 781130
rect 674944 779714 674972 781102
rect 675404 780844 675432 781374
rect 675312 780422 675432 780450
rect 675312 780314 675340 780422
rect 675128 780286 675340 780314
rect 675404 780300 675432 780422
rect 675128 780026 675156 780286
rect 675116 780020 675168 780026
rect 675116 779962 675168 779968
rect 675758 779920 675814 779929
rect 675758 779855 675814 779864
rect 674944 779686 675156 779714
rect 675772 779686 675800 779855
rect 675128 778478 675156 779686
rect 675312 779062 675432 779090
rect 675312 778598 675340 779062
rect 675404 779008 675432 779062
rect 675300 778592 675352 778598
rect 675300 778534 675352 778540
rect 675128 778450 675418 778478
rect 675116 778388 675168 778394
rect 675116 778330 675168 778336
rect 675128 776642 675156 778330
rect 675404 777322 675432 777852
rect 675312 777294 675432 777322
rect 675312 777034 675340 777294
rect 675300 777028 675352 777034
rect 675300 776970 675352 776976
rect 675128 776614 675418 776642
rect 675128 776002 675340 776030
rect 675128 775742 675156 776002
rect 675312 775962 675340 776002
rect 675404 775962 675432 776016
rect 675312 775934 675432 775962
rect 675116 775736 675168 775742
rect 675116 775678 675168 775684
rect 675024 775600 675076 775606
rect 674944 775548 675024 775554
rect 674944 775542 675076 775548
rect 674944 775526 675064 775542
rect 674944 774194 674972 775526
rect 675128 775322 675418 775350
rect 675128 774314 675156 775322
rect 675116 774308 675168 774314
rect 675116 774250 675168 774256
rect 674944 774166 675340 774194
rect 675312 774058 675340 774166
rect 675404 774058 675432 774180
rect 675312 774030 675432 774058
rect 674852 770026 675340 770054
rect 675312 750734 675340 770026
rect 674852 750706 675340 750734
rect 674852 742257 674880 750706
rect 675024 745272 675076 745278
rect 674944 745220 675024 745226
rect 674944 745214 675076 745220
rect 674944 745198 675064 745214
rect 674944 743322 674972 745198
rect 675312 743974 675432 744002
rect 675312 743866 675340 743974
rect 675128 743850 675340 743866
rect 675404 743852 675432 743974
rect 675116 743844 675340 743850
rect 675168 743838 675340 743844
rect 675116 743786 675168 743792
rect 674944 743294 675418 743322
rect 675404 742529 675432 742696
rect 675390 742520 675446 742529
rect 675390 742455 675446 742464
rect 674838 742248 674894 742257
rect 674838 742183 674894 742192
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 674944 742002 675340 742030
rect 675404 742016 675432 742070
rect 674944 741962 674972 742002
rect 674760 741934 674972 741962
rect 674760 734174 674788 741934
rect 675312 740166 675418 740194
rect 675312 739242 675340 740166
rect 675036 739214 675340 739242
rect 675036 736658 675064 739214
rect 675404 739158 675432 739636
rect 675392 739152 675444 739158
rect 675392 739094 675444 739100
rect 675404 738682 675432 739024
rect 675392 738676 675444 738682
rect 675392 738618 675444 738624
rect 675220 738330 675418 738358
rect 675220 738177 675248 738330
rect 675206 738168 675262 738177
rect 675206 738103 675262 738112
rect 675300 736976 675352 736982
rect 675300 736918 675352 736924
rect 675036 736630 675156 736658
rect 675128 736409 675156 736630
rect 674930 736400 674986 736409
rect 674930 736335 674986 736344
rect 675114 736400 675170 736409
rect 675114 736335 675170 736344
rect 674760 734146 674880 734174
rect 674656 727932 674708 727938
rect 674656 727874 674708 727880
rect 674852 727818 674880 734146
rect 674668 727790 674880 727818
rect 674668 727326 674696 727790
rect 674944 727682 674972 736335
rect 675312 735333 675340 736918
rect 675482 736128 675538 736137
rect 675482 736063 675538 736072
rect 675496 735896 675524 736063
rect 675312 735305 675418 735333
rect 675298 735040 675354 735049
rect 675036 734998 675298 735026
rect 675036 729858 675064 734998
rect 675298 734975 675354 734984
rect 675208 734868 675260 734874
rect 675208 734810 675260 734816
rect 675220 734754 675248 734810
rect 675128 734726 675248 734754
rect 675128 733428 675156 734726
rect 675312 734658 675418 734686
rect 675312 734330 675340 734658
rect 675300 734324 675352 734330
rect 675300 734266 675352 734272
rect 675482 734224 675538 734233
rect 675312 734168 675482 734174
rect 675312 734159 675538 734168
rect 675312 734146 675524 734159
rect 675312 733650 675340 734146
rect 675496 733825 675524 734031
rect 675482 733816 675538 733825
rect 675482 733751 675538 733760
rect 675300 733644 675352 733650
rect 675300 733586 675352 733592
rect 675312 733465 675418 733493
rect 675312 733428 675340 733465
rect 675128 733400 675340 733428
rect 675300 733304 675352 733310
rect 675300 733246 675352 733252
rect 675312 732034 675340 733246
rect 675758 733000 675814 733009
rect 675758 732935 675814 732944
rect 675772 732836 675800 732935
rect 675312 732006 675432 732034
rect 675404 731612 675432 732006
rect 675220 730986 675418 731014
rect 675220 730522 675248 730986
rect 675208 730516 675260 730522
rect 675208 730458 675260 730464
rect 675220 730337 675418 730365
rect 675220 729978 675248 730337
rect 675208 729972 675260 729978
rect 675208 729914 675260 729920
rect 675036 729830 675156 729858
rect 675128 727802 675156 729830
rect 675312 729150 675418 729178
rect 675312 728686 675340 729150
rect 675300 728680 675352 728686
rect 675300 728622 675352 728628
rect 675758 728376 675814 728385
rect 675758 728311 675814 728320
rect 675116 727796 675168 727802
rect 675116 727738 675168 727744
rect 674944 727666 675064 727682
rect 674944 727660 675076 727666
rect 674944 727654 675024 727660
rect 675024 727602 675076 727608
rect 674840 727456 674892 727462
rect 674840 727398 674892 727404
rect 674656 727320 674708 727326
rect 674656 727262 674708 727268
rect 674380 726640 674432 726646
rect 674380 726582 674432 726588
rect 674852 723217 674880 727398
rect 675024 727320 675076 727326
rect 675024 727262 675076 727268
rect 674838 723208 674894 723217
rect 674838 723143 674894 723152
rect 674024 722078 674144 722106
rect 673920 722016 673972 722022
rect 673920 721958 673972 721964
rect 674116 721857 674144 722078
rect 674102 721848 674158 721857
rect 673920 721812 673972 721818
rect 674102 721783 674158 721792
rect 673920 721754 673972 721760
rect 673932 720594 673960 721754
rect 675036 721721 675064 727262
rect 675772 721750 675800 728311
rect 675942 728104 675998 728113
rect 675942 728039 675998 728048
rect 675956 721750 675984 728039
rect 683304 727932 683356 727938
rect 683304 727874 683356 727880
rect 677324 727796 677376 727802
rect 677324 727738 677376 727744
rect 675760 721744 675812 721750
rect 675022 721712 675078 721721
rect 675760 721686 675812 721692
rect 675944 721744 675996 721750
rect 675944 721686 675996 721692
rect 675022 721647 675078 721656
rect 675760 721268 675812 721274
rect 675760 721210 675812 721216
rect 675944 721268 675996 721274
rect 675944 721210 675996 721216
rect 675772 720866 675800 721210
rect 675956 720866 675984 721210
rect 675760 720860 675812 720866
rect 675760 720802 675812 720808
rect 675944 720860 675996 720866
rect 675944 720802 675996 720808
rect 673920 720588 673972 720594
rect 673920 720530 673972 720536
rect 675760 720520 675812 720526
rect 675760 720462 675812 720468
rect 675944 720520 675996 720526
rect 675944 720462 675996 720468
rect 673920 720452 673972 720458
rect 673920 720394 673972 720400
rect 673932 717618 673960 720394
rect 673840 717590 673960 717618
rect 675772 717614 675800 720462
rect 675956 717614 675984 720462
rect 673840 712994 673868 717590
rect 675680 717586 675800 717614
rect 675864 717586 675984 717614
rect 674288 716508 674340 716514
rect 674288 716450 674340 716456
rect 674300 716394 674328 716450
rect 674024 716366 674328 716394
rect 674024 716310 674052 716366
rect 674012 716304 674064 716310
rect 674012 716246 674064 716252
rect 674012 715760 674064 715766
rect 674010 715728 674012 715737
rect 674064 715728 674066 715737
rect 674010 715663 674066 715672
rect 674012 715352 674064 715358
rect 674010 715320 674012 715329
rect 674064 715320 674066 715329
rect 674010 715255 674066 715264
rect 674010 715048 674066 715057
rect 674010 714983 674012 714992
rect 674064 714983 674066 714992
rect 674012 714954 674064 714960
rect 674288 714944 674340 714950
rect 674024 714892 674288 714898
rect 674024 714886 674340 714892
rect 674024 714882 674328 714886
rect 674012 714876 674328 714882
rect 674064 714870 674328 714876
rect 674012 714818 674064 714824
rect 674012 714536 674064 714542
rect 674010 714504 674012 714513
rect 674064 714504 674066 714513
rect 674010 714439 674066 714448
rect 674012 713720 674064 713726
rect 674010 713688 674012 713697
rect 674064 713688 674066 713697
rect 674010 713623 674066 713632
rect 674010 713280 674066 713289
rect 674010 713215 674012 713224
rect 674064 713215 674066 713224
rect 674012 713186 674064 713192
rect 673840 712966 674604 712994
rect 673748 712830 674512 712858
rect 674010 712464 674066 712473
rect 674010 712399 674012 712408
rect 674064 712399 674066 712408
rect 674012 712370 674064 712376
rect 674012 710048 674064 710054
rect 674010 710016 674012 710025
rect 674064 710016 674066 710025
rect 674010 709951 674066 709960
rect 674012 709640 674064 709646
rect 674010 709608 674012 709617
rect 674064 709608 674066 709617
rect 674010 709543 674066 709552
rect 674288 709572 674340 709578
rect 674288 709514 674340 709520
rect 674300 709458 674328 709514
rect 674024 709430 674328 709458
rect 674024 709374 674052 709430
rect 674012 709368 674064 709374
rect 674012 709310 674064 709316
rect 673656 708886 673960 708914
rect 673932 707954 673960 708886
rect 674288 708008 674340 708014
rect 674288 707954 674340 707956
rect 673932 707950 674340 707954
rect 673932 707926 674328 707950
rect 674484 707606 674512 712830
rect 674576 707954 674604 712966
rect 675680 712065 675708 717586
rect 675666 712056 675722 712065
rect 675666 711991 675722 712000
rect 675864 711249 675892 717586
rect 676034 716544 676090 716553
rect 676034 716479 676036 716488
rect 676088 716479 676090 716488
rect 676036 716450 676088 716456
rect 676034 716136 676090 716145
rect 676034 716071 676090 716080
rect 676048 714950 676076 716071
rect 676036 714944 676088 714950
rect 676036 714886 676088 714892
rect 677336 712094 677364 727738
rect 676220 712088 676272 712094
rect 676220 712030 676272 712036
rect 677324 712088 677376 712094
rect 677324 712030 677376 712036
rect 675850 711240 675906 711249
rect 675850 711175 675906 711184
rect 676034 710832 676090 710841
rect 676232 710818 676260 712030
rect 683316 711657 683344 727874
rect 683488 726640 683540 726646
rect 683488 726582 683540 726588
rect 683302 711648 683358 711657
rect 683302 711583 683358 711592
rect 676090 710790 676260 710818
rect 676034 710767 676090 710776
rect 676034 710424 676090 710433
rect 676034 710359 676090 710368
rect 676048 709578 676076 710359
rect 676036 709572 676088 709578
rect 676036 709514 676088 709520
rect 683500 708393 683528 726582
rect 684130 726472 684186 726481
rect 684130 726407 684186 726416
rect 684144 708801 684172 726407
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684130 708792 684186 708801
rect 684130 708727 684186 708736
rect 683486 708384 683542 708393
rect 683486 708319 683542 708328
rect 675852 708008 675904 708014
rect 674576 707926 674696 707954
rect 675852 707950 675904 707956
rect 674472 707600 674524 707606
rect 674472 707542 674524 707548
rect 674668 707198 674696 707926
rect 674656 707192 674708 707198
rect 674656 707134 674708 707140
rect 675864 706761 675892 707950
rect 676036 707600 676088 707606
rect 676034 707568 676036 707577
rect 676088 707568 676090 707577
rect 676034 707503 676090 707512
rect 676036 707192 676088 707198
rect 676034 707160 676036 707169
rect 676088 707160 676090 707169
rect 676034 707095 676090 707104
rect 675850 706752 675906 706761
rect 675850 706687 675906 706696
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 674012 705424 674064 705430
rect 674064 705372 674328 705378
rect 674012 705366 674328 705372
rect 674024 705362 674328 705366
rect 683132 705362 683160 705463
rect 674024 705356 674340 705362
rect 674024 705350 674288 705356
rect 674288 705298 674340 705304
rect 683120 705356 683172 705362
rect 683120 705298 683172 705304
rect 673564 705166 673684 705194
rect 673460 701480 673512 701486
rect 673460 701422 673512 701428
rect 673656 701162 673684 705166
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 703866 676076 705055
rect 674012 703860 674064 703866
rect 674288 703860 674340 703866
rect 674064 703820 674288 703848
rect 674012 703802 674064 703808
rect 674288 703802 674340 703808
rect 676036 703860 676088 703866
rect 676036 703802 676088 703808
rect 673920 701480 673972 701486
rect 673564 701134 673684 701162
rect 673840 701428 673920 701434
rect 673840 701422 673972 701428
rect 673840 701406 673960 701422
rect 673288 698266 673408 698294
rect 673182 697232 673238 697241
rect 673182 697167 673238 697176
rect 672906 687848 672962 687857
rect 672906 687783 672962 687792
rect 672722 669488 672778 669497
rect 672722 669423 672778 669432
rect 672540 665440 672592 665446
rect 672540 665382 672592 665388
rect 672722 651400 672778 651409
rect 672722 651335 672778 651344
rect 672356 619064 672408 619070
rect 672356 619006 672408 619012
rect 672354 603800 672410 603809
rect 672354 603735 672410 603744
rect 672368 527202 672396 603735
rect 672538 597408 672594 597417
rect 672538 597343 672594 597352
rect 672552 527406 672580 597343
rect 672736 576609 672764 651335
rect 672920 618225 672948 687783
rect 673196 619449 673224 697167
rect 673182 619440 673238 619449
rect 673182 619375 673238 619384
rect 672906 618216 672962 618225
rect 672906 618151 672962 618160
rect 673090 604208 673146 604217
rect 673090 604143 673146 604152
rect 672722 576600 672778 576609
rect 672722 576535 672778 576544
rect 672906 553344 672962 553353
rect 672906 553279 672962 553288
rect 672724 535016 672776 535022
rect 672722 534984 672724 534993
rect 672776 534984 672778 534993
rect 672722 534919 672778 534928
rect 672722 533488 672778 533497
rect 672722 533423 672778 533432
rect 672540 527400 672592 527406
rect 672540 527342 672592 527348
rect 672356 527196 672408 527202
rect 672356 527138 672408 527144
rect 672736 490113 672764 533423
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672630 489696 672686 489705
rect 672630 489631 672686 489640
rect 672172 455864 672224 455870
rect 672172 455806 672224 455812
rect 672000 455122 672120 455138
rect 672000 455116 672132 455122
rect 672000 455110 672080 455116
rect 672080 455058 672132 455064
rect 672448 453960 672500 453966
rect 672446 453928 672448 453937
rect 672500 453928 672502 453937
rect 672446 453863 672502 453872
rect 60002 430672 60058 430681
rect 60002 430607 60058 430616
rect 45834 427408 45890 427417
rect 45834 427343 45890 427352
rect 45664 427230 45784 427258
rect 45558 426864 45614 426873
rect 45558 426799 45614 426808
rect 44914 423192 44970 423201
rect 44914 423127 44970 423136
rect 44928 402937 44956 423127
rect 45098 421560 45154 421569
rect 45098 421495 45154 421504
rect 45112 406745 45140 421495
rect 45282 421152 45338 421161
rect 45282 421087 45338 421096
rect 45296 408105 45324 421087
rect 45282 408096 45338 408105
rect 45282 408031 45338 408040
rect 45098 406736 45154 406745
rect 45098 406671 45154 406680
rect 45282 405648 45338 405657
rect 45282 405583 45338 405592
rect 45296 402966 45324 405583
rect 45284 402960 45336 402966
rect 44914 402928 44970 402937
rect 45284 402902 45336 402908
rect 44914 402863 44970 402872
rect 44638 386472 44694 386481
rect 44638 386407 44694 386416
rect 44270 385656 44326 385665
rect 44270 385591 44326 385600
rect 45098 385248 45154 385257
rect 45098 385183 45154 385192
rect 44362 379128 44418 379137
rect 44362 379063 44418 379072
rect 44178 376272 44234 376281
rect 44178 376207 44234 376216
rect 44192 359666 44220 376207
rect 44376 364177 44404 379063
rect 44546 378720 44602 378729
rect 44546 378655 44602 378664
rect 44362 364168 44418 364177
rect 44362 364103 44418 364112
rect 44560 361593 44588 378655
rect 44730 377904 44786 377913
rect 44730 377839 44786 377848
rect 44744 364857 44772 377839
rect 44914 377496 44970 377505
rect 44914 377431 44970 377440
rect 44730 364848 44786 364857
rect 44730 364783 44786 364792
rect 44928 364334 44956 377431
rect 45112 369854 45140 385183
rect 45572 384033 45600 426799
rect 45756 418154 45784 427230
rect 46018 424008 46074 424017
rect 46018 423943 46074 423952
rect 45756 418126 45876 418154
rect 45848 384849 45876 418126
rect 46032 400217 46060 423943
rect 53838 407824 53894 407833
rect 53838 407759 53894 407768
rect 53852 404326 53880 407759
rect 53840 404320 53892 404326
rect 53840 404262 53892 404268
rect 51080 400240 51132 400246
rect 46018 400208 46074 400217
rect 51080 400182 51132 400188
rect 46018 400143 46074 400152
rect 51092 395729 51120 400182
rect 60016 400110 60044 430607
rect 61382 429312 61438 429321
rect 61382 429247 61438 429256
rect 60004 400104 60056 400110
rect 60004 400046 60056 400052
rect 61396 398313 61424 429247
rect 63130 427136 63186 427145
rect 63130 427071 63186 427080
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400616 62174 400625
rect 62118 400551 62174 400560
rect 62132 400246 62160 400551
rect 62120 400240 62172 400246
rect 63144 400217 63172 427071
rect 657542 403336 657598 403345
rect 657542 403271 657598 403280
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 62120 400182 62172 400188
rect 63130 400208 63186 400217
rect 63130 400143 63186 400152
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 61382 398304 61438 398313
rect 61382 398239 61438 398248
rect 51078 395720 51134 395729
rect 51078 395655 51134 395664
rect 61382 386472 61438 386481
rect 61382 386407 61438 386416
rect 45834 384840 45890 384849
rect 45834 384775 45890 384784
rect 46018 384432 46074 384441
rect 46018 384367 46074 384376
rect 45558 384024 45614 384033
rect 45558 383959 45614 383968
rect 45650 383616 45706 383625
rect 45650 383551 45706 383560
rect 45282 381440 45338 381449
rect 45282 381375 45338 381384
rect 45296 369854 45324 381375
rect 44836 364306 44956 364334
rect 45020 369826 45140 369854
rect 45204 369826 45324 369854
rect 44546 361584 44602 361593
rect 44546 361519 44602 361528
rect 44192 359650 44680 359666
rect 44192 359644 44692 359650
rect 44192 359638 44640 359644
rect 44640 359586 44692 359592
rect 44836 359514 44864 364306
rect 44824 359508 44876 359514
rect 44824 359450 44876 359456
rect 44822 355192 44878 355201
rect 44822 355127 44878 355136
rect 44638 354920 44694 354929
rect 44638 354855 44694 354864
rect 44652 354754 44680 354855
rect 44836 354754 44864 355127
rect 44640 354748 44692 354754
rect 44640 354690 44692 354696
rect 44824 354748 44876 354754
rect 44824 354690 44876 354696
rect 43732 354606 43944 354634
rect 44008 354606 44895 354634
rect 43916 354498 43944 354606
rect 43916 354482 44772 354498
rect 44867 354482 44895 354606
rect 43916 354476 44784 354482
rect 43916 354470 44732 354476
rect 44732 354418 44784 354424
rect 44855 354476 44907 354482
rect 44855 354418 44907 354424
rect 43258 353696 43314 353705
rect 43258 353631 43314 353640
rect 42338 353016 42394 353025
rect 42338 352951 42394 352960
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35808 344616 35860 344622
rect 35808 344558 35860 344564
rect 39856 344616 39908 344622
rect 39856 344558 39908 344564
rect 35820 344321 35848 344558
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 35622 343904 35678 343913
rect 35622 343839 35678 343848
rect 35636 343670 35664 343839
rect 35624 343664 35676 343670
rect 35624 343606 35676 343612
rect 35806 343496 35862 343505
rect 35806 343431 35862 343440
rect 35820 342242 35848 343431
rect 35808 342236 35860 342242
rect 35808 342178 35860 342184
rect 39868 341873 39896 344558
rect 40406 343904 40462 343913
rect 40406 343839 40462 343848
rect 40040 343664 40092 343670
rect 40040 343606 40092 343612
rect 35806 341864 35862 341873
rect 35806 341799 35862 341808
rect 39670 341864 39726 341873
rect 39670 341799 39726 341808
rect 39854 341864 39910 341873
rect 39854 341799 39910 341808
rect 35820 341562 35848 341799
rect 35808 341556 35860 341562
rect 35808 341498 35860 341504
rect 35808 341080 35860 341086
rect 35806 341048 35808 341057
rect 35860 341048 35862 341057
rect 35806 340983 35862 340992
rect 39684 340241 39712 341799
rect 40052 341442 40080 343606
rect 40222 342272 40278 342281
rect 40222 342207 40224 342216
rect 40276 342207 40278 342216
rect 40224 342178 40276 342184
rect 40420 341578 40448 343839
rect 45020 342553 45048 369826
rect 45204 343369 45232 369826
rect 45374 362944 45430 362953
rect 45374 362879 45430 362888
rect 45388 360194 45416 362879
rect 45376 360188 45428 360194
rect 45376 360130 45428 360136
rect 45376 359644 45428 359650
rect 45296 359592 45376 359598
rect 45296 359586 45428 359592
rect 45296 359570 45416 359586
rect 45296 353818 45324 359570
rect 45468 359508 45520 359514
rect 45468 359450 45520 359456
rect 45296 353790 45343 353818
rect 45315 353530 45343 353790
rect 45303 353524 45355 353530
rect 45303 353466 45355 353472
rect 45480 353274 45508 359450
rect 45434 353258 45508 353274
rect 45422 353252 45508 353258
rect 45474 353246 45508 353252
rect 45422 353194 45474 353200
rect 45190 343360 45246 343369
rect 45190 343295 45246 343304
rect 45006 342544 45062 342553
rect 45006 342479 45062 342488
rect 45466 342272 45522 342281
rect 45466 342207 45468 342216
rect 45520 342207 45522 342216
rect 45468 342178 45520 342184
rect 40236 341562 40448 341578
rect 40224 341556 40448 341562
rect 40276 341550 40448 341556
rect 40224 341498 40276 341504
rect 40052 341414 40540 341442
rect 40512 341306 40540 341414
rect 42246 341320 42302 341329
rect 40512 341278 42246 341306
rect 42246 341255 42302 341264
rect 40132 341080 40184 341086
rect 40130 341048 40132 341057
rect 40184 341048 40186 341057
rect 40130 340983 40186 340992
rect 45664 340785 45692 383551
rect 45834 353968 45890 353977
rect 45834 353903 45836 353912
rect 45888 353903 45890 353912
rect 45836 353874 45888 353880
rect 45836 353728 45888 353734
rect 45834 353696 45836 353705
rect 45888 353696 45890 353705
rect 45834 353631 45890 353640
rect 46032 343913 46060 384367
rect 47122 383208 47178 383217
rect 47122 383143 47178 383152
rect 46938 382392 46994 382401
rect 46938 382327 46994 382336
rect 46570 363216 46626 363225
rect 46570 363151 46626 363160
rect 46584 361554 46612 363151
rect 46572 361548 46624 361554
rect 46572 361490 46624 361496
rect 46952 353025 46980 382327
rect 47136 354385 47164 383143
rect 51724 357468 51776 357474
rect 51724 357410 51776 357416
rect 47122 354376 47178 354385
rect 47122 354311 47178 354320
rect 51736 353297 51764 357410
rect 61396 356017 61424 386407
rect 63406 385928 63462 385937
rect 63406 385863 63462 385872
rect 62946 381848 63002 381857
rect 62946 381783 63002 381792
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62118 357776 62174 357785
rect 62118 357711 62174 357720
rect 62132 357474 62160 357711
rect 62120 357468 62172 357474
rect 62120 357410 62172 357416
rect 61382 356008 61438 356017
rect 61382 355943 61438 355952
rect 62960 354521 62988 381783
rect 63420 357377 63448 385863
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 395312 652262 395321
rect 652206 395247 652262 395256
rect 652220 373969 652248 395247
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 654796 371006 654824 382871
rect 657556 373998 657584 403271
rect 672644 401713 672672 489631
rect 672920 482361 672948 553279
rect 673104 528873 673132 604143
rect 673090 528864 673146 528873
rect 673090 528799 673146 528808
rect 672906 482352 672962 482361
rect 672906 482287 672962 482296
rect 673380 456006 673408 698266
rect 673564 687585 673592 701134
rect 673840 700890 673868 701406
rect 674024 701282 674328 701298
rect 674012 701276 674340 701282
rect 674064 701270 674288 701276
rect 674012 701218 674064 701224
rect 674288 701218 674340 701224
rect 675116 701276 675168 701282
rect 675116 701218 675168 701224
rect 674012 701072 674064 701078
rect 674288 701072 674340 701078
rect 674064 701020 674288 701026
rect 674012 701014 674340 701020
rect 674024 700998 674328 701014
rect 673840 700862 673960 700890
rect 673736 696992 673788 696998
rect 673734 696960 673736 696969
rect 673788 696960 673790 696969
rect 673734 696895 673790 696904
rect 673734 690160 673790 690169
rect 673734 690095 673736 690104
rect 673788 690095 673790 690104
rect 673736 690066 673788 690072
rect 673736 688832 673788 688838
rect 673734 688800 673736 688809
rect 673788 688800 673790 688809
rect 673734 688735 673790 688744
rect 673734 688120 673790 688129
rect 673734 688055 673790 688064
rect 673550 687576 673606 687585
rect 673550 687511 673606 687520
rect 673550 671392 673606 671401
rect 673550 671327 673606 671336
rect 673564 670750 673592 671327
rect 673552 670744 673604 670750
rect 673552 670686 673604 670692
rect 673550 670576 673606 670585
rect 673550 670511 673606 670520
rect 673564 669526 673592 670511
rect 673552 669520 673604 669526
rect 673552 669462 673604 669468
rect 673550 668944 673606 668953
rect 673550 668879 673606 668888
rect 673564 668234 673592 668879
rect 673552 668228 673604 668234
rect 673552 668170 673604 668176
rect 673550 667312 673606 667321
rect 673550 667247 673606 667256
rect 673564 666602 673592 667247
rect 673552 666596 673604 666602
rect 673552 666538 673604 666544
rect 673550 666360 673606 666369
rect 673550 666295 673606 666304
rect 673564 665446 673592 666295
rect 673552 665440 673604 665446
rect 673552 665382 673604 665388
rect 673552 626000 673604 626006
rect 673550 625968 673552 625977
rect 673604 625968 673606 625977
rect 673550 625903 673606 625912
rect 673748 621014 673776 688055
rect 673932 671673 673960 700862
rect 675128 698337 675156 701218
rect 675392 701072 675444 701078
rect 675392 701014 675444 701020
rect 675404 698875 675432 701014
rect 675128 698309 675418 698337
rect 675128 697666 675418 697694
rect 675128 697241 675156 697666
rect 675114 697232 675170 697241
rect 675114 697167 675170 697176
rect 675220 697054 675432 697082
rect 675220 697049 675248 697054
rect 675128 697021 675248 697049
rect 675404 697035 675432 697054
rect 675128 696697 675156 697021
rect 675298 696960 675354 696969
rect 675298 696895 675354 696904
rect 675114 696688 675170 696697
rect 675114 696623 675170 696632
rect 675312 695722 675340 696895
rect 675312 695694 675524 695722
rect 675298 695464 675354 695473
rect 675298 695399 675354 695408
rect 675312 695042 675340 695399
rect 675496 695195 675524 695694
rect 675312 695014 675432 695042
rect 675404 694620 675432 695014
rect 675404 693530 675432 694008
rect 674472 693524 674524 693530
rect 674472 693466 674524 693472
rect 675392 693524 675444 693530
rect 675392 693466 675444 693472
rect 674288 693048 674340 693054
rect 674288 692990 674340 692996
rect 674102 689480 674158 689489
rect 674102 689415 674158 689424
rect 673918 671664 673974 671673
rect 673918 671599 673974 671608
rect 673920 671152 673972 671158
rect 673920 671094 673972 671100
rect 673932 670993 673960 671094
rect 673918 670984 673974 670993
rect 673918 670919 673974 670928
rect 673918 670168 673974 670177
rect 673918 670103 673920 670112
rect 673972 670103 673974 670112
rect 673920 670074 673972 670080
rect 673918 669760 673974 669769
rect 673918 669695 673974 669704
rect 673932 669390 673960 669695
rect 673920 669384 673972 669390
rect 673920 669326 673972 669332
rect 673920 668568 673972 668574
rect 673918 668536 673920 668545
rect 673972 668536 673974 668545
rect 673918 668471 673974 668480
rect 673918 668128 673974 668137
rect 673918 668063 673974 668072
rect 673932 667962 673960 668063
rect 673920 667956 673972 667962
rect 673920 667898 673972 667904
rect 673918 667720 673974 667729
rect 673918 667655 673974 667664
rect 673932 666942 673960 667655
rect 673920 666936 673972 666942
rect 673920 666878 673972 666884
rect 673918 666088 673974 666097
rect 673918 666023 673920 666032
rect 673972 666023 673974 666032
rect 673920 665994 673972 666000
rect 673918 665272 673974 665281
rect 673918 665207 673920 665216
rect 673972 665207 673974 665216
rect 673920 665178 673972 665184
rect 673918 664864 673974 664873
rect 673918 664799 673974 664808
rect 673932 664494 673960 664799
rect 673920 664488 673972 664494
rect 673920 664430 673972 664436
rect 673918 664048 673974 664057
rect 673918 663983 673920 663992
rect 673972 663983 673974 663992
rect 673920 663954 673972 663960
rect 673918 662008 673974 662017
rect 673918 661943 673920 661952
rect 673972 661943 673974 661952
rect 673920 661914 673972 661920
rect 673920 661632 673972 661638
rect 673918 661600 673920 661609
rect 673972 661600 673974 661609
rect 673918 661535 673974 661544
rect 673918 661192 673974 661201
rect 673918 661127 673920 661136
rect 673972 661127 673974 661136
rect 673920 661098 673972 661104
rect 673918 660240 673974 660249
rect 673918 660175 673920 660184
rect 673972 660175 673974 660184
rect 673920 660146 673972 660152
rect 673918 659968 673974 659977
rect 673918 659903 673974 659912
rect 673932 659734 673960 659903
rect 673920 659728 673972 659734
rect 673920 659670 673972 659676
rect 673918 655616 673974 655625
rect 673918 655551 673920 655560
rect 673972 655551 673974 655560
rect 673920 655522 673972 655528
rect 674116 654134 674144 689415
rect 674300 688129 674328 692990
rect 674286 688120 674342 688129
rect 674286 688055 674342 688064
rect 674484 683114 674512 693466
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 675128 693314 675340 693342
rect 675404 693328 675432 693382
rect 675128 693054 675156 693314
rect 675116 693048 675168 693054
rect 675116 692990 675168 692996
rect 675128 690866 675418 690894
rect 675128 690441 675156 690866
rect 675114 690432 675170 690441
rect 675114 690367 675170 690376
rect 674930 690160 674986 690169
rect 674930 690095 674986 690104
rect 674944 688922 674972 690095
rect 675404 689897 675432 690336
rect 675390 689888 675446 689897
rect 675390 689823 675446 689832
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689489 675156 689642
rect 675114 689480 675170 689489
rect 675114 689415 675170 689424
rect 675114 689208 675170 689217
rect 675114 689143 675170 689152
rect 675128 689058 675156 689143
rect 675128 689030 675418 689058
rect 674944 688894 675156 688922
rect 674930 688800 674986 688809
rect 674930 688735 674986 688744
rect 674654 687576 674710 687585
rect 674654 687511 674710 687520
rect 674668 683114 674696 687511
rect 674944 686678 674972 688735
rect 675128 688514 675156 688894
rect 675128 688486 675340 688514
rect 675312 688378 675340 688486
rect 675404 688378 675432 688500
rect 675312 688350 675432 688378
rect 675114 687848 675170 687857
rect 675170 687806 675418 687834
rect 675114 687783 675170 687792
rect 674944 686650 675248 686678
rect 675220 686610 675248 686650
rect 675404 686610 675432 686664
rect 675220 686582 675432 686610
rect 675482 686488 675538 686497
rect 675482 686423 675538 686432
rect 674930 686216 674986 686225
rect 674930 686151 674986 686160
rect 674392 683086 674512 683114
rect 674576 683086 674696 683114
rect 674944 683114 674972 686151
rect 675496 685984 675524 686423
rect 675482 685672 675538 685681
rect 675482 685607 675538 685616
rect 675114 685400 675170 685409
rect 675496 685372 675524 685607
rect 675114 685335 675170 685344
rect 675128 684162 675156 685335
rect 675128 684134 675418 684162
rect 674944 683086 675340 683114
rect 674116 654106 674328 654134
rect 674010 648408 674066 648417
rect 674010 648343 674066 648352
rect 674024 647986 674052 648343
rect 673472 620986 673776 621014
rect 673840 647958 674052 647986
rect 673472 619562 673500 620986
rect 673642 620664 673698 620673
rect 673642 620599 673698 620608
rect 673656 619682 673684 620599
rect 673644 619676 673696 619682
rect 673644 619618 673696 619624
rect 673472 619534 673592 619562
rect 673564 617409 673592 619534
rect 673550 617400 673606 617409
rect 673550 617335 673606 617344
rect 673840 601694 673868 647958
rect 674010 647320 674066 647329
rect 674010 647255 674012 647264
rect 674064 647255 674066 647264
rect 674012 647226 674064 647232
rect 674102 644328 674158 644337
rect 674102 644263 674158 644272
rect 674116 643226 674144 644263
rect 674116 643198 674236 643226
rect 674012 643136 674064 643142
rect 674010 643104 674012 643113
rect 674064 643104 674066 643113
rect 674010 643039 674066 643048
rect 674208 640334 674236 643198
rect 674116 640306 674236 640334
rect 674116 630674 674144 640306
rect 674300 636886 674328 654106
rect 674392 649994 674420 683086
rect 674576 682446 674604 683086
rect 674564 682440 674616 682446
rect 674564 682382 674616 682388
rect 674746 671664 674802 671673
rect 674746 671599 674802 671608
rect 674760 663513 674788 671599
rect 675312 666913 675340 683086
rect 683212 682440 683264 682446
rect 683212 682382 683264 682388
rect 681002 679008 681058 679017
rect 681002 678943 681058 678952
rect 675298 666904 675354 666913
rect 675298 666839 675354 666848
rect 681016 665825 681044 678943
rect 681002 665816 681058 665825
rect 681002 665751 681058 665760
rect 674930 664048 674986 664057
rect 674930 663983 674932 663992
rect 674984 663983 674986 663992
rect 676220 664012 676272 664018
rect 674932 663954 674984 663960
rect 676220 663954 676272 663960
rect 676232 663785 676260 663954
rect 676218 663776 676274 663785
rect 676218 663711 676274 663720
rect 674746 663504 674802 663513
rect 674746 663439 674802 663448
rect 683224 662969 683252 682382
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683210 662960 683266 662969
rect 683210 662895 683266 662904
rect 674562 660240 674618 660249
rect 674562 660175 674618 660184
rect 674576 659870 674604 660175
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 683132 659870 683160 660039
rect 674564 659864 674616 659870
rect 674564 659806 674616 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 674852 653126 675340 653154
rect 674392 649966 674512 649994
rect 674484 647234 674512 649966
rect 674852 647234 674880 653126
rect 675312 653018 675340 653126
rect 675404 653018 675432 653140
rect 675312 652990 675432 653018
rect 675312 652582 675432 652610
rect 675312 652474 675340 652582
rect 675128 652446 675340 652474
rect 675404 652460 675432 652582
rect 675128 652225 675156 652446
rect 675114 652216 675170 652225
rect 675114 652151 675170 652160
rect 675128 651834 675418 651862
rect 675128 651409 675156 651834
rect 675114 651400 675170 651409
rect 675114 651335 675170 651344
rect 674392 647206 674512 647234
rect 674760 647206 674880 647234
rect 674944 649998 675340 650026
rect 674392 637574 674420 647206
rect 674760 644881 674788 647206
rect 674746 644872 674802 644881
rect 674746 644807 674802 644816
rect 674944 643618 674972 649998
rect 675312 649994 675340 649998
rect 675404 649994 675432 650012
rect 675312 649966 675432 649994
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675404 648417 675432 648788
rect 675390 648408 675446 648417
rect 675390 648343 675446 648352
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675114 647320 675170 647329
rect 675114 647255 675170 647264
rect 675128 645674 675156 647255
rect 675128 645646 675418 645674
rect 675128 645102 675418 645130
rect 674932 643612 674984 643618
rect 674932 643554 674984 643560
rect 675128 643550 675156 645102
rect 675312 644461 675418 644489
rect 675312 644337 675340 644461
rect 675298 644328 675354 644337
rect 675298 644263 675354 644272
rect 675312 643810 675418 643838
rect 675116 643544 675168 643550
rect 675116 643486 675168 643492
rect 674932 643476 674984 643482
rect 674932 643418 674984 643424
rect 674748 643340 674800 643346
rect 674748 643282 674800 643288
rect 674564 642796 674616 642802
rect 674564 642738 674616 642744
rect 674392 637546 674512 637574
rect 674288 636880 674340 636886
rect 674288 636822 674340 636828
rect 674116 630646 674328 630674
rect 674300 627910 674328 630646
rect 674288 627904 674340 627910
rect 674288 627846 674340 627852
rect 674010 626376 674066 626385
rect 674010 626311 674066 626320
rect 674024 625734 674052 626311
rect 674012 625728 674064 625734
rect 674012 625670 674064 625676
rect 674010 625560 674066 625569
rect 674010 625495 674066 625504
rect 674024 625190 674052 625495
rect 674012 625184 674064 625190
rect 674012 625126 674064 625132
rect 674010 624744 674066 624753
rect 674010 624679 674012 624688
rect 674064 624679 674066 624688
rect 674012 624650 674064 624656
rect 674012 624368 674064 624374
rect 674010 624336 674012 624345
rect 674064 624336 674066 624345
rect 674010 624271 674066 624280
rect 674010 623928 674066 623937
rect 674010 623863 674012 623872
rect 674064 623863 674066 623872
rect 674012 623834 674064 623840
rect 674012 623552 674064 623558
rect 674010 623520 674012 623529
rect 674064 623520 674066 623529
rect 674010 623455 674066 623464
rect 674010 623112 674066 623121
rect 674010 623047 674012 623056
rect 674064 623047 674066 623056
rect 674012 623018 674064 623024
rect 674010 622296 674066 622305
rect 674010 622231 674012 622240
rect 674064 622231 674066 622240
rect 674012 622202 674064 622208
rect 674012 621784 674064 621790
rect 674012 621726 674064 621732
rect 674024 621489 674052 621726
rect 674010 621480 674066 621489
rect 674010 621415 674066 621424
rect 674012 621104 674064 621110
rect 674010 621072 674012 621081
rect 674064 621072 674066 621081
rect 674010 621007 674066 621016
rect 674484 621014 674512 637546
rect 674208 620986 674512 621014
rect 674012 620288 674064 620294
rect 674012 620230 674064 620236
rect 674024 619857 674052 620230
rect 674010 619848 674066 619857
rect 674010 619783 674066 619792
rect 674012 619064 674064 619070
rect 674010 619032 674012 619041
rect 674064 619032 674066 619041
rect 674010 618967 674066 618976
rect 674208 618633 674236 620986
rect 674380 620900 674432 620906
rect 674380 620842 674432 620848
rect 674194 618624 674250 618633
rect 674194 618559 674250 618568
rect 674010 616992 674066 617001
rect 674010 616927 674012 616936
rect 674064 616927 674066 616936
rect 674012 616898 674064 616904
rect 674012 616616 674064 616622
rect 674010 616584 674012 616593
rect 674064 616584 674066 616593
rect 674010 616519 674066 616528
rect 674012 615528 674064 615534
rect 674010 615496 674012 615505
rect 674064 615496 674066 615505
rect 674010 615431 674066 615440
rect 674010 614952 674066 614961
rect 674010 614887 674012 614896
rect 674064 614887 674066 614896
rect 674012 614858 674064 614864
rect 674010 611416 674066 611425
rect 674010 611351 674012 611360
rect 674064 611351 674066 611360
rect 674012 611322 674064 611328
rect 673840 601666 674052 601694
rect 673826 600400 673882 600409
rect 673826 600335 673828 600344
rect 673880 600335 673882 600344
rect 673828 600306 673880 600312
rect 673642 599856 673698 599865
rect 673642 599791 673698 599800
rect 673656 582374 673684 599791
rect 673828 599480 673880 599486
rect 673826 599448 673828 599457
rect 673880 599448 673882 599457
rect 673826 599383 673882 599392
rect 673826 599176 673882 599185
rect 673826 599111 673882 599120
rect 673840 582374 673868 599111
rect 674024 591433 674052 601666
rect 674194 598632 674250 598641
rect 674194 598567 674250 598576
rect 674010 591424 674066 591433
rect 674010 591359 674066 591368
rect 673472 582346 673684 582374
rect 673748 582346 673868 582374
rect 674208 582374 674236 598567
rect 674392 591326 674420 620842
rect 674380 591320 674432 591326
rect 674380 591262 674432 591268
rect 674208 582346 674328 582374
rect 673472 567194 673500 582346
rect 673748 567194 673776 582346
rect 674010 581088 674066 581097
rect 674300 581074 674328 582346
rect 674576 581346 674604 642738
rect 674760 621014 674788 643282
rect 674944 642649 674972 643418
rect 675114 643104 675170 643113
rect 675114 643039 675170 643048
rect 674852 642621 674972 642649
rect 674852 637650 674880 642621
rect 675128 641458 675156 643039
rect 675312 642802 675340 643810
rect 675482 643512 675538 643521
rect 675482 643447 675538 643456
rect 675496 643280 675524 643447
rect 675300 642796 675352 642802
rect 675300 642738 675352 642744
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675404 640665 675432 640795
rect 675390 640656 675446 640665
rect 675390 640591 675446 640600
rect 675298 640384 675354 640393
rect 675128 640342 675298 640370
rect 674852 637622 674972 637650
rect 674944 631417 674972 637622
rect 674930 631408 674986 631417
rect 674930 631343 674986 631352
rect 675128 630674 675156 640342
rect 675298 640319 675354 640328
rect 675220 640138 675418 640166
rect 675220 637574 675248 640138
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675220 637546 675340 637574
rect 675036 630646 675156 630674
rect 675036 629785 675064 630646
rect 675022 629776 675078 629785
rect 675022 629711 675078 629720
rect 675312 629218 675340 637546
rect 683304 636880 683356 636886
rect 683304 636822 683356 636828
rect 683946 636848 684002 636857
rect 675220 629190 675340 629218
rect 674930 625968 674986 625977
rect 674930 625903 674986 625912
rect 674944 625734 674972 625903
rect 674932 625728 674984 625734
rect 674932 625670 674984 625676
rect 675220 621014 675248 629190
rect 675392 627904 675444 627910
rect 675392 627846 675444 627852
rect 674668 620986 674788 621014
rect 674944 620986 675248 621014
rect 674668 592034 674696 620986
rect 674944 611354 674972 620986
rect 675404 620906 675432 627846
rect 676496 625728 676548 625734
rect 676494 625696 676496 625705
rect 676548 625696 676550 625705
rect 676494 625631 676550 625640
rect 675392 620900 675444 620906
rect 675392 620842 675444 620848
rect 683316 617953 683344 636822
rect 683946 636783 684002 636792
rect 683960 622033 683988 636783
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683946 622024 684002 622033
rect 683946 621959 684002 621968
rect 683302 617944 683358 617953
rect 683302 617879 683358 617888
rect 675116 615528 675168 615534
rect 675114 615496 675116 615505
rect 683120 615528 683172 615534
rect 675168 615496 675170 615505
rect 675114 615431 675170 615440
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 683118 615431 683174 615440
rect 674852 611326 674972 611354
rect 675114 611416 675170 611425
rect 675114 611351 675170 611360
rect 674852 604761 674880 611326
rect 675128 608682 675156 611351
rect 675128 608654 675418 608682
rect 675114 608288 675170 608297
rect 675114 608223 675170 608232
rect 675128 608138 675156 608223
rect 675128 608110 675418 608138
rect 675128 607465 675418 607493
rect 675128 607345 675156 607465
rect 675114 607336 675170 607345
rect 675114 607271 675170 607280
rect 675036 606818 675418 606846
rect 674838 604752 674894 604761
rect 674838 604687 674894 604696
rect 674840 604580 674892 604586
rect 674840 604522 674892 604528
rect 674852 592034 674880 604522
rect 675036 603922 675064 606818
rect 675312 604982 675418 605010
rect 675312 604586 675340 604982
rect 675300 604580 675352 604586
rect 675300 604522 675352 604528
rect 675404 604217 675432 604452
rect 675390 604208 675446 604217
rect 675390 604143 675446 604152
rect 674944 603894 675064 603922
rect 675312 603894 675432 603922
rect 674944 598934 674972 603894
rect 675114 603800 675170 603809
rect 675312 603786 675340 603894
rect 675170 603758 675340 603786
rect 675404 603772 675432 603894
rect 675114 603735 675170 603744
rect 675128 603146 675418 603174
rect 675128 602993 675156 603146
rect 675114 602984 675170 602993
rect 675114 602919 675170 602928
rect 675312 600766 675432 600794
rect 675114 600672 675170 600681
rect 675312 600658 675340 600766
rect 675170 600630 675340 600658
rect 675404 600644 675432 600766
rect 675114 600607 675170 600616
rect 675298 600400 675354 600409
rect 675298 600335 675354 600344
rect 675114 599448 675170 599457
rect 675114 599383 675170 599392
rect 674944 598906 675064 598934
rect 675036 595270 675064 598906
rect 675128 596442 675156 599383
rect 675312 598278 675340 600335
rect 675496 599865 675524 600100
rect 675482 599856 675538 599865
rect 675482 599791 675538 599800
rect 675496 599185 675524 599488
rect 675482 599176 675538 599185
rect 675482 599111 675538 599120
rect 675496 598641 675524 598808
rect 675482 598632 675538 598641
rect 675482 598567 675538 598576
rect 675312 598250 675418 598278
rect 675404 597417 675432 597652
rect 675390 597408 675446 597417
rect 675390 597343 675446 597352
rect 675128 596414 675418 596442
rect 675404 595513 675432 595816
rect 675390 595504 675446 595513
rect 675390 595439 675446 595448
rect 675024 595264 675076 595270
rect 675024 595206 675076 595212
rect 675036 595122 675418 595150
rect 674668 592006 674788 592034
rect 674852 592006 674972 592034
rect 674576 581318 674696 581346
rect 674300 581046 674512 581074
rect 674010 581023 674012 581032
rect 674064 581023 674066 581032
rect 674012 580994 674064 581000
rect 674012 580440 674064 580446
rect 674064 580388 674328 580394
rect 674012 580382 674328 580388
rect 674024 580366 674328 580382
rect 674300 580310 674328 580366
rect 674012 580304 674064 580310
rect 674010 580272 674012 580281
rect 674288 580304 674340 580310
rect 674064 580272 674066 580281
rect 674288 580246 674340 580252
rect 674010 580207 674066 580216
rect 674288 580168 674340 580174
rect 674024 580116 674288 580122
rect 674024 580110 674340 580116
rect 674024 580094 674328 580110
rect 674024 579698 674052 580094
rect 674012 579692 674064 579698
rect 674012 579634 674064 579640
rect 674024 579290 674328 579306
rect 674012 579284 674340 579290
rect 674064 579278 674288 579284
rect 674012 579226 674064 579232
rect 674288 579226 674340 579232
rect 674012 579080 674064 579086
rect 674010 579048 674012 579057
rect 674064 579048 674066 579057
rect 674010 578983 674066 578992
rect 674288 578468 674340 578474
rect 674288 578410 674340 578416
rect 674300 578354 674328 578410
rect 674024 578338 674328 578354
rect 674012 578332 674328 578338
rect 674064 578326 674328 578332
rect 674012 578274 674064 578280
rect 674012 578128 674064 578134
rect 674288 578128 674340 578134
rect 674064 578076 674288 578082
rect 674012 578070 674340 578076
rect 674024 578054 674328 578070
rect 674012 577856 674064 577862
rect 674064 577804 674328 577810
rect 674012 577798 674328 577804
rect 674024 577794 674328 577798
rect 674024 577788 674340 577794
rect 674024 577782 674288 577788
rect 674288 577730 674340 577736
rect 674288 577652 674340 577658
rect 674484 577640 674512 581046
rect 674668 579614 674696 581318
rect 674576 579586 674696 579614
rect 674576 577776 674604 579586
rect 674760 579442 674788 592006
rect 674944 584633 674972 592006
rect 675036 589274 675064 595122
rect 675208 595060 675260 595066
rect 675208 595002 675260 595008
rect 675220 589274 675248 595002
rect 675404 593609 675432 593980
rect 675390 593600 675446 593609
rect 675390 593535 675446 593544
rect 676034 592920 676090 592929
rect 676034 592855 676090 592864
rect 675484 591456 675536 591462
rect 675482 591424 675484 591433
rect 675536 591424 675538 591433
rect 675482 591359 675538 591368
rect 675036 589246 675156 589274
rect 675220 589246 675340 589274
rect 674930 584624 674986 584633
rect 674930 584559 674986 584568
rect 674760 579414 674880 579442
rect 674852 577930 674880 579414
rect 674840 577924 674892 577930
rect 674840 577866 674892 577872
rect 674576 577748 674880 577776
rect 674484 577612 674696 577640
rect 674288 577594 674340 577600
rect 674300 577538 674328 577594
rect 674024 577522 674328 577538
rect 674012 577516 674328 577522
rect 674064 577510 674328 577516
rect 674012 577458 674064 577464
rect 674010 577008 674066 577017
rect 674010 576943 674012 576952
rect 674064 576943 674066 576952
rect 674012 576914 674064 576920
rect 674288 576020 674340 576026
rect 674288 575962 674340 575968
rect 674300 575906 674328 575962
rect 674024 575878 674328 575906
rect 674024 575550 674052 575878
rect 674012 575544 674064 575550
rect 674012 575486 674064 575492
rect 674012 574592 674064 574598
rect 674010 574560 674012 574569
rect 674064 574560 674066 574569
rect 674010 574495 674066 574504
rect 674012 574320 674064 574326
rect 674010 574288 674012 574297
rect 674064 574288 674066 574297
rect 674010 574223 674066 574232
rect 674288 574184 674340 574190
rect 674024 574132 674288 574138
rect 674024 574126 674340 574132
rect 674024 574122 674328 574126
rect 674012 574116 674328 574122
rect 674064 574110 674328 574116
rect 674012 574058 674064 574064
rect 674012 573096 674064 573102
rect 674010 573064 674012 573073
rect 674064 573064 674066 573073
rect 674010 572999 674066 573008
rect 674288 572960 674340 572966
rect 674024 572908 674288 572914
rect 674024 572902 674340 572908
rect 674024 572886 674328 572902
rect 674024 572762 674052 572886
rect 674012 572756 674064 572762
rect 674012 572698 674064 572704
rect 674288 571940 674340 571946
rect 674288 571882 674340 571888
rect 674300 571826 674328 571882
rect 674024 571798 674328 571826
rect 674024 571470 674052 571798
rect 674012 571464 674064 571470
rect 674012 571406 674064 571412
rect 674288 570104 674340 570110
rect 674024 570052 674288 570058
rect 674024 570046 674340 570052
rect 674024 570030 674328 570046
rect 674024 569974 674052 570030
rect 674012 569968 674064 569974
rect 674012 569910 674064 569916
rect 674288 569288 674340 569294
rect 674288 569230 674340 569236
rect 674300 569106 674328 569230
rect 674024 569078 674328 569106
rect 674024 568614 674052 569078
rect 674012 568608 674064 568614
rect 674012 568550 674064 568556
rect 674668 567194 674696 577612
rect 674852 571305 674880 577748
rect 674838 571296 674894 571305
rect 674838 571231 674894 571240
rect 673472 567166 673684 567194
rect 673748 567166 674052 567194
rect 673656 528554 673684 567166
rect 673828 565888 673880 565894
rect 673826 565856 673828 565865
rect 673880 565856 673882 565865
rect 673826 565791 673882 565800
rect 673826 554840 673882 554849
rect 673826 554775 673828 554784
rect 673880 554775 673882 554784
rect 673828 554746 673880 554752
rect 673826 553752 673882 553761
rect 673826 553687 673828 553696
rect 673880 553687 673882 553696
rect 673828 553658 673880 553664
rect 674024 547913 674052 567166
rect 674116 567166 674696 567194
rect 674116 548162 674144 567166
rect 675128 563054 675156 589246
rect 675312 586265 675340 589246
rect 675298 586256 675354 586265
rect 675298 586191 675354 586200
rect 675484 577924 675536 577930
rect 675484 577866 675536 577872
rect 675496 571713 675524 577866
rect 675852 577788 675904 577794
rect 675852 577730 675904 577736
rect 675864 577425 675892 577730
rect 675850 577416 675906 577425
rect 675850 577351 675906 577360
rect 676048 575521 676076 592855
rect 683212 591456 683264 591462
rect 683212 591398 683264 591404
rect 682382 590608 682438 590617
rect 682382 590543 682438 590552
rect 676218 580544 676274 580553
rect 676218 580479 676274 580488
rect 676232 580174 676260 580479
rect 676404 580304 676456 580310
rect 676404 580246 676456 580252
rect 676220 580168 676272 580174
rect 676416 580145 676444 580246
rect 676220 580110 676272 580116
rect 676402 580136 676458 580145
rect 676402 580071 676458 580080
rect 676218 579320 676274 579329
rect 676218 579255 676220 579264
rect 676272 579255 676274 579264
rect 676220 579226 676272 579232
rect 676218 578504 676274 578513
rect 676218 578439 676220 578448
rect 676272 578439 676274 578448
rect 676220 578410 676272 578416
rect 676220 578128 676272 578134
rect 676218 578096 676220 578105
rect 676272 578096 676274 578105
rect 676218 578031 676274 578040
rect 676218 577688 676274 577697
rect 676218 577623 676220 577632
rect 676272 577623 676274 577632
rect 676220 577594 676272 577600
rect 682396 576065 682424 590543
rect 676218 576056 676274 576065
rect 676218 575991 676220 576000
rect 676272 575991 676274 576000
rect 682382 576056 682438 576065
rect 682382 575991 682438 576000
rect 676220 575962 676272 575968
rect 676034 575512 676090 575521
rect 676034 575447 676090 575456
rect 676218 574832 676274 574841
rect 676218 574767 676274 574776
rect 676232 574190 676260 574767
rect 676220 574184 676272 574190
rect 676220 574126 676272 574132
rect 683224 573617 683252 591398
rect 683396 591320 683448 591326
rect 683396 591262 683448 591268
rect 676218 573608 676274 573617
rect 676218 573543 676274 573552
rect 683210 573608 683266 573617
rect 683210 573543 683266 573552
rect 676232 572966 676260 573543
rect 676220 572960 676272 572966
rect 676220 572902 676272 572908
rect 683408 572801 683436 591262
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683394 572792 683450 572801
rect 683394 572727 683450 572736
rect 676218 571976 676274 571985
rect 676218 571911 676220 571920
rect 676272 571911 676274 571920
rect 676220 571882 676272 571888
rect 675482 571704 675538 571713
rect 675482 571639 675538 571648
rect 676218 570752 676274 570761
rect 676218 570687 676274 570696
rect 676232 570110 676260 570687
rect 676220 570104 676272 570110
rect 676220 570046 676272 570052
rect 676218 569528 676274 569537
rect 676218 569463 676274 569472
rect 676232 569294 676260 569463
rect 676220 569288 676272 569294
rect 676220 569230 676272 569236
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675404 563448 675432 565791
rect 675390 563136 675446 563145
rect 675390 563071 675446 563080
rect 674852 563026 675156 563054
rect 674472 559360 674524 559366
rect 674472 559302 674524 559308
rect 674288 558272 674340 558278
rect 674288 558214 674340 558220
rect 674300 554933 674328 558214
rect 674484 554933 674512 559302
rect 674656 557592 674708 557598
rect 674656 557534 674708 557540
rect 674208 554905 674328 554933
rect 674392 554905 674512 554933
rect 674208 550634 674236 554905
rect 674392 554826 674420 554905
rect 674300 554798 674420 554826
rect 674300 553394 674328 554798
rect 674472 554736 674524 554742
rect 674472 554678 674524 554684
rect 674300 553366 674420 553394
rect 674208 550606 674328 550634
rect 674116 548134 674236 548162
rect 674010 547904 674066 547913
rect 674010 547839 674066 547848
rect 674208 547754 674236 548134
rect 674024 547726 674236 547754
rect 674024 547641 674052 547726
rect 674010 547632 674066 547641
rect 674010 547567 674066 547576
rect 674300 540974 674328 550606
rect 673840 540946 674328 540974
rect 673840 534074 673868 540946
rect 674194 536072 674250 536081
rect 674194 536007 674250 536016
rect 674012 535696 674064 535702
rect 674010 535664 674012 535673
rect 674064 535664 674066 535673
rect 674010 535599 674066 535608
rect 674208 535514 674236 536007
rect 674024 535498 674236 535514
rect 674012 535492 674236 535498
rect 674064 535486 674236 535492
rect 674012 535434 674064 535440
rect 674010 535256 674066 535265
rect 674010 535191 674066 535200
rect 674024 534274 674052 535191
rect 674194 534440 674250 534449
rect 674194 534375 674250 534384
rect 674012 534268 674064 534274
rect 674012 534210 674064 534216
rect 674208 534154 674236 534375
rect 674024 534138 674236 534154
rect 674012 534132 674236 534138
rect 674064 534126 674236 534132
rect 674012 534074 674064 534080
rect 673472 528526 673684 528554
rect 673748 534046 673868 534074
rect 673472 527082 673500 528526
rect 673748 528374 673776 534046
rect 674010 533216 674066 533225
rect 674010 533151 674066 533160
rect 674024 532982 674052 533151
rect 674012 532976 674064 532982
rect 674012 532918 674064 532924
rect 674010 532808 674066 532817
rect 674010 532743 674012 532752
rect 674064 532743 674066 532752
rect 674012 532714 674064 532720
rect 674010 532400 674066 532409
rect 674010 532335 674066 532344
rect 674024 531758 674052 532335
rect 674194 531992 674250 532001
rect 674194 531927 674250 531936
rect 674012 531752 674064 531758
rect 674012 531694 674064 531700
rect 674208 531638 674236 531927
rect 674024 531610 674236 531638
rect 674024 531350 674052 531610
rect 674012 531344 674064 531350
rect 674012 531286 674064 531292
rect 674010 531176 674066 531185
rect 674010 531111 674066 531120
rect 674024 530534 674052 531111
rect 674194 530768 674250 530777
rect 674194 530703 674250 530712
rect 674012 530528 674064 530534
rect 674012 530470 674064 530476
rect 674012 530256 674064 530262
rect 674012 530198 674064 530204
rect 674024 530097 674052 530198
rect 674010 530088 674066 530097
rect 674010 530023 674066 530032
rect 674208 529938 674236 530703
rect 674024 529922 674236 529938
rect 674012 529916 674236 529922
rect 674064 529910 674236 529916
rect 674012 529858 674064 529864
rect 674194 529544 674250 529553
rect 674194 529479 674250 529488
rect 674010 529136 674066 529145
rect 674010 529071 674066 529080
rect 674024 528766 674052 529071
rect 674012 528760 674064 528766
rect 674012 528702 674064 528708
rect 674012 528624 674064 528630
rect 674208 528578 674236 529479
rect 674064 528572 674236 528578
rect 674012 528566 674236 528572
rect 674024 528550 674236 528566
rect 673748 528346 673868 528374
rect 673642 528184 673698 528193
rect 673642 528119 673698 528128
rect 673656 527202 673684 528119
rect 673644 527196 673696 527202
rect 673644 527138 673696 527144
rect 673472 527054 673592 527082
rect 673564 526833 673592 527054
rect 673550 526824 673606 526833
rect 673550 526759 673606 526768
rect 673840 499574 673868 528346
rect 674010 527912 674066 527921
rect 674010 527847 674066 527856
rect 674024 527406 674052 527847
rect 674012 527400 674064 527406
rect 674012 527342 674064 527348
rect 674392 509234 674420 553366
rect 673656 499546 673868 499574
rect 674300 509206 674420 509234
rect 673656 490634 673684 499546
rect 674300 494766 674328 509206
rect 674288 494760 674340 494766
rect 674288 494702 674340 494708
rect 673826 492144 673882 492153
rect 673826 492079 673882 492088
rect 673840 491366 673868 492079
rect 674012 491904 674064 491910
rect 674064 491852 674328 491858
rect 674012 491846 674328 491852
rect 674024 491842 674328 491846
rect 674024 491836 674340 491842
rect 674024 491830 674288 491836
rect 674288 491778 674340 491784
rect 674288 491700 674340 491706
rect 674288 491642 674340 491648
rect 674300 491586 674328 491642
rect 674024 491558 674328 491586
rect 674024 491502 674052 491558
rect 674012 491496 674064 491502
rect 674012 491438 674064 491444
rect 673828 491360 673880 491366
rect 673828 491302 673880 491308
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 673656 490606 674144 490634
rect 673920 489320 673972 489326
rect 673918 489288 673920 489297
rect 673972 489288 673974 489297
rect 673918 489223 673974 489232
rect 673920 488504 673972 488510
rect 673918 488472 673920 488481
rect 673972 488472 673974 488481
rect 673918 488407 673974 488416
rect 673918 486024 673974 486033
rect 673918 485959 673974 485968
rect 673932 485858 673960 485959
rect 673920 485852 673972 485858
rect 673920 485794 673972 485800
rect 674116 485774 674144 490606
rect 674116 485746 674236 485774
rect 674012 485648 674064 485654
rect 674010 485616 674012 485625
rect 674064 485616 674066 485625
rect 674010 485551 674066 485560
rect 674010 485208 674066 485217
rect 674010 485143 674066 485152
rect 674024 484430 674052 485143
rect 674012 484424 674064 484430
rect 674208 484401 674236 485746
rect 674012 484366 674064 484372
rect 674194 484392 674250 484401
rect 674194 484327 674250 484336
rect 674012 484016 674064 484022
rect 674010 483984 674012 483993
rect 674064 483984 674066 483993
rect 674010 483919 674066 483928
rect 674484 482769 674512 554678
rect 674668 483177 674696 557534
rect 674852 546514 674880 563026
rect 675404 562904 675432 563071
rect 675128 562278 675418 562306
rect 675128 561921 675156 562278
rect 675114 561912 675170 561921
rect 675114 561847 675170 561856
rect 675312 561734 675432 561762
rect 675312 561626 675340 561734
rect 674944 561598 675340 561626
rect 675404 561612 675432 561734
rect 674944 550634 674972 561598
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 675128 559762 675340 559790
rect 675404 559776 675432 559830
rect 675128 559366 675156 559762
rect 675116 559360 675168 559366
rect 675116 559302 675168 559308
rect 675128 559218 675418 559246
rect 675128 559065 675156 559218
rect 675114 559056 675170 559065
rect 675114 558991 675170 559000
rect 675404 558278 675432 558620
rect 675392 558272 675444 558278
rect 675392 558214 675444 558220
rect 675128 557926 675418 557954
rect 675128 557598 675156 557926
rect 675116 557592 675168 557598
rect 675116 557534 675168 557540
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675128 554905 675418 554933
rect 675128 554742 675156 554905
rect 675298 554840 675354 554849
rect 675298 554775 675354 554784
rect 675116 554736 675168 554742
rect 675116 554678 675168 554684
rect 675114 553752 675170 553761
rect 675114 553687 675170 553696
rect 675128 551253 675156 553687
rect 675312 553602 675340 554775
rect 675772 554033 675800 554268
rect 675758 554024 675814 554033
rect 675758 553959 675814 553968
rect 675220 553574 675340 553602
rect 675220 553093 675248 553574
rect 675404 553353 675432 553656
rect 675390 553344 675446 553353
rect 675390 553279 675446 553288
rect 675220 553065 675418 553093
rect 675312 552418 675418 552446
rect 675312 552129 675340 552418
rect 675298 552120 675354 552129
rect 675298 552055 675354 552064
rect 675128 551225 675418 551253
rect 674944 550606 675064 550634
rect 675036 550050 675064 550606
rect 675772 550361 675800 550596
rect 675758 550352 675814 550361
rect 675758 550287 675814 550296
rect 675024 550044 675076 550050
rect 675024 549986 675076 549992
rect 675128 549937 675418 549965
rect 675128 546922 675156 549937
rect 675300 549840 675352 549846
rect 675300 549782 675352 549788
rect 675312 547074 675340 549782
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675482 547904 675538 547913
rect 675482 547839 675538 547848
rect 675496 547194 675524 547839
rect 675666 547632 675722 547641
rect 675666 547567 675722 547576
rect 678242 547632 678298 547641
rect 678242 547567 678298 547576
rect 675484 547188 675536 547194
rect 675484 547130 675536 547136
rect 675312 547046 675432 547074
rect 675116 546916 675168 546922
rect 675116 546858 675168 546864
rect 675116 546712 675168 546718
rect 675116 546654 675168 546660
rect 674840 546508 674892 546514
rect 674840 546450 674892 546456
rect 675128 545578 675156 546654
rect 675036 545550 675156 545578
rect 675036 528554 675064 545550
rect 675404 541090 675432 547046
rect 675680 545766 675708 547567
rect 675668 545760 675720 545766
rect 675668 545702 675720 545708
rect 675574 545592 675630 545601
rect 675574 545527 675630 545536
rect 674944 528526 675064 528554
rect 675220 541062 675432 541090
rect 674654 483168 674710 483177
rect 674654 483103 674710 483112
rect 674470 482760 674526 482769
rect 674470 482695 674526 482704
rect 674944 480486 674972 528526
rect 675220 488510 675248 541062
rect 675588 540974 675616 545527
rect 675312 540946 675616 540974
rect 675312 518894 675340 540946
rect 678256 531865 678284 547567
rect 684316 547188 684368 547194
rect 684316 547130 684368 547136
rect 683486 547088 683542 547097
rect 683486 547023 683542 547032
rect 682382 546816 682438 546825
rect 682382 546751 682438 546760
rect 681004 546508 681056 546514
rect 681004 546450 681056 546456
rect 678242 531856 678298 531865
rect 678242 531791 678298 531800
rect 681016 525774 681044 546450
rect 682396 530641 682424 546751
rect 683304 545760 683356 545766
rect 683304 545702 683356 545708
rect 682382 530632 682438 530641
rect 682382 530567 682438 530576
rect 683316 526561 683344 545702
rect 683500 527377 683528 547023
rect 684328 527785 684356 547130
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 684314 527776 684370 527785
rect 684314 527711 684370 527720
rect 683486 527368 683542 527377
rect 683486 527303 683542 527312
rect 683302 526552 683358 526561
rect 683302 526487 683358 526496
rect 681004 525768 681056 525774
rect 681004 525710 681056 525716
rect 683120 525768 683172 525774
rect 683120 525710 683172 525716
rect 683302 525736 683358 525745
rect 683132 525337 683160 525710
rect 683302 525671 683358 525680
rect 683118 525328 683174 525337
rect 683118 525263 683174 525272
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 676864 518968 676916 518974
rect 676864 518910 676916 518916
rect 675312 518866 675708 518894
rect 675484 518696 675536 518702
rect 675484 518638 675536 518644
rect 675208 488504 675260 488510
rect 675208 488446 675260 488452
rect 674932 480480 674984 480486
rect 674932 480422 674984 480428
rect 675300 475244 675352 475250
rect 675300 475186 675352 475192
rect 673368 456000 673420 456006
rect 673368 455942 673420 455948
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673388 455194 673440 455200
rect 674288 455048 674340 455054
rect 673090 455016 673146 455025
rect 673090 454951 673146 454960
rect 674286 455016 674288 455025
rect 674340 455016 674342 455025
rect 674286 454951 674342 454960
rect 673104 454866 673132 454951
rect 673058 454850 673132 454866
rect 673046 454844 673132 454850
rect 673098 454838 673132 454844
rect 673046 454786 673098 454792
rect 674288 454776 674340 454782
rect 672906 454744 672962 454753
rect 672906 454679 672908 454688
rect 672960 454679 672962 454688
rect 674286 454744 674288 454753
rect 674340 454744 674342 454753
rect 674286 454679 674342 454688
rect 672908 454650 672960 454656
rect 674288 454504 674340 454510
rect 672814 454472 672870 454481
rect 672814 454407 672816 454416
rect 672868 454407 672870 454416
rect 674286 454472 674288 454481
rect 674340 454472 674342 454481
rect 674286 454407 674342 454416
rect 672816 454378 672868 454384
rect 675312 453937 675340 475186
rect 675496 455054 675524 518638
rect 675680 503878 675708 518866
rect 675668 503872 675720 503878
rect 675668 503814 675720 503820
rect 675852 491836 675904 491842
rect 675852 491778 675904 491784
rect 675864 491337 675892 491778
rect 676034 491736 676090 491745
rect 676034 491671 676036 491680
rect 676088 491671 676090 491680
rect 676036 491642 676088 491648
rect 675850 491328 675906 491337
rect 675850 491263 675906 491272
rect 675850 490512 675906 490521
rect 675850 490447 675906 490456
rect 675864 485774 675892 490447
rect 676036 488504 676088 488510
rect 676036 488446 676088 488452
rect 676048 487665 676076 488446
rect 676034 487656 676090 487665
rect 676034 487591 676090 487600
rect 675864 485746 675984 485774
rect 675666 480720 675722 480729
rect 675666 480655 675722 480664
rect 675484 455048 675536 455054
rect 675484 454990 675536 454996
rect 675680 454510 675708 480655
rect 675668 454504 675720 454510
rect 675668 454446 675720 454452
rect 675298 453928 675354 453937
rect 675298 453863 675354 453872
rect 675956 447817 675984 485746
rect 676876 454782 676904 518910
rect 677888 518838 677916 524447
rect 683316 518974 683344 525671
rect 683304 518968 683356 518974
rect 683304 518910 683356 518916
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 678244 503872 678296 503878
rect 678244 503814 678296 503820
rect 678256 486849 678284 503814
rect 683578 503704 683634 503713
rect 683578 503639 683634 503648
rect 683212 494760 683264 494766
rect 683212 494702 683264 494708
rect 678242 486840 678298 486849
rect 678242 486775 678298 486784
rect 683224 486441 683252 494702
rect 683592 487257 683620 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 487248 683634 487257
rect 683578 487183 683634 487192
rect 683210 486432 683266 486441
rect 683210 486367 683266 486376
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 680372 475250 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480486 683160 481063
rect 683120 480480 683172 480486
rect 683120 480422 683172 480428
rect 680360 475244 680412 475250
rect 680360 475186 680412 475192
rect 676864 454776 676916 454782
rect 676864 454718 676916 454724
rect 675942 447808 675998 447817
rect 675942 447743 675998 447752
rect 676034 410544 676090 410553
rect 676034 410479 676090 410488
rect 674564 403300 674616 403306
rect 674564 403242 674616 403248
rect 673182 402112 673238 402121
rect 673182 402047 673238 402056
rect 672630 401704 672686 401713
rect 672630 401639 672686 401648
rect 672906 401296 672962 401305
rect 672906 401231 672962 401240
rect 671986 397216 672042 397225
rect 671986 397151 672042 397160
rect 669226 393816 669282 393825
rect 669226 393751 669282 393760
rect 657544 373992 657596 373998
rect 657544 373934 657596 373940
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 654782 358592 654838 358601
rect 654782 358527 654838 358536
rect 63406 357368 63462 357377
rect 63406 357303 63462 357312
rect 652022 356688 652078 356697
rect 652022 356623 652078 356632
rect 62946 354512 63002 354521
rect 62946 354447 63002 354456
rect 51722 353288 51778 353297
rect 51722 353223 51778 353232
rect 46938 353016 46994 353025
rect 46938 352951 46994 352960
rect 46018 343904 46074 343913
rect 46018 343839 46074 343848
rect 63132 342236 63184 342242
rect 63132 342178 63184 342184
rect 62946 341728 63002 341737
rect 62946 341663 63002 341672
rect 62762 341456 62818 341465
rect 62762 341391 62818 341400
rect 45650 340776 45706 340785
rect 45650 340711 45706 340720
rect 39670 340232 39726 340241
rect 39670 340167 39726 340176
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35544 339658 35572 339759
rect 35532 339652 35584 339658
rect 35532 339594 35584 339600
rect 35820 339522 35848 339759
rect 37096 339652 37148 339658
rect 37096 339594 37148 339600
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37108 336569 37136 339594
rect 38844 339516 38896 339522
rect 38844 339458 38896 339464
rect 37094 336560 37150 336569
rect 37094 336495 37150 336504
rect 38856 335753 38884 339458
rect 46938 339280 46994 339289
rect 46938 339215 46994 339224
rect 45558 338872 45614 338881
rect 45558 338807 45614 338816
rect 45374 337920 45430 337929
rect 45374 337855 45430 337864
rect 45388 337770 45416 337855
rect 45388 337742 45508 337770
rect 35806 335744 35862 335753
rect 35806 335679 35862 335688
rect 38842 335744 38898 335753
rect 38842 335679 38898 335688
rect 35820 335374 35848 335679
rect 35808 335368 35860 335374
rect 35808 335310 35860 335316
rect 39856 335368 39908 335374
rect 39856 335310 39908 335316
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35820 334150 35848 334455
rect 35808 334144 35860 334150
rect 35808 334086 35860 334092
rect 39868 332489 39896 335310
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 44362 334656 44418 334665
rect 44362 334591 44418 334600
rect 40316 334144 40368 334150
rect 40316 334086 40368 334092
rect 40328 332897 40356 334086
rect 40314 332888 40370 332897
rect 40314 332823 40370 332832
rect 42890 332888 42946 332897
rect 42890 332823 42946 332832
rect 39854 332480 39910 332489
rect 39854 332415 39910 332424
rect 42430 327040 42486 327049
rect 42430 326975 42486 326984
rect 42444 326278 42472 326975
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42656 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42182 321898 42472 321926
rect 42076 321201 42104 321368
rect 42062 321192 42118 321201
rect 42062 321127 42118 321136
rect 42168 320521 42196 320725
rect 42154 320512 42210 320521
rect 42154 320447 42210 320456
rect 42076 319977 42104 320076
rect 41878 319968 41934 319977
rect 41878 319903 41934 319912
rect 42062 319968 42118 319977
rect 42062 319903 42118 319912
rect 41892 319532 41920 319903
rect 42444 319433 42472 321898
rect 42628 320793 42656 323734
rect 42904 321201 42932 332823
rect 43074 332480 43130 332489
rect 43074 332415 43130 332424
rect 42890 321192 42946 321201
rect 42890 321127 42946 321136
rect 42614 320784 42670 320793
rect 42614 320719 42670 320728
rect 43088 320521 43116 332415
rect 43074 320512 43130 320521
rect 43074 320447 43130 320456
rect 44192 319977 44220 334591
rect 44376 322833 44404 334591
rect 45282 327040 45338 327049
rect 45480 327026 45508 337742
rect 45338 326998 45508 327026
rect 45282 326975 45338 326984
rect 44362 322824 44418 322833
rect 44362 322759 44418 322768
rect 44178 319968 44234 319977
rect 44178 319903 44234 319912
rect 42430 319424 42486 319433
rect 42430 319359 42486 319368
rect 42246 319016 42302 319025
rect 42246 318951 42302 318960
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42260 316418 42288 318951
rect 42182 316390 42288 316418
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 45572 315489 45600 338807
rect 42154 315480 42210 315489
rect 42154 315415 42210 315424
rect 45558 315480 45614 315489
rect 45558 315415 45614 315424
rect 42168 315180 42196 315415
rect 42062 313712 42118 313721
rect 42062 313647 42118 313656
rect 42076 313344 42104 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42168 312174 42288 312202
rect 42168 312052 42196 312174
rect 42260 312066 42288 312174
rect 42260 312038 42472 312066
rect 42076 309097 42104 311508
rect 42444 310457 42472 312038
rect 46952 310457 46980 339215
rect 51722 334112 51778 334121
rect 51722 334047 51778 334056
rect 50342 333160 50398 333169
rect 50342 333095 50398 333104
rect 42430 310448 42486 310457
rect 42430 310383 42486 310392
rect 46938 310448 46994 310457
rect 46938 310383 46994 310392
rect 42062 309088 42118 309097
rect 42062 309023 42118 309032
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 35622 300928 35678 300937
rect 35622 300863 35678 300872
rect 35636 298790 35664 300863
rect 46202 300520 46258 300529
rect 46202 300455 46258 300464
rect 44362 299704 44418 299713
rect 44362 299639 44418 299648
rect 35806 298888 35862 298897
rect 35806 298823 35862 298832
rect 35624 298784 35676 298790
rect 35624 298726 35676 298732
rect 35820 298314 35848 298823
rect 41604 298784 41656 298790
rect 41786 298752 41842 298761
rect 41656 298732 41786 298738
rect 41604 298726 41786 298732
rect 41616 298710 41786 298726
rect 41786 298687 41842 298696
rect 35808 298308 35860 298314
rect 35808 298250 35860 298256
rect 41604 298308 41656 298314
rect 41604 298250 41656 298256
rect 41616 296562 41644 298250
rect 44178 297256 44234 297265
rect 44178 297191 44234 297200
rect 41786 296576 41842 296585
rect 41616 296534 41786 296562
rect 41786 296511 41842 296520
rect 42798 296576 42854 296585
rect 42798 296511 42854 296520
rect 35438 296440 35494 296449
rect 35438 296375 35494 296384
rect 35452 295526 35480 296375
rect 35622 296032 35678 296041
rect 35622 295967 35678 295976
rect 35440 295520 35492 295526
rect 35440 295462 35492 295468
rect 35636 295390 35664 295967
rect 35808 295656 35860 295662
rect 35806 295624 35808 295633
rect 40684 295656 40736 295662
rect 35860 295624 35862 295633
rect 40684 295598 40736 295604
rect 35806 295559 35862 295568
rect 40040 295520 40092 295526
rect 40040 295462 40092 295468
rect 35624 295384 35676 295390
rect 35624 295326 35676 295332
rect 35806 295216 35862 295225
rect 35806 295151 35862 295160
rect 33782 294808 33838 294817
rect 33782 294743 33838 294752
rect 32402 294400 32458 294409
rect 32402 294335 32458 294344
rect 32416 284889 32444 294335
rect 33796 286346 33824 294743
rect 35820 294302 35848 295151
rect 35808 294296 35860 294302
rect 35808 294238 35860 294244
rect 35806 293176 35862 293185
rect 35806 293111 35862 293120
rect 35820 292942 35848 293111
rect 35808 292936 35860 292942
rect 35808 292878 35860 292884
rect 35806 292768 35862 292777
rect 35806 292703 35862 292712
rect 35820 292602 35848 292703
rect 35808 292596 35860 292602
rect 35808 292538 35860 292544
rect 39212 292596 39264 292602
rect 39212 292538 39264 292544
rect 35806 291136 35862 291145
rect 35806 291071 35862 291080
rect 35622 290320 35678 290329
rect 35622 290255 35678 290264
rect 35636 289134 35664 290255
rect 35820 289950 35848 291071
rect 35808 289944 35860 289950
rect 35808 289886 35860 289892
rect 35624 289128 35676 289134
rect 35624 289070 35676 289076
rect 39224 288969 39252 292538
rect 40052 291378 40080 295462
rect 40040 291372 40092 291378
rect 40040 291314 40092 291320
rect 39210 288960 39266 288969
rect 39210 288895 39266 288904
rect 33784 286340 33836 286346
rect 33784 286282 33836 286288
rect 32402 284880 32458 284889
rect 32402 284815 32458 284824
rect 40696 284345 40724 295598
rect 41604 295384 41656 295390
rect 41656 295361 41828 295372
rect 41656 295352 41842 295361
rect 41656 295344 41786 295352
rect 41604 295326 41656 295332
rect 41786 295287 41842 295296
rect 41696 294296 41748 294302
rect 41696 294238 41748 294244
rect 41328 292868 41380 292874
rect 41328 292810 41380 292816
rect 41340 291122 41368 292810
rect 41708 292574 41736 294238
rect 41708 292546 42472 292574
rect 42246 291952 42302 291961
rect 42246 291887 42302 291896
rect 41696 291372 41748 291378
rect 41696 291314 41748 291320
rect 41708 291258 41736 291314
rect 41708 291242 42104 291258
rect 41708 291236 42116 291242
rect 41708 291230 42064 291236
rect 42064 291178 42116 291184
rect 41786 291136 41842 291145
rect 41340 291094 41786 291122
rect 41786 291071 41842 291080
rect 41696 289944 41748 289950
rect 41748 289892 42104 289898
rect 41696 289886 42104 289892
rect 41708 289882 42104 289886
rect 41708 289876 42116 289882
rect 41708 289870 42064 289876
rect 42064 289818 42116 289824
rect 42260 289241 42288 291887
rect 42246 289232 42302 289241
rect 42246 289167 42302 289176
rect 41696 289128 41748 289134
rect 41748 289076 42380 289082
rect 41696 289070 42380 289076
rect 41708 289054 42380 289070
rect 41696 286340 41748 286346
rect 41696 286282 41748 286288
rect 41708 286226 41736 286282
rect 41708 286198 42288 286226
rect 40682 284336 40738 284345
rect 40682 284271 40738 284280
rect 42260 283059 42288 286198
rect 42182 283031 42288 283059
rect 42352 281874 42380 289054
rect 42182 281846 42380 281874
rect 42248 281784 42300 281790
rect 42248 281726 42300 281732
rect 42260 281330 42288 281726
rect 42168 281302 42288 281330
rect 42168 281180 42196 281302
rect 42444 281058 42472 292546
rect 42616 291236 42668 291242
rect 42616 291178 42668 291184
rect 42628 281790 42656 291178
rect 42616 281784 42668 281790
rect 42616 281726 42668 281732
rect 42444 281030 42656 281058
rect 42182 280554 42472 280582
rect 42248 280152 42300 280158
rect 42248 280094 42300 280100
rect 42260 279426 42288 280094
rect 42168 279398 42288 279426
rect 42168 279344 42196 279398
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42182 278718 42288 278746
rect 41786 278488 41842 278497
rect 41786 278423 41842 278432
rect 41800 278188 41828 278423
rect 42062 277808 42118 277817
rect 42062 277743 42118 277752
rect 42076 277508 42104 277743
rect 42260 277394 42288 278718
rect 42430 278695 42486 278704
rect 42260 277366 42472 277394
rect 41786 277128 41842 277137
rect 41786 277063 41842 277072
rect 41800 276896 41828 277063
rect 42248 276820 42300 276826
rect 42248 276762 42300 276768
rect 42260 276570 42288 276762
rect 42444 276706 42472 277366
rect 42628 276826 42656 281030
rect 42616 276820 42668 276826
rect 42616 276762 42668 276768
rect 42444 276678 42656 276706
rect 42076 276542 42288 276570
rect 42076 276352 42104 276542
rect 42628 275913 42656 276678
rect 42614 275904 42670 275913
rect 42614 275839 42670 275848
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273170 42196 273224
rect 42338 273184 42394 273193
rect 42168 273142 42338 273170
rect 42338 273119 42394 273128
rect 42430 272912 42486 272921
rect 42430 272847 42486 272856
rect 42444 272558 42472 272847
rect 42182 272530 42472 272558
rect 41970 272368 42026 272377
rect 41970 272303 42026 272312
rect 41984 272000 42012 272303
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 41878 270056 41934 270065
rect 41878 269991 41934 270000
rect 41892 269521 41920 269991
rect 42156 269068 42208 269074
rect 42156 269010 42208 269016
rect 42168 268872 42196 269010
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 42168 266257 42196 268328
rect 42154 266248 42210 266257
rect 42154 266183 42210 266192
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42812 255921 42840 296511
rect 43166 295352 43222 295361
rect 43166 295287 43222 295296
rect 42982 291136 43038 291145
rect 42982 291071 43038 291080
rect 42996 280158 43024 291071
rect 42984 280152 43036 280158
rect 42984 280094 43036 280100
rect 43180 269074 43208 295287
rect 43352 289876 43404 289882
rect 43352 289818 43404 289824
rect 43364 282914 43392 289818
rect 43626 288960 43682 288969
rect 43626 288895 43682 288904
rect 43364 282886 43484 282914
rect 43168 269068 43220 269074
rect 43168 269010 43220 269016
rect 35806 255912 35862 255921
rect 35806 255847 35862 255856
rect 39762 255912 39818 255921
rect 39762 255847 39818 255856
rect 42798 255912 42854 255921
rect 42798 255847 42854 255856
rect 35820 255406 35848 255847
rect 39776 255406 39804 255847
rect 35808 255400 35860 255406
rect 35808 255342 35860 255348
rect 39764 255400 39816 255406
rect 39764 255342 39816 255348
rect 35808 254108 35860 254114
rect 35808 254050 35860 254056
rect 39212 254108 39264 254114
rect 39212 254050 39264 254056
rect 35820 253881 35848 254050
rect 35806 253872 35862 253881
rect 35806 253807 35862 253816
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35636 252618 35664 253399
rect 39224 253065 39252 254050
rect 43456 253934 43484 282886
rect 43640 277817 43668 288895
rect 43626 277808 43682 277817
rect 43626 277743 43682 277752
rect 44192 254946 44220 297191
rect 44376 256873 44404 299639
rect 44822 298072 44878 298081
rect 44822 298007 44878 298016
rect 44546 293584 44602 293593
rect 44546 293519 44602 293528
rect 44560 273193 44588 293519
rect 44546 273184 44602 273193
rect 44546 273119 44602 273128
rect 44362 256864 44418 256873
rect 44362 256799 44418 256808
rect 44638 256456 44694 256465
rect 44638 256391 44694 256400
rect 44100 254918 44220 254946
rect 44100 254561 44128 254918
rect 44270 254824 44326 254833
rect 44270 254759 44326 254768
rect 44086 254552 44142 254561
rect 44086 254487 44142 254496
rect 43272 253906 43484 253934
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 39210 253056 39266 253065
rect 39210 252991 39266 253000
rect 42798 253056 42854 253065
rect 42798 252991 42854 253000
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 41420 252748 41472 252754
rect 41420 252690 41472 252696
rect 35624 252612 35676 252618
rect 35624 252554 35676 252560
rect 40316 252612 40368 252618
rect 40316 252554 40368 252560
rect 40328 252249 40356 252554
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 40314 252240 40370 252249
rect 40314 252175 40370 252184
rect 35820 251394 35848 252175
rect 35808 251388 35860 251394
rect 35808 251330 35860 251336
rect 41432 251174 41460 252690
rect 41708 251394 41920 251410
rect 41696 251388 41920 251394
rect 41748 251382 41920 251388
rect 41696 251330 41748 251336
rect 41892 251174 41920 251382
rect 41432 251146 41736 251174
rect 41892 251146 42472 251174
rect 35806 250608 35862 250617
rect 35806 250543 35862 250552
rect 35820 249966 35848 250543
rect 35808 249960 35860 249966
rect 35808 249902 35860 249908
rect 39672 249960 39724 249966
rect 39672 249902 39724 249908
rect 39684 249393 39712 249902
rect 35806 249384 35862 249393
rect 35806 249319 35862 249328
rect 39670 249384 39726 249393
rect 39670 249319 39726 249328
rect 35820 248674 35848 249319
rect 35808 248668 35860 248674
rect 35808 248610 35860 248616
rect 41512 248668 41564 248674
rect 41512 248610 41564 248616
rect 41524 247761 41552 248610
rect 41708 248554 41736 251146
rect 41708 248526 42380 248554
rect 35622 247752 35678 247761
rect 35622 247687 35678 247696
rect 41510 247752 41566 247761
rect 41510 247687 41566 247696
rect 35636 247110 35664 247687
rect 35808 247240 35860 247246
rect 35808 247182 35860 247188
rect 41696 247240 41748 247246
rect 41696 247182 41748 247188
rect 35624 247104 35676 247110
rect 35624 247046 35676 247052
rect 35820 246945 35848 247182
rect 39856 247104 39908 247110
rect 39856 247046 39908 247052
rect 35806 246936 35862 246945
rect 35806 246871 35862 246880
rect 39868 245585 39896 247046
rect 39854 245576 39910 245585
rect 39854 245511 39910 245520
rect 41708 244274 41736 247182
rect 41708 244246 42288 244274
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 42260 238754 42288 244246
rect 42168 238726 42288 238754
rect 42168 238649 42196 238726
rect 42352 238014 42380 248526
rect 42182 237986 42380 238014
rect 42444 237425 42472 251146
rect 42430 237416 42486 237425
rect 42430 237351 42486 237360
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42430 234560 42486 234569
rect 42430 234495 42486 234504
rect 42444 234342 42472 234495
rect 42182 234314 42472 234342
rect 42182 233667 42472 233695
rect 42154 233336 42210 233345
rect 42154 233271 42210 233280
rect 42168 233104 42196 233271
rect 42444 232665 42472 233667
rect 42430 232656 42486 232665
rect 42430 232591 42486 232600
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 41786 230480 41842 230489
rect 41786 230415 41842 230424
rect 42432 230444 42484 230450
rect 41800 229976 41828 230415
rect 42432 230386 42484 230392
rect 42444 229378 42472 230386
rect 42182 229350 42472 229378
rect 41970 228984 42026 228993
rect 41970 228919 42026 228928
rect 41984 228820 42012 228919
rect 42432 227724 42484 227730
rect 42432 227666 42484 227672
rect 42444 226998 42472 227666
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42472 226318
rect 42246 226128 42302 226137
rect 42246 226063 42302 226072
rect 42260 225706 42288 226063
rect 42182 225678 42288 225706
rect 42168 223553 42196 225148
rect 42444 224913 42472 226290
rect 42614 225584 42670 225593
rect 42614 225519 42670 225528
rect 42430 224904 42486 224913
rect 42430 224839 42486 224848
rect 42154 223544 42210 223553
rect 42154 223479 42210 223488
rect 42628 219434 42656 225519
rect 41708 219406 42656 219434
rect 35806 217968 35862 217977
rect 35806 217903 35862 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35820 214713 35848 217903
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 41708 213994 41736 219406
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 35438 212256 35494 212265
rect 35438 212191 35494 212200
rect 35452 211206 35480 212191
rect 42812 211857 42840 252991
rect 42982 252240 43038 252249
rect 42982 252175 43038 252184
rect 42996 251174 43024 252175
rect 42904 251146 43024 251174
rect 43272 251174 43300 253906
rect 43272 251146 43484 251174
rect 42904 244274 42932 251146
rect 43074 249384 43130 249393
rect 43074 249319 43130 249328
rect 42904 244246 43024 244274
rect 42996 227730 43024 244246
rect 43088 238754 43116 249319
rect 43088 238726 43208 238754
rect 43180 230450 43208 238726
rect 43168 230444 43220 230450
rect 43168 230386 43220 230392
rect 42984 227724 43036 227730
rect 42984 227666 43036 227672
rect 35622 211848 35678 211857
rect 35622 211783 35678 211792
rect 39578 211848 39634 211857
rect 39578 211783 39634 211792
rect 42798 211848 42854 211857
rect 42798 211783 42854 211792
rect 35636 211342 35664 211783
rect 39592 211614 39620 211783
rect 35808 211608 35860 211614
rect 35808 211550 35860 211556
rect 39580 211608 39632 211614
rect 39580 211550 39632 211556
rect 35820 211449 35848 211550
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35624 211336 35676 211342
rect 35624 211278 35676 211284
rect 41696 211336 41748 211342
rect 41696 211278 41748 211284
rect 35440 211200 35492 211206
rect 35440 211142 35492 211148
rect 41328 211200 41380 211206
rect 41328 211142 41380 211148
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209846 35848 210151
rect 35808 209840 35860 209846
rect 35808 209782 35860 209788
rect 40316 209840 40368 209846
rect 40316 209782 40368 209788
rect 35622 208992 35678 209001
rect 35622 208927 35678 208936
rect 35636 208418 35664 208927
rect 35806 208584 35862 208593
rect 35806 208519 35808 208528
rect 35860 208519 35862 208528
rect 35808 208490 35860 208496
rect 35624 208412 35676 208418
rect 35624 208354 35676 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 208185 40080 208354
rect 40038 208176 40094 208185
rect 40038 208111 40094 208120
rect 35806 207768 35862 207777
rect 35806 207703 35862 207712
rect 35820 207194 35848 207703
rect 35808 207188 35860 207194
rect 35808 207130 35860 207136
rect 35806 206136 35862 206145
rect 35806 206071 35862 206080
rect 35820 205834 35848 206071
rect 35808 205828 35860 205834
rect 35808 205770 35860 205776
rect 40328 205737 40356 209782
rect 40684 208548 40736 208554
rect 40684 208490 40736 208496
rect 40696 206961 40724 208490
rect 41144 207188 41196 207194
rect 41144 207130 41196 207136
rect 40682 206952 40738 206961
rect 40682 206887 40738 206896
rect 41156 206145 41184 207130
rect 41340 206553 41368 211142
rect 41708 207777 41736 211278
rect 41694 207768 41750 207777
rect 41694 207703 41750 207712
rect 42890 206952 42946 206961
rect 42890 206887 42946 206896
rect 41326 206544 41382 206553
rect 41326 206479 41382 206488
rect 41142 206136 41198 206145
rect 41142 206071 41198 206080
rect 40684 205828 40736 205834
rect 40684 205770 40736 205776
rect 40314 205728 40370 205737
rect 40314 205663 40370 205672
rect 35806 204912 35862 204921
rect 35806 204847 35862 204856
rect 35820 204678 35848 204847
rect 35808 204672 35860 204678
rect 35808 204614 35860 204620
rect 35806 204504 35862 204513
rect 35806 204439 35862 204448
rect 35820 204338 35848 204439
rect 35808 204332 35860 204338
rect 35808 204274 35860 204280
rect 28538 203688 28594 203697
rect 28538 203623 28594 203632
rect 28552 199345 28580 203623
rect 40696 203289 40724 205770
rect 41696 204536 41748 204542
rect 41694 204504 41696 204513
rect 41748 204504 41750 204513
rect 41694 204439 41750 204448
rect 41696 204332 41748 204338
rect 41696 204274 41748 204280
rect 41708 204105 41736 204274
rect 41694 204096 41750 204105
rect 41694 204031 41750 204040
rect 40682 203280 40738 203289
rect 40682 203215 40738 203224
rect 28538 199336 28594 199345
rect 28538 199271 28594 199280
rect 42246 199336 42302 199345
rect 42246 199271 42302 199280
rect 42062 197024 42118 197033
rect 42062 196959 42118 196968
rect 42076 196656 42104 196959
rect 42260 195786 42288 199271
rect 42168 195758 42288 195786
rect 42168 195432 42196 195758
rect 41878 195256 41934 195265
rect 41878 195191 41934 195200
rect 41892 194820 41920 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 41786 193216 41842 193225
rect 41786 193151 41842 193160
rect 41800 192984 41828 193151
rect 42076 191593 42104 191760
rect 42062 191584 42118 191593
rect 42062 191519 42118 191528
rect 42168 191026 42196 191148
rect 42260 191026 42288 194919
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42904 190454 42932 206887
rect 43166 206136 43222 206145
rect 43166 206071 43222 206080
rect 43180 205634 43208 206071
rect 43180 205606 43300 205634
rect 43074 203280 43130 203289
rect 43074 203215 43130 203224
rect 43088 202874 43116 203215
rect 43088 202846 43208 202874
rect 43180 190454 43208 202846
rect 42430 190431 42486 190440
rect 42628 190426 42932 190454
rect 42996 190426 43208 190454
rect 42628 190074 42656 190426
rect 42536 190046 42656 190074
rect 42536 189938 42564 190046
rect 42182 189910 42564 189938
rect 42996 187490 43024 190426
rect 42536 187462 43024 187490
rect 42536 187459 42564 187462
rect 42182 187431 42564 187459
rect 42430 186824 42486 186833
rect 42182 186782 42430 186810
rect 42430 186759 42486 186768
rect 41786 186416 41842 186425
rect 41786 186351 41842 186360
rect 41800 186184 41828 186351
rect 41786 186008 41842 186017
rect 41786 185943 41842 185952
rect 41800 185605 41828 185943
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 43272 183546 43300 205606
rect 42536 183518 43300 183546
rect 42536 183138 42564 183518
rect 42182 183110 42564 183138
rect 42182 182463 42472 182491
rect 42076 179353 42104 181900
rect 42444 180713 42472 182463
rect 42430 180704 42486 180713
rect 42430 180639 42486 180648
rect 42062 179344 42118 179353
rect 42062 179279 42118 179288
rect 43456 44198 43484 251146
rect 43810 247752 43866 247761
rect 43810 247687 43866 247696
rect 43626 245576 43682 245585
rect 43626 245511 43682 245520
rect 43640 44334 43668 245511
rect 43824 234569 43852 247687
rect 43810 234560 43866 234569
rect 43810 234495 43866 234504
rect 44284 212129 44312 254759
rect 44454 251968 44510 251977
rect 44454 251903 44510 251912
rect 44468 233345 44496 251903
rect 44454 233336 44510 233345
rect 44454 233271 44510 233280
rect 44652 213761 44680 256391
rect 44836 255241 44864 298007
rect 45006 293992 45062 294001
rect 45006 293927 45062 293936
rect 45020 272921 45048 293927
rect 46216 292466 46244 300455
rect 46204 292460 46256 292466
rect 46204 292402 46256 292408
rect 48962 289912 49018 289921
rect 48962 289847 49018 289856
rect 46204 285728 46256 285734
rect 46204 285670 46256 285676
rect 45006 272912 45062 272921
rect 45006 272847 45062 272856
rect 46216 258097 46244 285670
rect 47768 280356 47820 280362
rect 47768 280298 47820 280304
rect 46202 258088 46258 258097
rect 46202 258023 46258 258032
rect 45558 255640 45614 255649
rect 45558 255575 45614 255584
rect 44822 255232 44878 255241
rect 44822 255167 44878 255176
rect 44822 252784 44878 252793
rect 44822 252719 44878 252728
rect 44836 226137 44864 252719
rect 45190 251560 45246 251569
rect 45190 251495 45246 251504
rect 45006 249112 45062 249121
rect 45006 249047 45062 249056
rect 45020 231849 45048 249047
rect 45204 240145 45232 251495
rect 45190 240136 45246 240145
rect 45190 240071 45246 240080
rect 45006 231840 45062 231849
rect 45006 231775 45062 231784
rect 44822 226128 44878 226137
rect 44822 226063 44878 226072
rect 44638 213752 44694 213761
rect 44638 213687 44694 213696
rect 45572 212945 45600 255575
rect 45926 251152 45982 251161
rect 45926 251087 45982 251096
rect 45742 248704 45798 248713
rect 45742 248639 45798 248648
rect 45756 232665 45784 248639
rect 45742 232656 45798 232665
rect 45742 232591 45798 232600
rect 45940 224913 45968 251087
rect 46110 248296 46166 248305
rect 46110 248231 46166 248240
rect 46124 235929 46152 248231
rect 47582 246664 47638 246673
rect 47582 246599 47638 246608
rect 46110 235920 46166 235929
rect 46110 235855 46166 235864
rect 45926 224904 45982 224913
rect 45926 224839 45982 224848
rect 45558 212936 45614 212945
rect 45558 212871 45614 212880
rect 44270 212120 44326 212129
rect 44270 212055 44326 212064
rect 46938 209672 46994 209681
rect 46938 209607 46994 209616
rect 44362 208448 44418 208457
rect 44362 208383 44418 208392
rect 44178 207224 44234 207233
rect 44178 207159 44234 207168
rect 43994 204504 44050 204513
rect 43994 204439 44050 204448
rect 43810 204096 43866 204105
rect 43810 204031 43866 204040
rect 43824 45218 43852 204031
rect 44008 191593 44036 204439
rect 43994 191584 44050 191593
rect 43994 191519 44050 191528
rect 44192 186833 44220 207159
rect 44376 197033 44404 208383
rect 44638 205320 44694 205329
rect 44638 205255 44694 205264
rect 44362 197024 44418 197033
rect 44362 196959 44418 196968
rect 44652 190505 44680 205255
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44638 190496 44694 190505
rect 44638 190431 44694 190440
rect 44178 186824 44234 186833
rect 44178 186759 44234 186768
rect 44836 74534 44864 204711
rect 46202 203552 46258 203561
rect 46202 203487 46258 203496
rect 44836 74506 45508 74534
rect 45480 49026 45508 74506
rect 46216 51746 46244 203487
rect 46952 180713 46980 209607
rect 46938 180704 46994 180713
rect 46938 180639 46994 180648
rect 47596 53106 47624 246599
rect 47780 214985 47808 280298
rect 47766 214976 47822 214985
rect 47766 214911 47822 214920
rect 47766 213344 47822 213353
rect 47766 213279 47822 213288
rect 47780 190505 47808 213279
rect 47950 210896 48006 210905
rect 47950 210831 48006 210840
rect 47964 195922 47992 210831
rect 48778 206544 48834 206553
rect 48778 206479 48834 206488
rect 47964 195894 48360 195922
rect 48332 194449 48360 195894
rect 48318 194440 48374 194449
rect 48318 194375 48374 194384
rect 48792 192409 48820 206479
rect 48778 192400 48834 192409
rect 48778 192335 48834 192344
rect 47766 190496 47822 190505
rect 47766 190431 47822 190440
rect 48976 53242 49004 289847
rect 49146 247480 49202 247489
rect 49146 247415 49202 247424
rect 48964 53236 49016 53242
rect 48964 53178 49016 53184
rect 47584 53100 47636 53106
rect 47584 53042 47636 53048
rect 46204 51740 46256 51746
rect 46204 51682 46256 51688
rect 49160 50386 49188 247415
rect 49514 207768 49570 207777
rect 49514 207703 49570 207712
rect 49528 196489 49556 207703
rect 49514 196480 49570 196489
rect 49514 196415 49570 196424
rect 50356 51882 50384 333095
rect 50526 290728 50582 290737
rect 50526 290663 50582 290672
rect 50540 53378 50568 290663
rect 50712 218884 50764 218890
rect 50712 218826 50764 218832
rect 50724 179353 50752 218826
rect 50710 179344 50766 179353
rect 50710 179279 50766 179288
rect 50528 53372 50580 53378
rect 50528 53314 50580 53320
rect 50344 51876 50396 51882
rect 50344 51818 50396 51824
rect 49148 50380 49200 50386
rect 49148 50322 49200 50328
rect 51736 49162 51764 334047
rect 53838 320784 53894 320793
rect 53838 320719 53894 320728
rect 53102 319424 53158 319433
rect 53102 319359 53158 319368
rect 53116 315994 53144 319359
rect 53852 317422 53880 320719
rect 53840 317416 53892 317422
rect 62120 317416 62172 317422
rect 53840 317358 53892 317364
rect 62118 317384 62120 317393
rect 62172 317384 62174 317393
rect 62118 317319 62174 317328
rect 62118 316024 62174 316033
rect 53104 315988 53156 315994
rect 62118 315959 62120 315968
rect 53104 315930 53156 315936
rect 62172 315959 62174 315968
rect 62120 315930 62172 315936
rect 62118 314800 62174 314809
rect 59912 314764 59964 314770
rect 62118 314735 62120 314744
rect 59912 314706 59964 314712
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 59924 309097 59952 314706
rect 62776 311817 62804 341391
rect 62960 313041 62988 341663
rect 63144 314129 63172 342178
rect 651380 328296 651432 328302
rect 651380 328238 651432 328244
rect 651392 328137 651420 328238
rect 651378 328128 651434 328137
rect 651378 328063 651434 328072
rect 652036 326913 652064 356623
rect 652390 352608 652446 352617
rect 652390 352543 652446 352552
rect 652404 329769 652432 352543
rect 653402 338736 653458 338745
rect 653402 338671 653458 338680
rect 652390 329760 652446 329769
rect 652390 329695 652446 329704
rect 652022 326904 652078 326913
rect 652022 326839 652078 326848
rect 651378 325680 651434 325689
rect 653416 325650 653444 338671
rect 654796 328302 654824 358527
rect 658922 346488 658978 346497
rect 658922 346423 658978 346432
rect 654784 328296 654836 328302
rect 654784 328238 654836 328244
rect 651378 325615 651380 325624
rect 651432 325615 651434 325624
rect 653404 325644 653456 325650
rect 651380 325586 651432 325592
rect 653404 325586 653456 325592
rect 63130 314120 63186 314129
rect 63130 314055 63186 314064
rect 653402 313304 653458 313313
rect 653402 313239 653458 313248
rect 62946 313032 63002 313041
rect 62946 312967 63002 312976
rect 62762 311808 62818 311817
rect 62762 311743 62818 311752
rect 652298 309904 652354 309913
rect 652298 309839 652354 309848
rect 59910 309088 59966 309097
rect 59910 309023 59966 309032
rect 651380 303544 651432 303550
rect 651380 303486 651432 303492
rect 651392 303385 651420 303486
rect 651378 303376 651434 303385
rect 651378 303311 651434 303320
rect 652312 302161 652340 309839
rect 653416 303550 653444 313239
rect 653404 303544 653456 303550
rect 653404 303486 653456 303492
rect 652298 302152 652354 302161
rect 652298 302087 652354 302096
rect 53102 301336 53158 301345
rect 53102 301271 53158 301280
rect 53116 291174 53144 301271
rect 654782 300928 654838 300937
rect 654782 300863 654838 300872
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 62762 298752 62818 298761
rect 62762 298687 62818 298696
rect 651470 298752 651526 298761
rect 651470 298687 651526 298696
rect 62118 295488 62174 295497
rect 58624 295452 58676 295458
rect 62118 295423 62120 295432
rect 58624 295394 58676 295400
rect 62172 295423 62174 295432
rect 62120 295394 62172 295400
rect 57244 294092 57296 294098
rect 57244 294034 57296 294040
rect 54484 292596 54536 292602
rect 54484 292538 54536 292544
rect 53104 291168 53156 291174
rect 53104 291110 53156 291116
rect 54496 266257 54524 292538
rect 55864 288516 55916 288522
rect 55864 288458 55916 288464
rect 54482 266248 54538 266257
rect 54482 266183 54538 266192
rect 55876 223553 55904 288458
rect 57256 275913 57284 294034
rect 58636 278769 58664 295394
rect 62118 294128 62174 294137
rect 62118 294063 62120 294072
rect 62172 294063 62174 294072
rect 62120 294034 62172 294040
rect 62302 292768 62358 292777
rect 62302 292703 62358 292712
rect 62316 292602 62344 292703
rect 62304 292596 62356 292602
rect 62304 292538 62356 292544
rect 62118 292496 62174 292505
rect 62118 292431 62120 292440
rect 62172 292431 62174 292440
rect 62120 292402 62172 292408
rect 62120 291168 62172 291174
rect 62120 291110 62172 291116
rect 62132 291009 62160 291110
rect 62118 291000 62174 291009
rect 62118 290935 62174 290944
rect 62776 289785 62804 298687
rect 651484 298178 651512 298687
rect 651472 298172 651524 298178
rect 651472 298114 651524 298120
rect 651470 297528 651526 297537
rect 651470 297463 651526 297472
rect 651484 297090 651512 297463
rect 651472 297084 651524 297090
rect 651472 297026 651524 297032
rect 652666 296848 652722 296857
rect 652666 296783 652722 296792
rect 652680 296002 652708 296783
rect 652668 295996 652720 296002
rect 652668 295938 652720 295944
rect 652390 295352 652446 295361
rect 652390 295287 652446 295296
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651470 293040 651526 293049
rect 651470 292975 651526 292984
rect 651484 292602 651512 292975
rect 651472 292596 651524 292602
rect 651472 292538 651524 292544
rect 652206 291544 652262 291553
rect 652206 291479 652262 291488
rect 651470 290456 651526 290465
rect 651470 290391 651526 290400
rect 651484 289882 651512 290391
rect 651472 289876 651524 289882
rect 651472 289818 651524 289824
rect 62762 289776 62818 289785
rect 62762 289711 62818 289720
rect 651470 289232 651526 289241
rect 651470 289167 651526 289176
rect 62118 288552 62174 288561
rect 62118 288487 62120 288496
rect 62172 288487 62174 288496
rect 62120 288458 62172 288464
rect 651484 288454 651512 289167
rect 652022 288552 652078 288561
rect 652022 288487 652078 288496
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651470 287464 651526 287473
rect 651470 287399 651526 287408
rect 63130 287192 63186 287201
rect 63130 287127 63186 287136
rect 62118 285968 62174 285977
rect 62118 285903 62174 285912
rect 62132 285734 62160 285903
rect 62120 285728 62172 285734
rect 62120 285670 62172 285676
rect 62118 284472 62174 284481
rect 60004 284436 60056 284442
rect 62118 284407 62120 284416
rect 60004 284378 60056 284384
rect 62172 284407 62174 284416
rect 62120 284378 62172 284384
rect 58622 278760 58678 278769
rect 58622 278695 58678 278704
rect 57242 275904 57298 275913
rect 57242 275839 57298 275848
rect 60016 256737 60044 284378
rect 62762 283248 62818 283257
rect 62762 283183 62818 283192
rect 62118 280936 62174 280945
rect 62118 280871 62174 280880
rect 61382 280392 61438 280401
rect 62132 280362 62160 280871
rect 61382 280327 61438 280336
rect 62120 280356 62172 280362
rect 60002 256728 60058 256737
rect 60002 256663 60058 256672
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 55862 223544 55918 223553
rect 55862 223479 55918 223488
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 60648 227452 60700 227458
rect 60648 227394 60700 227400
rect 58992 225616 59044 225622
rect 58992 225558 59044 225564
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217274 59032 225558
rect 59360 221468 59412 221474
rect 59360 221410 59412 221416
rect 59372 218074 59400 221410
rect 59820 218748 59872 218754
rect 59820 218690 59872 218696
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218690
rect 60660 217274 60688 227394
rect 61396 219434 61424 280327
rect 62120 280298 62172 280304
rect 61660 228540 61712 228546
rect 61660 228482 61712 228488
rect 61304 219406 61424 219434
rect 61304 217977 61332 219406
rect 61672 218210 61700 228482
rect 62028 225208 62080 225214
rect 62028 225150 62080 225156
rect 61660 218204 61712 218210
rect 61660 218146 61712 218152
rect 62040 218074 62068 225150
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 62028 218068 62080 218074
rect 62028 218010 62080 218016
rect 61290 217968 61346 217977
rect 61290 217903 61346 217912
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218962
rect 62776 218890 62804 283183
rect 62946 282160 63002 282169
rect 62946 282095 63002 282104
rect 62960 225593 62988 282095
rect 63144 267073 63172 287127
rect 651484 287094 651512 287399
rect 651472 287088 651524 287094
rect 651472 287030 651524 287036
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 651470 283384 651526 283393
rect 651470 283319 651526 283328
rect 651484 282946 651512 283319
rect 651472 282940 651524 282946
rect 651472 282882 651524 282888
rect 651470 280936 651526 280945
rect 651470 280871 651526 280880
rect 651484 280226 651512 280871
rect 651472 280220 651524 280226
rect 651472 280162 651524 280168
rect 65904 273970 65932 278052
rect 67100 274378 67128 278052
rect 67088 274372 67140 274378
rect 67088 274314 67140 274320
rect 65892 273964 65944 273970
rect 65892 273906 65944 273912
rect 68204 271182 68232 278052
rect 69400 272542 69428 278052
rect 69388 272536 69440 272542
rect 69388 272478 69440 272484
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269958 70624 278052
rect 71792 275330 71820 278052
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 272678 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272672 73028 272678
rect 72976 272614 73028 272620
rect 75380 271318 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76748 274712 76800 274718
rect 76748 274654 76800 274660
rect 75368 271312 75420 271318
rect 75368 271254 75420 271260
rect 70584 269952 70636 269958
rect 70584 269894 70636 269900
rect 76760 269822 76788 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76748 269816 76800 269822
rect 76748 269758 76800 269764
rect 78876 269550 78904 278052
rect 80072 277394 80100 278052
rect 80072 277366 80192 277394
rect 80164 269958 80192 277366
rect 81268 275466 81296 278052
rect 81256 275460 81308 275466
rect 81256 275402 81308 275408
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 79968 269952 80020 269958
rect 79968 269894 80020 269900
rect 80152 269952 80204 269958
rect 80152 269894 80204 269900
rect 78864 269544 78916 269550
rect 78864 269486 78916 269492
rect 79980 267170 80008 269894
rect 84120 269074 84148 278038
rect 85500 270094 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 270088 85540 270094
rect 85488 270030 85540 270036
rect 84108 269068 84160 269074
rect 84108 269010 84160 269016
rect 86236 267442 86264 275538
rect 87156 271454 87184 278052
rect 87144 271448 87196 271454
rect 87144 271390 87196 271396
rect 88352 270366 88380 278052
rect 89456 278038 89562 278066
rect 89456 274242 89484 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89444 274236 89496 274242
rect 89444 274178 89496 274184
rect 88340 270360 88392 270366
rect 88340 270302 88392 270308
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 79968 267164 80020 267170
rect 79968 267106 80020 267112
rect 63130 267064 63186 267073
rect 90376 267034 90404 274654
rect 92400 268394 92428 278038
rect 93044 275738 93072 278052
rect 93032 275732 93084 275738
rect 93032 275674 93084 275680
rect 94240 271590 94268 278052
rect 95436 274378 95464 278052
rect 96632 274582 96660 278052
rect 97842 278038 97948 278066
rect 96620 274576 96672 274582
rect 96620 274518 96672 274524
rect 95884 274508 95936 274514
rect 95884 274450 95936 274456
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 271584 94280 271590
rect 94228 271526 94280 271532
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 95896 267578 95924 274450
rect 97920 270230 97948 278038
rect 99024 272950 99052 278052
rect 100128 275874 100156 278052
rect 100116 275868 100168 275874
rect 100116 275810 100168 275816
rect 101324 273086 101352 278052
rect 101312 273080 101364 273086
rect 101312 273022 101364 273028
rect 99012 272944 99064 272950
rect 99012 272886 99064 272892
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 102520 268530 102548 278052
rect 103716 274786 103744 278052
rect 104926 278038 105216 278066
rect 103704 274780 103756 274786
rect 103704 274722 103756 274728
rect 104808 274780 104860 274786
rect 104808 274722 104860 274728
rect 102508 268524 102560 268530
rect 102508 268466 102560 268472
rect 95884 267572 95936 267578
rect 95884 267514 95936 267520
rect 104820 267306 104848 274722
rect 105188 274514 105216 278038
rect 105176 274508 105228 274514
rect 105176 274450 105228 274456
rect 106108 271726 106136 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 271862 108436 278052
rect 109618 278038 110276 278066
rect 108396 271856 108448 271862
rect 108396 271798 108448 271804
rect 106096 271720 106148 271726
rect 106096 271662 106148 271668
rect 110248 268666 110276 278038
rect 110800 275058 110828 278052
rect 110788 275052 110840 275058
rect 110788 274994 110840 275000
rect 111996 268938 112024 278052
rect 113206 278038 113496 278066
rect 113468 273834 113496 278038
rect 113456 273828 113508 273834
rect 113456 273770 113508 273776
rect 114388 273222 114416 278052
rect 115506 278038 115888 278066
rect 114376 273216 114428 273222
rect 114376 273158 114428 273164
rect 111984 268932 112036 268938
rect 111984 268874 112036 268880
rect 115860 268802 115888 278038
rect 116688 271046 116716 278052
rect 117884 274650 117912 278052
rect 117688 274644 117740 274650
rect 117688 274586 117740 274592
rect 117872 274644 117924 274650
rect 117872 274586 117924 274592
rect 116676 271040 116728 271046
rect 116676 270982 116728 270988
rect 115848 268796 115900 268802
rect 115848 268738 115900 268744
rect 110236 268660 110288 268666
rect 110236 268602 110288 268608
rect 117700 267714 117728 274586
rect 119080 272270 119108 278052
rect 120276 272406 120304 278052
rect 121486 278038 121684 278066
rect 120264 272400 120316 272406
rect 120264 272342 120316 272348
rect 119068 272264 119120 272270
rect 119068 272206 119120 272212
rect 121460 270360 121512 270366
rect 121460 270302 121512 270308
rect 117688 267708 117740 267714
rect 117688 267650 117740 267656
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 63130 266999 63186 267008
rect 90364 267028 90416 267034
rect 90364 266970 90416 266976
rect 121472 266898 121500 270302
rect 121656 269278 121684 278038
rect 122484 278038 122590 278066
rect 122484 270366 122512 278038
rect 123772 273698 123800 278052
rect 123760 273692 123812 273698
rect 123760 273634 123812 273640
rect 124968 270910 124996 278052
rect 126178 278038 126928 278066
rect 124956 270904 125008 270910
rect 124956 270846 125008 270852
rect 122472 270360 122524 270366
rect 122472 270302 122524 270308
rect 126900 269686 126928 278038
rect 127360 270774 127388 278052
rect 127348 270768 127400 270774
rect 127348 270710 127400 270716
rect 126888 269680 126940 269686
rect 126888 269622 126940 269628
rect 121644 269272 121696 269278
rect 121644 269214 121696 269220
rect 128556 268258 128584 278052
rect 129476 278038 129674 278066
rect 129476 270502 129504 278038
rect 130856 272134 130884 278052
rect 132052 274922 132080 278052
rect 133262 278038 133828 278066
rect 132040 274916 132092 274922
rect 132040 274858 132092 274864
rect 130844 272128 130896 272134
rect 130844 272070 130896 272076
rect 129464 270496 129516 270502
rect 129464 270438 129516 270444
rect 133800 269550 133828 278038
rect 134444 273562 134472 278052
rect 134432 273556 134484 273562
rect 134432 273498 134484 273504
rect 135640 273426 135668 278052
rect 136836 274786 136864 278052
rect 136824 274780 136876 274786
rect 136824 274722 136876 274728
rect 137652 274780 137704 274786
rect 137652 274722 137704 274728
rect 136824 273964 136876 273970
rect 136824 273906 136876 273912
rect 135628 273420 135680 273426
rect 135628 273362 135680 273368
rect 130384 269544 130436 269550
rect 130384 269486 130436 269492
rect 133788 269544 133840 269550
rect 133788 269486 133840 269492
rect 128544 268252 128596 268258
rect 128544 268194 128596 268200
rect 121460 266892 121512 266898
rect 121460 266834 121512 266840
rect 130396 266762 130424 269486
rect 130384 266756 130436 266762
rect 130384 266698 130436 266704
rect 136836 264330 136864 273906
rect 137664 269074 137692 274722
rect 137940 270638 137968 278052
rect 139136 275194 139164 278052
rect 140346 278038 140728 278066
rect 139124 275188 139176 275194
rect 139124 275130 139176 275136
rect 139400 272536 139452 272542
rect 139400 272478 139452 272484
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137928 270632 137980 270638
rect 137928 270574 137980 270580
rect 137468 269068 137520 269074
rect 137468 269010 137520 269016
rect 137652 269068 137704 269074
rect 137652 269010 137704 269016
rect 137480 266626 137508 269010
rect 138112 267572 138164 267578
rect 138112 267514 138164 267520
rect 137468 266620 137520 266626
rect 137468 266562 137520 266568
rect 136836 264302 137310 264330
rect 138124 264316 138152 267514
rect 138492 264330 138520 271118
rect 139412 264330 139440 272478
rect 140700 269414 140728 278038
rect 141056 275324 141108 275330
rect 141056 275266 141108 275272
rect 140688 269408 140740 269414
rect 140688 269350 140740 269356
rect 140596 267164 140648 267170
rect 140596 267106 140648 267112
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140608 264316 140636 267106
rect 141068 264330 141096 275266
rect 141528 272542 141556 278052
rect 142160 272672 142212 272678
rect 142160 272614 142212 272620
rect 141516 272536 141568 272542
rect 141516 272478 141568 272484
rect 142172 264330 142200 272614
rect 142724 271318 142752 278052
rect 143920 274786 143948 278052
rect 143908 274780 143960 274786
rect 143908 274722 143960 274728
rect 144368 274780 144420 274786
rect 144368 274722 144420 274728
rect 142712 271312 142764 271318
rect 142712 271254 142764 271260
rect 144184 271312 144236 271318
rect 144184 271254 144236 271260
rect 142712 271176 142764 271182
rect 142712 271118 142764 271124
rect 142724 264330 142752 271118
rect 143908 269816 143960 269822
rect 143908 269758 143960 269764
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143920 264316 143948 269758
rect 144196 267170 144224 271254
rect 144380 269822 144408 274722
rect 145116 274106 145144 278052
rect 145564 275460 145616 275466
rect 145564 275402 145616 275408
rect 145104 274100 145156 274106
rect 145104 274042 145156 274048
rect 145104 273964 145156 273970
rect 145104 273906 145156 273912
rect 144368 269816 144420 269822
rect 144368 269758 144420 269764
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 144184 267164 144236 267170
rect 144184 267106 144236 267112
rect 144748 264316 144776 267378
rect 144920 266892 144972 266898
rect 144920 266834 144972 266840
rect 144932 266490 144960 266834
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 273906
rect 145380 266892 145432 266898
rect 145380 266834 145432 266840
rect 145392 266626 145420 266834
rect 145576 266626 145604 275402
rect 146220 275330 146248 278052
rect 146208 275324 146260 275330
rect 146208 275266 146260 275272
rect 146944 275188 146996 275194
rect 146944 275130 146996 275136
rect 146956 274786 146984 275130
rect 146944 274780 146996 274786
rect 146944 274722 146996 274728
rect 147416 273970 147444 278052
rect 147404 273964 147456 273970
rect 147404 273906 147456 273912
rect 146944 273420 146996 273426
rect 146944 273362 146996 273368
rect 146392 269952 146444 269958
rect 146392 269894 146444 269900
rect 145380 266620 145432 266626
rect 145380 266562 145432 266568
rect 145564 266620 145616 266626
rect 145564 266562 145616 266568
rect 145116 264302 145590 264330
rect 146404 264316 146432 269894
rect 146956 267442 146984 273362
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 146944 267436 146996 267442
rect 146944 267378 146996 267384
rect 147220 266756 147272 266762
rect 147220 266698 147272 266704
rect 147232 264316 147260 266698
rect 148048 266620 148100 266626
rect 148048 266562 148100 266568
rect 148060 264316 148088 266562
rect 148428 264330 148456 272750
rect 148612 271182 148640 278052
rect 149808 275194 149836 278052
rect 151018 278038 151768 278066
rect 149796 275188 149848 275194
rect 149796 275130 149848 275136
rect 149704 275052 149756 275058
rect 149704 274994 149756 275000
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149428 270088 149480 270094
rect 149428 270030 149480 270036
rect 149440 264330 149468 270030
rect 149716 266762 149744 274994
rect 151740 268258 151768 278038
rect 152004 274236 152056 274242
rect 152004 274178 152056 274184
rect 150440 268252 150492 268258
rect 150440 268194 150492 268200
rect 151728 268252 151780 268258
rect 151728 268194 151780 268200
rect 150452 267578 150480 268194
rect 150440 267572 150492 267578
rect 150440 267514 150492 267520
rect 151360 267028 151412 267034
rect 151360 266970 151412 266976
rect 150532 266892 150584 266898
rect 150532 266834 150584 266840
rect 149704 266756 149756 266762
rect 149704 266698 149756 266704
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266834
rect 151372 264316 151400 266970
rect 152016 265674 152044 274178
rect 152200 272678 152228 278052
rect 153396 275058 153424 278052
rect 154316 278038 154514 278066
rect 153384 275052 153436 275058
rect 153384 274994 153436 275000
rect 152188 272672 152240 272678
rect 152188 272614 152240 272620
rect 152188 271448 152240 271454
rect 152188 271390 152240 271396
rect 152004 265668 152056 265674
rect 152004 265610 152056 265616
rect 152200 264316 152228 271390
rect 154316 271318 154344 278038
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 275052 154540 275058
rect 154488 274994 154540 275000
rect 154304 271312 154356 271318
rect 154304 271254 154356 271260
rect 154500 267034 154528 274994
rect 154776 267734 154804 275538
rect 155696 274242 155724 278052
rect 155960 275732 156012 275738
rect 155960 275674 156012 275680
rect 155684 274236 155736 274242
rect 155684 274178 155736 274184
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 154684 267706 154804 267734
rect 154488 267028 154540 267034
rect 154488 266970 154540 266976
rect 153844 266484 153896 266490
rect 153844 266426 153896 266432
rect 152740 265668 152792 265674
rect 152740 265610 152792 265616
rect 152752 264330 152780 265610
rect 152752 264302 153042 264330
rect 153856 264316 153884 266426
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 155972 265674 156000 275674
rect 156892 275602 156920 278052
rect 156880 275596 156932 275602
rect 156880 275538 156932 275544
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 156144 271584 156196 271590
rect 156144 271526 156196 271532
rect 155960 265668 156012 265674
rect 155960 265610 156012 265616
rect 156156 264330 156184 271526
rect 156788 265668 156840 265674
rect 156788 265610 156840 265616
rect 156800 264330 156828 265610
rect 157628 264330 157656 274314
rect 158088 272814 158116 278052
rect 158076 272808 158128 272814
rect 158076 272750 158128 272756
rect 159284 271454 159312 278052
rect 160480 275466 160508 278052
rect 161584 275874 161612 278052
rect 162124 276004 162176 276010
rect 162124 275946 162176 275952
rect 161388 275868 161440 275874
rect 161388 275810 161440 275816
rect 161572 275868 161624 275874
rect 161572 275810 161624 275816
rect 161756 275868 161808 275874
rect 161756 275810 161808 275816
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161400 273170 161428 275810
rect 161768 275754 161796 275810
rect 161676 275726 161796 275754
rect 161676 275058 161704 275726
rect 161848 275460 161900 275466
rect 161848 275402 161900 275408
rect 161860 275058 161888 275402
rect 161664 275052 161716 275058
rect 161664 274994 161716 275000
rect 161848 275052 161900 275058
rect 161848 274994 161900 275000
rect 161400 273142 161612 273170
rect 160192 273080 160244 273086
rect 160192 273022 160244 273028
rect 159272 271448 159324 271454
rect 159272 271390 159324 271396
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 156156 264302 156354 264330
rect 156800 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159640 267708 159692 267714
rect 159640 267650 159692 267656
rect 159652 264316 159680 267650
rect 160204 265674 160232 273022
rect 160376 272944 160428 272950
rect 160376 272886 160428 272892
rect 160192 265668 160244 265674
rect 160192 265610 160244 265616
rect 160388 264330 160416 272886
rect 161584 267734 161612 273142
rect 161584 267706 161704 267734
rect 161020 265668 161072 265674
rect 161020 265610 161072 265616
rect 161032 264330 161060 265610
rect 161676 264330 161704 267706
rect 162136 266422 162164 275946
rect 162780 272950 162808 278052
rect 163976 277394 164004 278052
rect 165186 278038 165476 278066
rect 163976 277366 164096 277394
rect 164068 275738 164096 277366
rect 163136 275732 163188 275738
rect 163136 275674 163188 275680
rect 164056 275732 164108 275738
rect 164056 275674 164108 275680
rect 162768 272944 162820 272950
rect 162768 272886 162820 272892
rect 162952 268524 163004 268530
rect 162952 268466 163004 268472
rect 162124 266416 162176 266422
rect 162124 266358 162176 266364
rect 160388 264302 160494 264330
rect 161032 264302 161322 264330
rect 161676 264302 162150 264330
rect 162964 264316 162992 268466
rect 163148 268122 163176 275674
rect 163320 274508 163372 274514
rect 163320 274450 163372 274456
rect 163136 268116 163188 268122
rect 163136 268058 163188 268064
rect 163332 264330 163360 274450
rect 164976 271720 165028 271726
rect 164976 271662 165028 271668
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 163332 264302 163806 264330
rect 164620 264316 164648 267242
rect 164988 264330 165016 271662
rect 165448 269958 165476 278038
rect 166368 274378 166396 278052
rect 167000 275868 167052 275874
rect 167000 275810 167052 275816
rect 166356 274372 166408 274378
rect 166356 274314 166408 274320
rect 165896 271856 165948 271862
rect 165896 271798 165948 271804
rect 165436 269952 165488 269958
rect 165436 269894 165488 269900
rect 165908 264330 165936 271798
rect 167012 268666 167040 275810
rect 167564 274922 167592 278052
rect 167552 274916 167604 274922
rect 167552 274858 167604 274864
rect 168760 274514 168788 278052
rect 169878 278038 170168 278066
rect 169024 274916 169076 274922
rect 169024 274858 169076 274864
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 167828 269272 167880 269278
rect 167828 269214 167880 269220
rect 167000 268660 167052 268666
rect 167000 268602 167052 268608
rect 167644 268388 167696 268394
rect 167644 268330 167696 268336
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167656 264330 167684 268330
rect 167840 267714 167868 269214
rect 168748 268932 168800 268938
rect 168748 268874 168800 268880
rect 168012 268388 168064 268394
rect 168012 268330 168064 268336
rect 168024 268122 168052 268330
rect 168012 268116 168064 268122
rect 168012 268058 168064 268064
rect 167828 267708 167880 267714
rect 167828 267650 167880 267656
rect 167656 264302 167946 264330
rect 168760 264316 168788 268874
rect 169036 267306 169064 274858
rect 169944 273828 169996 273834
rect 169944 273770 169996 273776
rect 169024 267300 169076 267306
rect 169024 267242 169076 267248
rect 169576 266756 169628 266762
rect 169576 266698 169628 266704
rect 169588 264316 169616 266698
rect 169956 264330 169984 273770
rect 170140 271590 170168 278038
rect 171060 275738 171088 278052
rect 171048 275732 171100 275738
rect 171048 275674 171100 275680
rect 171600 273216 171652 273222
rect 171600 273158 171652 273164
rect 170128 271584 170180 271590
rect 170128 271526 170180 271532
rect 171232 268524 171284 268530
rect 171232 268466 171284 268472
rect 169956 264302 170430 264330
rect 171244 264316 171272 268466
rect 171612 264330 171640 273158
rect 172256 273086 172284 278052
rect 173466 278038 173756 278066
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 173256 272264 173308 272270
rect 173256 272206 173308 272212
rect 172520 271040 172572 271046
rect 172520 270982 172572 270988
rect 172532 264330 172560 270982
rect 173268 264330 173296 272206
rect 173728 270094 173756 278038
rect 174648 274854 174676 278052
rect 174636 274848 174688 274854
rect 174636 274790 174688 274796
rect 174452 274780 174504 274786
rect 174452 274722 174504 274728
rect 174176 274644 174228 274650
rect 174176 274586 174228 274592
rect 173716 270088 173768 270094
rect 173716 270030 173768 270036
rect 174188 264330 174216 274586
rect 174464 272270 174492 274722
rect 175280 272400 175332 272406
rect 175280 272342 175332 272348
rect 174452 272264 174504 272270
rect 174452 272206 174504 272212
rect 175292 264330 175320 272342
rect 175752 271726 175780 278052
rect 175924 275052 175976 275058
rect 175924 274994 175976 275000
rect 175936 273834 175964 274994
rect 175924 273828 175976 273834
rect 175924 273770 175976 273776
rect 175740 271720 175792 271726
rect 175740 271662 175792 271668
rect 176200 270360 176252 270366
rect 176200 270302 176252 270308
rect 171612 264302 172086 264330
rect 172532 264302 172914 264330
rect 173268 264302 173742 264330
rect 174188 264302 174570 264330
rect 175292 264302 175398 264330
rect 176212 264316 176240 270302
rect 176948 268530 176976 278052
rect 178144 275874 178172 278052
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 273692 177540 273698
rect 177488 273634 177540 273640
rect 176936 268524 176988 268530
rect 176936 268466 176988 268472
rect 177028 267708 177080 267714
rect 177028 267650 177080 267656
rect 177040 264316 177068 267650
rect 177500 264330 177528 273634
rect 178684 270904 178736 270910
rect 178684 270846 178736 270852
rect 178316 269680 178368 269686
rect 178316 269622 178368 269628
rect 178328 264330 178356 269622
rect 178696 266422 178724 270846
rect 179340 270230 179368 278052
rect 180550 278038 180748 278066
rect 181746 278038 182036 278066
rect 179880 270768 179932 270774
rect 179880 270710 179932 270716
rect 179328 270224 179380 270230
rect 179328 270166 179380 270172
rect 178684 266416 178736 266422
rect 178684 266358 178736 266364
rect 179512 266416 179564 266422
rect 179512 266358 179564 266364
rect 177500 264302 177882 264330
rect 178328 264302 178710 264330
rect 179524 264316 179552 266358
rect 179892 264330 179920 270710
rect 180720 270366 180748 278038
rect 181168 270496 181220 270502
rect 181168 270438 181220 270444
rect 180708 270360 180760 270366
rect 180708 270302 180760 270308
rect 179892 264302 180366 264330
rect 181180 264316 181208 270438
rect 182008 267714 182036 278038
rect 182732 274848 182784 274854
rect 182732 274790 182784 274796
rect 182456 272128 182508 272134
rect 182456 272070 182508 272076
rect 181996 267708 182048 267714
rect 181996 267650 182048 267656
rect 181996 267572 182048 267578
rect 181996 267514 182048 267520
rect 182008 264316 182036 267514
rect 182468 264330 182496 272070
rect 182744 267714 182772 274790
rect 182928 274650 182956 278052
rect 182916 274644 182968 274650
rect 182916 274586 182968 274592
rect 184124 273222 184152 278052
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185124 273556 185176 273562
rect 185124 273498 185176 273504
rect 184112 273216 184164 273222
rect 184112 273158 184164 273164
rect 183652 269544 183704 269550
rect 183652 269486 183704 269492
rect 182732 267708 182784 267714
rect 182732 267650 182784 267656
rect 182468 264302 182850 264330
rect 183664 264316 183692 269486
rect 184480 268660 184532 268666
rect 184480 268602 184532 268608
rect 184492 264316 184520 268602
rect 185136 264330 185164 273498
rect 186424 269550 186452 278052
rect 187344 278038 187634 278066
rect 186412 269544 186464 269550
rect 186412 269486 186464 269492
rect 186136 269068 186188 269074
rect 186136 269010 186188 269016
rect 185136 264302 185334 264330
rect 186148 264316 186176 269010
rect 187344 268666 187372 278038
rect 188816 271862 188844 278052
rect 189080 275324 189132 275330
rect 189080 275266 189132 275272
rect 189092 272542 189120 275266
rect 190012 275058 190040 278052
rect 191222 278038 191512 278066
rect 192418 278038 192800 278066
rect 193522 278038 193628 278066
rect 190000 275052 190052 275058
rect 190000 274994 190052 275000
rect 189080 272536 189132 272542
rect 189080 272478 189132 272484
rect 189172 272400 189224 272406
rect 189172 272342 189224 272348
rect 188804 271856 188856 271862
rect 188804 271798 188856 271804
rect 187700 270632 187752 270638
rect 187700 270574 187752 270580
rect 187332 268660 187384 268666
rect 187332 268602 187384 268608
rect 186964 267436 187016 267442
rect 186964 267378 187016 267384
rect 186976 264316 187004 267378
rect 187712 264330 187740 270574
rect 188620 269408 188672 269414
rect 188620 269350 188672 269356
rect 187712 264302 187818 264330
rect 188632 264316 188660 269350
rect 189184 265674 189212 272342
rect 189356 272264 189408 272270
rect 189356 272206 189408 272212
rect 189172 265668 189224 265674
rect 189172 265610 189224 265616
rect 189368 264330 189396 272206
rect 191484 271998 191512 278038
rect 191748 275188 191800 275194
rect 191748 275130 191800 275136
rect 191472 271992 191524 271998
rect 191472 271934 191524 271940
rect 191760 270502 191788 275130
rect 192392 274100 192444 274106
rect 192392 274042 192444 274048
rect 191748 270496 191800 270502
rect 191748 270438 191800 270444
rect 190828 269816 190880 269822
rect 190828 269758 190880 269764
rect 189908 265668 189960 265674
rect 189908 265610 189960 265616
rect 189920 264330 189948 265610
rect 190840 264330 190868 269758
rect 191932 267164 191984 267170
rect 191932 267106 191984 267112
rect 189368 264302 189474 264330
rect 189920 264302 190302 264330
rect 190840 264302 191130 264330
rect 191944 264316 191972 267106
rect 192404 264330 192432 274042
rect 192576 271856 192628 271862
rect 192576 271798 192628 271804
rect 192588 267170 192616 271798
rect 192772 271046 192800 278038
rect 193404 273964 193456 273970
rect 193404 273906 193456 273912
rect 192760 271040 192812 271046
rect 192760 270982 192812 270988
rect 192576 267164 192628 267170
rect 192576 267106 192628 267112
rect 193416 264330 193444 273906
rect 193600 272406 193628 278038
rect 194704 272542 194732 278052
rect 195900 273970 195928 278052
rect 195888 273964 195940 273970
rect 195888 273906 195940 273912
rect 194048 272536 194100 272542
rect 194048 272478 194100 272484
rect 194692 272536 194744 272542
rect 194692 272478 194744 272484
rect 193588 272400 193640 272406
rect 193588 272342 193640 272348
rect 194060 264330 194088 272478
rect 197096 271182 197124 278052
rect 198292 274106 198320 278052
rect 198740 275460 198792 275466
rect 198740 275402 198792 275408
rect 198280 274100 198332 274106
rect 198280 274042 198332 274048
rect 197544 272672 197596 272678
rect 197544 272614 197596 272620
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 197084 271176 197136 271182
rect 197084 271118 197136 271124
rect 194796 264330 194824 271118
rect 196900 270496 196952 270502
rect 196900 270438 196952 270444
rect 196072 268252 196124 268258
rect 196072 268194 196124 268200
rect 192404 264302 192786 264330
rect 193416 264302 193614 264330
rect 194060 264302 194442 264330
rect 194796 264302 195270 264330
rect 196084 264316 196112 268194
rect 196912 264316 196940 270438
rect 197556 264330 197584 272614
rect 198096 271312 198148 271318
rect 198096 271254 198148 271260
rect 198108 264330 198136 271254
rect 198752 267850 198780 275402
rect 199488 272678 199516 278052
rect 200592 277394 200620 278052
rect 200500 277366 200620 277394
rect 200120 274236 200172 274242
rect 200120 274178 200172 274184
rect 199476 272672 199528 272678
rect 199476 272614 199528 272620
rect 198740 267844 198792 267850
rect 198740 267786 198792 267792
rect 199384 267028 199436 267034
rect 199384 266970 199436 266976
rect 197556 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 266970
rect 200132 264330 200160 274178
rect 200500 269686 200528 277366
rect 200672 272808 200724 272814
rect 200672 272750 200724 272756
rect 200488 269680 200540 269686
rect 200488 269622 200540 269628
rect 200684 264330 200712 272750
rect 201788 270502 201816 278052
rect 202328 271448 202380 271454
rect 202328 271390 202380 271396
rect 201776 270496 201828 270502
rect 201776 270438 201828 270444
rect 201868 267844 201920 267850
rect 201868 267786 201920 267792
rect 200132 264302 200238 264330
rect 200684 264302 201066 264330
rect 201880 264316 201908 267786
rect 202340 264330 202368 271390
rect 202984 269822 203012 278052
rect 203904 278038 204194 278066
rect 202972 269816 203024 269822
rect 202972 269758 203024 269764
rect 203904 268394 203932 278038
rect 205376 274242 205404 278052
rect 206376 275596 206428 275602
rect 206376 275538 206428 275544
rect 205364 274236 205416 274242
rect 205364 274178 205416 274184
rect 204260 273828 204312 273834
rect 204260 273770 204312 273776
rect 204076 269544 204128 269550
rect 204076 269486 204128 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 203892 268388 203944 268394
rect 203892 268330 203944 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204088 266898 204116 269486
rect 204076 266892 204128 266898
rect 204076 266834 204128 266840
rect 204272 264330 204300 273770
rect 204720 272944 204772 272950
rect 204720 272886 204772 272892
rect 204732 264330 204760 272886
rect 206008 269952 206060 269958
rect 206008 269894 206060 269900
rect 204272 264302 204378 264330
rect 204732 264302 205206 264330
rect 206020 264316 206048 269894
rect 206388 264330 206416 275538
rect 206572 273834 206600 278052
rect 207768 274378 207796 278052
rect 208492 274508 208544 274514
rect 208492 274450 208544 274456
rect 207296 274372 207348 274378
rect 207296 274314 207348 274320
rect 207756 274372 207808 274378
rect 207756 274314 207808 274320
rect 206560 273828 206612 273834
rect 206560 273770 206612 273776
rect 207308 264330 207336 274314
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208504 264316 208532 274450
rect 208872 272814 208900 278052
rect 208860 272808 208912 272814
rect 208860 272750 208912 272756
rect 209780 271584 209832 271590
rect 209780 271526 209832 271532
rect 209320 267300 209372 267306
rect 209320 267242 209372 267248
rect 209332 264316 209360 267242
rect 209792 264330 209820 271526
rect 210068 269958 210096 278052
rect 211264 277394 211292 278052
rect 212276 278038 212474 278066
rect 211264 277366 211384 277394
rect 211068 275732 211120 275738
rect 211068 275674 211120 275680
rect 210608 273080 210660 273086
rect 210608 273022 210660 273028
rect 210056 269952 210108 269958
rect 210056 269894 210108 269900
rect 210620 264330 210648 273022
rect 211080 271810 211108 275674
rect 211080 271782 211200 271810
rect 211172 267734 211200 271782
rect 211356 268802 211384 277366
rect 212276 271318 212304 278038
rect 213000 271720 213052 271726
rect 213000 271662 213052 271668
rect 212264 271312 212316 271318
rect 212264 271254 212316 271260
rect 212632 270088 212684 270094
rect 212632 270030 212684 270036
rect 211344 268796 211396 268802
rect 211344 268738 211396 268744
rect 211172 267706 211384 267734
rect 211356 264330 211384 267706
rect 209792 264302 210174 264330
rect 210620 264302 211002 264330
rect 211356 264302 211830 264330
rect 212644 264316 212672 270030
rect 213012 264330 213040 271662
rect 213656 271454 213684 278052
rect 214852 275466 214880 278052
rect 215970 278038 216536 278066
rect 214840 275460 214892 275466
rect 214840 275402 214892 275408
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 214104 270224 214156 270230
rect 214104 270166 214156 270172
rect 214116 266558 214144 270166
rect 214288 267708 214340 267714
rect 214288 267650 214340 267656
rect 214104 266552 214156 266558
rect 214104 266494 214156 266500
rect 213012 264302 213486 264330
rect 214300 264316 214328 267650
rect 214576 266694 214604 274586
rect 215300 270360 215352 270366
rect 215300 270302 215352 270308
rect 215116 268524 215168 268530
rect 215116 268466 215168 268472
rect 214564 266688 214616 266694
rect 214564 266630 214616 266636
rect 215128 264316 215156 268466
rect 215312 266422 215340 270302
rect 216508 270094 216536 278038
rect 217152 275874 217180 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 217140 275868 217192 275874
rect 217140 275810 217192 275816
rect 216496 270088 216548 270094
rect 216496 270030 216548 270036
rect 215944 266552 215996 266558
rect 215944 266494 215996 266500
rect 215300 266416 215352 266422
rect 215300 266358 215352 266364
rect 215956 264316 215984 266494
rect 216692 264330 216720 275810
rect 218348 275330 218376 278052
rect 218336 275324 218388 275330
rect 218336 275266 218388 275272
rect 218704 275052 218756 275058
rect 218704 274994 218756 275000
rect 218716 267306 218744 274994
rect 218888 273216 218940 273222
rect 218888 273158 218940 273164
rect 218704 267300 218756 267306
rect 218704 267242 218756 267248
rect 218900 267034 218928 273158
rect 219544 272950 219572 278052
rect 220464 278038 220754 278066
rect 219532 272944 219584 272950
rect 219532 272886 219584 272892
rect 219440 268660 219492 268666
rect 219440 268602 219492 268608
rect 219256 267572 219308 267578
rect 219256 267514 219308 267520
rect 218888 267028 218940 267034
rect 218888 266970 218940 266976
rect 218428 266688 218480 266694
rect 218428 266630 218480 266636
rect 217600 266416 217652 266422
rect 217600 266358 217652 266364
rect 216692 264302 216798 264330
rect 217612 264316 217640 266358
rect 218440 264316 218468 266630
rect 219268 264316 219296 267514
rect 219452 266422 219480 268602
rect 220464 268530 220492 278038
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220452 268524 220504 268530
rect 220452 268466 220504 268472
rect 220084 267028 220136 267034
rect 220084 266970 220136 266976
rect 219440 266416 219492 266422
rect 219440 266358 219492 266364
rect 220096 264316 220124 266970
rect 220912 266892 220964 266898
rect 220912 266834 220964 266840
rect 220924 264316 220952 266834
rect 221292 264330 221320 275946
rect 221936 275602 221964 278052
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 223132 271590 223160 278052
rect 224040 275868 224092 275874
rect 224040 275810 224092 275816
rect 224052 273086 224080 275810
rect 224236 275738 224264 278052
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 224040 273080 224092 273086
rect 224040 273022 224092 273028
rect 224224 272400 224276 272406
rect 224224 272342 224276 272348
rect 223120 271584 223172 271590
rect 223120 271526 223172 271532
rect 223488 268796 223540 268802
rect 223488 268738 223540 268744
rect 223500 267306 223528 268738
rect 223028 267300 223080 267306
rect 223028 267242 223080 267248
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 222568 266416 222620 266422
rect 222568 266358 222620 266364
rect 221292 264302 221766 264330
rect 222580 264316 222608 266358
rect 223040 264330 223068 267242
rect 223948 267164 224000 267170
rect 223948 267106 224000 267112
rect 223960 264330 223988 267106
rect 224236 266422 224264 272342
rect 225432 271862 225460 278052
rect 225052 271856 225104 271862
rect 225052 271798 225104 271804
rect 225420 271856 225472 271862
rect 225420 271798 225472 271804
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 223040 264302 223422 264330
rect 223960 264302 224250 264330
rect 225064 264316 225092 271798
rect 225512 271040 225564 271046
rect 225512 270982 225564 270988
rect 225524 264330 225552 270982
rect 226628 270230 226656 278052
rect 227824 274514 227852 278052
rect 227812 274508 227864 274514
rect 227812 274450 227864 274456
rect 229020 273970 229048 278052
rect 229192 274100 229244 274106
rect 229192 274042 229244 274048
rect 227904 273964 227956 273970
rect 227904 273906 227956 273912
rect 229008 273964 229060 273970
rect 229008 273906 229060 273912
rect 227168 272536 227220 272542
rect 227168 272478 227220 272484
rect 226616 270224 226668 270230
rect 226616 270166 226668 270172
rect 226892 269680 226944 269686
rect 226892 269622 226944 269628
rect 226904 266626 226932 269622
rect 226892 266620 226944 266626
rect 226892 266562 226944 266568
rect 226708 266416 226760 266422
rect 226708 266358 226760 266364
rect 225524 264302 225906 264330
rect 226720 264316 226748 266358
rect 227180 264330 227208 272478
rect 227916 264330 227944 273906
rect 229204 273850 229232 274042
rect 229112 273822 229232 273850
rect 228364 271856 228416 271862
rect 228364 271798 228416 271804
rect 228376 267034 228404 271798
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 265674 229140 273822
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230572 272672 230624 272678
rect 230572 272614 230624 272620
rect 229284 271176 229336 271182
rect 229284 271118 229336 271124
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 229100 265668 229152 265674
rect 229100 265610 229152 265616
rect 229296 265554 229324 271118
rect 229652 265668 229704 265674
rect 229652 265610 229704 265616
rect 229204 265526 229324 265554
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229204 264316 229232 265526
rect 229664 264330 229692 265610
rect 230584 264330 230612 272614
rect 231688 268394 231716 278038
rect 232516 275874 232544 278052
rect 232504 275868 232556 275874
rect 232504 275810 232556 275816
rect 232780 275732 232832 275738
rect 232780 275674 232832 275680
rect 232228 270496 232280 270502
rect 232228 270438 232280 270444
rect 230756 268388 230808 268394
rect 230756 268330 230808 268336
rect 231676 268388 231728 268394
rect 231676 268330 231728 268336
rect 230768 266762 230796 268330
rect 230756 266756 230808 266762
rect 230756 266698 230808 266704
rect 231676 266620 231728 266626
rect 231676 266562 231728 266568
rect 229664 264302 230046 264330
rect 230584 264302 230874 264330
rect 231688 264316 231716 266562
rect 232240 264330 232268 270438
rect 232792 270366 232820 275674
rect 233712 272678 233740 278052
rect 233884 274372 233936 274378
rect 233884 274314 233936 274320
rect 233700 272672 233752 272678
rect 233700 272614 233752 272620
rect 232780 270360 232832 270366
rect 232780 270302 232832 270308
rect 233332 269816 233384 269822
rect 233332 269758 233384 269764
rect 232240 264302 232530 264330
rect 233344 264316 233372 269758
rect 233896 266422 233924 274314
rect 234712 274236 234764 274242
rect 234712 274178 234764 274184
rect 234160 266756 234212 266762
rect 234160 266698 234212 266704
rect 233884 266416 233936 266422
rect 233884 266358 233936 266364
rect 234172 264316 234200 266698
rect 234724 264330 234752 274178
rect 234908 274106 234936 278052
rect 236104 275738 236132 278052
rect 236092 275732 236144 275738
rect 236092 275674 236144 275680
rect 236644 275460 236696 275466
rect 236644 275402 236696 275408
rect 234896 274100 234948 274106
rect 234896 274042 234948 274048
rect 235448 273828 235500 273834
rect 235448 273770 235500 273776
rect 235460 264330 235488 273770
rect 236656 267442 236684 275402
rect 237300 274242 237328 278052
rect 237288 274236 237340 274242
rect 237288 274178 237340 274184
rect 237380 272808 237432 272814
rect 237380 272750 237432 272756
rect 236644 267436 236696 267442
rect 236644 267378 236696 267384
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 234724 264302 235014 264330
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237392 264330 237420 272750
rect 238496 272542 238524 278052
rect 239404 275596 239456 275602
rect 239404 275538 239456 275544
rect 239416 275346 239444 275538
rect 239600 275466 239628 278052
rect 240810 278038 241468 278066
rect 239864 275868 239916 275874
rect 239864 275810 239916 275816
rect 239588 275460 239640 275466
rect 239588 275402 239640 275408
rect 239416 275318 239536 275346
rect 238484 272536 238536 272542
rect 238484 272478 238536 272484
rect 239312 271312 239364 271318
rect 239312 271254 239364 271260
rect 238300 269952 238352 269958
rect 238300 269894 238352 269900
rect 237392 264302 237498 264330
rect 238312 264316 238340 269894
rect 239324 267734 239352 271254
rect 239508 267734 239536 275318
rect 239876 271726 239904 275810
rect 239864 271720 239916 271726
rect 239864 271662 239916 271668
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 239324 267706 239444 267734
rect 239508 267706 239628 267734
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 239140 264316 239168 267242
rect 239416 264466 239444 267706
rect 239600 266422 239628 267706
rect 239588 266416 239640 266422
rect 239588 266358 239640 266364
rect 239416 264438 239536 264466
rect 239508 264330 239536 264438
rect 240428 264330 240456 271390
rect 241440 269822 241468 278038
rect 241992 269958 242020 278052
rect 243188 275602 243216 278052
rect 244398 278038 244688 278066
rect 243176 275596 243228 275602
rect 243176 275538 243228 275544
rect 243084 275324 243136 275330
rect 243084 275266 243136 275272
rect 242440 270088 242492 270094
rect 242440 270030 242492 270036
rect 241980 269952 242032 269958
rect 241980 269894 242032 269900
rect 241428 269816 241480 269822
rect 241428 269758 241480 269764
rect 241612 267436 241664 267442
rect 241612 267378 241664 267384
rect 239508 264302 239982 264330
rect 240428 264302 240810 264330
rect 241624 264316 241652 267378
rect 242452 264316 242480 270030
rect 243096 265674 243124 275266
rect 243268 273080 243320 273086
rect 243268 273022 243320 273028
rect 243084 265668 243136 265674
rect 243084 265610 243136 265616
rect 243280 264316 243308 273022
rect 244464 272944 244516 272950
rect 244464 272886 244516 272892
rect 243820 265668 243872 265674
rect 243820 265610 243872 265616
rect 243832 264330 243860 265610
rect 244476 264330 244504 272886
rect 244660 271318 244688 278038
rect 244648 271312 244700 271318
rect 244648 271254 244700 271260
rect 245580 268666 245608 278052
rect 246790 278038 246988 278066
rect 247894 278038 248368 278066
rect 245568 268660 245620 268666
rect 245568 268602 245620 268608
rect 245752 268524 245804 268530
rect 245752 268466 245804 268472
rect 243832 264302 244122 264330
rect 244476 264302 244950 264330
rect 245764 264316 245792 268466
rect 246960 267170 246988 278038
rect 247224 271584 247276 271590
rect 247224 271526 247276 271532
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 271526
rect 247868 270360 247920 270366
rect 247868 270302 247920 270308
rect 247880 264330 247908 270302
rect 248340 270094 248368 278038
rect 248880 274508 248932 274514
rect 248880 274450 248932 274456
rect 248328 270088 248380 270094
rect 248328 270030 248380 270036
rect 248892 266558 248920 274450
rect 249076 274378 249104 278052
rect 249064 274372 249116 274378
rect 249064 274314 249116 274320
rect 250272 271454 250300 278052
rect 250444 273964 250496 273970
rect 250444 273906 250496 273912
rect 250260 271448 250312 271454
rect 250260 271390 250312 271396
rect 249892 270224 249944 270230
rect 249892 270166 249944 270172
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 248880 266552 248932 266558
rect 248880 266494 248932 266500
rect 247236 264302 247434 264330
rect 247880 264302 248262 264330
rect 249076 264316 249104 266834
rect 249904 264316 249932 270166
rect 250456 266422 250484 273906
rect 251468 272950 251496 278052
rect 251916 275460 251968 275466
rect 251916 275402 251968 275408
rect 251456 272944 251508 272950
rect 251456 272886 251508 272892
rect 251732 271176 251784 271182
rect 251732 271118 251784 271124
rect 251744 267734 251772 271118
rect 251928 267734 251956 275402
rect 252664 272814 252692 278052
rect 253388 275732 253440 275738
rect 253388 275674 253440 275680
rect 252652 272808 252704 272814
rect 252652 272750 252704 272756
rect 253204 268388 253256 268394
rect 253204 268330 253256 268336
rect 251744 267706 251864 267734
rect 251928 267706 252048 267734
rect 250720 266552 250772 266558
rect 250720 266494 250772 266500
rect 250444 266416 250496 266422
rect 250444 266358 250496 266364
rect 250732 264316 250760 266494
rect 251548 266416 251600 266422
rect 251548 266358 251600 266364
rect 251560 264316 251588 266358
rect 251836 264330 251864 267706
rect 252020 266762 252048 267706
rect 252008 266756 252060 266762
rect 252008 266698 252060 266704
rect 251836 264302 252402 264330
rect 253216 264316 253244 268330
rect 253400 266422 253428 275674
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 272672 253992 272678
rect 253940 272614 253992 272620
rect 253388 266416 253440 266422
rect 253388 266358 253440 266364
rect 253952 265674 253980 272614
rect 254124 271720 254176 271726
rect 254124 271662 254176 271668
rect 253940 265668 253992 265674
rect 253940 265610 253992 265616
rect 254136 265554 254164 271662
rect 254964 271182 254992 278052
rect 255320 275596 255372 275602
rect 255320 275538 255372 275544
rect 255332 274106 255360 275538
rect 256160 275330 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275324 256200 275330
rect 256148 275266 256200 275272
rect 258356 274712 258408 274718
rect 258356 274654 258408 274660
rect 256976 274236 257028 274242
rect 256976 274178 257028 274184
rect 255320 274100 255372 274106
rect 255320 274042 255372 274048
rect 255412 273964 255464 273970
rect 255412 273906 255464 273912
rect 254952 271176 255004 271182
rect 254952 271118 255004 271124
rect 254492 265668 254544 265674
rect 254492 265610 254544 265616
rect 254044 265526 254164 265554
rect 254044 264316 254072 265526
rect 254504 264330 254532 265610
rect 255424 264330 255452 273906
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 254504 264302 254886 264330
rect 255424 264302 255714 264330
rect 256528 264316 256556 266358
rect 256988 264330 257016 274178
rect 258080 272536 258132 272542
rect 258080 272478 258132 272484
rect 258092 264330 258120 272478
rect 258368 268394 258396 274654
rect 258552 273970 258580 278052
rect 258540 273964 258592 273970
rect 258540 273906 258592 273912
rect 259748 270230 259776 278052
rect 260958 278038 261248 278066
rect 261220 274106 261248 278038
rect 261956 278038 262062 278066
rect 261024 274100 261076 274106
rect 261024 274042 261076 274048
rect 261208 274100 261260 274106
rect 261208 274042 261260 274048
rect 259736 270224 259788 270230
rect 259736 270166 259788 270172
rect 260380 269952 260432 269958
rect 260380 269894 260432 269900
rect 259828 269816 259880 269822
rect 259828 269758 259880 269764
rect 258356 268388 258408 268394
rect 258356 268330 258408 268336
rect 259000 266756 259052 266762
rect 259000 266698 259052 266704
rect 256988 264302 257370 264330
rect 258092 264302 258198 264330
rect 259012 264316 259040 266698
rect 259840 264316 259868 269758
rect 260392 264330 260420 269894
rect 261036 264330 261064 274042
rect 261956 269822 261984 278038
rect 262864 275596 262916 275602
rect 262864 275538 262916 275544
rect 262220 271312 262272 271318
rect 262220 271254 262272 271260
rect 261944 269816 261996 269822
rect 261944 269758 261996 269764
rect 262232 264330 262260 271254
rect 262876 270366 262904 275538
rect 263244 275466 263272 278052
rect 263232 275460 263284 275466
rect 263232 275402 263284 275408
rect 264440 272406 264468 278052
rect 265256 274372 265308 274378
rect 265256 274314 265308 274320
rect 264428 272400 264480 272406
rect 264428 272342 264480 272348
rect 262864 270360 262916 270366
rect 262864 270302 262916 270308
rect 264796 270088 264848 270094
rect 264796 270030 264848 270036
rect 263140 268660 263192 268666
rect 263140 268602 263192 268608
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262232 264302 262338 264330
rect 263152 264316 263180 268602
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263980 264316 264008 267106
rect 264808 264316 264836 270030
rect 265268 264330 265296 274314
rect 265636 271454 265664 278052
rect 266832 272678 266860 278052
rect 268028 274718 268056 278052
rect 268660 275324 268712 275330
rect 268660 275266 268712 275272
rect 268016 274712 268068 274718
rect 268016 274654 268068 274660
rect 267004 272944 267056 272950
rect 267004 272886 267056 272892
rect 266820 272672 266872 272678
rect 266820 272614 266872 272620
rect 265624 271448 265676 271454
rect 265624 271390 265676 271396
rect 266452 271312 266504 271318
rect 266452 271254 266504 271260
rect 265268 264302 265650 264330
rect 266464 264316 266492 271254
rect 267016 264330 267044 272886
rect 267924 272536 267976 272542
rect 267924 272478 267976 272484
rect 267936 264330 267964 272478
rect 268672 271930 268700 275266
rect 269224 275126 269252 278052
rect 269212 275120 269264 275126
rect 269212 275062 269264 275068
rect 268660 271924 268712 271930
rect 268660 271866 268712 271872
rect 270328 271182 270356 278052
rect 271524 272814 271552 278052
rect 272432 274712 272484 274718
rect 272432 274654 272484 274660
rect 272064 273964 272116 273970
rect 272064 273906 272116 273912
rect 271512 272808 271564 272814
rect 271512 272750 271564 272756
rect 270500 271924 270552 271930
rect 270500 271866 270552 271872
rect 269304 271176 269356 271182
rect 269304 271118 269356 271124
rect 270316 271176 270368 271182
rect 270316 271118 270368 271124
rect 268936 268388 268988 268394
rect 268936 268330 268988 268336
rect 267016 264302 267306 264330
rect 267936 264302 268134 264330
rect 268948 264316 268976 268330
rect 269316 264330 269344 271118
rect 270512 264330 270540 271866
rect 271420 270224 271472 270230
rect 271420 270166 271472 270172
rect 269316 264302 269790 264330
rect 270512 264302 270618 264330
rect 271432 264316 271460 270166
rect 272076 264330 272104 273906
rect 272444 269278 272472 274654
rect 272720 273970 272748 278052
rect 273260 275460 273312 275466
rect 273260 275402 273312 275408
rect 272708 273964 272760 273970
rect 272708 273906 272760 273912
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 272432 269272 272484 269278
rect 272432 269214 272484 269220
rect 272076 264302 272274 264330
rect 273088 264316 273116 269894
rect 273272 269006 273300 275402
rect 273916 275330 273944 278052
rect 273904 275324 273956 275330
rect 273904 275266 273956 275272
rect 274916 275120 274968 275126
rect 274916 275062 274968 275068
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269000 273312 269006
rect 273260 268942 273312 268948
rect 273548 264330 273576 274042
rect 274732 269816 274784 269822
rect 274732 269758 274784 269764
rect 273548 264302 273930 264330
rect 274744 264316 274772 269758
rect 274928 269142 274956 275062
rect 275112 274106 275140 278052
rect 276322 278038 276704 278066
rect 275100 274100 275152 274106
rect 275100 274042 275152 274048
rect 276020 272400 276072 272406
rect 276020 272342 276072 272348
rect 274916 269136 274968 269142
rect 274916 269078 274968 269084
rect 275560 269000 275612 269006
rect 275560 268942 275612 268948
rect 275572 264316 275600 268942
rect 276032 264330 276060 272342
rect 276676 271318 276704 278038
rect 277504 275670 277532 278052
rect 277492 275664 277544 275670
rect 277492 275606 277544 275612
rect 278608 273154 278636 278052
rect 279818 278038 280108 278066
rect 278596 273148 278648 273154
rect 278596 273090 278648 273096
rect 277584 272672 277636 272678
rect 277584 272614 277636 272620
rect 276848 271448 276900 271454
rect 276848 271390 276900 271396
rect 276664 271312 276716 271318
rect 276664 271254 276716 271260
rect 276860 264330 276888 271390
rect 277596 264330 277624 272614
rect 280080 269822 280108 278038
rect 280344 272808 280396 272814
rect 280344 272750 280396 272756
rect 280068 269816 280120 269822
rect 280068 269758 280120 269764
rect 278872 269272 278924 269278
rect 278872 269214 278924 269220
rect 276032 264302 276414 264330
rect 276860 264302 277242 264330
rect 277596 264302 278070 264330
rect 278884 264316 278912 269214
rect 279700 269136 279752 269142
rect 279700 269078 279752 269084
rect 279712 264316 279740 269078
rect 280356 265674 280384 272750
rect 281000 272678 281028 278052
rect 282196 274310 282224 278052
rect 282920 275324 282972 275330
rect 282920 275266 282972 275272
rect 282184 274304 282236 274310
rect 282184 274246 282236 274252
rect 281816 273964 281868 273970
rect 281816 273906 281868 273912
rect 280988 272672 281040 272678
rect 280988 272614 281040 272620
rect 280528 271176 280580 271182
rect 280528 271118 280580 271124
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 280540 264316 280568 271118
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281828 264330 281856 273906
rect 282932 264330 282960 275266
rect 283392 274718 283420 278052
rect 284588 275874 284616 278052
rect 284576 275868 284628 275874
rect 284576 275810 284628 275816
rect 284300 275664 284352 275670
rect 284300 275606 284352 275612
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283472 274100 283524 274106
rect 283472 274042 283524 274048
rect 283484 264330 283512 274042
rect 284312 265674 284340 275606
rect 285692 275466 285720 278052
rect 286888 275602 286916 278052
rect 286876 275596 286928 275602
rect 286876 275538 286928 275544
rect 285680 275460 285732 275466
rect 285680 275402 285732 275408
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274922 289308 278052
rect 290096 275868 290148 275874
rect 290096 275810 290148 275816
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 287704 274304 287756 274310
rect 287704 274246 287756 274252
rect 285864 273148 285916 273154
rect 285864 273090 285916 273096
rect 284484 271312 284536 271318
rect 284484 271254 284536 271260
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271254
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 285876 264330 285904 273090
rect 286324 272672 286376 272678
rect 286324 272614 286376 272620
rect 286336 266898 286364 272614
rect 287152 269816 287204 269822
rect 287152 269758 287204 269764
rect 286324 266892 286376 266898
rect 286324 266834 286376 266840
rect 281000 264302 281382 264330
rect 281828 264302 282210 264330
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 285876 264302 286350 264330
rect 287164 264316 287192 269758
rect 287716 266422 287744 274246
rect 287980 266892 288032 266898
rect 287980 266834 288032 266840
rect 287704 266416 287756 266422
rect 287704 266358 287756 266364
rect 287992 264316 288020 266834
rect 288808 266416 288860 266422
rect 288808 266358 288860 266364
rect 288820 264316 288848 266358
rect 289188 264330 289216 274654
rect 290108 264330 290136 275810
rect 290476 275262 290504 278052
rect 291672 275466 291700 278052
rect 291844 275596 291896 275602
rect 291844 275538 291896 275544
rect 291200 275460 291252 275466
rect 291200 275402 291252 275408
rect 291660 275460 291712 275466
rect 291660 275402 291712 275408
rect 290464 275256 290516 275262
rect 290464 275198 290516 275204
rect 291212 264330 291240 275402
rect 291856 264330 291884 275538
rect 292672 275052 292724 275058
rect 292672 274994 292724 275000
rect 292684 264330 292712 274994
rect 292868 274718 292896 278052
rect 293972 274990 294000 278052
rect 294144 275256 294196 275262
rect 294144 275198 294196 275204
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 293408 274916 293460 274922
rect 293408 274858 293460 274864
rect 292856 274712 292908 274718
rect 292856 274654 292908 274660
rect 293420 264330 293448 274858
rect 294156 264330 294184 275198
rect 295168 274854 295196 278052
rect 295432 275460 295484 275466
rect 295432 275402 295484 275408
rect 295156 274848 295208 274854
rect 295156 274790 295208 274796
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291212 264302 291318 264330
rect 291856 264302 292146 264330
rect 292684 264302 292974 264330
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295444 264316 295472 275402
rect 296364 274718 296392 278052
rect 297560 275398 297588 278052
rect 297548 275392 297600 275398
rect 297548 275334 297600 275340
rect 298756 275262 298784 278052
rect 299952 275398 299980 278052
rect 300964 278038 301070 278066
rect 302266 278038 302464 278066
rect 299572 275392 299624 275398
rect 299572 275334 299624 275340
rect 299940 275392 299992 275398
rect 299940 275334 299992 275340
rect 298744 275256 298796 275262
rect 298744 275198 298796 275204
rect 296812 274984 296864 274990
rect 296812 274926 296864 274932
rect 295800 274712 295852 274718
rect 295800 274654 295852 274660
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 295812 264330 295840 274654
rect 296824 264330 296852 274926
rect 297456 274848 297508 274854
rect 297456 274790 297508 274796
rect 297468 264330 297496 274790
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298388 264330 298416 274654
rect 295812 264302 296286 264330
rect 296824 264302 297114 264330
rect 297468 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 275334
rect 300032 275256 300084 275262
rect 300032 275198 300084 275204
rect 300044 264330 300072 275198
rect 300964 266422 300992 278038
rect 301136 275392 301188 275398
rect 301136 275334 301188 275340
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 301148 264330 301176 275334
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 301148 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 277394 310560 278052
rect 310992 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 318826 278038 319024 278066
rect 310532 277366 310652 277394
rect 310624 266694 310652 277366
rect 310612 266688 310664 266694
rect 310612 266630 310664 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310992 266422 311020 278038
rect 311912 266558 311940 278038
rect 312360 266688 312412 266694
rect 312360 266630 312412 266636
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 310980 266416 311032 266422
rect 310980 266358 311032 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312372 264330 312400 266630
rect 312820 266552 312872 266558
rect 312820 266494 312872 266500
rect 312018 264302 312400 264330
rect 312832 264316 312860 266494
rect 313292 266422 313320 278038
rect 314476 267028 314528 267034
rect 314476 266970 314528 266976
rect 313648 266892 313700 266898
rect 313648 266834 313700 266840
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 266834
rect 314488 264316 314516 266970
rect 314672 266694 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266688 314712 266694
rect 314660 266630 314712 266636
rect 315316 264316 315344 267378
rect 316052 266558 316080 278038
rect 317432 266898 317460 278038
rect 318708 273284 318760 273290
rect 318708 273226 318760 273232
rect 318720 267734 318748 273226
rect 318628 267706 318748 267734
rect 317788 267164 317840 267170
rect 317788 267106 317840 267112
rect 317420 266892 317472 266898
rect 317420 266834 317472 266840
rect 316960 266688 317012 266694
rect 316960 266630 317012 266636
rect 316040 266552 316092 266558
rect 316040 266494 316092 266500
rect 316408 266552 316460 266558
rect 316408 266494 316460 266500
rect 316420 264330 316448 266494
rect 316158 264302 316448 264330
rect 316972 264316 317000 266630
rect 317800 264316 317828 267106
rect 318628 264316 318656 267706
rect 318996 267034 319024 278038
rect 319180 278038 320022 278066
rect 320192 278038 321218 278066
rect 321572 278038 322414 278066
rect 322952 278038 323518 278066
rect 319180 267442 319208 278038
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319168 267436 319220 267442
rect 319168 267378 319220 267384
rect 318984 267028 319036 267034
rect 318984 266970 319036 266976
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321572 266694 321600 278038
rect 322756 272672 322808 272678
rect 322756 272614 322808 272620
rect 321928 266892 321980 266898
rect 321928 266834 321980 266840
rect 321560 266688 321612 266694
rect 321560 266630 321612 266636
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 266834
rect 322768 264316 322796 272614
rect 322952 267170 322980 278038
rect 324044 273964 324096 273970
rect 324044 273906 324096 273912
rect 322940 267164 322992 267170
rect 322940 267106 322992 267112
rect 324056 264330 324084 273906
rect 324700 273290 324728 278052
rect 325712 278038 325910 278066
rect 325332 274236 325384 274242
rect 325332 274178 325384 274184
rect 324688 273284 324740 273290
rect 324688 273226 324740 273232
rect 325344 266422 325372 274178
rect 325516 272536 325568 272542
rect 325516 272478 325568 272484
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 272478
rect 325712 269142 325740 278038
rect 326436 271312 326488 271318
rect 326436 271254 326488 271260
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 271254
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 327540 273284 327592 273290
rect 327540 273226 327592 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327552 266898 327580 273226
rect 329472 273080 329524 273086
rect 329472 273022 329524 273028
rect 327724 270088 327776 270094
rect 327724 270030 327776 270036
rect 327540 266892 327592 266898
rect 327540 266834 327592 266840
rect 327736 264316 327764 270030
rect 329484 266422 329512 273022
rect 330588 272678 330616 278052
rect 331784 273970 331812 278052
rect 332980 274242 333008 278052
rect 333796 274372 333848 274378
rect 333796 274314 333848 274320
rect 332968 274236 333020 274242
rect 332968 274178 333020 274184
rect 332324 274100 332376 274106
rect 332324 274042 332376 274048
rect 331772 273964 331824 273970
rect 331772 273906 331824 273912
rect 331956 273964 332008 273970
rect 331956 273906 332008 273912
rect 330576 272672 330628 272678
rect 330576 272614 330628 272620
rect 329656 271448 329708 271454
rect 329656 271390 329708 271396
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 329472 266416 329524 266422
rect 329472 266358 329524 266364
rect 328564 264316 328592 266358
rect 329668 264330 329696 271390
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 330208 266416 330260 266422
rect 330208 266358 330260 266364
rect 329406 264302 329696 264330
rect 330220 264316 330248 266358
rect 331048 264316 331076 267706
rect 331968 266422 331996 273906
rect 331956 266416 332008 266422
rect 331956 266358 332008 266364
rect 332336 264330 332364 274042
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 274314
rect 334176 272542 334204 278052
rect 335372 274666 335400 278052
rect 335096 274638 335400 274666
rect 335556 278038 336582 278066
rect 336752 278038 337778 278066
rect 334164 272536 334216 272542
rect 334164 272478 334216 272484
rect 335096 271318 335124 274638
rect 335268 272944 335320 272950
rect 335268 272886 335320 272892
rect 335084 271312 335136 271318
rect 335084 271254 335136 271260
rect 335084 269952 335136 269958
rect 335084 269894 335136 269900
rect 334348 266416 334400 266422
rect 334348 266358 334400 266364
rect 333546 264302 333836 264330
rect 334360 264316 334388 266358
rect 335096 264330 335124 269894
rect 335280 266422 335308 272886
rect 335556 269822 335584 278038
rect 336372 272808 336424 272814
rect 336372 272750 336424 272756
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 335268 266416 335320 266422
rect 335268 266358 335320 266364
rect 336384 264330 336412 272750
rect 336752 270094 336780 278038
rect 338868 273086 338896 278052
rect 338856 273080 338908 273086
rect 338856 273022 338908 273028
rect 338028 272672 338080 272678
rect 338028 272614 338080 272620
rect 336740 270088 336792 270094
rect 336740 270030 336792 270036
rect 336832 269816 336884 269822
rect 336832 269758 336884 269764
rect 335096 264302 335202 264330
rect 336030 264302 336412 264330
rect 336844 264316 336872 269758
rect 338040 264330 338068 272614
rect 340064 271454 340092 278052
rect 341260 273970 341288 278052
rect 341248 273964 341300 273970
rect 341248 273906 341300 273912
rect 342076 273964 342128 273970
rect 342076 273906 342128 273912
rect 340052 271448 340104 271454
rect 340052 271390 340104 271396
rect 340604 271448 340656 271454
rect 340604 271390 340656 271396
rect 339408 271312 339460 271318
rect 339408 271254 339460 271260
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337686 264302 338068 264330
rect 338500 264316 338528 268466
rect 339420 267734 339448 271254
rect 339328 267706 339448 267734
rect 339328 264316 339356 267706
rect 340616 264330 340644 271390
rect 340972 267572 341024 267578
rect 340972 267514 341024 267520
rect 340170 264302 340644 264330
rect 340984 264316 341012 267514
rect 342088 264330 342116 273906
rect 342456 271182 342484 278052
rect 343456 274236 343508 274242
rect 343456 274178 343508 274184
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 342628 266688 342680 266694
rect 342628 266630 342680 266636
rect 341826 264302 342116 264330
rect 342640 264316 342668 266630
rect 343468 264316 343496 274178
rect 343652 274106 343680 278052
rect 343836 278038 344862 278066
rect 343640 274100 343692 274106
rect 343640 274042 343692 274048
rect 343836 266898 343864 278038
rect 345952 274378 345980 278052
rect 346872 278038 347162 278066
rect 347792 278038 348358 278066
rect 345940 274372 345992 274378
rect 345940 274314 345992 274320
rect 346872 272950 346900 278038
rect 347044 274372 347096 274378
rect 347044 274314 347096 274320
rect 346860 272944 346912 272950
rect 346860 272886 346912 272892
rect 344652 272536 344704 272542
rect 344652 272478 344704 272484
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272478
rect 345112 270224 345164 270230
rect 345112 270166 345164 270172
rect 344310 264302 344692 264330
rect 345124 264316 345152 270166
rect 345940 270088 345992 270094
rect 345940 270030 345992 270036
rect 345952 264316 345980 270030
rect 347056 266694 347084 274314
rect 347596 271176 347648 271182
rect 347596 271118 347648 271124
rect 347044 266688 347096 266694
rect 347044 266630 347096 266636
rect 347412 266552 347464 266558
rect 347412 266494 347464 266500
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 346780 264316 346808 266358
rect 347424 264330 347452 266494
rect 347608 266422 347636 271118
rect 347792 269958 347820 278038
rect 349540 272814 349568 278052
rect 350552 278038 350750 278066
rect 350356 274100 350408 274106
rect 350356 274042 350408 274048
rect 349804 273080 349856 273086
rect 349804 273022 349856 273028
rect 349528 272808 349580 272814
rect 349528 272750 349580 272756
rect 347780 269952 347832 269958
rect 347780 269894 347832 269900
rect 348424 268388 348476 268394
rect 348424 268330 348476 268336
rect 347596 266416 347648 266422
rect 347596 266358 347648 266364
rect 347424 264302 347622 264330
rect 348436 264316 348464 268330
rect 349816 266558 349844 273022
rect 350080 267436 350132 267442
rect 350080 267378 350132 267384
rect 349804 266552 349856 266558
rect 349804 266494 349856 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 267378
rect 350368 266422 350396 274042
rect 350552 269822 350580 278038
rect 350724 274712 350776 274718
rect 350724 274654 350776 274660
rect 350540 269816 350592 269822
rect 350540 269758 350592 269764
rect 350736 268530 350764 274654
rect 351932 272678 351960 278052
rect 353128 274718 353156 278052
rect 353116 274712 353168 274718
rect 353116 274654 353168 274660
rect 352564 272808 352616 272814
rect 352564 272750 352616 272756
rect 351920 272672 351972 272678
rect 351920 272614 351972 272620
rect 351736 269952 351788 269958
rect 351736 269894 351788 269900
rect 350724 268524 350776 268530
rect 350724 268466 350776 268472
rect 350908 266552 350960 266558
rect 350908 266494 350960 266500
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 266494
rect 351748 264316 351776 269894
rect 352576 266558 352604 272750
rect 353944 271720 353996 271726
rect 353944 271662 353996 271668
rect 353392 267300 353444 267306
rect 353392 267242 353444 267248
rect 352564 266552 352616 266558
rect 352564 266494 352616 266500
rect 352564 266416 352616 266422
rect 352564 266358 352616 266364
rect 352576 264316 352604 266358
rect 353404 264316 353432 267242
rect 353956 266422 353984 271662
rect 354232 271318 354260 278052
rect 355152 278038 355442 278066
rect 354496 272672 354548 272678
rect 354496 272614 354548 272620
rect 354220 271312 354272 271318
rect 354220 271254 354272 271260
rect 353944 266416 353996 266422
rect 353944 266358 353996 266364
rect 354508 264330 354536 272614
rect 355152 271454 355180 278038
rect 356624 271862 356652 278052
rect 357820 273970 357848 278052
rect 358084 274508 358136 274514
rect 358084 274450 358136 274456
rect 357808 273964 357860 273970
rect 357808 273906 357860 273912
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271448 355192 271454
rect 355140 271390 355192 271396
rect 355048 269816 355100 269822
rect 355048 269758 355100 269764
rect 354246 264302 354536 264330
rect 355060 264316 355088 269758
rect 355336 267578 355364 271798
rect 357164 271584 357216 271590
rect 357164 271526 357216 271532
rect 355324 267572 355376 267578
rect 355324 267514 355376 267520
rect 355876 267028 355928 267034
rect 355876 266970 355928 266976
rect 355888 264316 355916 266970
rect 357176 264330 357204 271526
rect 358096 267442 358124 274450
rect 359016 274378 359044 278052
rect 359004 274372 359056 274378
rect 359004 274314 359056 274320
rect 360212 274242 360240 278052
rect 361212 275324 361264 275330
rect 361212 275266 361264 275272
rect 360200 274236 360252 274242
rect 360200 274178 360252 274184
rect 360108 273964 360160 273970
rect 360108 273906 360160 273912
rect 358728 271448 358780 271454
rect 358728 271390 358780 271396
rect 358084 267436 358136 267442
rect 358084 267378 358136 267384
rect 357532 266552 357584 266558
rect 357532 266494 357584 266500
rect 356730 264302 357204 264330
rect 357544 264316 357572 266494
rect 358740 264330 358768 271390
rect 359832 268524 359884 268530
rect 359832 268466 359884 268472
rect 359648 266756 359700 266762
rect 359648 266698 359700 266704
rect 359188 266416 359240 266422
rect 359188 266358 359240 266364
rect 358386 264302 358768 264330
rect 359200 264316 359228 266358
rect 359660 264330 359688 266698
rect 359844 266558 359872 268466
rect 359832 266552 359884 266558
rect 359832 266494 359884 266500
rect 360120 266422 360148 273906
rect 360108 266416 360160 266422
rect 360108 266358 360160 266364
rect 361224 264330 361252 275266
rect 361408 272542 361436 278052
rect 361592 278038 362526 278066
rect 362972 278038 363722 278066
rect 364536 278038 364918 278066
rect 361396 272536 361448 272542
rect 361396 272478 361448 272484
rect 361592 270230 361620 278038
rect 362776 272944 362828 272950
rect 362776 272886 362828 272892
rect 361580 270224 361632 270230
rect 361580 270166 361632 270172
rect 362500 267572 362552 267578
rect 362500 267514 362552 267520
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 359660 264302 360042 264330
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 267514
rect 362788 266422 362816 272886
rect 362972 270094 363000 278038
rect 363788 272536 363840 272542
rect 363788 272478 363840 272484
rect 362960 270088 363012 270094
rect 362960 270030 363012 270036
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 272478
rect 364536 271182 364564 278038
rect 364984 274236 365036 274242
rect 364984 274178 365036 274184
rect 364524 271176 364576 271182
rect 364524 271118 364576 271124
rect 364156 270224 364208 270230
rect 364156 270166 364208 270172
rect 363354 264302 363828 264330
rect 364168 264316 364196 270166
rect 364996 267306 365024 274178
rect 366100 273086 366128 278052
rect 367112 278038 367310 278066
rect 366364 273216 366416 273222
rect 366364 273158 366416 273164
rect 366088 273080 366140 273086
rect 366088 273022 366140 273028
rect 365444 271312 365496 271318
rect 365444 271254 365496 271260
rect 364984 267300 365036 267306
rect 364984 267242 365036 267248
rect 365456 264330 365484 271254
rect 365812 267164 365864 267170
rect 365812 267106 365864 267112
rect 365010 264302 365484 264330
rect 365824 264316 365852 267106
rect 366376 266762 366404 273158
rect 366916 271176 366968 271182
rect 366916 271118 366968 271124
rect 366364 266756 366416 266762
rect 366364 266698 366416 266704
rect 366928 264330 366956 271118
rect 367112 268394 367140 278038
rect 368492 274106 368520 278052
rect 369596 274514 369624 278052
rect 369584 274508 369636 274514
rect 369584 274450 369636 274456
rect 369308 274372 369360 274378
rect 369308 274314 369360 274320
rect 368480 274100 368532 274106
rect 368480 274042 368532 274048
rect 369124 274100 369176 274106
rect 369124 274042 369176 274048
rect 367468 270360 367520 270366
rect 367468 270302 367520 270308
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 366666 264302 366956 264330
rect 367480 264316 367508 270302
rect 369136 267578 369164 274042
rect 369124 267572 369176 267578
rect 369124 267514 369176 267520
rect 369124 266552 369176 266558
rect 369124 266494 369176 266500
rect 368296 266416 368348 266422
rect 368296 266358 368348 266364
rect 368308 264316 368336 266358
rect 369136 264316 369164 266494
rect 369320 266422 369348 274314
rect 370792 272814 370820 278052
rect 371252 278038 372002 278066
rect 372816 278038 373198 278066
rect 370780 272808 370832 272814
rect 370780 272750 370832 272756
rect 369952 270088 370004 270094
rect 369952 270030 370004 270036
rect 369964 266558 369992 270030
rect 371252 269958 371280 278038
rect 372816 271726 372844 278038
rect 373264 274372 373316 274378
rect 373264 274314 373316 274320
rect 372804 271720 372856 271726
rect 372804 271662 372856 271668
rect 371240 269952 371292 269958
rect 371240 269894 371292 269900
rect 372436 269952 372488 269958
rect 372436 269894 372488 269900
rect 372160 268388 372212 268394
rect 372160 268330 372212 268336
rect 370780 267572 370832 267578
rect 370780 267514 370832 267520
rect 369952 266552 370004 266558
rect 369952 266494 370004 266500
rect 369308 266416 369360 266422
rect 369308 266358 369360 266364
rect 369952 266416 370004 266422
rect 369952 266358 370004 266364
rect 369964 264316 369992 266358
rect 370792 264316 370820 267514
rect 371608 267436 371660 267442
rect 371608 267378 371660 267384
rect 371620 264316 371648 267378
rect 372172 266422 372200 268330
rect 372160 266416 372212 266422
rect 372160 266358 372212 266364
rect 372448 264316 372476 269894
rect 373276 267442 373304 274314
rect 374380 274242 374408 278052
rect 374368 274236 374420 274242
rect 374368 274178 374420 274184
rect 374644 273352 374696 273358
rect 374644 273294 374696 273300
rect 373264 267436 373316 267442
rect 373264 267378 373316 267384
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373276 264316 373304 267242
rect 374656 267034 374684 273294
rect 375196 272808 375248 272814
rect 375196 272750 375248 272756
rect 374644 267028 374696 267034
rect 374644 266970 374696 266976
rect 374920 266552 374972 266558
rect 374920 266494 374972 266500
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 266494
rect 375208 266422 375236 272750
rect 375576 272678 375604 278052
rect 376786 278038 376984 278066
rect 375564 272672 375616 272678
rect 375564 272614 375616 272620
rect 376576 271856 376628 271862
rect 376576 271798 376628 271804
rect 375748 267028 375800 267034
rect 375748 266970 375800 266976
rect 375196 266416 375248 266422
rect 375196 266358 375248 266364
rect 375760 264316 375788 266970
rect 376588 264316 376616 271798
rect 376956 269822 376984 278038
rect 377876 273358 377904 278052
rect 377864 273352 377916 273358
rect 377864 273294 377916 273300
rect 377404 273080 377456 273086
rect 377404 273022 377456 273028
rect 376944 269816 376996 269822
rect 376944 269758 376996 269764
rect 377416 267578 377444 273022
rect 379072 271590 379100 278052
rect 379532 278038 380282 278066
rect 379336 274236 379388 274242
rect 379336 274178 379388 274184
rect 379060 271584 379112 271590
rect 379060 271526 379112 271532
rect 377680 269816 377732 269822
rect 377680 269758 377732 269764
rect 377404 267572 377456 267578
rect 377404 267514 377456 267520
rect 377692 264330 377720 269758
rect 378232 267708 378284 267714
rect 378232 267650 378284 267656
rect 377430 264302 377720 264330
rect 378244 264316 378272 267650
rect 379348 264330 379376 274178
rect 379532 268530 379560 278038
rect 381464 271454 381492 278052
rect 382660 273970 382688 278052
rect 382924 274644 382976 274650
rect 382924 274586 382976 274592
rect 382648 273964 382700 273970
rect 382648 273906 382700 273912
rect 382004 272672 382056 272678
rect 382004 272614 382056 272620
rect 381452 271448 381504 271454
rect 381452 271390 381504 271396
rect 381544 271040 381596 271046
rect 381544 270982 381596 270988
rect 379704 269068 379756 269074
rect 379704 269010 379756 269016
rect 379520 268524 379572 268530
rect 379520 268466 379572 268472
rect 379716 266558 379744 269010
rect 380716 267572 380768 267578
rect 380716 267514 380768 267520
rect 379704 266552 379756 266558
rect 379704 266494 379756 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379376 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267514
rect 381556 266422 381584 270982
rect 381544 266416 381596 266422
rect 381544 266358 381596 266364
rect 382016 264330 382044 272614
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 382936 267170 382964 274586
rect 383856 273222 383884 278052
rect 385052 275330 385080 278052
rect 385880 278038 386170 278066
rect 385040 275324 385092 275330
rect 385040 275266 385092 275272
rect 383844 273216 383896 273222
rect 383844 273158 383896 273164
rect 385880 272950 385908 278038
rect 386052 275460 386104 275466
rect 386052 275402 386104 275408
rect 385868 272944 385920 272950
rect 385868 272886 385920 272892
rect 384948 271720 385000 271726
rect 384948 271662 385000 271668
rect 384764 269680 384816 269686
rect 384764 269622 384816 269628
rect 383200 267436 383252 267442
rect 383200 267378 383252 267384
rect 382924 267164 382976 267170
rect 382924 267106 382976 267112
rect 383212 264316 383240 267378
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 269622
rect 384960 266422 384988 271662
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 386064 264330 386092 275402
rect 387352 274106 387380 278052
rect 387340 274100 387392 274106
rect 387340 274042 387392 274048
rect 387432 273964 387484 273970
rect 387432 273906 387484 273912
rect 387444 266422 387472 273906
rect 388548 272542 388576 278052
rect 389192 278038 389758 278066
rect 388536 272536 388588 272542
rect 388536 272478 388588 272484
rect 388996 272400 389048 272406
rect 388996 272342 389048 272348
rect 387616 271584 387668 271590
rect 387616 271526 387668 271532
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 387432 266416 387484 266422
rect 387432 266358 387484 266364
rect 384776 264302 384882 264330
rect 385710 264302 386092 264330
rect 386524 264316 386552 266358
rect 387628 264330 387656 271526
rect 388168 266756 388220 266762
rect 388168 266698 388220 266704
rect 387366 264302 387656 264330
rect 388180 264316 388208 266698
rect 389008 264316 389036 272342
rect 389192 270230 389220 278038
rect 390940 271318 390968 278052
rect 392136 274650 392164 278052
rect 392124 274644 392176 274650
rect 392124 274586 392176 274592
rect 392584 273692 392636 273698
rect 392584 273634 392636 273640
rect 390928 271312 390980 271318
rect 390928 271254 390980 271260
rect 391848 271312 391900 271318
rect 391848 271254 391900 271260
rect 389180 270224 389232 270230
rect 389180 270166 389232 270172
rect 390100 270224 390152 270230
rect 390100 270166 390152 270172
rect 389824 268796 389876 268802
rect 389824 268738 389876 268744
rect 389836 264316 389864 268738
rect 390112 267034 390140 270166
rect 390652 267164 390704 267170
rect 390652 267106 390704 267112
rect 390100 267028 390152 267034
rect 390100 266970 390152 266976
rect 390664 264316 390692 267106
rect 391860 264330 391888 271254
rect 392032 269544 392084 269550
rect 392032 269486 392084 269492
rect 392044 267306 392072 269486
rect 392596 267714 392624 273634
rect 393332 271182 393360 278052
rect 393516 278038 394450 278066
rect 393320 271176 393372 271182
rect 393320 271118 393372 271124
rect 393516 270366 393544 278038
rect 395632 274514 395660 278052
rect 396092 278038 396842 278066
rect 397472 278038 398038 278066
rect 395620 274508 395672 274514
rect 395620 274450 395672 274456
rect 394332 274100 394384 274106
rect 394332 274042 394384 274048
rect 393964 271448 394016 271454
rect 393964 271390 394016 271396
rect 393504 270360 393556 270366
rect 393504 270302 393556 270308
rect 392584 267708 392636 267714
rect 392584 267650 392636 267656
rect 392032 267300 392084 267306
rect 392032 267242 392084 267248
rect 393136 267028 393188 267034
rect 393136 266970 393188 266976
rect 392308 266892 392360 266898
rect 392308 266834 392360 266840
rect 391506 264302 391888 264330
rect 392320 264316 392348 266834
rect 393148 264316 393176 266970
rect 393976 266898 394004 271390
rect 393964 266892 394016 266898
rect 393964 266834 394016 266840
rect 394344 264330 394372 274042
rect 395620 270496 395672 270502
rect 395620 270438 395672 270444
rect 394792 266416 394844 266422
rect 394792 266358 394844 266364
rect 393990 264302 394372 264330
rect 394804 264316 394832 266358
rect 395632 264316 395660 270438
rect 396092 270094 396120 278038
rect 397276 272536 397328 272542
rect 397276 272478 397328 272484
rect 396080 270088 396132 270094
rect 396080 270030 396132 270036
rect 396172 268660 396224 268666
rect 396172 268602 396224 268608
rect 396184 266422 396212 268602
rect 397092 266756 397144 266762
rect 397092 266698 397144 266704
rect 396172 266416 396224 266422
rect 396172 266358 396224 266364
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 396460 264316 396488 266358
rect 397104 264330 397132 266698
rect 397288 266422 397316 272478
rect 397472 268394 397500 278038
rect 399220 273086 399248 278052
rect 400324 274378 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274372 400364 274378
rect 400312 274314 400364 274320
rect 400128 273828 400180 273834
rect 400128 273770 400180 273776
rect 399208 273080 399260 273086
rect 399208 273022 399260 273028
rect 399944 270088 399996 270094
rect 399944 270030 399996 270036
rect 397460 268388 397512 268394
rect 397460 268330 397512 268336
rect 398104 267708 398156 267714
rect 398104 267650 398156 267656
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 267650
rect 399956 267578 399984 270030
rect 399944 267572 399996 267578
rect 399944 267514 399996 267520
rect 400140 266422 400168 273770
rect 400508 269958 400536 278038
rect 401508 273216 401560 273222
rect 401508 273158 401560 273164
rect 400864 270360 400916 270366
rect 400864 270302 400916 270308
rect 400496 269952 400548 269958
rect 400496 269894 400548 269900
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 398944 264316 398972 266358
rect 400128 266280 400180 266286
rect 400128 266222 400180 266228
rect 400140 264330 400168 266222
rect 400876 264330 400904 270302
rect 401520 267734 401548 273158
rect 401704 269550 401732 278038
rect 403912 272814 403940 278052
rect 404372 278038 405122 278066
rect 405752 278038 406318 278066
rect 404176 274644 404228 274650
rect 404176 274586 404228 274592
rect 403900 272808 403952 272814
rect 403900 272750 403952 272756
rect 402612 271176 402664 271182
rect 402612 271118 402664 271124
rect 401876 269952 401928 269958
rect 401876 269894 401928 269900
rect 401692 269544 401744 269550
rect 401692 269486 401744 269492
rect 399786 264302 400168 264330
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401888 267442 401916 269894
rect 401876 267436 401928 267442
rect 401876 267378 401928 267384
rect 402624 264330 402652 271118
rect 403256 268524 403308 268530
rect 403256 268466 403308 268472
rect 403072 267300 403124 267306
rect 403072 267242 403124 267248
rect 402270 264302 402652 264330
rect 403084 264316 403112 267242
rect 403268 266422 403296 268466
rect 403256 266416 403308 266422
rect 403256 266358 403308 266364
rect 404188 264330 404216 274586
rect 404372 269074 404400 278038
rect 405752 270230 405780 278038
rect 406844 272944 406896 272950
rect 406844 272886 406896 272892
rect 405740 270224 405792 270230
rect 405740 270166 405792 270172
rect 404544 269544 404596 269550
rect 404544 269486 404596 269492
rect 404360 269068 404412 269074
rect 404360 269010 404412 269016
rect 404556 266626 404584 269486
rect 405556 267436 405608 267442
rect 405556 267378 405608 267384
rect 404544 266620 404596 266626
rect 404544 266562 404596 266568
rect 404728 266620 404780 266626
rect 404728 266562 404780 266568
rect 403926 264302 404216 264330
rect 404740 264316 404768 266562
rect 405568 264316 405596 267378
rect 406856 264330 406884 272886
rect 407500 271862 407528 278052
rect 408512 278038 408618 278066
rect 408224 273080 408276 273086
rect 408224 273022 408276 273028
rect 407488 271856 407540 271862
rect 407488 271798 407540 271804
rect 407764 271856 407816 271862
rect 407764 271798 407816 271804
rect 407776 266762 407804 271798
rect 408040 268388 408092 268394
rect 408040 268330 408092 268336
rect 407764 266756 407816 266762
rect 407764 266698 407816 266704
rect 407212 266416 407264 266422
rect 407212 266358 407264 266364
rect 406410 264302 406884 264330
rect 407224 264316 407252 266358
rect 408052 264316 408080 268330
rect 408236 266422 408264 273022
rect 408512 269822 408540 278038
rect 409236 274508 409288 274514
rect 409236 274450 409288 274456
rect 408500 269816 408552 269822
rect 408500 269758 408552 269764
rect 408224 266416 408276 266422
rect 408224 266358 408276 266364
rect 409248 264330 409276 274450
rect 409800 273698 409828 278052
rect 410996 274242 411024 278052
rect 411824 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 274236 411036 274242
rect 410984 274178 411036 274184
rect 409788 273692 409840 273698
rect 409788 273634 409840 273640
rect 411824 271046 411852 278038
rect 412272 272808 412324 272814
rect 412272 272750 412324 272756
rect 411812 271040 411864 271046
rect 411812 270982 411864 270988
rect 409696 270224 409748 270230
rect 409696 270166 409748 270172
rect 408894 264302 409276 264330
rect 409708 264316 409736 270166
rect 410524 267572 410576 267578
rect 410524 267514 410576 267520
rect 410536 264316 410564 267514
rect 412284 266422 412312 272750
rect 412652 270094 412680 278038
rect 413468 274916 413520 274922
rect 413468 274858 413520 274864
rect 412640 270088 412692 270094
rect 412640 270030 412692 270036
rect 412456 269816 412508 269822
rect 412456 269758 412508 269764
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 411364 264316 411392 266358
rect 412468 264330 412496 269758
rect 412640 268116 412692 268122
rect 412640 268058 412692 268064
rect 412652 266626 412680 268058
rect 412640 266620 412692 266626
rect 412640 266562 412692 266568
rect 413480 264330 413508 274858
rect 413836 274372 413888 274378
rect 413836 274314 413888 274320
rect 412206 264302 412496 264330
rect 413034 264302 413508 264330
rect 413848 264316 413876 274314
rect 414584 272678 414612 278052
rect 415412 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 272672 414624 272678
rect 414572 272614 414624 272620
rect 414480 271040 414532 271046
rect 414480 270982 414532 270988
rect 414492 267714 414520 270982
rect 414664 270088 414716 270094
rect 414664 270030 414716 270036
rect 414480 267708 414532 267714
rect 414480 267650 414532 267656
rect 414676 264316 414704 270030
rect 415412 268938 415440 278038
rect 416412 275324 416464 275330
rect 416412 275266 416464 275272
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 416424 266422 416452 275266
rect 416596 274236 416648 274242
rect 416596 274178 416648 274184
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 415504 264316 415532 266358
rect 416608 264330 416636 274178
rect 416792 269958 416820 278038
rect 418080 271726 418108 278052
rect 418264 278038 419290 278066
rect 418068 271720 418120 271726
rect 418068 271662 418120 271668
rect 417424 270904 417476 270910
rect 417424 270846 417476 270852
rect 416780 269952 416832 269958
rect 416780 269894 416832 269900
rect 417148 269952 417200 269958
rect 417148 269894 417200 269900
rect 416346 264302 416636 264330
rect 417160 264316 417188 269894
rect 417436 267170 417464 270846
rect 418264 269686 418292 278038
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420644 275052 420696 275058
rect 420644 274994 420696 275000
rect 419172 272672 419224 272678
rect 419172 272614 419224 272620
rect 418252 269680 418304 269686
rect 418252 269622 418304 269628
rect 417424 267164 417476 267170
rect 417424 267106 417476 267112
rect 417976 267164 418028 267170
rect 417976 267106 418028 267112
rect 417988 264316 418016 267106
rect 419184 264330 419212 272614
rect 420184 271720 420236 271726
rect 420184 271662 420236 271668
rect 419632 268252 419684 268258
rect 419632 268194 419684 268200
rect 418830 264302 419212 264330
rect 419644 264316 419672 268194
rect 420196 267034 420224 271662
rect 420184 267028 420236 267034
rect 420184 266970 420236 266976
rect 420656 264330 420684 274994
rect 421668 273970 421696 278052
rect 421656 273964 421708 273970
rect 421656 273906 421708 273912
rect 421840 273964 421892 273970
rect 421840 273906 421892 273912
rect 421852 267734 421880 273906
rect 422864 271590 422892 278052
rect 423692 278038 423982 278066
rect 423404 275460 423456 275466
rect 423404 275402 423456 275408
rect 422852 271584 422904 271590
rect 422852 271526 422904 271532
rect 422944 270632 422996 270638
rect 422944 270574 422996 270580
rect 422116 269680 422168 269686
rect 422116 269622 422168 269628
rect 421760 267706 421880 267734
rect 421760 264330 421788 267706
rect 420486 264302 420684 264330
rect 421314 264302 421788 264330
rect 422128 264316 422156 269622
rect 422956 267306 422984 270574
rect 422944 267300 422996 267306
rect 422944 267242 422996 267248
rect 423416 264330 423444 275402
rect 423692 269550 423720 278038
rect 425164 272406 425192 278052
rect 425348 278038 426374 278066
rect 425152 272400 425204 272406
rect 425152 272342 425204 272348
rect 423680 269544 423732 269550
rect 423680 269486 423732 269492
rect 423956 269272 424008 269278
rect 423956 269214 424008 269220
rect 423772 267708 423824 267714
rect 423772 267650 423824 267656
rect 422970 264302 423444 264330
rect 423784 264316 423812 267650
rect 423968 267442 423996 269214
rect 425348 268802 425376 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426348 272128 426400 272134
rect 426348 272070 426400 272076
rect 425336 268796 425388 268802
rect 425336 268738 425388 268744
rect 426360 267734 426388 272070
rect 426268 267706 426388 267734
rect 423956 267436 424008 267442
rect 423956 267378 424008 267384
rect 424600 267300 424652 267306
rect 424600 267242 424652 267248
rect 424612 264316 424640 267242
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 267706
rect 427096 266422 427124 275130
rect 427556 270910 427584 278052
rect 428752 271318 428780 278052
rect 429948 271454 429976 278052
rect 430212 275596 430264 275602
rect 430212 275538 430264 275544
rect 429936 271448 429988 271454
rect 429936 271390 429988 271396
rect 428740 271312 428792 271318
rect 428740 271254 428792 271260
rect 427544 270904 427596 270910
rect 427544 270846 427596 270852
rect 427452 270768 427504 270774
rect 427452 270710 427504 270716
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270710
rect 429108 269408 429160 269414
rect 429108 269350 429160 269356
rect 429120 267578 429148 269350
rect 429108 267572 429160 267578
rect 429108 267514 429160 267520
rect 427912 266892 427964 266898
rect 427912 266834 427964 266840
rect 427110 264302 427492 264330
rect 427924 264316 427952 266834
rect 428740 266756 428792 266762
rect 428740 266698 428792 266704
rect 428752 264316 428780 266698
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275538
rect 431144 271726 431172 278052
rect 432248 274106 432276 278052
rect 433444 277394 433472 278052
rect 433352 277366 433472 277394
rect 433628 278038 434654 278066
rect 432236 274100 432288 274106
rect 432236 274042 432288 274048
rect 432604 274100 432656 274106
rect 432604 274042 432656 274048
rect 431132 271720 431184 271726
rect 431132 271662 431184 271668
rect 430396 270904 430448 270910
rect 430396 270846 430448 270852
rect 430408 266422 430436 270846
rect 432236 269544 432288 269550
rect 432236 269486 432288 269492
rect 432052 267436 432104 267442
rect 432052 267378 432104 267384
rect 431224 267028 431276 267034
rect 431224 266970 431276 266976
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 430224 264302 430422 264330
rect 431236 264316 431264 266970
rect 432064 264316 432092 267378
rect 432248 267170 432276 269486
rect 432236 267164 432288 267170
rect 432236 267106 432288 267112
rect 432616 267034 432644 274042
rect 433352 268666 433380 277366
rect 433628 270502 433656 278038
rect 435640 275732 435692 275738
rect 435640 275674 435692 275680
rect 434628 271720 434680 271726
rect 434628 271662 434680 271668
rect 433616 270496 433668 270502
rect 433616 270438 433668 270444
rect 433708 268932 433760 268938
rect 433708 268874 433760 268880
rect 433340 268660 433392 268666
rect 433340 268602 433392 268608
rect 432880 267164 432932 267170
rect 432880 267106 432932 267112
rect 432604 267028 432656 267034
rect 432604 266970 432656 266976
rect 432892 264316 432920 267106
rect 433720 264316 433748 268874
rect 434640 267734 434668 271662
rect 434548 267706 434668 267734
rect 434548 264316 434576 267706
rect 435652 264330 435680 275674
rect 435836 272542 435864 278052
rect 435824 272536 435876 272542
rect 435824 272478 435876 272484
rect 437032 271862 437060 278052
rect 438136 278038 438242 278066
rect 437020 271856 437072 271862
rect 437020 271798 437072 271804
rect 437204 271856 437256 271862
rect 437204 271798 437256 271804
rect 436192 269068 436244 269074
rect 436192 269010 436244 269016
rect 435390 264302 435680 264330
rect 436204 264316 436232 269010
rect 437216 264330 437244 271798
rect 438136 271046 438164 278038
rect 439332 273834 439360 278052
rect 440252 278038 440542 278066
rect 439320 273828 439372 273834
rect 439320 273770 439372 273776
rect 438768 272536 438820 272542
rect 438768 272478 438820 272484
rect 438124 271040 438176 271046
rect 438124 270982 438176 270988
rect 438308 271040 438360 271046
rect 438308 270982 438360 270988
rect 438320 264330 438348 270982
rect 438780 267734 438808 272478
rect 439964 271584 440016 271590
rect 439964 271526 440016 271532
rect 437046 264302 437244 264330
rect 437874 264302 438348 264330
rect 438688 267706 438808 267734
rect 438688 264316 438716 267706
rect 439976 264330 440004 271526
rect 440252 268530 440280 278038
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273692 440936 273698
rect 440884 273634 440936 273640
rect 440240 268524 440292 268530
rect 440240 268466 440292 268472
rect 440896 267714 440924 273634
rect 441632 270366 441660 277366
rect 442264 273828 442316 273834
rect 442264 273770 442316 273776
rect 441620 270360 441672 270366
rect 441620 270302 441672 270308
rect 441160 268796 441212 268802
rect 441160 268738 441212 268744
rect 440884 267708 440936 267714
rect 440884 267650 440936 267656
rect 440332 266620 440384 266626
rect 440332 266562 440384 266568
rect 439530 264302 440004 264330
rect 440344 264316 440372 266562
rect 441172 264316 441200 268738
rect 442276 266762 442304 273770
rect 442920 273222 442948 278052
rect 442908 273216 442960 273222
rect 442908 273158 442960 273164
rect 442908 271448 442960 271454
rect 442908 271390 442960 271396
rect 442724 266892 442776 266898
rect 442724 266834 442776 266840
rect 442264 266756 442316 266762
rect 442264 266698 442316 266704
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 266834
rect 442920 266422 442948 271390
rect 444116 271182 444144 278052
rect 445024 275868 445076 275874
rect 445024 275810 445076 275816
rect 444104 271176 444156 271182
rect 444104 271118 444156 271124
rect 443644 268660 443696 268666
rect 443644 268602 443696 268608
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 442736 264302 442842 264330
rect 443656 264316 443684 268602
rect 445036 266626 445064 275810
rect 445312 270638 445340 278052
rect 446508 274650 446536 278052
rect 447152 278038 447626 278066
rect 448532 278038 448822 278066
rect 446496 274644 446548 274650
rect 446496 274586 446548 274592
rect 446404 273556 446456 273562
rect 446404 273498 446456 273504
rect 445668 271312 445720 271318
rect 445668 271254 445720 271260
rect 445300 270632 445352 270638
rect 445300 270574 445352 270580
rect 445300 267572 445352 267578
rect 445300 267514 445352 267520
rect 445024 266620 445076 266626
rect 445024 266562 445076 266568
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 444484 264316 444512 266358
rect 445312 264316 445340 267514
rect 445680 266422 445708 271254
rect 446416 267306 446444 273498
rect 446956 272264 447008 272270
rect 446956 272206 447008 272212
rect 446404 267300 446456 267306
rect 446404 267242 446456 267248
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446128 266416 446180 266422
rect 446128 266358 446180 266364
rect 446140 264316 446168 266358
rect 446968 264316 446996 272206
rect 447152 268122 447180 278038
rect 447784 271992 447836 271998
rect 447784 271934 447836 271940
rect 447140 268116 447192 268122
rect 447140 268058 447192 268064
rect 447796 266422 447824 271934
rect 448532 269278 448560 278038
rect 450004 272950 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 450544 274644 450596 274650
rect 450544 274586 450596 274592
rect 449992 272944 450044 272950
rect 449992 272886 450044 272892
rect 449716 272400 449768 272406
rect 449716 272342 449768 272348
rect 448520 269272 448572 269278
rect 448520 269214 448572 269220
rect 448612 268524 448664 268530
rect 448612 268466 448664 268472
rect 448152 267300 448204 267306
rect 448152 267242 448204 267248
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 448164 264330 448192 267242
rect 447810 264302 448192 264330
rect 448624 264316 448652 268466
rect 449728 264330 449756 272342
rect 450268 267708 450320 267714
rect 450268 267650 450320 267656
rect 449466 264302 449756 264330
rect 450280 264316 450308 267650
rect 450556 267034 450584 274586
rect 450832 273086 450860 278038
rect 450820 273080 450872 273086
rect 450820 273022 450872 273028
rect 451188 273080 451240 273086
rect 451188 273022 451240 273028
rect 451200 267734 451228 273022
rect 451384 268394 451412 278038
rect 453592 274514 453620 278052
rect 454052 278038 454710 278066
rect 455432 278038 455906 278066
rect 453580 274508 453632 274514
rect 453580 274450 453632 274456
rect 453764 274508 453816 274514
rect 453764 274450 453816 274456
rect 453776 273358 453804 274450
rect 453304 273352 453356 273358
rect 453304 273294 453356 273300
rect 453764 273352 453816 273358
rect 453764 273294 453816 273300
rect 452292 273216 452344 273222
rect 452292 273158 452344 273164
rect 451372 268388 451424 268394
rect 451372 268330 451424 268336
rect 451108 267706 451228 267734
rect 450544 267028 450596 267034
rect 450544 266970 450596 266976
rect 451108 264316 451136 267706
rect 452304 264330 452332 273158
rect 453316 267442 453344 273294
rect 453580 270496 453632 270502
rect 453580 270438 453632 270444
rect 453304 267436 453356 267442
rect 453304 267378 453356 267384
rect 452752 266620 452804 266626
rect 452752 266562 452804 266568
rect 451950 264302 452332 264330
rect 452764 264316 452792 266562
rect 453592 264316 453620 270438
rect 454052 270230 454080 278038
rect 454408 276004 454460 276010
rect 454408 275946 454460 275952
rect 454420 275738 454448 275946
rect 454408 275732 454460 275738
rect 454408 275674 454460 275680
rect 455236 272944 455288 272950
rect 455236 272886 455288 272892
rect 454040 270224 454092 270230
rect 454040 270166 454092 270172
rect 455052 267028 455104 267034
rect 455052 266970 455104 266976
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455064 264330 455092 266970
rect 455248 266422 455276 272886
rect 455432 269414 455460 278038
rect 457088 272814 457116 278052
rect 457444 276004 457496 276010
rect 457444 275946 457496 275952
rect 457076 272808 457128 272814
rect 457076 272750 457128 272756
rect 456064 270360 456116 270366
rect 456064 270302 456116 270308
rect 455420 269408 455472 269414
rect 455420 269350 455472 269356
rect 455236 266416 455288 266422
rect 455236 266358 455288 266364
rect 455064 264302 455262 264330
rect 456076 264316 456104 270302
rect 457456 267306 457484 275946
rect 458088 272944 458140 272950
rect 458088 272886 458140 272892
rect 457444 267300 457496 267306
rect 457444 267242 457496 267248
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456904 264316 456932 266358
rect 457732 264316 457760 266698
rect 458100 266422 458128 272886
rect 458284 269822 458312 278052
rect 459480 274922 459508 278052
rect 459468 274916 459520 274922
rect 459468 274858 459520 274864
rect 460676 274378 460704 278052
rect 460952 278038 461886 278066
rect 460664 274372 460716 274378
rect 460664 274314 460716 274320
rect 460020 273420 460072 273426
rect 460020 273362 460072 273368
rect 459468 271176 459520 271182
rect 459468 271118 459520 271124
rect 458548 270224 458600 270230
rect 458548 270166 458600 270172
rect 458272 269816 458324 269822
rect 458272 269758 458324 269764
rect 458088 266416 458140 266422
rect 458088 266358 458140 266364
rect 458560 264316 458588 270166
rect 459480 267734 459508 271118
rect 459388 267706 459508 267734
rect 459388 264316 459416 267706
rect 460032 267170 460060 273362
rect 460952 270094 460980 278038
rect 462976 275330 463004 278052
rect 462964 275324 463016 275330
rect 462964 275266 463016 275272
rect 463148 275324 463200 275330
rect 463148 275266 463200 275272
rect 462226 272368 462282 272377
rect 462226 272303 462282 272312
rect 460940 270088 460992 270094
rect 460940 270030 460992 270036
rect 461400 270088 461452 270094
rect 461400 270030 461452 270036
rect 460204 267436 460256 267442
rect 460204 267378 460256 267384
rect 460020 267164 460072 267170
rect 460020 267106 460072 267112
rect 460216 264316 460244 267378
rect 461412 264330 461440 270030
rect 462240 264330 462268 272303
rect 463160 264330 463188 275266
rect 464172 274242 464200 278052
rect 465092 278038 465382 278066
rect 464160 274236 464212 274242
rect 464160 274178 464212 274184
rect 463332 272944 463384 272950
rect 463384 272892 463924 272898
rect 463332 272886 463924 272892
rect 463344 272870 463924 272886
rect 463896 272814 463924 272870
rect 463884 272808 463936 272814
rect 463884 272750 463936 272756
rect 465092 269958 465120 278038
rect 466564 277394 466592 278052
rect 466472 277366 466592 277394
rect 467392 278038 467774 278066
rect 467944 278038 468970 278066
rect 465724 274372 465776 274378
rect 465724 274314 465776 274320
rect 465736 273426 465764 274314
rect 465724 273420 465776 273426
rect 465724 273362 465776 273368
rect 465080 269952 465132 269958
rect 465080 269894 465132 269900
rect 463516 269816 463568 269822
rect 463516 269758 463568 269764
rect 461058 264302 461440 264330
rect 461886 264302 462268 264330
rect 462714 264302 463188 264330
rect 463528 264316 463556 269758
rect 466472 269550 466500 277366
rect 467392 272678 467420 278038
rect 467564 273420 467616 273426
rect 467564 273362 467616 273368
rect 467380 272672 467432 272678
rect 467380 272614 467432 272620
rect 466460 269544 466512 269550
rect 466460 269486 466512 269492
rect 466000 269408 466052 269414
rect 466000 269350 466052 269356
rect 464344 268388 464396 268394
rect 464344 268330 464396 268336
rect 464356 264316 464384 268330
rect 465172 267164 465224 267170
rect 465172 267106 465224 267112
rect 465184 264316 465212 267106
rect 466012 264316 466040 269350
rect 466828 266416 466880 266422
rect 466828 266358 466880 266364
rect 466840 264316 466868 266358
rect 467576 264330 467604 273362
rect 467748 272672 467800 272678
rect 467748 272614 467800 272620
rect 467760 266422 467788 272614
rect 467944 268258 467972 278038
rect 470152 275058 470180 278052
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 469864 274780 469916 274786
rect 469864 274722 469916 274728
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467932 268252 467984 268258
rect 467932 268194 467984 268200
rect 467748 266416 467800 266422
rect 467748 266358 467800 266364
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 469876 266626 469904 274722
rect 471256 273970 471284 278052
rect 471992 278038 472466 278066
rect 473372 278038 473662 278066
rect 471612 276276 471664 276282
rect 471612 276218 471664 276224
rect 471244 273964 471296 273970
rect 471244 273906 471296 273912
rect 470416 272672 470468 272678
rect 470414 272640 470416 272649
rect 470600 272672 470652 272678
rect 470468 272640 470470 272649
rect 470414 272575 470470 272584
rect 470598 272640 470600 272649
rect 470652 272640 470654 272649
rect 470598 272575 470654 272584
rect 470428 272462 470824 272490
rect 470428 272377 470456 272462
rect 470414 272368 470470 272377
rect 470414 272303 470470 272312
rect 470796 272134 470824 272462
rect 470554 272128 470606 272134
rect 470784 272128 470836 272134
rect 470606 272076 470640 272082
rect 470554 272070 470640 272076
rect 470784 272070 470836 272076
rect 470566 272054 470640 272070
rect 470612 271969 470640 272054
rect 470598 271960 470654 271969
rect 470598 271895 470654 271904
rect 470968 269272 471020 269278
rect 470968 269214 471020 269220
rect 470140 267300 470192 267306
rect 470140 267242 470192 267248
rect 469864 266620 469916 266626
rect 469864 266562 469916 266568
rect 469312 265124 469364 265130
rect 469312 265066 469364 265072
rect 469324 264316 469352 265066
rect 470152 264316 470180 267242
rect 470980 264316 471008 269214
rect 471624 264330 471652 276218
rect 471992 269686 472020 278038
rect 473372 275466 473400 278038
rect 473360 275460 473412 275466
rect 473360 275402 473412 275408
rect 473360 274916 473412 274922
rect 473360 274858 473412 274864
rect 473372 269686 473400 274858
rect 474372 274236 474424 274242
rect 474372 274178 474424 274184
rect 471980 269680 472032 269686
rect 471980 269622 472032 269628
rect 472624 269680 472676 269686
rect 472624 269622 472676 269628
rect 473360 269680 473412 269686
rect 473360 269622 473412 269628
rect 471624 264302 471822 264330
rect 472636 264316 472664 269622
rect 474384 266422 474412 274178
rect 474844 273698 474872 278052
rect 476040 277394 476068 278052
rect 475948 277366 476068 277394
rect 475384 275868 475436 275874
rect 475384 275810 475436 275816
rect 475396 275466 475424 275810
rect 475384 275460 475436 275466
rect 475384 275402 475436 275408
rect 475752 273964 475804 273970
rect 475752 273906 475804 273912
rect 474832 273692 474884 273698
rect 474832 273634 474884 273640
rect 474648 269408 474700 269414
rect 474648 269350 474700 269356
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 474372 266416 474424 266422
rect 474372 266358 474424 266364
rect 473464 264316 473492 266358
rect 474660 264330 474688 269350
rect 475108 265260 475160 265266
rect 475108 265202 475160 265208
rect 474306 264302 474688 264330
rect 475120 264316 475148 265202
rect 475764 264330 475792 273906
rect 475948 273562 475976 277366
rect 477040 276412 477092 276418
rect 477040 276354 477092 276360
rect 476120 275052 476172 275058
rect 476120 274994 476172 275000
rect 475936 273556 475988 273562
rect 475936 273498 475988 273504
rect 476132 273426 476160 274994
rect 476120 273420 476172 273426
rect 476120 273362 476172 273368
rect 477052 264330 477080 276354
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 478064 271969 478092 278038
rect 478512 276548 478564 276554
rect 478512 276490 478564 276496
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 478524 266422 478552 276490
rect 478696 273420 478748 273426
rect 478696 273362 478748 273368
rect 477592 266416 477644 266422
rect 477592 266358 477644 266364
rect 478512 266416 478564 266422
rect 478512 266358 478564 266364
rect 475764 264302 475962 264330
rect 476790 264302 477080 264330
rect 477604 264316 477632 266358
rect 478708 264330 478736 273362
rect 479168 270774 479196 278038
rect 479524 275868 479576 275874
rect 479524 275810 479576 275816
rect 479156 270768 479208 270774
rect 479156 270710 479208 270716
rect 479536 266762 479564 275810
rect 480732 274650 480760 278052
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481928 273834 481956 278052
rect 482836 277364 482888 277370
rect 482836 277306 482888 277312
rect 481916 273828 481968 273834
rect 481916 273770 481968 273776
rect 481364 273556 481416 273562
rect 481364 273498 481416 273504
rect 479524 266756 479576 266762
rect 479524 266698 479576 266704
rect 480076 265532 480128 265538
rect 480076 265474 480128 265480
rect 479248 265396 479300 265402
rect 479248 265338 479300 265344
rect 478446 264302 478736 264330
rect 479260 264316 479288 265338
rect 480088 264316 480116 265474
rect 481376 264330 481404 273498
rect 482560 266552 482612 266558
rect 482560 266494 482612 266500
rect 481732 266416 481784 266422
rect 481732 266358 481784 266364
rect 480930 264302 481404 264330
rect 481744 264316 481772 266358
rect 482572 264316 482600 266494
rect 482848 266422 482876 277306
rect 483124 270910 483152 278052
rect 484320 275602 484348 278052
rect 484308 275596 484360 275602
rect 484308 275538 484360 275544
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 485228 275460 485280 275466
rect 485228 275402 485280 275408
rect 485056 275194 485084 275402
rect 485044 275188 485096 275194
rect 485044 275130 485096 275136
rect 485240 275058 485268 275402
rect 485228 275052 485280 275058
rect 485228 274994 485280 275000
rect 485516 274106 485544 278052
rect 485688 277228 485740 277234
rect 485688 277170 485740 277176
rect 485504 274100 485556 274106
rect 485504 274042 485556 274048
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483112 270904 483164 270910
rect 483112 270846 483164 270852
rect 484320 266422 484348 273634
rect 485228 271720 485280 271726
rect 485228 271662 485280 271668
rect 485412 271720 485464 271726
rect 485412 271662 485464 271668
rect 485240 271046 485268 271662
rect 485228 271040 485280 271046
rect 485228 270982 485280 270988
rect 485424 269770 485452 271662
rect 485056 269742 485452 269770
rect 485056 266558 485084 269742
rect 485700 267734 485728 277170
rect 486620 274514 486648 278052
rect 486608 274508 486660 274514
rect 486608 274450 486660 274456
rect 487816 274378 487844 278052
rect 488552 278038 489026 278066
rect 488356 274644 488408 274650
rect 488356 274586 488408 274592
rect 487804 274372 487856 274378
rect 487804 274314 487856 274320
rect 487068 273828 487120 273834
rect 487068 273770 487120 273776
rect 486884 270768 486936 270774
rect 486884 270710 486936 270716
rect 485424 267706 485728 267734
rect 485044 266552 485096 266558
rect 485044 266494 485096 266500
rect 482836 266416 482888 266422
rect 482836 266358 482888 266364
rect 483388 266416 483440 266422
rect 483388 266358 483440 266364
rect 484308 266416 484360 266422
rect 484308 266358 484360 266364
rect 483400 264316 483428 266358
rect 484216 266280 484268 266286
rect 484216 266222 484268 266228
rect 484228 264316 484256 266222
rect 485424 264330 485452 267706
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 485070 264302 485452 264330
rect 485884 264316 485912 266358
rect 486896 264330 486924 270710
rect 487080 266422 487108 273770
rect 487068 266416 487120 266422
rect 487068 266358 487120 266364
rect 487528 266212 487580 266218
rect 487528 266154 487580 266160
rect 486726 264302 486924 264330
rect 487540 264316 487568 266154
rect 488368 264316 488396 274586
rect 488552 268938 488580 278038
rect 489918 272776 489974 272785
rect 489918 272711 489974 272720
rect 489932 272626 489960 272711
rect 489886 272598 489960 272626
rect 489886 272542 489914 272598
rect 489874 272536 489926 272542
rect 489874 272478 489926 272484
rect 490012 272536 490064 272542
rect 490012 272478 490064 272484
rect 490024 272218 490052 272478
rect 489886 272190 490052 272218
rect 489886 272134 489914 272190
rect 489874 272128 489926 272134
rect 489874 272070 489926 272076
rect 490012 272128 490064 272134
rect 490012 272070 490064 272076
rect 490024 271726 490052 272070
rect 490012 271720 490064 271726
rect 490012 271662 490064 271668
rect 490208 271046 490236 278052
rect 491404 275194 491432 278052
rect 491772 278038 492614 278066
rect 491392 275188 491444 275194
rect 491392 275130 491444 275136
rect 491208 274100 491260 274106
rect 491208 274042 491260 274048
rect 490196 271040 490248 271046
rect 490196 270982 490248 270988
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 268932 488592 268938
rect 488540 268874 488592 268880
rect 489656 264330 489684 270574
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 491220 264330 491248 274042
rect 491772 269074 491800 278038
rect 493324 275188 493376 275194
rect 493324 275130 493376 275136
rect 492404 275052 492456 275058
rect 492404 274994 492456 275000
rect 492416 270910 492444 274994
rect 492404 270904 492456 270910
rect 492404 270846 492456 270852
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491760 269068 491812 269074
rect 491760 269010 491812 269016
rect 492600 266490 492628 270846
rect 493336 266898 493364 275130
rect 493704 271862 493732 278052
rect 494900 275058 494928 278052
rect 495728 278038 496110 278066
rect 495072 277092 495124 277098
rect 495072 277034 495124 277040
rect 494888 275052 494940 275058
rect 494888 274994 494940 275000
rect 493692 271856 493744 271862
rect 493692 271798 493744 271804
rect 493600 268252 493652 268258
rect 493600 268194 493652 268200
rect 493324 266892 493376 266898
rect 493324 266834 493376 266840
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492588 266484 492640 266490
rect 492588 266426 492640 266432
rect 490866 264302 491248 264330
rect 491680 264316 491708 266426
rect 492496 266076 492548 266082
rect 492496 266018 492548 266024
rect 492508 264316 492536 266018
rect 493612 264330 493640 268194
rect 495084 267734 495112 277034
rect 495728 272785 495756 278038
rect 495714 272776 495770 272785
rect 495714 272711 495770 272720
rect 496544 271856 496596 271862
rect 496544 271798 496596 271804
rect 495256 271040 495308 271046
rect 495256 270982 495308 270988
rect 494992 267706 495112 267734
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 493350 264302 493640 264330
rect 494164 264316 494192 266426
rect 494992 264316 495020 267706
rect 495268 266490 495296 270982
rect 495808 268116 495860 268122
rect 495808 268058 495860 268064
rect 495256 266484 495308 266490
rect 495256 266426 495308 266432
rect 495820 264316 495848 268058
rect 496556 264330 496584 271798
rect 497292 271590 497320 278052
rect 498488 275738 498516 278052
rect 499684 277394 499712 278052
rect 499592 277366 499712 277394
rect 498476 275732 498528 275738
rect 498476 275674 498528 275680
rect 497464 275188 497516 275194
rect 497464 275130 497516 275136
rect 497280 271584 497332 271590
rect 497280 271526 497332 271532
rect 497476 267578 497504 275130
rect 499304 271584 499356 271590
rect 499304 271526 499356 271532
rect 498292 269068 498344 269074
rect 498292 269010 498344 269016
rect 497464 267572 497516 267578
rect 497464 267514 497516 267520
rect 497464 266892 497516 266898
rect 497464 266834 497516 266840
rect 496556 264302 496662 264330
rect 497476 264316 497504 266834
rect 498304 264316 498332 269010
rect 499316 264330 499344 271526
rect 499592 268802 499620 277366
rect 500880 271454 500908 278052
rect 501604 275596 501656 275602
rect 501604 275538 501656 275544
rect 500868 271448 500920 271454
rect 500868 271390 500920 271396
rect 500776 268932 500828 268938
rect 500776 268874 500828 268880
rect 499580 268796 499632 268802
rect 499580 268738 499632 268744
rect 499948 266620 500000 266626
rect 499948 266562 500000 266568
rect 499146 264302 499344 264330
rect 499960 264316 499988 266562
rect 500788 264316 500816 268874
rect 501616 267714 501644 275538
rect 501984 275058 502012 278052
rect 502352 278038 503194 278066
rect 501972 275052 502024 275058
rect 501972 274994 502024 275000
rect 501972 271720 502024 271726
rect 501972 271662 502024 271668
rect 501604 267708 501656 267714
rect 501604 267650 501656 267656
rect 501984 264330 502012 271662
rect 502352 268666 502380 278038
rect 503444 275052 503496 275058
rect 503444 274994 503496 275000
rect 502340 268660 502392 268666
rect 502340 268602 502392 268608
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268602
rect 503456 266490 503484 274994
rect 504376 271318 504404 278052
rect 505572 275194 505600 278052
rect 505560 275188 505612 275194
rect 505560 275130 505612 275136
rect 506768 271998 506796 278052
rect 507964 277394 507992 278052
rect 507964 277366 508084 277394
rect 507860 275732 507912 275738
rect 507860 275674 507912 275680
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506756 271992 506808 271998
rect 506756 271934 506808 271940
rect 507124 271992 507176 271998
rect 507124 271934 507176 271940
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 504364 271312 504416 271318
rect 504364 271254 504416 271260
rect 504824 267572 504876 267578
rect 504824 267514 504876 267520
rect 503444 266484 503496 266490
rect 503444 266426 503496 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 267514
rect 505020 266490 505048 271390
rect 505744 268796 505796 268802
rect 505744 268738 505796 268744
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 504836 264302 504942 264330
rect 505756 264316 505784 268738
rect 507136 266762 507164 271934
rect 507504 267734 507532 275130
rect 507872 274242 507900 275674
rect 507860 274236 507912 274242
rect 507860 274178 507912 274184
rect 508056 272270 508084 277366
rect 509068 276010 509096 278052
rect 509252 278038 510278 278066
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 508596 274372 508648 274378
rect 508596 274314 508648 274320
rect 508044 272264 508096 272270
rect 508044 272206 508096 272212
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 507124 266756 507176 266762
rect 507124 266698 507176 266704
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 508608 264330 508636 274314
rect 509056 269544 509108 269550
rect 509056 269486 509108 269492
rect 508254 264302 508636 264330
rect 509068 264316 509096 269486
rect 509252 268530 509280 278038
rect 511460 272406 511488 278052
rect 511632 276956 511684 276962
rect 511632 276898 511684 276904
rect 511448 272400 511500 272406
rect 511448 272342 511500 272348
rect 509240 268524 509292 268530
rect 509240 268466 509292 268472
rect 511644 267734 511672 276898
rect 512656 275602 512684 278052
rect 512644 275596 512696 275602
rect 512644 275538 512696 275544
rect 511816 274236 511868 274242
rect 511816 274178 511868 274184
rect 511552 267706 511672 267734
rect 509884 266756 509936 266762
rect 509884 266698 509936 266704
rect 509896 264316 509924 266698
rect 510712 266620 510764 266626
rect 510712 266562 510764 266568
rect 510724 264316 510752 266562
rect 511552 264316 511580 267706
rect 511828 266626 511856 274178
rect 513852 273086 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 273080 513892 273086
rect 513840 273022 513892 273028
rect 512644 272400 512696 272406
rect 512644 272342 512696 272348
rect 512656 267034 512684 272342
rect 513196 268524 513248 268530
rect 513196 268466 513248 268472
rect 512644 267028 512696 267034
rect 512644 266970 512696 266976
rect 511816 266620 511868 266626
rect 511816 266562 511868 266568
rect 512368 265940 512420 265946
rect 512368 265882 512420 265888
rect 512380 264316 512408 265882
rect 513208 264316 513236 268466
rect 514496 264330 514524 276762
rect 515048 273222 515076 278052
rect 515404 275596 515456 275602
rect 515404 275538 515456 275544
rect 515036 273216 515088 273222
rect 515036 273158 515088 273164
rect 515220 273216 515272 273222
rect 515220 273158 515272 273164
rect 515232 272406 515260 273158
rect 515220 272400 515272 272406
rect 515220 272342 515272 272348
rect 514852 267708 514904 267714
rect 514852 267650 514904 267656
rect 514050 264302 514524 264330
rect 514864 264316 514892 267650
rect 515416 267442 515444 275538
rect 516244 274786 516272 278052
rect 516796 278038 517362 278066
rect 516232 274780 516284 274786
rect 516232 274722 516284 274728
rect 516796 270502 516824 278038
rect 517152 276004 517204 276010
rect 517152 275946 517204 275952
rect 516784 270496 516836 270502
rect 516784 270438 516836 270444
rect 515404 267436 515456 267442
rect 515404 267378 515456 267384
rect 516508 266620 516560 266626
rect 516508 266562 516560 266568
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266562
rect 517164 264330 517192 275946
rect 518544 272950 518572 278052
rect 518716 276684 518768 276690
rect 518716 276626 518768 276632
rect 518532 272944 518584 272950
rect 518532 272886 518584 272892
rect 517336 272400 517388 272406
rect 517336 272342 517388 272348
rect 517348 266626 517376 272342
rect 517520 270496 517572 270502
rect 517520 270438 517572 270444
rect 517532 267734 517560 270438
rect 518728 267734 518756 276626
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 517532 267706 517744 267734
rect 517520 267572 517572 267578
rect 517520 267514 517572 267520
rect 517532 266626 517560 267514
rect 517716 266898 517744 267706
rect 518544 267706 518756 267734
rect 517704 266892 517756 266898
rect 517704 266834 517756 266840
rect 517336 266620 517388 266626
rect 517336 266562 517388 266568
rect 517520 266620 517572 266626
rect 517520 266562 517572 266568
rect 518544 264330 518572 267706
rect 519820 267436 519872 267442
rect 519820 267378 519872 267384
rect 518992 266892 519044 266898
rect 518992 266834 519044 266840
rect 517164 264302 517362 264330
rect 518190 264302 518572 264330
rect 519004 264316 519032 266834
rect 519832 264316 519860 267378
rect 520108 266898 520136 272206
rect 520292 270366 520320 278038
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520280 270360 520332 270366
rect 520280 270302 520332 270308
rect 520096 266892 520148 266898
rect 520096 266834 520148 266840
rect 520648 265668 520700 265674
rect 520648 265610 520700 265616
rect 520660 264316 520688 265610
rect 521488 264316 521516 273158
rect 522132 272814 522160 278052
rect 523328 275874 523356 278052
rect 524432 278038 524538 278066
rect 525352 278038 525642 278066
rect 523316 275868 523368 275874
rect 523316 275810 523368 275816
rect 524144 275868 524196 275874
rect 524144 275810 524196 275816
rect 524156 272814 524184 275810
rect 522120 272808 522172 272814
rect 522120 272750 522172 272756
rect 522764 272808 522816 272814
rect 522764 272750 522816 272756
rect 524144 272808 524196 272814
rect 524144 272750 524196 272756
rect 522776 264330 522804 272750
rect 523868 271176 523920 271182
rect 523866 271144 523868 271153
rect 524052 271176 524104 271182
rect 523920 271144 523922 271153
rect 524052 271118 524104 271124
rect 523866 271079 523922 271088
rect 523132 270224 523184 270230
rect 523132 270166 523184 270172
rect 522330 264302 522804 264330
rect 523144 264316 523172 270166
rect 524064 267734 524092 271118
rect 524432 270366 524460 278038
rect 525352 271153 525380 278038
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 526444 274780 526496 274786
rect 526444 274722 526496 274728
rect 525338 271144 525394 271153
rect 525338 271079 525394 271088
rect 524420 270360 524472 270366
rect 524420 270302 524472 270308
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 523972 267706 524092 267734
rect 523972 264316 524000 267706
rect 524788 267028 524840 267034
rect 524788 266970 524840 266976
rect 524800 264316 524828 266970
rect 525628 264316 525656 270302
rect 526456 267170 526484 274722
rect 526812 273080 526864 273086
rect 526812 273022 526864 273028
rect 526444 267164 526496 267170
rect 526444 267106 526496 267112
rect 526824 264330 526852 273022
rect 527192 270094 527220 278038
rect 528192 275596 528244 275602
rect 528192 275538 528244 275544
rect 527180 270088 527232 270094
rect 527180 270030 527232 270036
rect 528204 266898 528232 275538
rect 529216 272542 529244 278052
rect 530412 275330 530440 278052
rect 531332 278038 531622 278066
rect 530400 275324 530452 275330
rect 530400 275266 530452 275272
rect 529848 272944 529900 272950
rect 529848 272886 529900 272892
rect 529204 272536 529256 272542
rect 529204 272478 529256 272484
rect 528376 270088 528428 270094
rect 528376 270030 528428 270036
rect 527272 266892 527324 266898
rect 527272 266834 527324 266840
rect 528192 266892 528244 266898
rect 528192 266834 528244 266840
rect 526470 264302 526852 264330
rect 527284 264316 527312 266834
rect 528388 264330 528416 270030
rect 529664 267572 529716 267578
rect 529664 267514 529716 267520
rect 528928 266892 528980 266898
rect 528928 266834 528980 266840
rect 528126 264302 528416 264330
rect 528940 264316 528968 266834
rect 529676 264330 529704 267514
rect 529860 266898 529888 272886
rect 530398 270192 530454 270201
rect 530398 270127 530454 270136
rect 530412 269686 530440 270127
rect 531332 269822 531360 278038
rect 532332 275324 532384 275330
rect 532332 275266 532384 275272
rect 531964 269952 532016 269958
rect 531964 269894 532016 269900
rect 531320 269816 531372 269822
rect 531320 269758 531372 269764
rect 531976 269686 532004 269894
rect 530400 269680 530452 269686
rect 530400 269622 530452 269628
rect 530584 269680 530636 269686
rect 530584 269622 530636 269628
rect 531964 269680 532016 269686
rect 531964 269622 532016 269628
rect 529848 266892 529900 266898
rect 529848 266834 529900 266840
rect 529676 264302 529782 264330
rect 530596 264316 530624 269622
rect 532344 267734 532372 275266
rect 532516 272808 532568 272814
rect 532516 272750 532568 272756
rect 532252 267706 532372 267734
rect 531412 266892 531464 266898
rect 531412 266834 531464 266840
rect 531424 264316 531452 266834
rect 532252 264316 532280 267706
rect 532528 266898 532556 272750
rect 532712 268394 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 533712 272536 533764 272542
rect 533712 272478 533764 272484
rect 533528 270360 533580 270366
rect 533528 270302 533580 270308
rect 533160 270224 533212 270230
rect 533160 270166 533212 270172
rect 533172 269686 533200 270166
rect 533540 269958 533568 270302
rect 533528 269952 533580 269958
rect 533528 269894 533580 269900
rect 533160 269680 533212 269686
rect 533160 269622 533212 269628
rect 532700 268388 532752 268394
rect 532700 268330 532752 268336
rect 532516 266892 532568 266898
rect 532516 266834 532568 266840
rect 533068 266892 533120 266898
rect 533068 266834 533120 266840
rect 533080 264316 533108 266834
rect 533724 264330 533752 272478
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266898 534028 269894
rect 534736 267306 534764 274722
rect 536300 272678 536328 278052
rect 537496 275466 537524 278052
rect 538508 278038 538706 278066
rect 537484 275460 537536 275466
rect 537484 275402 537536 275408
rect 537300 275324 537352 275330
rect 537300 275266 537352 275272
rect 537576 275324 537628 275330
rect 537576 275266 537628 275272
rect 537944 275324 537996 275330
rect 537944 275266 537996 275272
rect 537312 275097 537340 275266
rect 537298 275088 537354 275097
rect 537298 275023 537354 275032
rect 536748 274508 536800 274514
rect 536748 274450 536800 274456
rect 536288 272672 536340 272678
rect 536288 272614 536340 272620
rect 536564 272672 536616 272678
rect 536564 272614 536616 272620
rect 534724 267300 534776 267306
rect 534724 267242 534776 267248
rect 534724 267164 534776 267170
rect 534724 267106 534776 267112
rect 533988 266892 534040 266898
rect 533988 266834 534040 266840
rect 533724 264302 533922 264330
rect 534736 264316 534764 267106
rect 535552 266892 535604 266898
rect 535552 266834 535604 266840
rect 535564 264316 535592 266834
rect 536576 264330 536604 272614
rect 536760 266898 536788 274450
rect 536748 266892 536800 266898
rect 536748 266834 536800 266840
rect 537588 264330 537616 275266
rect 537956 274786 537984 275266
rect 538126 275088 538182 275097
rect 538126 275023 538182 275032
rect 538140 274786 538168 275023
rect 537944 274780 537996 274786
rect 537944 274722 537996 274728
rect 538128 274780 538180 274786
rect 538128 274722 538180 274728
rect 537760 269952 537812 269958
rect 537758 269920 537760 269929
rect 537944 269952 537996 269958
rect 537812 269920 537814 269929
rect 537944 269894 537996 269900
rect 538310 269920 538366 269929
rect 537758 269855 537814 269864
rect 536406 264302 536604 264330
rect 537234 264302 537616 264330
rect 537956 264330 537984 269894
rect 538310 269855 538366 269864
rect 538324 269414 538352 269855
rect 538508 269822 538536 278038
rect 539888 277394 539916 278052
rect 539888 277366 540008 277394
rect 539322 273728 539378 273737
rect 539322 273663 539378 273672
rect 538496 269816 538548 269822
rect 538496 269758 538548 269764
rect 538680 269816 538732 269822
rect 538680 269758 538732 269764
rect 538128 269408 538180 269414
rect 538128 269350 538180 269356
rect 538312 269408 538364 269414
rect 538692 269362 538720 269758
rect 538312 269350 538364 269356
rect 538140 269226 538168 269350
rect 538508 269334 538720 269362
rect 538508 269226 538536 269334
rect 538140 269198 538536 269226
rect 539336 264330 539364 273663
rect 539692 266892 539744 266898
rect 539692 266834 539744 266840
rect 537956 264302 538062 264330
rect 538890 264302 539364 264330
rect 539704 264316 539732 266834
rect 539980 265130 540008 277366
rect 540992 275330 541020 278052
rect 541176 278038 542202 278066
rect 540980 275324 541032 275330
rect 540980 275266 541032 275272
rect 541176 269362 541204 278038
rect 543384 276282 543412 278052
rect 543372 276276 543424 276282
rect 543372 276218 543424 276224
rect 543004 275324 543056 275330
rect 543004 275266 543056 275272
rect 542266 274816 542322 274825
rect 543016 274786 543044 275266
rect 544580 274922 544608 278052
rect 545776 275738 545804 278052
rect 546512 278038 546986 278066
rect 547892 278038 548090 278066
rect 545764 275732 545816 275738
rect 545764 275674 545816 275680
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 543186 274816 543242 274825
rect 542266 274751 542322 274760
rect 543004 274780 543056 274786
rect 540624 269334 541204 269362
rect 540624 269278 540652 269334
rect 540612 269272 540664 269278
rect 540612 269214 540664 269220
rect 540796 269272 540848 269278
rect 540796 269214 540848 269220
rect 539968 265124 540020 265130
rect 539968 265066 540020 265072
rect 540808 264330 540836 269214
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 540546 264302 540836 264330
rect 541360 264316 541388 268330
rect 542280 267734 542308 274751
rect 543186 274751 543188 274760
rect 543004 274722 543056 274728
rect 543240 274751 543242 274760
rect 543188 274722 543240 274728
rect 543188 269952 543240 269958
rect 543188 269894 543240 269900
rect 542820 269816 542872 269822
rect 542820 269758 542872 269764
rect 542832 269090 542860 269758
rect 543200 269278 543228 269894
rect 543188 269272 543240 269278
rect 543188 269214 543240 269220
rect 546512 269210 546540 278038
rect 547510 274000 547566 274009
rect 547510 273935 547512 273944
rect 547564 273935 547566 273944
rect 547696 273964 547748 273970
rect 547512 273906 547564 273912
rect 547696 273906 547748 273912
rect 547708 273737 547736 273906
rect 547694 273728 547750 273737
rect 547694 273663 547750 273672
rect 543372 269204 543424 269210
rect 543372 269146 543424 269152
rect 546500 269204 546552 269210
rect 546500 269146 546552 269152
rect 543384 269090 543412 269146
rect 542832 269062 543412 269090
rect 542188 267706 542308 267734
rect 542188 264316 542216 267706
rect 543004 267300 543056 267306
rect 543004 267242 543056 267248
rect 543016 264316 543044 267242
rect 547892 265266 547920 278038
rect 549272 274009 549300 278052
rect 550468 276418 550496 278052
rect 551664 276554 551692 278052
rect 552492 278038 552874 278066
rect 553412 278038 554070 278066
rect 554792 278038 555266 278066
rect 551652 276548 551704 276554
rect 551652 276490 551704 276496
rect 550456 276412 550508 276418
rect 550456 276354 550508 276360
rect 549258 274000 549314 274009
rect 549258 273935 549314 273944
rect 549902 273728 549958 273737
rect 549902 273663 549958 273672
rect 549916 266490 549944 273663
rect 552492 273426 552520 278038
rect 552846 273728 552902 273737
rect 552664 273692 552716 273698
rect 552846 273663 552848 273672
rect 552664 273634 552716 273640
rect 552900 273663 552902 273672
rect 552848 273634 552900 273640
rect 552676 273426 552704 273634
rect 552480 273420 552532 273426
rect 552480 273362 552532 273368
rect 552664 273420 552716 273426
rect 552664 273362 552716 273368
rect 549904 266484 549956 266490
rect 549904 266426 549956 266432
rect 553412 265402 553440 278038
rect 554792 265538 554820 278038
rect 556356 273562 556384 278052
rect 557552 277370 557580 278052
rect 557540 277364 557592 277370
rect 557540 277306 557592 277312
rect 556344 273556 556396 273562
rect 556344 273498 556396 273504
rect 556804 273556 556856 273562
rect 556804 273498 556856 273504
rect 556816 266626 556844 273498
rect 558748 272134 558776 278052
rect 559944 273426 559972 278052
rect 560496 278038 561154 278066
rect 559932 273420 559984 273426
rect 559932 273362 559984 273368
rect 558736 272128 558788 272134
rect 558736 272070 558788 272076
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 560496 266354 560524 278038
rect 562336 277234 562364 278052
rect 562324 277228 562376 277234
rect 562324 277170 562376 277176
rect 562600 273828 562652 273834
rect 562600 273770 562652 273776
rect 562612 273714 562640 273770
rect 562244 273698 562640 273714
rect 563440 273698 563468 278052
rect 562232 273692 562640 273698
rect 562284 273686 562640 273692
rect 563428 273692 563480 273698
rect 562232 273634 562284 273640
rect 563428 273634 563480 273640
rect 563704 273692 563756 273698
rect 563704 273634 563756 273640
rect 563716 266762 563744 273634
rect 564636 270774 564664 278052
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 563704 266756 563756 266762
rect 563704 266698 563756 266704
rect 560484 266348 560536 266354
rect 560484 266290 560536 266296
rect 565832 266218 565860 278052
rect 567028 274650 567056 278052
rect 567016 274644 567068 274650
rect 567016 274586 567068 274592
rect 568224 270638 568252 278052
rect 569420 271998 569448 278052
rect 569972 278038 570630 278066
rect 569972 274106 570000 278038
rect 569960 274100 570012 274106
rect 569960 274042 570012 274048
rect 569408 271992 569460 271998
rect 569408 271934 569460 271940
rect 571720 270910 571748 278052
rect 572732 278038 572930 278066
rect 571984 274100 572036 274106
rect 571984 274042 572036 274048
rect 571996 273834 572024 274042
rect 571984 273828 572036 273834
rect 571984 273770 572036 273776
rect 571708 270904 571760 270910
rect 571708 270846 571760 270852
rect 571984 270904 572036 270910
rect 571984 270846 572036 270852
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 571996 267714 572024 270846
rect 571984 267708 572036 267714
rect 571984 267650 572036 267656
rect 565820 266212 565872 266218
rect 565820 266154 565872 266160
rect 572732 266082 572760 278038
rect 574112 268258 574140 278052
rect 575308 271046 575336 278052
rect 576504 277098 576532 278052
rect 576872 278038 577714 278066
rect 578528 278038 578910 278066
rect 579632 278038 580014 278066
rect 581012 278038 581210 278066
rect 576492 277092 576544 277098
rect 576492 277034 576544 277040
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 574100 268252 574152 268258
rect 574100 268194 574152 268200
rect 576872 268122 576900 278038
rect 578528 271862 578556 278038
rect 578516 271856 578568 271862
rect 578516 271798 578568 271804
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 268116 576912 268122
rect 576860 268058 576912 268064
rect 578896 267442 578924 271798
rect 579632 270502 579660 278038
rect 579620 270496 579672 270502
rect 579620 270438 579672 270444
rect 581012 269074 581040 278038
rect 582392 271590 582420 278052
rect 583588 274106 583616 278052
rect 583772 278038 584798 278066
rect 583576 274100 583628 274106
rect 583576 274042 583628 274048
rect 582380 271584 582432 271590
rect 582380 271526 582432 271532
rect 581644 270496 581696 270502
rect 581644 270438 581696 270444
rect 581656 269414 581684 270438
rect 581644 269408 581696 269414
rect 581644 269350 581696 269356
rect 581000 269068 581052 269074
rect 581000 269010 581052 269016
rect 583772 268938 583800 278038
rect 585980 271726 586008 278052
rect 587084 275058 587112 278052
rect 587912 278038 588294 278066
rect 587072 275052 587124 275058
rect 587072 274994 587124 275000
rect 585968 271720 586020 271726
rect 585968 271662 586020 271668
rect 585784 271584 585836 271590
rect 585784 271526 585836 271532
rect 583760 268932 583812 268938
rect 583760 268874 583812 268880
rect 585796 267578 585824 271526
rect 587912 268666 587940 278038
rect 589476 271454 589504 278052
rect 590672 273562 590700 278052
rect 590856 278038 591882 278066
rect 590660 273556 590712 273562
rect 590660 273498 590712 273504
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 590856 268802 590884 278038
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 595088 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 595088 274378 595116 278038
rect 595076 274372 595128 274378
rect 595076 274314 595128 274320
rect 595444 274372 595496 274378
rect 595444 274314 595496 274320
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 590844 268796 590896 268802
rect 590844 268738 590896 268744
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 585784 267572 585836 267578
rect 585784 267514 585836 267520
rect 578884 267436 578936 267442
rect 578884 267378 578936 267384
rect 595456 266898 595484 274314
rect 596192 269550 596220 278038
rect 597756 273834 597784 278052
rect 598952 274242 598980 278052
rect 600148 276962 600176 278052
rect 600332 278038 601358 278066
rect 601712 278038 602462 278066
rect 600136 276956 600188 276962
rect 600136 276898 600188 276904
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 597744 273828 597796 273834
rect 597744 273770 597796 273776
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 595444 266892 595496 266898
rect 595444 266834 595496 266840
rect 572720 266076 572772 266082
rect 572720 266018 572772 266024
rect 600332 265946 600360 278038
rect 601712 268530 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 270910 604868 278052
rect 605852 278038 606050 278066
rect 604828 270904 604880 270910
rect 604828 270846 604880 270852
rect 601700 268524 601752 268530
rect 601700 268466 601752 268472
rect 600320 265940 600372 265946
rect 600320 265882 600372 265888
rect 605852 265810 605880 278038
rect 607232 272406 607260 278052
rect 608428 276010 608456 278052
rect 609624 276690 609652 278052
rect 609612 276684 609664 276690
rect 609612 276626 609664 276632
rect 608416 276004 608468 276010
rect 608416 275946 608468 275952
rect 607220 272400 607272 272406
rect 607220 272342 607272 272348
rect 610728 272270 610756 278052
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611924 271862 611952 278052
rect 612752 278038 613134 278066
rect 611912 271856 611964 271862
rect 611912 271798 611964 271804
rect 612004 271312 612056 271318
rect 612004 271254 612056 271260
rect 612016 267034 612044 271254
rect 612004 267028 612056 267034
rect 612004 266970 612056 266976
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 612752 265674 612780 278038
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 616156 278038 616722 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 616156 269686 616184 278038
rect 617812 271182 617840 278052
rect 618640 278038 619022 278066
rect 619652 278038 620218 278066
rect 618640 271318 618668 278038
rect 618628 271312 618680 271318
rect 618628 271254 618680 271260
rect 618904 271312 618956 271318
rect 618904 271254 618956 271260
rect 617800 271176 617852 271182
rect 617800 271118 617852 271124
rect 616144 269680 616196 269686
rect 616144 269622 616196 269628
rect 618916 267170 618944 271254
rect 619652 270230 619680 278038
rect 621400 273086 621428 278052
rect 622596 275602 622624 278052
rect 623806 278038 624004 278066
rect 622584 275596 622636 275602
rect 622584 275538 622636 275544
rect 621388 273080 621440 273086
rect 621388 273022 621440 273028
rect 620284 270496 620336 270502
rect 620284 270438 620336 270444
rect 619640 270224 619692 270230
rect 619640 270166 619692 270172
rect 620296 270094 620324 270438
rect 623976 270230 624004 278038
rect 624988 272950 625016 278052
rect 624976 272944 625028 272950
rect 624976 272886 625028 272892
rect 626092 271590 626120 278052
rect 626552 278038 627302 278066
rect 626080 271584 626132 271590
rect 626080 271526 626132 271532
rect 625804 271176 625856 271182
rect 625804 271118 625856 271124
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 620284 270088 620336 270094
rect 620284 270030 620336 270036
rect 625816 267306 625844 271118
rect 626552 270366 626580 278038
rect 628484 272814 628512 278052
rect 629680 275330 629708 278052
rect 630692 278038 630890 278066
rect 629668 275324 629720 275330
rect 629668 275266 629720 275272
rect 628472 272808 628524 272814
rect 628472 272750 628524 272756
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 630692 270094 630720 278038
rect 632072 272542 632100 278052
rect 632060 272536 632112 272542
rect 632060 272478 632112 272484
rect 633268 271318 633296 278052
rect 634372 274514 634400 278052
rect 634360 274508 634412 274514
rect 634360 274450 634412 274456
rect 635568 272678 635596 278052
rect 636764 275466 636792 278052
rect 637592 278038 637974 278066
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 635556 272672 635608 272678
rect 635556 272614 635608 272620
rect 633256 271312 633308 271318
rect 633256 271254 633308 271260
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 637592 269822 637620 278038
rect 639156 273970 639184 278052
rect 640352 274378 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 274372 640392 274378
rect 640340 274314 640392 274320
rect 639144 273964 639196 273970
rect 639144 273906 639196 273912
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 641732 268394 641760 278038
rect 643848 274786 643876 278052
rect 643836 274780 643888 274786
rect 643836 274722 643888 274728
rect 645044 271182 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271176 645084 271182
rect 645032 271118 645084 271124
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 625804 267300 625856 267306
rect 625804 267242 625856 267248
rect 618904 267164 618956 267170
rect 618904 267106 618956 267112
rect 612740 265668 612792 265674
rect 612740 265610 612792 265616
rect 554780 265532 554832 265538
rect 554780 265474 554832 265480
rect 553400 265396 553452 265402
rect 553400 265338 553452 265344
rect 547880 265260 547932 265266
rect 547880 265202 547932 265208
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 645872 261526 645900 278038
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 560944 259480 560996 259486
rect 560944 259422 560996 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553490 255640 553546 255649
rect 553490 255575 553492 255584
rect 553544 255575 553546 255584
rect 555424 255604 555476 255610
rect 553492 255546 553544 255552
rect 555424 255546 555476 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 554136 251194 554188 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 137928 231328 137980 231334
rect 137928 231270 137980 231276
rect 91744 231192 91796 231198
rect 91744 231134 91796 231140
rect 86224 229900 86276 229906
rect 86224 229842 86276 229848
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227724 64840 227730
rect 64788 227666 64840 227672
rect 62946 225584 63002 225593
rect 62946 225519 63002 225528
rect 64604 220380 64656 220386
rect 64604 220322 64656 220328
rect 64616 219434 64644 220322
rect 64800 219434 64828 227666
rect 66168 225752 66220 225758
rect 66168 225694 66220 225700
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 63132 219156 63184 219162
rect 63132 219098 63184 219104
rect 62764 218884 62816 218890
rect 62764 218826 62816 218832
rect 63144 217138 63172 219098
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 225694
rect 67272 218204 67324 218210
rect 67272 218146 67324 218152
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 66444 218068 66496 218074
rect 66444 218010 66496 218016
rect 64708 217246 64782 217274
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218010
rect 67284 217138 67312 218146
rect 67560 218074 67588 228618
rect 68296 218210 68324 229706
rect 82084 229628 82136 229634
rect 82084 229570 82136 229576
rect 72424 226160 72476 226166
rect 72424 226102 72476 226108
rect 68928 224256 68980 224262
rect 68928 224198 68980 224204
rect 68744 223168 68796 223174
rect 68744 223110 68796 223116
rect 68284 218204 68336 218210
rect 68284 218146 68336 218152
rect 68756 218074 68784 223110
rect 67548 218068 67600 218074
rect 67548 218010 67600 218016
rect 68100 218068 68152 218074
rect 68100 218010 68152 218016
rect 68744 218068 68796 218074
rect 68744 218010 68796 218016
rect 68112 217138 68140 218010
rect 68940 217274 68968 224198
rect 71412 222896 71464 222902
rect 71412 222838 71464 222844
rect 69756 220244 69808 220250
rect 69756 220186 69808 220192
rect 69768 217274 69796 220186
rect 70584 219156 70636 219162
rect 70584 219098 70636 219104
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219098
rect 71424 217274 71452 222838
rect 72436 219026 72464 226102
rect 76564 225888 76616 225894
rect 76564 225830 76616 225836
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220108 73120 220114
rect 73068 220050 73120 220056
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220050
rect 73724 218074 73752 224334
rect 75828 223032 75880 223038
rect 75828 222974 75880 222980
rect 73896 221604 73948 221610
rect 73896 221546 73948 221552
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221546
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 222974
rect 76380 220652 76432 220658
rect 76380 220594 76432 220600
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220594
rect 76576 218210 76604 225830
rect 79968 224664 80020 224670
rect 79968 224606 80020 224612
rect 78588 222760 78640 222766
rect 78588 222702 78640 222708
rect 77208 219020 77260 219026
rect 77208 218962 77260 218968
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218962
rect 78600 218074 78628 222702
rect 79692 220516 79744 220522
rect 79692 220458 79744 220464
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220458
rect 79980 218074 80008 224606
rect 81348 223440 81400 223446
rect 81348 223382 81400 223388
rect 80520 220856 80572 220862
rect 80520 220798 80572 220804
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 220798
rect 81360 217274 81388 223382
rect 82096 221610 82124 229570
rect 86236 229094 86264 229842
rect 86144 229066 86264 229094
rect 83464 226024 83516 226030
rect 83464 225966 83516 225972
rect 82084 221604 82136 221610
rect 82084 221546 82136 221552
rect 83004 220992 83056 220998
rect 83004 220934 83056 220940
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220934
rect 83476 218074 83504 225966
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 85304 223304 85356 223310
rect 85304 223246 85356 223252
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 85316 218074 85344 223246
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224470
rect 86144 220862 86172 229066
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 222624 88024 222630
rect 87972 222566 88024 222572
rect 86316 221604 86368 221610
rect 86316 221546 86368 221552
rect 86132 220856 86184 220862
rect 86132 220798 86184 220804
rect 86328 217274 86356 221546
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 222566
rect 88260 218074 88288 227802
rect 89628 227180 89680 227186
rect 89628 227122 89680 227128
rect 89444 224800 89496 224806
rect 89444 224742 89496 224748
rect 89456 218074 89484 224742
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227122
rect 91284 222012 91336 222018
rect 91284 221954 91336 221960
rect 90456 218068 90508 218074
rect 90456 218010 90508 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 218010
rect 91296 217274 91324 221954
rect 91756 218074 91784 231134
rect 128268 231056 128320 231062
rect 128268 230998 128320 231004
rect 97908 230920 97960 230926
rect 97908 230862 97960 230868
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 93768 228812 93820 228818
rect 93768 228754 93820 228760
rect 93780 218074 93808 228754
rect 95252 227866 95280 230114
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96436 227316 96488 227322
rect 96436 227258 96488 227264
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94596 221876 94648 221882
rect 94596 221818 94648 221824
rect 91744 218068 91796 218074
rect 91744 218010 91796 218016
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92066 217252 92118 217258
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92066 217194 92118 217200
rect 92078 216988 92106 217194
rect 92952 217138 92980 218010
rect 93768 217456 93820 217462
rect 93768 217398 93820 217404
rect 93780 217138 93808 217398
rect 94608 217274 94636 221818
rect 96264 218074 96292 224878
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217246 94636 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217246
rect 95436 217138 95464 218010
rect 96448 217274 96476 227258
rect 97724 221740 97776 221746
rect 97724 221682 97776 221688
rect 97736 219434 97764 221682
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 218010
rect 97828 217274 97856 219406
rect 97920 218090 97948 230862
rect 110328 230784 110380 230790
rect 110328 230726 110380 230732
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 229084 100720 229090
rect 100668 229026 100720 229032
rect 99288 223576 99340 223582
rect 99288 223518 99340 223524
rect 98552 222760 98604 222766
rect 98552 222702 98604 222708
rect 98564 222494 98592 222702
rect 98552 222488 98604 222494
rect 98552 222430 98604 222436
rect 97920 218074 98040 218090
rect 99300 218074 99328 223518
rect 100392 218612 100444 218618
rect 100392 218554 100444 218560
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218554
rect 100680 218074 100708 229026
rect 102152 227458 102180 229434
rect 106188 229084 106240 229090
rect 106188 229026 106240 229032
rect 102140 227452 102192 227458
rect 102140 227394 102192 227400
rect 103428 227452 103480 227458
rect 103428 227394 103480 227400
rect 102048 224120 102100 224126
rect 102048 224062 102100 224068
rect 101220 220788 101272 220794
rect 101220 220730 101272 220736
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217274 101260 220730
rect 102060 217274 102088 224062
rect 103440 218074 103468 227394
rect 106004 223984 106056 223990
rect 106004 223926 106056 223932
rect 104532 221332 104584 221338
rect 104532 221274 104584 221280
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217246 101260 217274
rect 102014 217246 102088 217274
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217246
rect 102014 216988 102042 217246
rect 102888 217138 102916 218010
rect 103704 217592 103756 217598
rect 103704 217534 103756 217540
rect 103716 217138 103744 217534
rect 104544 217274 104572 221274
rect 105820 219496 105872 219502
rect 105820 219438 105872 219444
rect 105832 218618 105860 219438
rect 105820 218612 105872 218618
rect 105820 218554 105872 218560
rect 106016 218074 106044 223926
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 229026
rect 110144 227588 110196 227594
rect 110144 227530 110196 227536
rect 106924 226500 106976 226506
rect 106924 226442 106976 226448
rect 106936 219298 106964 226442
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 107844 219972 107896 219978
rect 107844 219914 107896 219920
rect 106924 219292 106976 219298
rect 106924 219234 106976 219240
rect 107016 218612 107068 218618
rect 107016 218554 107068 218560
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218554
rect 107856 217274 107884 219914
rect 108684 217274 108712 223790
rect 110156 218074 110184 227530
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217274 110368 230726
rect 118608 230648 118660 230654
rect 118608 230590 118660 230596
rect 111064 229356 111116 229362
rect 111064 229298 111116 229304
rect 111076 227730 111104 229298
rect 112812 228268 112864 228274
rect 112812 228210 112864 228216
rect 111064 227724 111116 227730
rect 111064 227666 111116 227672
rect 111984 222148 112036 222154
rect 111984 222090 112036 222096
rect 111156 221196 111208 221202
rect 111156 221138 111208 221144
rect 111168 217274 111196 221138
rect 111996 217274 112024 222090
rect 112824 217274 112852 228210
rect 117228 227724 117280 227730
rect 117228 227666 117280 227672
rect 115296 223712 115348 223718
rect 115296 223654 115348 223660
rect 114468 219836 114520 219842
rect 114468 219778 114520 219784
rect 113640 219292 113692 219298
rect 113640 219234 113692 219240
rect 109466 217110 109540 217138
rect 110294 217246 110368 217274
rect 111122 217246 111196 217274
rect 111950 217246 112024 217274
rect 112778 217246 112852 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 216988 111150 217246
rect 111950 216988 111978 217246
rect 112778 216988 112806 217246
rect 113652 217138 113680 219234
rect 114480 217274 114508 219778
rect 115308 217274 115336 223654
rect 117240 218074 117268 227666
rect 118424 222488 118476 222494
rect 118424 222430 118476 222436
rect 118436 219434 118464 222430
rect 118436 219406 118556 219434
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 117976 218346 118004 219098
rect 117964 218340 118016 218346
rect 117964 218282 118016 218288
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117780 218068 117832 218074
rect 117780 218010 117832 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 115262 217246 115336 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115262 216988 115290 217246
rect 116136 217138 116164 218010
rect 116952 217728 117004 217734
rect 116952 217670 117004 217676
rect 116964 217138 116992 217670
rect 117792 217138 117820 218010
rect 118528 217274 118556 219406
rect 118620 218090 118648 230590
rect 126888 230036 126940 230042
rect 126888 229978 126940 229984
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 118620 218074 118740 218090
rect 120000 218074 120028 228074
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 226296 122616 226302
rect 122564 226238 122616 226244
rect 121092 219700 121144 219706
rect 121092 219642 121144 219648
rect 120264 218476 120316 218482
rect 120264 218418 120316 218424
rect 118620 218068 118752 218074
rect 118620 218062 118700 218068
rect 118700 218010 118752 218016
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 118528 217246 118602 217274
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217138 120304 218418
rect 121104 217274 121132 219642
rect 122576 218074 122604 226238
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 226850
rect 123496 218346 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225480 125284 225486
rect 125232 225422 125284 225428
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123484 218340 123536 218346
rect 123484 218282 123536 218288
rect 123576 218204 123628 218210
rect 123576 218146 123628 218152
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 218146
rect 124416 217274 124444 221002
rect 125244 217274 125272 225422
rect 126520 222624 126572 222630
rect 126520 222566 126572 222572
rect 126532 222358 126560 222566
rect 126520 222352 126572 222358
rect 126520 222294 126572 222300
rect 126716 218074 126744 227938
rect 126060 218068 126112 218074
rect 126060 218010 126112 218016
rect 126704 218068 126756 218074
rect 126704 218010 126756 218016
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218010
rect 126900 217274 126928 229978
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 127808 219972 127860 219978
rect 127808 219914 127860 219920
rect 127636 219706 127664 219914
rect 127624 219700 127676 219706
rect 127624 219642 127676 219648
rect 127820 219570 127848 219914
rect 127808 219564 127860 219570
rect 127808 219506 127860 219512
rect 128280 218074 128308 230998
rect 130384 230444 130436 230450
rect 130384 230386 130436 230392
rect 129556 226772 129608 226778
rect 129556 226714 129608 226720
rect 129372 225344 129424 225350
rect 129372 225286 129424 225292
rect 129384 218074 129412 225286
rect 127716 218068 127768 218074
rect 127716 218010 127768 218016
rect 128268 218068 128320 218074
rect 128268 218010 128320 218016
rect 128544 218068 128596 218074
rect 128544 218010 128596 218016
rect 129372 218068 129424 218074
rect 129372 218010 129424 218016
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218010
rect 128556 217138 128584 218010
rect 129568 217274 129596 226714
rect 130396 225214 130424 230386
rect 133788 230308 133840 230314
rect 133788 230250 133840 230256
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 130384 225208 130436 225214
rect 130384 225150 130436 225156
rect 132408 225072 132460 225078
rect 132408 225014 132460 225020
rect 132420 218346 132448 225014
rect 132592 219156 132644 219162
rect 132592 219098 132644 219104
rect 131856 218340 131908 218346
rect 131856 218282 131908 218288
rect 132408 218340 132460 218346
rect 132408 218282 132460 218288
rect 130200 218068 130252 218074
rect 130200 218010 130252 218016
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218010
rect 131028 217864 131080 217870
rect 131028 217806 131080 217812
rect 131040 217138 131068 217806
rect 131868 217138 131896 218282
rect 132604 218226 132632 219098
rect 132512 218198 132632 218226
rect 132512 218074 132540 218198
rect 133524 218074 133552 227802
rect 133800 219434 133828 230250
rect 136548 226636 136600 226642
rect 136548 226578 136600 226584
rect 135076 225208 135128 225214
rect 135076 225150 135128 225156
rect 134340 219564 134392 219570
rect 134340 219506 134392 219512
rect 133708 219406 133828 219434
rect 132500 218068 132552 218074
rect 132500 218010 132552 218016
rect 132684 218068 132736 218074
rect 132684 218010 132736 218016
rect 133512 218068 133564 218074
rect 133512 218010 133564 218016
rect 132696 217138 132724 218010
rect 133708 217274 133736 219406
rect 134352 217274 134380 219506
rect 130166 217110 130240 217138
rect 130994 217110 131068 217138
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 225150
rect 136560 218074 136588 226578
rect 137940 219434 137968 231270
rect 140042 229120 140098 229129
rect 140042 229055 140098 229064
rect 139306 228304 139362 228313
rect 139306 228239 139362 228248
rect 139124 222352 139176 222358
rect 139124 222294 139176 222300
rect 137664 219406 137968 219434
rect 136824 218340 136876 218346
rect 136824 218282 136876 218288
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 136548 218068 136600 218074
rect 136548 218010 136600 218016
rect 135088 217246 135162 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217110
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218010
rect 136836 217138 136864 218282
rect 137664 217274 137692 219406
rect 139136 218074 139164 222294
rect 138480 218068 138532 218074
rect 138480 218010 138532 218016
rect 139124 218068 139176 218074
rect 139124 218010 139176 218016
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 218010
rect 139320 217274 139348 228239
rect 140056 219026 140084 229055
rect 141160 228410 141188 231676
rect 141344 231662 141818 231690
rect 142172 231662 142462 231690
rect 142816 231662 143106 231690
rect 141148 228404 141200 228410
rect 141148 228346 141200 228352
rect 141148 226160 141200 226166
rect 141146 226128 141148 226137
rect 141200 226128 141202 226137
rect 141146 226063 141202 226072
rect 141344 221474 141372 231662
rect 142172 227050 142200 231662
rect 142434 230480 142490 230489
rect 142434 230415 142436 230424
rect 142488 230415 142490 230424
rect 142620 230444 142672 230450
rect 142436 230386 142488 230392
rect 142620 230386 142672 230392
rect 142632 229770 142660 230386
rect 142620 229764 142672 229770
rect 142620 229706 142672 229712
rect 142816 228698 142844 231662
rect 142988 229084 143040 229090
rect 142988 229026 143040 229032
rect 143448 229084 143500 229090
rect 143448 229026 143500 229032
rect 142632 228670 142844 228698
rect 143000 228682 143028 229026
rect 142988 228676 143040 228682
rect 142632 228546 142660 228670
rect 142988 228618 143040 228624
rect 142620 228540 142672 228546
rect 142620 228482 142672 228488
rect 142988 228540 143040 228546
rect 142988 228482 143040 228488
rect 143000 228313 143028 228482
rect 142986 228304 143042 228313
rect 142986 228239 143042 228248
rect 142160 227044 142212 227050
rect 142160 226986 142212 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141516 226160 141568 226166
rect 141516 226102 141568 226108
rect 141528 225622 141556 226102
rect 141516 225616 141568 225622
rect 141516 225558 141568 225564
rect 141792 225616 141844 225622
rect 141792 225558 141844 225564
rect 141332 221468 141384 221474
rect 141332 221410 141384 221416
rect 140778 220416 140834 220425
rect 140778 220351 140834 220360
rect 140792 219706 140820 220351
rect 140780 219700 140832 219706
rect 140780 219642 140832 219648
rect 140964 219700 141016 219706
rect 140964 219642 141016 219648
rect 140044 219020 140096 219026
rect 140044 218962 140096 218968
rect 139492 218340 139544 218346
rect 139492 218282 139544 218288
rect 140136 218340 140188 218346
rect 140136 218282 140188 218288
rect 139504 218074 139532 218282
rect 139492 218068 139544 218074
rect 139492 218010 139544 218016
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218282
rect 140976 217274 141004 219642
rect 141804 217274 141832 225558
rect 142250 220416 142306 220425
rect 141976 220380 142028 220386
rect 142250 220351 142306 220360
rect 141976 220322 142028 220328
rect 141988 219745 142016 220322
rect 142264 220250 142292 220351
rect 142252 220244 142304 220250
rect 142252 220186 142304 220192
rect 141974 219736 142030 219745
rect 141974 219671 142030 219680
rect 142436 218884 142488 218890
rect 142436 218826 142488 218832
rect 142448 218618 142476 218826
rect 143276 218618 143304 226986
rect 142436 218612 142488 218618
rect 142436 218554 142488 218560
rect 142620 218612 142672 218618
rect 142620 218554 142672 218560
rect 143264 218612 143316 218618
rect 143264 218554 143316 218560
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218554
rect 143460 217274 143488 229026
rect 143736 218754 143764 231676
rect 144104 231662 144394 231690
rect 144104 230489 144132 231662
rect 144090 230480 144146 230489
rect 144090 230415 144146 230424
rect 143998 229528 144054 229537
rect 143998 229463 144000 229472
rect 144052 229463 144054 229472
rect 144184 229492 144236 229498
rect 144000 229434 144052 229440
rect 144184 229434 144236 229440
rect 144196 219745 144224 229434
rect 145024 226166 145052 231676
rect 145392 231662 145682 231690
rect 146326 231662 146616 231690
rect 145392 229537 145420 231662
rect 146208 231600 146260 231606
rect 146208 231542 146260 231548
rect 146220 230450 146248 231542
rect 146208 230444 146260 230450
rect 146208 230386 146260 230392
rect 145378 229528 145434 229537
rect 145378 229463 145434 229472
rect 146206 229392 146262 229401
rect 146206 229327 146262 229336
rect 146220 229090 146248 229327
rect 146208 229084 146260 229090
rect 146208 229026 146260 229032
rect 146392 229084 146444 229090
rect 146392 229026 146444 229032
rect 146404 228970 146432 229026
rect 145944 228942 146432 228970
rect 145944 228546 145972 228942
rect 145932 228540 145984 228546
rect 145932 228482 145984 228488
rect 146116 228540 146168 228546
rect 146116 228482 146168 228488
rect 145012 226160 145064 226166
rect 145196 226160 145248 226166
rect 145012 226102 145064 226108
rect 145194 226128 145196 226137
rect 145248 226128 145250 226137
rect 145194 226063 145250 226072
rect 145930 222320 145986 222329
rect 145930 222255 145986 222264
rect 144642 220688 144698 220697
rect 144642 220623 144698 220632
rect 144656 220386 144684 220623
rect 144644 220380 144696 220386
rect 144644 220322 144696 220328
rect 144828 220380 144880 220386
rect 144828 220322 144880 220328
rect 144182 219736 144238 219745
rect 144182 219671 144238 219680
rect 143724 218748 143776 218754
rect 143724 218690 143776 218696
rect 144840 218618 144868 220322
rect 145944 218618 145972 222255
rect 144276 218612 144328 218618
rect 144276 218554 144328 218560
rect 144828 218612 144880 218618
rect 144828 218554 144880 218560
rect 145104 218612 145156 218618
rect 145104 218554 145156 218560
rect 145932 218612 145984 218618
rect 145932 218554 145984 218560
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144288 217138 144316 218554
rect 145116 217138 145144 218554
rect 146128 217274 146156 228482
rect 146588 226506 146616 231662
rect 146760 231464 146812 231470
rect 146760 231406 146812 231412
rect 146576 226500 146628 226506
rect 146576 226442 146628 226448
rect 146772 226166 146800 231406
rect 146956 229498 146984 231676
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 147232 231470 147260 231662
rect 147220 231464 147272 231470
rect 147220 231406 147272 231412
rect 147634 230444 147686 230450
rect 147634 230386 147686 230392
rect 147646 230194 147674 230386
rect 147324 230166 147674 230194
rect 147128 229560 147180 229566
rect 147128 229502 147180 229508
rect 146944 229492 146996 229498
rect 146944 229434 146996 229440
rect 147140 229129 147168 229502
rect 147126 229120 147182 229129
rect 147126 229055 147182 229064
rect 146760 226160 146812 226166
rect 146760 226102 146812 226108
rect 147324 224954 147352 230166
rect 147968 229809 147996 231662
rect 147586 229800 147642 229809
rect 147954 229800 148010 229809
rect 147586 229735 147642 229744
rect 147772 229764 147824 229770
rect 147600 229362 147628 229735
rect 147954 229735 148010 229744
rect 147772 229706 147824 229712
rect 147784 229650 147812 229706
rect 147784 229634 148180 229650
rect 147784 229628 148192 229634
rect 147784 229622 148140 229628
rect 148140 229570 148192 229576
rect 147770 229392 147826 229401
rect 147588 229356 147640 229362
rect 147770 229327 147772 229336
rect 147588 229298 147640 229304
rect 147824 229327 147826 229336
rect 147772 229298 147824 229304
rect 148888 228410 148916 231676
rect 149532 230450 149560 231676
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 151004 231662 151478 231690
rect 149520 230444 149572 230450
rect 149520 230386 149572 230392
rect 148876 228404 148928 228410
rect 148876 228346 148928 228352
rect 148968 226160 149020 226166
rect 148968 226102 149020 226108
rect 146588 224926 147352 224954
rect 146588 223174 146616 224926
rect 147678 223408 147734 223417
rect 147678 223343 147734 223352
rect 147692 223258 147720 223343
rect 147646 223230 147720 223258
rect 147646 223174 147674 223230
rect 146576 223168 146628 223174
rect 146576 223110 146628 223116
rect 146760 223168 146812 223174
rect 146760 223110 146812 223116
rect 147634 223168 147686 223174
rect 147634 223110 147686 223116
rect 147772 223168 147824 223174
rect 147772 223110 147824 223116
rect 146772 222494 146800 223110
rect 147784 223009 147812 223110
rect 147310 223000 147366 223009
rect 147310 222935 147366 222944
rect 147770 223000 147826 223009
rect 147770 222935 147826 222944
rect 146760 222488 146812 222494
rect 146760 222430 146812 222436
rect 147128 222352 147180 222358
rect 147126 222320 147128 222329
rect 147180 222320 147182 222329
rect 147126 222255 147182 222264
rect 147324 219434 147352 222935
rect 147588 221468 147640 221474
rect 147588 221410 147640 221416
rect 147128 219428 147352 219434
rect 147180 219406 147352 219428
rect 147128 219370 147180 219376
rect 146760 218748 146812 218754
rect 146760 218690 146812 218696
rect 144242 217110 144316 217138
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 144242 216988 144270 217110
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218690
rect 147600 217274 147628 221410
rect 148980 219434 149008 226102
rect 149808 225758 149836 231662
rect 150544 231606 150572 231662
rect 150532 231600 150584 231606
rect 150532 231542 150584 231548
rect 150346 229256 150402 229265
rect 150346 229191 150402 229200
rect 150072 226500 150124 226506
rect 150072 226442 150124 226448
rect 149796 225752 149848 225758
rect 149796 225694 149848 225700
rect 150084 224954 150112 226442
rect 150360 224954 150388 229191
rect 151004 224954 151032 231662
rect 151176 229356 151228 229362
rect 151176 229298 151228 229304
rect 151188 225842 151216 229298
rect 149992 224926 150112 224954
rect 150176 224926 150388 224954
rect 150912 224926 151032 224954
rect 151096 225814 151216 225842
rect 149242 220960 149298 220969
rect 149242 220895 149298 220904
rect 149256 220658 149284 220895
rect 149244 220652 149296 220658
rect 149244 220594 149296 220600
rect 149428 220652 149480 220658
rect 149428 220594 149480 220600
rect 149440 220250 149468 220594
rect 149428 220244 149480 220250
rect 149428 220186 149480 220192
rect 149992 219434 150020 224926
rect 148416 219428 148468 219434
rect 148416 219370 148468 219376
rect 148968 219428 149020 219434
rect 148968 219370 149020 219376
rect 149244 219428 149296 219434
rect 149244 219370 149296 219376
rect 149980 219428 150032 219434
rect 149980 219370 150032 219376
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 219370
rect 149256 217138 149284 219370
rect 150176 217274 150204 224926
rect 150912 220697 150940 224926
rect 151096 220930 151124 225814
rect 151268 225752 151320 225758
rect 151268 225694 151320 225700
rect 151280 224954 151308 225694
rect 151280 224926 151676 224954
rect 151084 220924 151136 220930
rect 151084 220866 151136 220872
rect 150898 220688 150954 220697
rect 150898 220623 150954 220632
rect 150900 220244 150952 220250
rect 150900 220186 150952 220192
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150204 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150912 217138 150940 220186
rect 151648 217274 151676 224926
rect 152108 222902 152136 231676
rect 152464 231328 152516 231334
rect 152464 231270 152516 231276
rect 152476 230518 152504 231270
rect 152464 230512 152516 230518
rect 152464 230454 152516 230460
rect 152464 228676 152516 228682
rect 152464 228618 152516 228624
rect 152476 228410 152504 228618
rect 152464 228404 152516 228410
rect 152464 228346 152516 228352
rect 152752 224262 152780 231676
rect 153396 229226 153424 231676
rect 153580 231662 154054 231690
rect 154698 231662 154988 231690
rect 153384 229220 153436 229226
rect 153384 229162 153436 229168
rect 153108 228676 153160 228682
rect 153108 228618 153160 228624
rect 152740 224256 152792 224262
rect 152740 224198 152792 224204
rect 152278 223408 152334 223417
rect 152278 223343 152334 223352
rect 152292 222902 152320 223343
rect 152096 222896 152148 222902
rect 152096 222838 152148 222844
rect 152280 222896 152332 222902
rect 152280 222838 152332 222844
rect 152186 222728 152242 222737
rect 152186 222663 152242 222672
rect 152200 218890 152228 222663
rect 153120 219434 153148 228618
rect 153580 220114 153608 231662
rect 153844 229356 153896 229362
rect 153844 229298 153896 229304
rect 153568 220108 153620 220114
rect 153568 220050 153620 220056
rect 152556 219428 152608 219434
rect 152556 219370 152608 219376
rect 153108 219428 153160 219434
rect 153108 219370 153160 219376
rect 152372 219292 152424 219298
rect 152372 219234 152424 219240
rect 152384 218890 152412 219234
rect 152188 218884 152240 218890
rect 152188 218826 152240 218832
rect 152372 218884 152424 218890
rect 152372 218826 152424 218832
rect 151648 217246 151722 217274
rect 150866 217110 150940 217138
rect 150866 216988 150894 217110
rect 151694 216988 151722 217246
rect 152568 217138 152596 219370
rect 153856 219298 153884 229298
rect 154960 223038 154988 231662
rect 155328 224398 155356 231676
rect 155500 231600 155552 231606
rect 155500 231542 155552 231548
rect 155316 224392 155368 224398
rect 155316 224334 155368 224340
rect 154948 223032 155000 223038
rect 154948 222974 155000 222980
rect 155132 223032 155184 223038
rect 155132 222974 155184 222980
rect 155144 222737 155172 222974
rect 155512 222902 155540 231542
rect 155776 231328 155828 231334
rect 155776 231270 155828 231276
rect 155788 229226 155816 231270
rect 155972 229634 156000 231676
rect 156156 231662 156630 231690
rect 156984 231662 157274 231690
rect 155960 229628 156012 229634
rect 155960 229570 156012 229576
rect 155776 229220 155828 229226
rect 155776 229162 155828 229168
rect 155776 224256 155828 224262
rect 155776 224198 155828 224204
rect 155500 222896 155552 222902
rect 155500 222838 155552 222844
rect 155130 222728 155186 222737
rect 155130 222663 155186 222672
rect 155040 220924 155092 220930
rect 155040 220866 155092 220872
rect 154212 220108 154264 220114
rect 154212 220050 154264 220056
rect 153200 219292 153252 219298
rect 153200 219234 153252 219240
rect 153844 219292 153896 219298
rect 153844 219234 153896 219240
rect 153212 219026 153240 219234
rect 153200 219020 153252 219026
rect 153200 218962 153252 218968
rect 153384 219020 153436 219026
rect 153384 218962 153436 218968
rect 153396 217138 153424 218962
rect 154224 217274 154252 220050
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155052 217138 155080 220866
rect 155788 217274 155816 224198
rect 156156 220969 156184 231662
rect 156984 231606 157012 231662
rect 156972 231600 157024 231606
rect 156972 231542 157024 231548
rect 156604 231464 156656 231470
rect 156604 231406 156656 231412
rect 156616 229362 156644 231406
rect 157294 230172 157346 230178
rect 157294 230114 157346 230120
rect 157432 230172 157484 230178
rect 157432 230114 157484 230120
rect 156786 229936 156842 229945
rect 156786 229871 156788 229880
rect 156840 229871 156842 229880
rect 156788 229842 156840 229848
rect 157306 229786 157334 230114
rect 157444 229945 157472 230114
rect 157430 229936 157486 229945
rect 157430 229871 157486 229880
rect 157306 229758 157656 229786
rect 157340 229628 157392 229634
rect 157340 229570 157392 229576
rect 156604 229356 156656 229362
rect 156604 229298 156656 229304
rect 156880 229084 156932 229090
rect 156880 229026 156932 229032
rect 156892 228857 156920 229026
rect 156878 228848 156934 228857
rect 156878 228783 156934 228792
rect 156878 227488 156934 227497
rect 156878 227423 156934 227432
rect 156892 227186 156920 227423
rect 156880 227180 156932 227186
rect 156880 227122 156932 227128
rect 157352 224398 157380 229570
rect 157628 229226 157656 229758
rect 157616 229220 157668 229226
rect 157616 229162 157668 229168
rect 157524 229084 157576 229090
rect 157524 229026 157576 229032
rect 157536 228857 157564 229026
rect 157522 228848 157578 228857
rect 157522 228783 157578 228792
rect 157904 225894 157932 231676
rect 158548 229906 158576 231676
rect 158916 231662 159206 231690
rect 158536 229900 158588 229906
rect 158536 229842 158588 229848
rect 157892 225888 157944 225894
rect 157892 225830 157944 225836
rect 156696 224392 156748 224398
rect 156696 224334 156748 224340
rect 157340 224392 157392 224398
rect 157340 224334 157392 224340
rect 156142 220960 156198 220969
rect 156142 220895 156198 220904
rect 155788 217246 155862 217274
rect 155006 217110 155080 217138
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 224334
rect 157248 223440 157300 223446
rect 157246 223408 157248 223417
rect 157432 223440 157484 223446
rect 157300 223408 157302 223417
rect 157246 223343 157302 223352
rect 157430 223408 157432 223417
rect 157484 223408 157486 223417
rect 157430 223343 157486 223352
rect 157524 223032 157576 223038
rect 157524 222974 157576 222980
rect 157536 217138 157564 222974
rect 158350 221640 158406 221649
rect 158350 221575 158406 221584
rect 158364 217138 158392 221575
rect 158916 220522 158944 231662
rect 159362 229392 159418 229401
rect 159362 229327 159364 229336
rect 159416 229327 159418 229336
rect 159364 229298 159416 229304
rect 159836 223446 159864 231676
rect 160006 228168 160062 228177
rect 160006 228103 160062 228112
rect 159824 223440 159876 223446
rect 159824 223382 159876 223388
rect 158904 220516 158956 220522
rect 158904 220458 158956 220464
rect 160020 219434 160048 228103
rect 160192 227180 160244 227186
rect 160192 227122 160244 227128
rect 160204 224262 160232 227122
rect 160480 224670 160508 231676
rect 161124 230178 161152 231676
rect 161768 231334 161796 231676
rect 161756 231328 161808 231334
rect 161756 231270 161808 231276
rect 161112 230172 161164 230178
rect 161112 230114 161164 230120
rect 160468 224664 160520 224670
rect 160468 224606 160520 224612
rect 161664 224392 161716 224398
rect 161664 224334 161716 224340
rect 160192 224256 160244 224262
rect 160192 224198 160244 224204
rect 160834 220416 160890 220425
rect 160834 220351 160890 220360
rect 159180 219428 159232 219434
rect 159180 219370 159232 219376
rect 160008 219428 160060 219434
rect 160008 219370 160060 219376
rect 159192 217138 159220 219370
rect 160008 219292 160060 219298
rect 160008 219234 160060 219240
rect 160020 217138 160048 219234
rect 160848 217138 160876 220351
rect 161676 217138 161704 224334
rect 162124 223440 162176 223446
rect 162124 223382 162176 223388
rect 162136 218890 162164 223382
rect 162412 223310 162440 231676
rect 163056 226030 163084 231676
rect 163700 231470 163728 231676
rect 163688 231464 163740 231470
rect 163688 231406 163740 231412
rect 163964 229900 164016 229906
rect 163964 229842 164016 229848
rect 163044 226024 163096 226030
rect 163044 225966 163096 225972
rect 162400 223304 162452 223310
rect 162400 223246 162452 223252
rect 163976 219434 164004 229842
rect 164344 221610 164372 231676
rect 164988 222766 165016 231676
rect 165160 224664 165212 224670
rect 165160 224606 165212 224612
rect 164976 222760 165028 222766
rect 164976 222702 165028 222708
rect 164514 221640 164570 221649
rect 164332 221604 164384 221610
rect 164514 221575 164516 221584
rect 164332 221546 164384 221552
rect 164568 221575 164570 221584
rect 164516 221546 164568 221552
rect 164148 220516 164200 220522
rect 164148 220458 164200 220464
rect 163320 219428 163372 219434
rect 163320 219370 163372 219376
rect 163964 219428 164016 219434
rect 163964 219370 164016 219376
rect 162124 218884 162176 218890
rect 162124 218826 162176 218832
rect 162492 218884 162544 218890
rect 162492 218826 162544 218832
rect 161940 218748 161992 218754
rect 161940 218690 161992 218696
rect 161952 218482 161980 218690
rect 161940 218476 161992 218482
rect 161940 218418 161992 218424
rect 162504 217138 162532 218826
rect 163332 217138 163360 219370
rect 164160 217138 164188 220458
rect 165172 217274 165200 224606
rect 165632 224534 165660 231676
rect 166276 229226 166304 231676
rect 166552 231662 166934 231690
rect 167196 231662 167578 231690
rect 166264 229220 166316 229226
rect 166264 229162 166316 229168
rect 166552 227497 166580 231662
rect 166998 229256 167054 229265
rect 166998 229191 167054 229200
rect 166814 228984 166870 228993
rect 167012 228954 167040 229191
rect 166814 228919 166870 228928
rect 167000 228948 167052 228954
rect 166828 228818 166856 228919
rect 167000 228890 167052 228896
rect 166816 228812 166868 228818
rect 166816 228754 166868 228760
rect 166954 228812 167006 228818
rect 166954 228754 167006 228760
rect 166966 228698 166994 228754
rect 166828 228670 166994 228698
rect 166828 228410 166856 228670
rect 166816 228404 166868 228410
rect 166816 228346 166868 228352
rect 166954 228404 167006 228410
rect 166954 228346 167006 228352
rect 166966 228290 166994 228346
rect 166828 228262 166994 228290
rect 166828 228177 166856 228262
rect 166814 228168 166870 228177
rect 166814 228103 166870 228112
rect 166538 227488 166594 227497
rect 166538 227423 166594 227432
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165988 224392 166040 224398
rect 165988 224334 166040 224340
rect 165620 222760 165672 222766
rect 165620 222702 165672 222708
rect 165632 218618 165660 222702
rect 165804 218748 165856 218754
rect 165804 218690 165856 218696
rect 165620 218612 165672 218618
rect 165620 218554 165672 218560
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217110 158392 217138
rect 159146 217110 159220 217138
rect 159974 217110 160048 217138
rect 160802 217110 160876 217138
rect 161630 217110 161704 217138
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 164114 217110 164188 217138
rect 164942 217246 165200 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217110
rect 159146 216988 159174 217110
rect 159974 216988 160002 217110
rect 160802 216988 160830 217110
rect 161630 216988 161658 217110
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217110
rect 164942 216988 164970 217246
rect 165816 217138 165844 218690
rect 166000 218210 166028 224334
rect 167196 222018 167224 231662
rect 167366 229256 167422 229265
rect 167366 229191 167368 229200
rect 167420 229191 167422 229200
rect 167368 229162 167420 229168
rect 167366 228984 167422 228993
rect 167366 228919 167368 228928
rect 167420 228919 167422 228928
rect 167368 228890 167420 228896
rect 168208 224806 168236 231676
rect 168852 231198 168880 231676
rect 168840 231192 168892 231198
rect 168840 231134 168892 231140
rect 169496 228954 169524 231676
rect 169864 231662 170154 231690
rect 170324 231662 170798 231690
rect 169484 228948 169536 228954
rect 169484 228890 169536 228896
rect 169482 227352 169538 227361
rect 169482 227287 169484 227296
rect 169536 227287 169538 227296
rect 169484 227258 169536 227264
rect 169668 225888 169720 225894
rect 169668 225830 169720 225836
rect 168196 224800 168248 224806
rect 168196 224742 168248 224748
rect 168288 224256 168340 224262
rect 168288 224198 168340 224204
rect 167184 222012 167236 222018
rect 167184 221954 167236 221960
rect 167460 222012 167512 222018
rect 167460 221954 167512 221960
rect 166998 220960 167054 220969
rect 166998 220895 167054 220904
rect 167012 220810 167040 220895
rect 166966 220794 167040 220810
rect 166954 220788 167040 220794
rect 166368 220748 166856 220776
rect 166368 220658 166396 220748
rect 166828 220674 166856 220748
rect 167006 220782 167040 220788
rect 167184 220788 167236 220794
rect 166954 220730 167006 220736
rect 167184 220730 167236 220736
rect 167196 220674 167224 220730
rect 166356 220652 166408 220658
rect 166356 220594 166408 220600
rect 166540 220652 166592 220658
rect 166828 220646 167224 220674
rect 166540 220594 166592 220600
rect 166552 220425 166580 220594
rect 166908 220516 166960 220522
rect 166908 220458 166960 220464
rect 167092 220516 167144 220522
rect 167092 220458 167144 220464
rect 166538 220416 166594 220425
rect 166538 220351 166594 220360
rect 166920 220289 166948 220458
rect 167104 220289 167132 220458
rect 166906 220280 166962 220289
rect 166906 220215 166962 220224
rect 167090 220280 167146 220289
rect 167090 220215 167146 220224
rect 166632 218612 166684 218618
rect 166632 218554 166684 218560
rect 165988 218204 166040 218210
rect 165988 218146 166040 218152
rect 166644 217138 166672 218554
rect 167472 217138 167500 221954
rect 168300 217138 168328 224198
rect 169680 219298 169708 225830
rect 169864 221882 169892 231662
rect 169852 221876 169904 221882
rect 169852 221818 169904 221824
rect 169116 219292 169168 219298
rect 169116 219234 169168 219240
rect 169668 219292 169720 219298
rect 169668 219234 169720 219240
rect 169128 217138 169156 219234
rect 169760 218884 169812 218890
rect 169760 218826 169812 218832
rect 169944 218884 169996 218890
rect 169944 218826 169996 218832
rect 169574 218512 169630 218521
rect 169772 218482 169800 218826
rect 169574 218447 169576 218456
rect 169628 218447 169630 218456
rect 169760 218476 169812 218482
rect 169576 218418 169628 218424
rect 169760 218418 169812 218424
rect 169956 217138 169984 218826
rect 170324 217326 170352 231662
rect 171048 229764 171100 229770
rect 171048 229706 171100 229712
rect 171060 218890 171088 229706
rect 171230 227624 171286 227633
rect 171230 227559 171286 227568
rect 171244 227458 171272 227559
rect 171232 227452 171284 227458
rect 171232 227394 171284 227400
rect 171428 226930 171456 231676
rect 171704 231662 172086 231690
rect 171704 227361 171732 231662
rect 172150 227624 172206 227633
rect 172150 227559 172206 227568
rect 172164 227458 172192 227559
rect 172152 227452 172204 227458
rect 172152 227394 172204 227400
rect 171690 227352 171746 227361
rect 171690 227287 171746 227296
rect 171600 227180 171652 227186
rect 171600 227122 171652 227128
rect 171244 226902 171456 226930
rect 171048 218884 171100 218890
rect 171048 218826 171100 218832
rect 170772 218068 170824 218074
rect 170772 218010 170824 218016
rect 170312 217320 170364 217326
rect 170312 217262 170364 217268
rect 170784 217138 170812 218010
rect 171244 217462 171272 226902
rect 171612 225894 171640 227122
rect 171600 225888 171652 225894
rect 171600 225830 171652 225836
rect 171784 225888 171836 225894
rect 171784 225830 171836 225836
rect 171796 224954 171824 225830
rect 171428 224926 171824 224954
rect 171428 218210 171456 224926
rect 171968 224800 172020 224806
rect 171968 224742 172020 224748
rect 172152 224800 172204 224806
rect 172152 224742 172204 224748
rect 171600 224528 171652 224534
rect 171600 224470 171652 224476
rect 171612 224126 171640 224470
rect 171980 224398 172008 224742
rect 171784 224392 171836 224398
rect 171784 224334 171836 224340
rect 171968 224392 172020 224398
rect 171968 224334 172020 224340
rect 171796 224126 171824 224334
rect 171600 224120 171652 224126
rect 171600 224062 171652 224068
rect 171784 224120 171836 224126
rect 171784 224062 171836 224068
rect 171784 223440 171836 223446
rect 171784 223382 171836 223388
rect 171796 222902 171824 223382
rect 171784 222896 171836 222902
rect 171784 222838 171836 222844
rect 171600 221740 171652 221746
rect 171600 221682 171652 221688
rect 171612 221202 171640 221682
rect 171784 221604 171836 221610
rect 171784 221546 171836 221552
rect 171796 221202 171824 221546
rect 171600 221196 171652 221202
rect 171600 221138 171652 221144
rect 171784 221196 171836 221202
rect 171784 221138 171836 221144
rect 172164 219298 172192 224742
rect 172716 221882 172744 231676
rect 172992 231662 173374 231690
rect 172992 224942 173020 231662
rect 174004 230926 174032 231676
rect 174280 231662 174662 231690
rect 175306 231662 175596 231690
rect 173992 230920 174044 230926
rect 173992 230862 174044 230868
rect 174280 229226 174308 231662
rect 174268 229220 174320 229226
rect 174268 229162 174320 229168
rect 173346 228848 173402 228857
rect 173346 228783 173402 228792
rect 174818 228848 174874 228857
rect 174818 228783 174820 228792
rect 172980 224936 173032 224942
rect 172980 224878 173032 224884
rect 172888 222896 172940 222902
rect 172888 222838 172940 222844
rect 172704 221876 172756 221882
rect 172704 221818 172756 221824
rect 171600 219292 171652 219298
rect 171600 219234 171652 219240
rect 172152 219292 172204 219298
rect 172152 219234 172204 219240
rect 172428 219292 172480 219298
rect 172428 219234 172480 219240
rect 171416 218204 171468 218210
rect 171416 218146 171468 218152
rect 171232 217456 171284 217462
rect 171232 217398 171284 217404
rect 171612 217138 171640 219234
rect 172440 217138 172468 219234
rect 172900 218521 172928 222838
rect 173360 219298 173388 228783
rect 174872 228783 174874 228792
rect 174820 228754 174872 228760
rect 174084 221876 174136 221882
rect 174084 221818 174136 221824
rect 173348 219292 173400 219298
rect 173348 219234 173400 219240
rect 172886 218512 172942 218521
rect 172886 218447 172942 218456
rect 173256 218204 173308 218210
rect 173256 218146 173308 218152
rect 173268 217138 173296 218146
rect 174096 217138 174124 221818
rect 174912 221740 174964 221746
rect 174912 221682 174964 221688
rect 174924 217138 174952 221682
rect 175568 220969 175596 231662
rect 175752 231662 175950 231690
rect 176304 231662 176594 231690
rect 175752 223582 175780 231662
rect 175740 223576 175792 223582
rect 175740 223518 175792 223524
rect 176304 223174 176332 231662
rect 176752 230172 176804 230178
rect 176752 230114 176804 230120
rect 176764 229094 176792 230114
rect 176672 229066 176792 229094
rect 176672 223530 176700 229066
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 177408 225026 177436 231662
rect 176488 223502 176700 223530
rect 177316 224998 177436 225026
rect 176292 223168 176344 223174
rect 176292 223110 176344 223116
rect 176488 221490 176516 223502
rect 176304 221462 176516 221490
rect 175554 220960 175610 220969
rect 175554 220895 175610 220904
rect 175740 218748 175792 218754
rect 175740 218690 175792 218696
rect 175752 217138 175780 218690
rect 176304 217274 176332 221462
rect 177316 221377 177344 224998
rect 177488 224936 177540 224942
rect 177488 224878 177540 224884
rect 176474 221368 176530 221377
rect 176474 221303 176476 221312
rect 176528 221303 176530 221312
rect 177302 221368 177358 221377
rect 177302 221303 177358 221312
rect 176476 221274 176528 221280
rect 177304 221196 177356 221202
rect 177304 221138 177356 221144
rect 176474 220824 176530 220833
rect 176474 220759 176476 220768
rect 176528 220759 176530 220768
rect 176614 220788 176666 220794
rect 176476 220730 176528 220736
rect 176614 220730 176666 220736
rect 176626 220674 176654 220730
rect 176488 220646 176654 220674
rect 176488 218074 176516 220646
rect 176476 218068 176528 218074
rect 176476 218010 176528 218016
rect 177316 217274 177344 221138
rect 177500 219162 177528 224878
rect 178512 224534 178540 231676
rect 178788 231662 179170 231690
rect 178500 224528 178552 224534
rect 178500 224470 178552 224476
rect 178788 219434 178816 231662
rect 179800 229094 179828 231676
rect 179984 231662 180458 231690
rect 179984 229094 180012 231662
rect 179708 229066 179828 229094
rect 179892 229066 180012 229094
rect 179708 228954 179736 229066
rect 179696 228948 179748 228954
rect 179696 228890 179748 228896
rect 178960 224800 179012 224806
rect 178960 224742 179012 224748
rect 179328 224800 179380 224806
rect 179328 224742 179380 224748
rect 178972 224534 179000 224742
rect 178960 224528 179012 224534
rect 178960 224470 179012 224476
rect 178420 219406 178816 219434
rect 177488 219156 177540 219162
rect 177488 219098 177540 219104
rect 178224 218068 178276 218074
rect 178224 218010 178276 218016
rect 176304 217246 176562 217274
rect 177316 217246 177390 217274
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 168254 217110 168328 217138
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171566 217110 171640 217138
rect 172394 217110 172468 217138
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217110 174952 217138
rect 175706 217110 175780 217138
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217110
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217110
rect 172394 216988 172422 217110
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217110
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 216988 177390 217246
rect 178236 217138 178264 218010
rect 178420 217598 178448 219406
rect 179052 219156 179104 219162
rect 179052 219098 179104 219104
rect 178408 217592 178460 217598
rect 178408 217534 178460 217540
rect 179064 217138 179092 219098
rect 179340 218074 179368 224742
rect 179892 220833 179920 229066
rect 180064 228948 180116 228954
rect 180064 228890 180116 228896
rect 179878 220824 179934 220833
rect 179878 220759 179934 220768
rect 180076 218890 180104 228890
rect 181088 223990 181116 231676
rect 181352 227452 181404 227458
rect 181352 227394 181404 227400
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 180524 220788 180576 220794
rect 180524 220730 180576 220736
rect 180708 220788 180760 220794
rect 180708 220730 180760 220736
rect 180536 220153 180564 220730
rect 180522 220144 180578 220153
rect 180522 220079 180578 220088
rect 180064 218884 180116 218890
rect 180064 218826 180116 218832
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 179328 218068 179380 218074
rect 179328 218010 179380 218016
rect 179892 217138 179920 218146
rect 180720 217274 180748 220730
rect 181168 218748 181220 218754
rect 181168 218690 181220 218696
rect 181180 218346 181208 218690
rect 181364 218482 181392 227394
rect 181732 223446 181760 231676
rect 182376 227594 182404 231676
rect 182652 231662 183034 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181720 223440 181772 223446
rect 181720 223382 181772 223388
rect 181996 223168 182048 223174
rect 181996 223110 182048 223116
rect 181352 218476 181404 218482
rect 181352 218418 181404 218424
rect 182008 218346 182036 223110
rect 182652 221610 182680 231662
rect 183664 223854 183692 231676
rect 184308 230790 184336 231676
rect 184296 230784 184348 230790
rect 184296 230726 184348 230732
rect 184664 229220 184716 229226
rect 184664 229162 184716 229168
rect 183652 223848 183704 223854
rect 183652 223790 183704 223796
rect 184388 223848 184440 223854
rect 184388 223790 184440 223796
rect 183192 223576 183244 223582
rect 183192 223518 183244 223524
rect 182640 221604 182692 221610
rect 182640 221546 182692 221552
rect 182364 219292 182416 219298
rect 182364 219234 182416 219240
rect 181168 218340 181220 218346
rect 181168 218282 181220 218288
rect 181536 218340 181588 218346
rect 181536 218282 181588 218288
rect 181996 218340 182048 218346
rect 181996 218282 182048 218288
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181548 217138 181576 218282
rect 182376 217138 182404 219234
rect 183204 217274 183232 223518
rect 184400 218754 184428 223790
rect 184676 223582 184704 229162
rect 184952 228274 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184940 228268 184992 228274
rect 184940 228210 184992 228216
rect 184664 223576 184716 223582
rect 184664 223518 184716 223524
rect 184848 223440 184900 223446
rect 184848 223382 184900 223388
rect 184662 221776 184718 221785
rect 184662 221711 184718 221720
rect 184676 219434 184704 221711
rect 184676 219406 184796 219434
rect 184388 218748 184440 218754
rect 184388 218690 184440 218696
rect 184020 218340 184072 218346
rect 184020 218282 184072 218288
rect 181502 217110 181576 217138
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 181502 216988 181530 217110
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218282
rect 184768 217274 184796 219406
rect 184860 218362 184888 223382
rect 185136 219842 185164 231662
rect 185400 227588 185452 227594
rect 185400 227530 185452 227536
rect 185412 226914 185440 227530
rect 185584 227316 185636 227322
rect 185584 227258 185636 227264
rect 185596 226914 185624 227258
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185872 222154 185900 231662
rect 186136 227452 186188 227458
rect 186136 227394 186188 227400
rect 185860 222148 185912 222154
rect 185860 222090 185912 222096
rect 185766 221776 185822 221785
rect 185766 221711 185768 221720
rect 185820 221711 185822 221720
rect 185768 221682 185820 221688
rect 185860 221332 185912 221338
rect 185860 221274 185912 221280
rect 185872 221218 185900 221274
rect 185320 221202 185900 221218
rect 185308 221196 185900 221202
rect 185360 221190 185900 221196
rect 185308 221138 185360 221144
rect 185766 220144 185822 220153
rect 185766 220079 185822 220088
rect 185780 219978 185808 220079
rect 185768 219972 185820 219978
rect 185768 219914 185820 219920
rect 185124 219836 185176 219842
rect 185124 219778 185176 219784
rect 184860 218346 184980 218362
rect 186148 218346 186176 227394
rect 186884 223310 186912 231676
rect 187528 227730 187556 231676
rect 188172 230654 188200 231676
rect 188160 230648 188212 230654
rect 188160 230590 188212 230596
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 187700 227724 187752 227730
rect 187700 227666 187752 227672
rect 187712 227458 187740 227666
rect 187700 227452 187752 227458
rect 187700 227394 187752 227400
rect 188816 223718 188844 231676
rect 189092 231662 189474 231690
rect 189092 229094 189120 231662
rect 189092 229066 189304 229094
rect 188804 223712 188856 223718
rect 188804 223654 188856 223660
rect 187332 223576 187384 223582
rect 187332 223518 187384 223524
rect 186872 223304 186924 223310
rect 186872 223246 186924 223252
rect 186504 218476 186556 218482
rect 186504 218418 186556 218424
rect 184860 218340 184992 218346
rect 184860 218334 184940 218340
rect 184940 218282 184992 218288
rect 185676 218340 185728 218346
rect 185676 218282 185728 218288
rect 186136 218340 186188 218346
rect 186136 218282 186188 218288
rect 184768 217246 184842 217274
rect 183986 217110 184060 217138
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218282
rect 186516 217138 186544 218418
rect 187344 217138 187372 223518
rect 188160 223304 188212 223310
rect 188160 223246 188212 223252
rect 188172 217138 188200 223246
rect 188988 218884 189040 218890
rect 188988 218826 189040 218832
rect 189000 217138 189028 218826
rect 189276 217734 189304 229066
rect 189724 228268 189776 228274
rect 189724 228210 189776 228216
rect 189736 219298 189764 228210
rect 190104 228138 190132 231676
rect 190656 231662 190762 231690
rect 190656 229094 190684 231662
rect 190472 229066 190684 229094
rect 190092 228132 190144 228138
rect 190092 228074 190144 228080
rect 189908 227452 189960 227458
rect 189908 227394 189960 227400
rect 189724 219292 189776 219298
rect 189724 219234 189776 219240
rect 189920 219178 189948 227394
rect 190472 219858 190500 229066
rect 191392 222630 191420 231676
rect 191564 223984 191616 223990
rect 191564 223926 191616 223932
rect 191380 222624 191432 222630
rect 191380 222566 191432 222572
rect 190644 219972 190696 219978
rect 190644 219914 190696 219920
rect 190104 219842 190500 219858
rect 190092 219836 190500 219842
rect 190144 219830 190500 219836
rect 190092 219778 190144 219784
rect 189644 219150 189948 219178
rect 189644 218754 189672 219150
rect 189632 218748 189684 218754
rect 189632 218690 189684 218696
rect 189816 218748 189868 218754
rect 189816 218690 189868 218696
rect 189264 217728 189316 217734
rect 189264 217670 189316 217676
rect 189828 217138 189856 218690
rect 190656 217138 190684 219914
rect 191576 217274 191604 223926
rect 192036 222766 192064 231676
rect 192680 227594 192708 231676
rect 192944 228132 192996 228138
rect 192944 228074 192996 228080
rect 192668 227588 192720 227594
rect 192668 227530 192720 227536
rect 192024 222760 192076 222766
rect 192024 222702 192076 222708
rect 192956 219298 192984 228074
rect 193324 221066 193352 231676
rect 193968 226302 193996 231676
rect 193956 226296 194008 226302
rect 193956 226238 194008 226244
rect 194140 226296 194192 226302
rect 194140 226238 194192 226244
rect 193956 222760 194008 222766
rect 193956 222702 194008 222708
rect 193312 221060 193364 221066
rect 193312 221002 193364 221008
rect 192300 219292 192352 219298
rect 192300 219234 192352 219240
rect 192944 219292 192996 219298
rect 192944 219234 192996 219240
rect 193128 219292 193180 219298
rect 193128 219234 193180 219240
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217110 187372 217138
rect 188126 217110 188200 217138
rect 188954 217110 189028 217138
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191604 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217110
rect 188126 216988 188154 217110
rect 188954 216988 188982 217110
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 219234
rect 193140 217138 193168 219234
rect 193968 217138 193996 222702
rect 194152 218890 194180 226238
rect 194612 224126 194640 231676
rect 195060 230648 195112 230654
rect 195060 230590 195112 230596
rect 195072 230042 195100 230590
rect 195060 230036 195112 230042
rect 195060 229978 195112 229984
rect 195256 229094 195284 231676
rect 195900 231062 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197464 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231056 195940 231062
rect 195888 230998 195940 231004
rect 195428 230036 195480 230042
rect 195428 229978 195480 229984
rect 195440 229094 195468 229978
rect 195164 229066 195284 229094
rect 195348 229066 195468 229094
rect 195164 228002 195192 229066
rect 195152 227996 195204 228002
rect 195152 227938 195204 227944
rect 194600 224120 194652 224126
rect 194600 224062 194652 224068
rect 194784 224120 194836 224126
rect 194784 224062 194836 224068
rect 194140 218884 194192 218890
rect 194140 218826 194192 218832
rect 194324 218884 194376 218890
rect 194324 218826 194376 218832
rect 194336 218482 194364 218826
rect 194324 218476 194376 218482
rect 194324 218418 194376 218424
rect 194796 217138 194824 224062
rect 195348 218754 195376 229066
rect 196176 225486 196204 231662
rect 196912 230654 196940 231662
rect 196900 230648 196952 230654
rect 196900 230590 196952 230596
rect 197464 226778 197492 231662
rect 198016 229094 198044 231662
rect 197740 229066 198044 229094
rect 197452 226772 197504 226778
rect 197452 226714 197504 226720
rect 196348 226024 196400 226030
rect 196348 225966 196400 225972
rect 196164 225480 196216 225486
rect 196164 225422 196216 225428
rect 196360 219609 196388 225966
rect 197176 222624 197228 222630
rect 197176 222566 197228 222572
rect 195886 219600 195942 219609
rect 195886 219535 195942 219544
rect 196346 219600 196402 219609
rect 196346 219535 196402 219544
rect 195900 219162 195928 219535
rect 195888 219156 195940 219162
rect 195888 219098 195940 219104
rect 195336 218748 195388 218754
rect 195336 218690 195388 218696
rect 195612 218748 195664 218754
rect 195612 218690 195664 218696
rect 195624 217138 195652 218690
rect 196440 218340 196492 218346
rect 196440 218282 196492 218288
rect 196452 217138 196480 218282
rect 197188 217274 197216 222566
rect 197740 217870 197768 229066
rect 198004 225480 198056 225486
rect 198004 225422 198056 225428
rect 198016 218754 198044 225422
rect 199120 225350 199148 231676
rect 199108 225344 199160 225350
rect 199108 225286 199160 225292
rect 199764 224942 199792 231676
rect 200408 227866 200436 231676
rect 200592 231662 201066 231690
rect 200592 229094 200620 231662
rect 200592 229066 200804 229094
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 227724 200080 227730
rect 200028 227666 200080 227672
rect 200040 225026 200068 227666
rect 200040 224998 200160 225026
rect 199752 224936 199804 224942
rect 199752 224878 199804 224884
rect 199936 224936 199988 224942
rect 199936 224878 199988 224884
rect 199948 224074 199976 224878
rect 200132 224754 200160 224998
rect 199856 224046 199976 224074
rect 200040 224726 200160 224754
rect 199856 223990 199884 224046
rect 199844 223984 199896 223990
rect 199844 223926 199896 223932
rect 200040 219298 200068 224726
rect 200396 222148 200448 222154
rect 200396 222090 200448 222096
rect 198188 219292 198240 219298
rect 198188 219234 198240 219240
rect 198924 219292 198976 219298
rect 198924 219234 198976 219240
rect 200028 219292 200080 219298
rect 200028 219234 200080 219240
rect 198200 218754 198228 219234
rect 198004 218748 198056 218754
rect 198004 218690 198056 218696
rect 198188 218748 198240 218754
rect 198188 218690 198240 218696
rect 198096 218476 198148 218482
rect 198096 218418 198148 218424
rect 197728 217864 197780 217870
rect 197728 217806 197780 217812
rect 197188 217246 197262 217274
rect 192266 217110 192340 217138
rect 193094 217110 193168 217138
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217110
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218418
rect 198936 217138 198964 219234
rect 199752 219156 199804 219162
rect 199752 219098 199804 219104
rect 199764 217138 199792 219098
rect 200408 218482 200436 222090
rect 200776 219570 200804 229066
rect 201696 225078 201724 231676
rect 202340 230314 202368 231676
rect 202998 231662 203196 231690
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202878 229120 202934 229129
rect 202878 229055 202880 229064
rect 202932 229055 202934 229064
rect 202880 229026 202932 229032
rect 203168 226642 203196 231662
rect 203628 230518 203656 231676
rect 203616 230512 203668 230518
rect 203616 230454 203668 230460
rect 203524 227860 203576 227866
rect 203524 227802 203576 227808
rect 203156 226636 203208 226642
rect 203156 226578 203208 226584
rect 203156 225616 203208 225622
rect 203156 225558 203208 225564
rect 203168 225350 203196 225558
rect 203156 225344 203208 225350
rect 203156 225286 203208 225292
rect 201684 225072 201736 225078
rect 201684 225014 201736 225020
rect 202604 225072 202656 225078
rect 202604 225014 202656 225020
rect 201408 223984 201460 223990
rect 201408 223926 201460 223932
rect 201132 219700 201184 219706
rect 201132 219642 201184 219648
rect 200764 219564 200816 219570
rect 200764 219506 200816 219512
rect 201144 219434 201172 219642
rect 200592 219406 201172 219434
rect 200396 218476 200448 218482
rect 200396 218418 200448 218424
rect 200592 217274 200620 219406
rect 201420 217274 201448 223926
rect 202420 220380 202472 220386
rect 202420 220322 202472 220328
rect 202432 219745 202460 220322
rect 202418 219736 202474 219745
rect 202418 219671 202474 219680
rect 202616 219434 202644 225014
rect 202788 220380 202840 220386
rect 202788 220322 202840 220328
rect 202800 219842 202828 220322
rect 202788 219836 202840 219842
rect 202788 219778 202840 219784
rect 203154 219736 203210 219745
rect 203154 219671 203156 219680
rect 203208 219671 203210 219680
rect 203156 219642 203208 219648
rect 202616 219406 202828 219434
rect 202604 219292 202656 219298
rect 202604 219234 202656 219240
rect 202616 218618 202644 219234
rect 202604 218612 202656 218618
rect 202604 218554 202656 218560
rect 202800 218482 202828 219406
rect 203536 219026 203564 227802
rect 204076 227044 204128 227050
rect 204076 226986 204128 226992
rect 204088 226642 204116 226986
rect 204076 226636 204128 226642
rect 204076 226578 204128 226584
rect 203892 225752 203944 225758
rect 203892 225694 203944 225700
rect 203524 219020 203576 219026
rect 203524 218962 203576 218968
rect 203064 218612 203116 218618
rect 203064 218554 203116 218560
rect 202236 218476 202288 218482
rect 202236 218418 202288 218424
rect 202788 218476 202840 218482
rect 202788 218418 202840 218424
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217246 200620 217274
rect 201374 217246 201448 217274
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217246
rect 201374 216988 201402 217246
rect 202248 217138 202276 218418
rect 203076 217138 203104 218554
rect 203904 217274 203932 225694
rect 204272 225214 204300 231676
rect 204720 229084 204772 229090
rect 204720 229026 204772 229032
rect 204732 228138 204760 229026
rect 204720 228132 204772 228138
rect 204720 228074 204772 228080
rect 204916 227882 204944 231676
rect 205192 231662 205574 231690
rect 205836 231662 206218 231690
rect 205192 229129 205220 231662
rect 205178 229120 205234 229129
rect 205178 229055 205234 229064
rect 205456 227996 205508 228002
rect 205456 227938 205508 227944
rect 204548 227854 204944 227882
rect 204548 225894 204576 227854
rect 204904 227724 204956 227730
rect 204904 227666 204956 227672
rect 204916 227458 204944 227666
rect 204720 227452 204772 227458
rect 204720 227394 204772 227400
rect 204904 227452 204956 227458
rect 204904 227394 204956 227400
rect 204732 226778 204760 227394
rect 204720 226772 204772 226778
rect 204720 226714 204772 226720
rect 204732 226358 205128 226386
rect 204536 225888 204588 225894
rect 204536 225830 204588 225836
rect 204732 225758 204760 226358
rect 205100 226302 205128 226358
rect 204904 226296 204956 226302
rect 204904 226238 204956 226244
rect 205088 226296 205140 226302
rect 205088 226238 205140 226244
rect 204916 225894 204944 226238
rect 204904 225888 204956 225894
rect 204904 225830 204956 225836
rect 204720 225752 204772 225758
rect 204720 225694 204772 225700
rect 204904 225752 204956 225758
rect 204904 225694 204956 225700
rect 204916 225486 204944 225694
rect 204904 225480 204956 225486
rect 204904 225422 204956 225428
rect 204260 225208 204312 225214
rect 204260 225150 204312 225156
rect 204536 225208 204588 225214
rect 204536 225150 204588 225156
rect 204548 219434 204576 225150
rect 204904 221468 204956 221474
rect 204904 221410 204956 221416
rect 205088 221468 205140 221474
rect 205088 221410 205140 221416
rect 204916 221202 204944 221410
rect 204904 221196 204956 221202
rect 204904 221138 204956 221144
rect 205100 221066 205128 221410
rect 205088 221060 205140 221066
rect 205088 221002 205140 221008
rect 204536 219428 204588 219434
rect 204536 219370 204588 219376
rect 204720 218476 204772 218482
rect 204720 218418 204772 218424
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218418
rect 205468 217274 205496 227938
rect 205836 219570 205864 231662
rect 206284 230444 206336 230450
rect 206284 230386 206336 230392
rect 205824 219564 205876 219570
rect 205824 219506 205876 219512
rect 206296 219434 206324 230386
rect 206848 222494 206876 231676
rect 207492 223854 207520 231676
rect 208136 226642 208164 231676
rect 208596 231662 208794 231690
rect 208124 226636 208176 226642
rect 208124 226578 208176 226584
rect 207480 223848 207532 223854
rect 207480 223790 207532 223796
rect 207664 223848 207716 223854
rect 207664 223790 207716 223796
rect 206836 222488 206888 222494
rect 206836 222430 206888 222436
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206204 219406 206324 219434
rect 206204 218618 206232 219406
rect 206376 219020 206428 219026
rect 206376 218962 206428 218968
rect 206192 218612 206244 218618
rect 206192 218554 206244 218560
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218962
rect 207216 217274 207244 219642
rect 207676 219298 207704 223790
rect 207848 222488 207900 222494
rect 207848 222430 207900 222436
rect 207664 219292 207716 219298
rect 207664 219234 207716 219240
rect 207860 218482 207888 222430
rect 208596 219570 208624 231662
rect 209424 225350 209452 231676
rect 210068 229498 210096 231676
rect 210424 230308 210476 230314
rect 210424 230250 210476 230256
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 209596 225480 209648 225486
rect 209596 225422 209648 225428
rect 209412 225344 209464 225350
rect 209412 225286 209464 225292
rect 209608 219586 209636 225422
rect 208584 219564 208636 219570
rect 208584 219506 208636 219512
rect 209516 219558 209636 219586
rect 208032 218612 208084 218618
rect 208032 218554 208084 218560
rect 207848 218476 207900 218482
rect 207848 218418 207900 218424
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 208044 217138 208072 218554
rect 209516 218482 209544 219558
rect 210436 219434 210464 230250
rect 210712 228546 210740 231676
rect 211172 231662 211370 231690
rect 210700 228540 210752 228546
rect 210700 228482 210752 228488
rect 210976 227860 211028 227866
rect 210976 227802 211028 227808
rect 209688 219428 209740 219434
rect 209688 219370 209740 219376
rect 210424 219428 210476 219434
rect 210424 219370 210476 219376
rect 208860 218476 208912 218482
rect 208860 218418 208912 218424
rect 209504 218476 209556 218482
rect 209504 218418 209556 218424
rect 208872 217138 208900 218418
rect 209700 217138 209728 219370
rect 210148 218612 210200 218618
rect 210148 218554 210200 218560
rect 210160 218346 210188 218554
rect 210148 218340 210200 218346
rect 210148 218282 210200 218288
rect 210332 218340 210384 218346
rect 210332 218282 210384 218288
rect 210344 218074 210372 218282
rect 210988 218074 211016 227802
rect 211172 221202 211200 231662
rect 212000 222358 212028 231676
rect 212356 229084 212408 229090
rect 212356 229026 212408 229032
rect 212368 228682 212396 229026
rect 212356 228676 212408 228682
rect 212356 228618 212408 228624
rect 212172 226636 212224 226642
rect 212172 226578 212224 226584
rect 211988 222352 212040 222358
rect 211988 222294 212040 222300
rect 211160 221196 211212 221202
rect 211160 221138 211212 221144
rect 211528 221196 211580 221202
rect 211528 221138 211580 221144
rect 211344 219292 211396 219298
rect 211344 219234 211396 219240
rect 210332 218068 210384 218074
rect 210332 218010 210384 218016
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 210528 217138 210556 218010
rect 211356 217138 211384 219234
rect 211540 218482 211568 221138
rect 211712 220108 211764 220114
rect 211712 220050 211764 220056
rect 211724 219570 211752 220050
rect 211712 219564 211764 219570
rect 211712 219506 211764 219512
rect 211528 218476 211580 218482
rect 211528 218418 211580 218424
rect 212184 217274 212212 226578
rect 212644 222902 212672 231676
rect 213288 226506 213316 231676
rect 213946 231662 214144 231690
rect 214116 229094 214144 231662
rect 213920 229084 213972 229090
rect 214116 229066 214328 229094
rect 214576 229090 214604 231676
rect 214748 230036 214800 230042
rect 214748 229978 214800 229984
rect 214760 229634 214788 229978
rect 214748 229628 214800 229634
rect 214748 229570 214800 229576
rect 215220 229362 215248 231676
rect 215208 229356 215260 229362
rect 215208 229298 215260 229304
rect 213920 229026 213972 229032
rect 213276 226500 213328 226506
rect 213276 226442 213328 226448
rect 213932 226250 213960 229026
rect 214104 227044 214156 227050
rect 214104 226986 214156 226992
rect 214116 226778 214144 226986
rect 214104 226772 214156 226778
rect 214104 226714 214156 226720
rect 213472 226222 213960 226250
rect 213472 226166 213500 226222
rect 213460 226160 213512 226166
rect 213460 226102 213512 226108
rect 213644 226160 213696 226166
rect 213644 226102 213696 226108
rect 213656 225894 213684 226102
rect 213644 225888 213696 225894
rect 213644 225830 213696 225836
rect 212632 222896 212684 222902
rect 212632 222838 212684 222844
rect 213184 222896 213236 222902
rect 213184 222838 213236 222844
rect 213000 219428 213052 219434
rect 213000 219370 213052 219376
rect 207998 217110 208072 217138
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217110 210556 217138
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 207998 216988 208026 217110
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217110
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 219370
rect 213196 218346 213224 222838
rect 213828 220244 213880 220250
rect 213828 220186 213880 220192
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 220186
rect 214300 220114 214328 229066
rect 214564 229084 214616 229090
rect 214564 229026 214616 229032
rect 214748 229084 214800 229090
rect 214748 229026 214800 229032
rect 214564 228404 214616 228410
rect 214564 228346 214616 228352
rect 214576 228138 214604 228346
rect 214564 228132 214616 228138
rect 214564 228074 214616 228080
rect 214760 228002 214788 229026
rect 215864 228546 215892 231676
rect 216048 231662 216522 231690
rect 215852 228540 215904 228546
rect 215852 228482 215904 228488
rect 214748 227996 214800 228002
rect 214748 227938 214800 227944
rect 214748 227588 214800 227594
rect 214748 227530 214800 227536
rect 214932 227588 214984 227594
rect 214932 227530 214984 227536
rect 214760 226914 214788 227530
rect 214748 226908 214800 226914
rect 214748 226850 214800 226856
rect 214944 226642 214972 227530
rect 214932 226636 214984 226642
rect 214932 226578 214984 226584
rect 215208 225208 215260 225214
rect 215208 225150 215260 225156
rect 214564 220380 214616 220386
rect 214564 220322 214616 220328
rect 214576 220114 214604 220322
rect 214288 220108 214340 220114
rect 214288 220050 214340 220056
rect 214564 220108 214616 220114
rect 214564 220050 214616 220056
rect 215220 218074 215248 225150
rect 216048 224954 216076 231662
rect 216220 228540 216272 228546
rect 216220 228482 216272 228488
rect 216232 224954 216260 228482
rect 216404 226500 216456 226506
rect 216404 226442 216456 226448
rect 216416 224954 216444 226442
rect 217152 225622 217180 231676
rect 217508 228132 217560 228138
rect 217508 228074 217560 228080
rect 217140 225616 217192 225622
rect 217140 225558 217192 225564
rect 215956 224926 216076 224954
rect 216140 224926 216260 224954
rect 216324 224926 216444 224954
rect 215956 219570 215984 224926
rect 215944 219564 215996 219570
rect 215944 219506 215996 219512
rect 216140 218074 216168 224926
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 216128 218068 216180 218074
rect 216128 218010 216180 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217274 216352 224926
rect 217140 220244 217192 220250
rect 217140 220186 217192 220192
rect 217152 217274 217180 220186
rect 217520 219434 217548 228074
rect 217796 227730 217824 231676
rect 218152 228812 218204 228818
rect 218152 228754 218204 228760
rect 218164 228410 218192 228754
rect 218152 228404 218204 228410
rect 218152 228346 218204 228352
rect 217784 227724 217836 227730
rect 217784 227666 217836 227672
rect 218440 226778 218468 231676
rect 218428 226772 218480 226778
rect 218428 226714 218480 226720
rect 219084 223038 219112 231676
rect 219636 231662 219742 231690
rect 219440 228132 219492 228138
rect 219440 228074 219492 228080
rect 219452 227730 219480 228074
rect 219440 227724 219492 227730
rect 219440 227666 219492 227672
rect 219438 227488 219494 227497
rect 219438 227423 219494 227432
rect 219452 227322 219480 227423
rect 219440 227316 219492 227322
rect 219440 227258 219492 227264
rect 219348 226772 219400 226778
rect 219348 226714 219400 226720
rect 219072 223032 219124 223038
rect 219072 222974 219124 222980
rect 218060 221060 218112 221066
rect 218060 221002 218112 221008
rect 217336 219406 217548 219434
rect 217336 218618 217364 219406
rect 218072 219298 218100 221002
rect 218060 219292 218112 219298
rect 218060 219234 218112 219240
rect 217324 218612 217376 218618
rect 217324 218554 217376 218560
rect 217968 218476 218020 218482
rect 217968 218418 218020 218424
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217246 216352 217274
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217246
rect 217106 216988 217134 217246
rect 217980 217138 218008 218418
rect 219360 218074 219388 226714
rect 219636 220930 219664 231662
rect 220084 230036 220136 230042
rect 220084 229978 220136 229984
rect 220096 229770 220124 229978
rect 220084 229764 220136 229770
rect 220084 229706 220136 229712
rect 220372 229498 220400 231676
rect 220360 229492 220412 229498
rect 220360 229434 220412 229440
rect 220636 229492 220688 229498
rect 220636 229434 220688 229440
rect 219900 228948 219952 228954
rect 219900 228890 219952 228896
rect 219912 228138 219940 228890
rect 220176 228540 220228 228546
rect 220176 228482 220228 228488
rect 219900 228132 219952 228138
rect 219900 228074 219952 228080
rect 220188 227882 220216 228482
rect 220096 227866 220216 227882
rect 220084 227860 220216 227866
rect 220136 227854 220216 227860
rect 220084 227802 220136 227808
rect 220452 227724 220504 227730
rect 220452 227666 220504 227672
rect 220464 227497 220492 227666
rect 220450 227488 220506 227497
rect 220450 227423 220506 227432
rect 219808 227316 219860 227322
rect 219808 227258 219860 227264
rect 219820 226914 219848 227258
rect 220268 227180 220320 227186
rect 220268 227122 220320 227128
rect 220280 226914 220308 227122
rect 219808 226908 219860 226914
rect 219808 226850 219860 226856
rect 220268 226908 220320 226914
rect 220268 226850 220320 226856
rect 220452 226636 220504 226642
rect 220452 226578 220504 226584
rect 220084 226160 220136 226166
rect 220084 226102 220136 226108
rect 220096 225894 220124 226102
rect 220084 225888 220136 225894
rect 220084 225830 220136 225836
rect 220084 225616 220136 225622
rect 220084 225558 220136 225564
rect 220096 225214 220124 225558
rect 220084 225208 220136 225214
rect 220084 225150 220136 225156
rect 219624 220924 219676 220930
rect 219624 220866 219676 220872
rect 219624 218612 219676 218618
rect 219624 218554 219676 218560
rect 218796 218068 218848 218074
rect 218796 218010 218848 218016
rect 219348 218068 219400 218074
rect 219348 218010 219400 218016
rect 218808 217138 218836 218010
rect 219636 217138 219664 218554
rect 220464 217274 220492 226578
rect 220648 226506 220676 229434
rect 221016 228002 221044 231676
rect 221292 231662 221674 231690
rect 222212 231662 222318 231690
rect 221004 227996 221056 228002
rect 221004 227938 221056 227944
rect 220636 226500 220688 226506
rect 220636 226442 220688 226448
rect 220636 222012 220688 222018
rect 220636 221954 220688 221960
rect 220820 222012 220872 222018
rect 220820 221954 220872 221960
rect 220648 220930 220676 221954
rect 220832 221474 220860 221954
rect 220820 221468 220872 221474
rect 220820 221410 220872 221416
rect 221004 221468 221056 221474
rect 221004 221410 221056 221416
rect 221016 221066 221044 221410
rect 221004 221060 221056 221066
rect 221004 221002 221056 221008
rect 220636 220924 220688 220930
rect 220636 220866 220688 220872
rect 221292 220658 221320 231662
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221280 220652 221332 220658
rect 221280 220594 221332 220600
rect 221844 218074 221872 226442
rect 222016 226160 222068 226166
rect 222016 226102 222068 226108
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 226102
rect 222212 222018 222240 231662
rect 222948 225350 222976 231676
rect 223592 227730 223620 231676
rect 223776 231662 224250 231690
rect 223580 227724 223632 227730
rect 223580 227666 223632 227672
rect 222936 225344 222988 225350
rect 222936 225286 222988 225292
rect 222200 222012 222252 222018
rect 222200 221954 222252 221960
rect 223488 220924 223540 220930
rect 223488 220866 223540 220872
rect 223500 218482 223528 220866
rect 223776 220658 223804 231662
rect 224592 227792 224644 227798
rect 224592 227734 224644 227740
rect 223764 220652 223816 220658
rect 223764 220594 223816 220600
rect 223764 220516 223816 220522
rect 223764 220458 223816 220464
rect 223488 218476 223540 218482
rect 223488 218418 223540 218424
rect 222936 218340 222988 218346
rect 222936 218282 222988 218288
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218282
rect 223776 217274 223804 220458
rect 224604 217274 224632 227734
rect 224880 224670 224908 231676
rect 225524 229906 225552 231676
rect 225512 229900 225564 229906
rect 225512 229842 225564 229848
rect 226168 229094 226196 231676
rect 225800 229066 226196 229094
rect 226536 231662 226826 231690
rect 227088 231662 227470 231690
rect 225800 228138 225828 229066
rect 225788 228132 225840 228138
rect 225788 228074 225840 228080
rect 225972 228132 226024 228138
rect 225972 228074 226024 228080
rect 225604 226772 225656 226778
rect 225604 226714 225656 226720
rect 224868 224664 224920 224670
rect 224868 224606 224920 224612
rect 225616 218210 225644 226714
rect 225984 219434 226012 228074
rect 226536 221066 226564 231662
rect 226708 227724 226760 227730
rect 226708 227666 226760 227672
rect 226720 226642 226748 227666
rect 226708 226636 226760 226642
rect 226708 226578 226760 226584
rect 227088 224398 227116 231662
rect 227536 224664 227588 224670
rect 227536 224606 227588 224612
rect 227076 224392 227128 224398
rect 227076 224334 227128 224340
rect 226524 221060 226576 221066
rect 226524 221002 226576 221008
rect 225984 219406 226196 219434
rect 225972 218476 226024 218482
rect 225972 218418 226024 218424
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217246 223804 217274
rect 224558 217246 224632 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217246
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218418
rect 226168 218074 226196 219406
rect 227548 218074 227576 224606
rect 228100 223854 228128 231676
rect 228744 227050 228772 231676
rect 229296 231662 229402 231690
rect 228732 227044 228784 227050
rect 228732 226986 228784 226992
rect 228916 227044 228968 227050
rect 228916 226986 228968 226992
rect 228928 226506 228956 226986
rect 228916 226500 228968 226506
rect 228916 226442 228968 226448
rect 228732 224392 228784 224398
rect 228732 224334 228784 224340
rect 228088 223848 228140 223854
rect 228088 223790 228140 223796
rect 227904 221060 227956 221066
rect 227904 221002 227956 221008
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227076 218068 227128 218074
rect 227076 218010 227128 218016
rect 227536 218068 227588 218074
rect 227536 218010 227588 218016
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227088 217138 227116 218010
rect 227916 217274 227944 221002
rect 228744 217274 228772 224334
rect 229296 220114 229324 231662
rect 230032 224262 230060 231676
rect 230676 230042 230704 231676
rect 230664 230036 230716 230042
rect 230664 229978 230716 229984
rect 230480 229900 230532 229906
rect 230480 229842 230532 229848
rect 230020 224256 230072 224262
rect 230492 224210 230520 229842
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230020 224198 230072 224204
rect 230400 224182 230520 224210
rect 229284 220108 229336 220114
rect 229284 220050 229336 220056
rect 230204 220108 230256 220114
rect 230204 220050 230256 220056
rect 230216 219434 230244 220050
rect 230216 219406 230336 219434
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 227042 217110 227116 217138
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217110
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230308 217274 230336 219406
rect 230400 218090 230428 224182
rect 231136 219434 231164 229434
rect 231320 228410 231348 231676
rect 231308 228404 231360 228410
rect 231308 228346 231360 228352
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231044 219406 231164 219434
rect 231044 218346 231072 219406
rect 231032 218340 231084 218346
rect 231032 218282 231084 218288
rect 230400 218074 230520 218090
rect 231688 218074 231716 224198
rect 231964 221882 231992 231676
rect 232608 224534 232636 231676
rect 233252 229094 233280 231676
rect 233896 229094 233924 231676
rect 233252 229066 233372 229094
rect 232596 224528 232648 224534
rect 232596 224470 232648 224476
rect 233148 224528 233200 224534
rect 233148 224470 233200 224476
rect 232136 222012 232188 222018
rect 232136 221954 232188 221960
rect 231952 221876 232004 221882
rect 231952 221818 232004 221824
rect 232148 221610 232176 221954
rect 232136 221604 232188 221610
rect 232136 221546 232188 221552
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 230400 218068 230532 218074
rect 230400 218062 230480 218068
rect 230480 218010 230532 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217138 232912 218282
rect 233160 218074 233188 224470
rect 233344 222902 233372 229066
rect 233712 229066 233924 229094
rect 234172 231662 234554 231690
rect 234724 231662 235198 231690
rect 234172 229094 234200 231662
rect 234172 229066 234292 229094
rect 233712 227186 233740 229066
rect 233884 228404 233936 228410
rect 233884 228346 233936 228352
rect 233896 227866 233924 228346
rect 233884 227860 233936 227866
rect 233884 227802 233936 227808
rect 233700 227180 233752 227186
rect 233700 227122 233752 227128
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 221876 233752 221882
rect 233700 221818 233752 221824
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221818
rect 234068 221468 234120 221474
rect 234068 221410 234120 221416
rect 234080 221066 234108 221410
rect 234264 221338 234292 229066
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234252 221332 234304 221338
rect 234252 221274 234304 221280
rect 234068 221060 234120 221066
rect 234068 221002 234120 221008
rect 234540 217274 234568 222838
rect 234724 222018 234752 231662
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 227180 235868 227186
rect 235816 227122 235868 227128
rect 234712 222012 234764 222018
rect 234712 221954 234764 221960
rect 235828 218074 235856 227122
rect 236472 226030 236500 231676
rect 236748 231662 237130 231690
rect 236460 226024 236512 226030
rect 236460 225966 236512 225972
rect 236748 220794 236776 231662
rect 237760 224806 237788 231676
rect 238404 226778 238432 231676
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238392 226772 238444 226778
rect 238392 226714 238444 226720
rect 237748 224800 237800 224806
rect 237748 224742 237800 224748
rect 237012 222352 237064 222358
rect 237012 222294 237064 222300
rect 236736 220788 236788 220794
rect 236736 220730 236788 220736
rect 236184 220652 236236 220658
rect 236184 220594 236236 220600
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217110 232912 217138
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217110
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217274 236224 220594
rect 237024 217274 237052 222294
rect 237840 221332 237892 221338
rect 237840 221274 237892 221280
rect 237852 217274 237880 221274
rect 235322 217110 235396 217138
rect 236150 217246 236224 217274
rect 236978 217246 237052 217274
rect 237806 217246 237880 217274
rect 238588 217274 238616 228754
rect 239048 228274 239076 231676
rect 239036 228268 239088 228274
rect 239036 228210 239088 228216
rect 239312 227860 239364 227866
rect 239312 227802 239364 227808
rect 239324 218890 239352 227802
rect 239692 223446 239720 231676
rect 239680 223440 239732 223446
rect 239680 223382 239732 223388
rect 240336 223174 240364 231676
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227322 241652 231676
rect 241612 227316 241664 227322
rect 241612 227258 241664 227264
rect 241152 226772 241204 226778
rect 241152 226714 241204 226720
rect 240324 223168 240376 223174
rect 240324 223110 240376 223116
rect 239496 219292 239548 219298
rect 239496 219234 239548 219240
rect 239312 218884 239364 218890
rect 239312 218826 239364 218832
rect 238588 217246 238662 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217246
rect 236978 216988 237006 217246
rect 237806 216988 237834 217246
rect 238634 216988 238662 217246
rect 239508 217138 239536 219234
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 226714
rect 242268 223582 242296 231676
rect 242926 231662 243124 231690
rect 242532 230036 242584 230042
rect 242532 229978 242584 229984
rect 242544 229094 242572 229978
rect 242544 229066 242756 229094
rect 242256 223576 242308 223582
rect 242256 223518 242308 223524
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 241980 218204 242032 218210
rect 241980 218146 242032 218152
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 218146
rect 242728 217274 242756 229066
rect 242900 225344 242952 225350
rect 242820 225292 242900 225298
rect 242820 225286 242952 225292
rect 242820 225270 242940 225286
rect 242820 218226 242848 225270
rect 243096 221746 243124 231662
rect 243556 227866 243584 231676
rect 243544 227860 243596 227866
rect 243544 227802 243596 227808
rect 244200 225894 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244188 225888 244240 225894
rect 244188 225830 244240 225836
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243084 221740 243136 221746
rect 243084 221682 243136 221688
rect 243728 221604 243780 221610
rect 243728 221546 243780 221552
rect 243740 221338 243768 221546
rect 243728 221332 243780 221338
rect 243728 221274 243780 221280
rect 243544 219156 243596 219162
rect 243544 219098 243596 219104
rect 242820 218210 242940 218226
rect 243556 218210 243584 219098
rect 242820 218204 242952 218210
rect 242820 218198 242900 218204
rect 242900 218146 242952 218152
rect 243544 218204 243596 218210
rect 243544 218146 243596 218152
rect 244108 218074 244136 223382
rect 244476 219978 244504 231662
rect 245120 223310 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229356 246540 229362
rect 246488 229298 246540 229304
rect 246304 227860 246356 227866
rect 246304 227802 246356 227808
rect 245476 223848 245528 223854
rect 245476 223790 245528 223796
rect 245108 223304 245160 223310
rect 245108 223246 245160 223252
rect 245292 223032 245344 223038
rect 245292 222974 245344 222980
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 245304 218074 245332 222974
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 245292 218068 245344 218074
rect 245292 218010 245344 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217138 244504 218010
rect 245488 217274 245516 223790
rect 246120 218884 246172 218890
rect 246120 218826 246172 218832
rect 243602 217110 243676 217138
rect 244430 217110 244504 217138
rect 245258 217246 245516 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 218826
rect 246316 218754 246344 227802
rect 246500 220658 246528 229298
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 247420 222766 247448 231676
rect 248064 224942 248092 231676
rect 248708 227866 248736 231676
rect 248984 231662 249366 231690
rect 248984 229094 249012 231662
rect 248892 229066 249012 229094
rect 248696 227860 248748 227866
rect 248696 227802 248748 227808
rect 248892 225758 248920 229066
rect 249064 227860 249116 227866
rect 249064 227802 249116 227808
rect 248880 225752 248932 225758
rect 248880 225694 248932 225700
rect 248052 224936 248104 224942
rect 248052 224878 248104 224884
rect 248328 224800 248380 224806
rect 248328 224742 248380 224748
rect 247408 222760 247460 222766
rect 247408 222702 247460 222708
rect 246488 220652 246540 220658
rect 246488 220594 246540 220600
rect 246948 220652 247000 220658
rect 246948 220594 247000 220600
rect 246304 218748 246356 218754
rect 246304 218690 246356 218696
rect 246960 217274 246988 220594
rect 248340 218074 248368 224742
rect 249076 218210 249104 227802
rect 249248 227316 249300 227322
rect 249248 227258 249300 227264
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249260 218074 249288 227258
rect 249432 223576 249484 223582
rect 249432 223518 249484 223524
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248328 218068 248380 218074
rect 248328 218010 248380 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 249248 218068 249300 218074
rect 249248 218010 249300 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217274 249472 223518
rect 249996 222630 250024 231676
rect 250640 224126 250668 231676
rect 251284 228002 251312 231676
rect 251272 227996 251324 228002
rect 251272 227938 251324 227944
rect 251928 227458 251956 231676
rect 252586 231662 252784 231690
rect 251916 227452 251968 227458
rect 251916 227394 251968 227400
rect 252468 226024 252520 226030
rect 252468 225966 252520 225972
rect 251088 225752 251140 225758
rect 251088 225694 251140 225700
rect 250628 224120 250680 224126
rect 250628 224062 250680 224068
rect 250904 223304 250956 223310
rect 250904 223246 250956 223252
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 250916 218074 250944 223246
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217246 249472 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217246
rect 250272 217138 250300 218010
rect 251100 217274 251128 225694
rect 252480 218074 252508 225966
rect 252756 219842 252784 231662
rect 252940 231662 253230 231690
rect 252940 222154 252968 231662
rect 253860 227866 253888 231676
rect 253848 227860 253900 227866
rect 253848 227802 253900 227808
rect 254504 225078 254532 231676
rect 254952 228268 255004 228274
rect 254952 228210 255004 228216
rect 254492 225072 254544 225078
rect 254492 225014 254544 225020
rect 252928 222148 252980 222154
rect 252928 222090 252980 222096
rect 253848 220924 253900 220930
rect 253848 220866 253900 220872
rect 253572 219972 253624 219978
rect 253572 219914 253624 219920
rect 252744 219836 252796 219842
rect 252744 219778 252796 219784
rect 252744 218748 252796 218754
rect 252744 218690 252796 218696
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218690
rect 253584 217274 253612 219914
rect 253860 219026 253888 220866
rect 254400 220788 254452 220794
rect 254400 220730 254452 220736
rect 253848 219020 253900 219026
rect 253848 218962 253900 218968
rect 254412 217274 254440 220730
rect 254964 219434 254992 228210
rect 255148 226302 255176 231676
rect 255136 226296 255188 226302
rect 255136 226238 255188 226244
rect 255792 223990 255820 231676
rect 256436 230450 256464 231676
rect 256424 230444 256476 230450
rect 256424 230386 256476 230392
rect 256516 229764 256568 229770
rect 256516 229706 256568 229712
rect 255780 223984 255832 223990
rect 255780 223926 255832 223932
rect 254964 219406 255176 219434
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 254366 217246 254440 217274
rect 255148 217274 255176 219406
rect 256528 218074 256556 229706
rect 257080 229090 257108 231676
rect 257264 231662 257738 231690
rect 257068 229084 257120 229090
rect 257068 229026 257120 229032
rect 257264 219706 257292 231662
rect 257896 229084 257948 229090
rect 257896 229026 257948 229032
rect 257712 228948 257764 228954
rect 257712 228890 257764 228896
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 255148 217246 255222 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254366 216988 254394 217246
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 228890
rect 257908 218074 257936 229026
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 258092 219434 258120 222090
rect 258644 220930 258672 231662
rect 259368 227452 259420 227458
rect 259368 227394 259420 227400
rect 258632 220924 258684 220930
rect 258632 220866 258684 220872
rect 258080 219428 258132 219434
rect 258080 219370 258132 219376
rect 259184 219020 259236 219026
rect 259184 218962 259236 218968
rect 257896 218068 257948 218074
rect 257896 218010 257948 218016
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259196 217274 259224 218962
rect 259380 218074 259408 227394
rect 259656 225486 259684 231676
rect 260300 228546 260328 231676
rect 260944 229094 260972 231676
rect 261588 230314 261616 231676
rect 261576 230308 261628 230314
rect 261576 230250 261628 230256
rect 260852 229066 260972 229094
rect 260288 228540 260340 228546
rect 260288 228482 260340 228488
rect 260656 226296 260708 226302
rect 260656 226238 260708 226244
rect 259644 225480 259696 225486
rect 259644 225422 259696 225428
rect 260668 219434 260696 226238
rect 260852 221202 260880 229066
rect 262232 227594 262260 231676
rect 262416 231662 262890 231690
rect 263152 231662 263534 231690
rect 263888 231662 264178 231690
rect 262220 227588 262272 227594
rect 262220 227530 262272 227536
rect 261852 225888 261904 225894
rect 261852 225830 261904 225836
rect 261024 222012 261076 222018
rect 261024 221954 261076 221960
rect 260840 221196 260892 221202
rect 260840 221138 260892 221144
rect 260668 219406 260788 219434
rect 260760 218074 260788 219406
rect 259368 218068 259420 218074
rect 259368 218010 259420 218016
rect 260196 218068 260248 218074
rect 260196 218010 260248 218016
rect 260748 218068 260800 218074
rect 260748 218010 260800 218016
rect 259196 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260208 217138 260236 218010
rect 261036 217274 261064 221954
rect 261864 217274 261892 225830
rect 262416 220386 262444 231662
rect 263152 221746 263180 231662
rect 263888 222154 263916 231662
rect 264244 230172 264296 230178
rect 264244 230114 264296 230120
rect 263876 222148 263928 222154
rect 263876 222090 263928 222096
rect 263140 221740 263192 221746
rect 263140 221682 263192 221688
rect 263508 221740 263560 221746
rect 263508 221682 263560 221688
rect 262404 220380 262456 220386
rect 262404 220322 262456 220328
rect 262680 220380 262732 220386
rect 262680 220322 262732 220328
rect 262692 217274 262720 220322
rect 263520 217274 263548 221682
rect 264256 220386 264284 230114
rect 264808 228682 264836 231676
rect 265176 231662 265466 231690
rect 264796 228676 264848 228682
rect 264796 228618 264848 228624
rect 264796 227588 264848 227594
rect 264796 227530 264848 227536
rect 264244 220380 264296 220386
rect 264244 220322 264296 220328
rect 264612 220380 264664 220386
rect 264612 220322 264664 220328
rect 264624 218618 264652 220322
rect 264612 218612 264664 218618
rect 264612 218554 264664 218560
rect 264808 218074 264836 227530
rect 265176 220250 265204 231662
rect 266096 225622 266124 231676
rect 266740 229634 266768 231676
rect 266728 229628 266780 229634
rect 266728 229570 266780 229576
rect 267384 226914 267412 231676
rect 268028 227730 268056 231676
rect 268212 231662 268686 231690
rect 268016 227724 268068 227730
rect 268016 227666 268068 227672
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 266084 225616 266136 225622
rect 266084 225558 266136 225564
rect 267004 225616 267056 225622
rect 267004 225558 267056 225564
rect 266268 224936 266320 224942
rect 266268 224878 266320 224884
rect 265164 220244 265216 220250
rect 265164 220186 265216 220192
rect 265992 218612 266044 218618
rect 265992 218554 266044 218560
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 260162 217110 260236 217138
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 262646 217246 262720 217274
rect 263474 217246 263548 217274
rect 260162 216988 260190 217110
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262646 216988 262674 217246
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 218554
rect 266280 218074 266308 224878
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266832 217274 266860 221274
rect 267016 218482 267044 225558
rect 268212 221066 268240 231662
rect 268936 228540 268988 228546
rect 268936 228482 268988 228488
rect 268200 221060 268252 221066
rect 268200 221002 268252 221008
rect 267648 220244 267700 220250
rect 267648 220186 267700 220192
rect 267004 218476 267056 218482
rect 267004 218418 267056 218424
rect 267660 217274 267688 220186
rect 268948 218074 268976 228482
rect 269316 220386 269344 231676
rect 269960 226166 269988 231676
rect 269948 226160 270000 226166
rect 269948 226102 270000 226108
rect 270224 226160 270276 226166
rect 270224 226102 270276 226108
rect 270040 222148 270092 222154
rect 270040 222090 270092 222096
rect 269304 220380 269356 220386
rect 269304 220322 269356 220328
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270052 217274 270080 222090
rect 270236 218074 270264 226102
rect 270604 220522 270632 231676
rect 271248 227050 271276 231676
rect 271892 229498 271920 231676
rect 271880 229492 271932 229498
rect 271880 229434 271932 229440
rect 272536 228138 272564 231676
rect 273180 229094 273208 231676
rect 272720 229066 273208 229094
rect 272524 228132 272576 228138
rect 272524 228074 272576 228080
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 220516 270644 220522
rect 270592 220458 270644 220464
rect 270776 219836 270828 219842
rect 270776 219778 270828 219784
rect 270788 218346 270816 219778
rect 270776 218340 270828 218346
rect 270776 218282 270828 218288
rect 270224 218068 270276 218074
rect 270224 218010 270276 218016
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 270052 217246 270126 217274
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272720 224754 272748 229066
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274272 228404 274324 228410
rect 274272 228346 274324 228352
rect 272352 224726 272748 224754
rect 272352 224670 272380 224726
rect 272340 224664 272392 224670
rect 272340 224606 272392 224612
rect 272524 224664 272576 224670
rect 272524 224606 272576 224612
rect 272340 224528 272392 224534
rect 272340 224470 272392 224476
rect 272352 224262 272380 224470
rect 272340 224256 272392 224262
rect 272340 224198 272392 224204
rect 272340 219156 272392 219162
rect 272340 219098 272392 219104
rect 272352 218618 272380 219098
rect 272340 218612 272392 218618
rect 272340 218554 272392 218560
rect 272536 218074 272564 224606
rect 273444 220380 273496 220386
rect 273444 220322 273496 220328
rect 272892 219428 272944 219434
rect 272892 219370 272944 219376
rect 272708 219292 272760 219298
rect 272708 219234 272760 219240
rect 272720 218618 272748 219234
rect 272708 218612 272760 218618
rect 272708 218554 272760 218560
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 272904 217274 272932 219370
rect 273456 217274 273484 220322
rect 274284 217274 274312 228346
rect 274468 225622 274496 231676
rect 274456 225616 274508 225622
rect 274456 225558 274508 225564
rect 275112 224534 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 224528 275152 224534
rect 275100 224470 275152 224476
rect 275100 224392 275152 224398
rect 275100 224334 275152 224340
rect 275112 217274 275140 224334
rect 275296 220114 275324 231662
rect 275652 230308 275704 230314
rect 275652 230250 275704 230256
rect 275664 229094 275692 230250
rect 275664 229066 275876 229094
rect 275284 220108 275336 220114
rect 275284 220050 275336 220056
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272582 217246 272932 217274
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 277044 229906 277072 231676
rect 277032 229900 277084 229906
rect 277032 229842 277084 229848
rect 276296 229628 276348 229634
rect 276296 229570 276348 229576
rect 276308 223582 276336 229570
rect 277688 224262 277716 231676
rect 277964 231662 278346 231690
rect 277676 224256 277728 224262
rect 277676 224198 277728 224204
rect 276296 223576 276348 223582
rect 276296 223518 276348 223524
rect 277964 221882 277992 231662
rect 278412 225616 278464 225622
rect 278412 225558 278464 225564
rect 277952 221876 278004 221882
rect 277952 221818 278004 221824
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 276756 220516 276808 220522
rect 276756 220458 276808 220464
rect 276768 217274 276796 220458
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276722 217246 276796 217274
rect 276722 216988 276750 217246
rect 277596 217138 277624 218010
rect 278424 217274 278452 225558
rect 278976 224126 279004 231676
rect 279160 231662 279634 231690
rect 278964 224120 279016 224126
rect 278964 224062 279016 224068
rect 278596 223576 278648 223582
rect 278596 223518 278648 223524
rect 278608 218074 278636 223518
rect 279160 219842 279188 231662
rect 280264 227186 280292 231676
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 279424 224052 279476 224058
rect 279424 223994 279476 224000
rect 279148 219836 279200 219842
rect 279148 219778 279200 219784
rect 279056 219292 279108 219298
rect 279056 219234 279108 219240
rect 279068 218890 279096 219234
rect 279056 218884 279108 218890
rect 279056 218826 279108 218832
rect 279240 218884 279292 218890
rect 279240 218826 279292 218832
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218826
rect 279436 218618 279464 223994
rect 280908 222358 280936 231676
rect 281356 227180 281408 227186
rect 281356 227122 281408 227128
rect 280896 222352 280948 222358
rect 280896 222294 280948 222300
rect 280068 221876 280120 221882
rect 280068 221818 280120 221824
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 280080 217274 280108 221818
rect 281368 219434 281396 227122
rect 281552 222902 281580 231676
rect 282196 229362 282224 231676
rect 282552 229900 282604 229906
rect 282552 229842 282604 229848
rect 282184 229356 282236 229362
rect 282184 229298 282236 229304
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282564 217274 282592 229842
rect 282840 228818 282868 231676
rect 282828 228812 282880 228818
rect 282828 228754 282880 228760
rect 283484 223174 283512 231676
rect 283760 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 282736 222896 282788 222902
rect 282736 222838 282788 222844
rect 282748 218074 282776 222838
rect 283760 221610 283788 231662
rect 284772 224058 284800 231676
rect 285048 231662 285430 231690
rect 285048 225350 285076 231662
rect 285496 228676 285548 228682
rect 285496 228618 285548 228624
rect 285036 225344 285088 225350
rect 285036 225286 285088 225292
rect 284760 224052 284812 224058
rect 284760 223994 284812 224000
rect 284208 222760 284260 222766
rect 284208 222702 284260 222708
rect 283748 221604 283800 221610
rect 283748 221546 283800 221552
rect 284024 221468 284076 221474
rect 284024 221410 284076 221416
rect 284036 219434 284064 221410
rect 284036 219406 284156 219434
rect 282736 218068 282788 218074
rect 282736 218010 282788 218016
rect 283380 218068 283432 218074
rect 283380 218010 283432 218016
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282592 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283392 217138 283420 218010
rect 284128 217274 284156 219406
rect 284220 218090 284248 222702
rect 284220 218074 284340 218090
rect 285508 218074 285536 228618
rect 286060 223446 286088 231676
rect 286704 226778 286732 231676
rect 287060 230444 287112 230450
rect 287060 230386 287112 230392
rect 286692 226772 286744 226778
rect 286692 226714 286744 226720
rect 287072 226166 287100 230386
rect 287348 230042 287376 231676
rect 287624 231662 288006 231690
rect 287336 230036 287388 230042
rect 287336 229978 287388 229984
rect 287060 226160 287112 226166
rect 287060 226102 287112 226108
rect 286324 224528 286376 224534
rect 286324 224470 286376 224476
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 286336 219298 286364 224470
rect 287624 223854 287652 231662
rect 288072 226160 288124 226166
rect 288072 226102 288124 226108
rect 287612 223848 287664 223854
rect 287612 223790 287664 223796
rect 286692 219836 286744 219842
rect 286692 219778 286744 219784
rect 286324 219292 286376 219298
rect 286324 219234 286376 219240
rect 285864 218884 285916 218890
rect 285864 218826 285916 218832
rect 284220 218068 284352 218074
rect 284220 218062 284300 218068
rect 284300 218010 284352 218016
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 283346 217110 283420 217138
rect 283346 216988 283374 217110
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 218826
rect 286704 217274 286732 219778
rect 288084 218074 288112 226102
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 288072 218068 288124 218074
rect 288072 218010 288124 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288636 220658 288664 231676
rect 288992 223304 289044 223310
rect 288992 223246 289044 223252
rect 288624 220652 288676 220658
rect 288624 220594 288676 220600
rect 289004 218482 289032 223246
rect 289280 223038 289308 231676
rect 289924 224534 289952 231676
rect 290568 227322 290596 231676
rect 290556 227316 290608 227322
rect 290556 227258 290608 227264
rect 291016 227316 291068 227322
rect 291016 227258 291068 227264
rect 289912 224528 289964 224534
rect 289912 224470 289964 224476
rect 290832 224528 290884 224534
rect 290832 224470 290884 224476
rect 289728 224256 289780 224262
rect 289728 224198 289780 224204
rect 289268 223032 289320 223038
rect 289268 222974 289320 222980
rect 288992 218476 289044 218482
rect 288992 218418 289044 218424
rect 289740 218074 289768 224198
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289728 218068 289780 218074
rect 289728 218010 289780 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224470
rect 291028 219434 291056 227258
rect 291212 223446 291240 231676
rect 291856 224806 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 293144 226030 293172 231676
rect 293328 231662 293802 231690
rect 293132 226024 293184 226030
rect 293132 225966 293184 225972
rect 291844 224800 291896 224806
rect 291844 224742 291896 224748
rect 291200 223440 291252 223446
rect 291200 223382 291252 223388
rect 291476 223032 291528 223038
rect 291476 222974 291528 222980
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291488 219026 291516 222974
rect 292488 220108 292540 220114
rect 292488 220050 292540 220056
rect 291660 219292 291712 219298
rect 291660 219234 291712 219240
rect 291476 219020 291528 219026
rect 291476 218962 291528 218968
rect 291672 218890 291700 219234
rect 291660 218884 291712 218890
rect 291660 218826 291712 218832
rect 291660 218748 291712 218754
rect 291660 218690 291712 218696
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291672 217138 291700 218690
rect 292500 217274 292528 220050
rect 293328 219978 293356 231662
rect 293776 227724 293828 227730
rect 293776 227666 293828 227672
rect 293316 219972 293368 219978
rect 293316 219914 293368 219920
rect 293788 218074 293816 227666
rect 294432 225758 294460 231676
rect 294420 225752 294472 225758
rect 294420 225694 294472 225700
rect 294880 224800 294932 224806
rect 294880 224742 294932 224748
rect 294892 219434 294920 224742
rect 295076 223310 295104 231676
rect 295720 228274 295748 231676
rect 296364 229090 296392 231676
rect 296824 231662 297022 231690
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296628 228812 296680 228818
rect 296628 228754 296680 228760
rect 295708 228268 295760 228274
rect 295708 228210 295760 228216
rect 296444 225752 296496 225758
rect 296444 225694 296496 225700
rect 295064 223304 295116 223310
rect 295064 223246 295116 223252
rect 296456 219434 296484 225694
rect 294892 219406 295012 219434
rect 296456 219406 296576 219434
rect 294144 219020 294196 219026
rect 294144 218962 294196 218968
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 291626 217110 291700 217138
rect 292454 217246 292528 217274
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218962
rect 294984 217274 295012 219406
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228754
rect 296824 220794 296852 231662
rect 297652 229770 297680 231676
rect 297640 229764 297692 229770
rect 297640 229706 297692 229712
rect 296996 229628 297048 229634
rect 296996 229570 297048 229576
rect 297008 224262 297036 229570
rect 298296 227458 298324 231676
rect 298284 227452 298336 227458
rect 298284 227394 298336 227400
rect 298940 226302 298968 231676
rect 299584 228954 299612 231676
rect 299572 228948 299624 228954
rect 299572 228890 299624 228896
rect 298928 226296 298980 226302
rect 298928 226238 298980 226244
rect 299388 226024 299440 226030
rect 299388 225966 299440 225972
rect 297364 225480 297416 225486
rect 297364 225422 297416 225428
rect 296996 224256 297048 224262
rect 296996 224198 297048 224204
rect 296812 220788 296864 220794
rect 296812 220730 296864 220736
rect 297376 219434 297404 225422
rect 299112 224256 299164 224262
rect 299112 224198 299164 224204
rect 297548 223372 297600 223378
rect 297548 223314 297600 223320
rect 297364 219428 297416 219434
rect 297364 219370 297416 219376
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297560 218890 297588 223314
rect 297548 218884 297600 218890
rect 297548 218826 297600 218832
rect 297456 218204 297508 218210
rect 297456 218146 297508 218152
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218146
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 298296 217138 298324 218010
rect 299124 217274 299152 224198
rect 299400 218074 299428 225966
rect 300228 223038 300256 231676
rect 300676 228948 300728 228954
rect 300676 228890 300728 228896
rect 300216 223032 300268 223038
rect 300216 222974 300268 222980
rect 300492 218612 300544 218618
rect 300492 218554 300544 218560
rect 299388 218068 299440 218074
rect 299388 218010 299440 218016
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299152 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 218554
rect 300688 218074 300716 228890
rect 300872 225894 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 300860 225888 300912 225894
rect 300860 225830 300912 225836
rect 301056 221746 301084 231662
rect 301700 222018 301728 231662
rect 302804 230178 302832 231676
rect 302792 230172 302844 230178
rect 302792 230114 302844 230120
rect 302884 230036 302936 230042
rect 302884 229978 302936 229984
rect 302148 229084 302200 229090
rect 302148 229026 302200 229032
rect 301688 222012 301740 222018
rect 301688 221954 301740 221960
rect 301044 221740 301096 221746
rect 301044 221682 301096 221688
rect 302160 218074 302188 229026
rect 302424 221604 302476 221610
rect 302424 221546 302476 221552
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 221546
rect 302896 218210 302924 229978
rect 303448 224942 303476 231676
rect 303816 231662 304106 231690
rect 303436 224936 303488 224942
rect 303436 224878 303488 224884
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302884 218204 302936 218210
rect 302884 218146 302936 218152
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304736 227594 304764 231676
rect 304724 227588 304776 227594
rect 304724 227530 304776 227536
rect 304264 224936 304316 224942
rect 304264 224878 304316 224884
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304080 219428 304132 219434
rect 304080 219370 304132 219376
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 219370
rect 304276 218482 304304 224878
rect 305380 223378 305408 231676
rect 306024 228546 306052 231676
rect 306392 231662 306682 231690
rect 306852 231662 307326 231690
rect 306012 228540 306064 228546
rect 306012 228482 306064 228488
rect 306196 227452 306248 227458
rect 306196 227394 306248 227400
rect 305368 223372 305420 223378
rect 305368 223314 305420 223320
rect 304908 220652 304960 220658
rect 304908 220594 304960 220600
rect 304264 218476 304316 218482
rect 304264 218418 304316 218424
rect 304920 217274 304948 220594
rect 306208 218074 306236 227394
rect 306392 222154 306420 231662
rect 306380 222148 306432 222154
rect 306380 222090 306432 222096
rect 306852 220250 306880 231662
rect 307956 230450 307984 231676
rect 307944 230444 307996 230450
rect 307944 230386 307996 230392
rect 308404 230444 308456 230450
rect 308404 230386 308456 230392
rect 308220 226296 308272 226302
rect 308220 226238 308272 226244
rect 307668 223304 307720 223310
rect 307668 223246 307720 223252
rect 306840 220244 306892 220250
rect 306840 220186 306892 220192
rect 307392 219156 307444 219162
rect 307392 219098 307444 219104
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 219098
rect 307680 218074 307708 223246
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308232 217274 308260 226238
rect 308416 219434 308444 230386
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 309244 220386 309272 231676
rect 309888 224670 309916 231676
rect 310336 227044 310388 227050
rect 310336 226986 310388 226992
rect 309876 224664 309928 224670
rect 309876 224606 309928 224612
rect 309232 220380 309284 220386
rect 309232 220322 309284 220328
rect 308956 220244 309008 220250
rect 308956 220186 309008 220192
rect 308404 219428 308456 219434
rect 308404 219370 308456 219376
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217246 308260 217274
rect 308968 217274 308996 220186
rect 310348 218074 310376 226986
rect 310532 225486 310560 231676
rect 310520 225480 310572 225486
rect 310520 225422 310572 225428
rect 311176 224398 311204 231676
rect 311360 231662 311834 231690
rect 311164 224392 311216 224398
rect 311164 224334 311216 224340
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310336 218068 310388 218074
rect 310336 218010 310388 218016
rect 308968 217246 309042 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217246
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 311360 220522 311388 231662
rect 312464 228410 312492 231676
rect 313108 230314 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230308 313148 230314
rect 313096 230250 313148 230256
rect 312636 230172 312688 230178
rect 312636 230114 312688 230120
rect 312452 228404 312504 228410
rect 312452 228346 312504 228352
rect 311532 224664 311584 224670
rect 311532 224606 311584 224612
rect 311348 220516 311400 220522
rect 311348 220458 311400 220464
rect 310980 219428 311032 219434
rect 310980 219370 311032 219376
rect 310992 218618 311020 219370
rect 311164 219020 311216 219026
rect 311164 218962 311216 218968
rect 311176 218618 311204 218962
rect 310980 218612 311032 218618
rect 310980 218554 311032 218560
rect 311164 218612 311216 218618
rect 311164 218554 311216 218560
rect 311544 217274 311572 224606
rect 312648 222154 312676 230114
rect 312912 225888 312964 225894
rect 312912 225830 312964 225836
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 225830
rect 313292 225622 313320 231662
rect 313936 229094 313964 231662
rect 313752 229066 313964 229094
rect 313280 225616 313332 225622
rect 313280 225558 313332 225564
rect 313188 222012 313240 222018
rect 313188 221954 313240 221960
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221954
rect 313752 221882 313780 229066
rect 313924 228540 313976 228546
rect 313924 228482 313976 228488
rect 313740 221876 313792 221882
rect 313740 221818 313792 221824
rect 313936 219298 313964 228482
rect 315040 223582 315068 231676
rect 315408 231662 315698 231690
rect 315408 229094 315436 231662
rect 315316 229066 315436 229094
rect 315316 224942 315344 229066
rect 315488 227588 315540 227594
rect 315488 227530 315540 227536
rect 315304 224936 315356 224942
rect 315304 224878 315356 224884
rect 315028 223576 315080 223582
rect 315028 223518 315080 223524
rect 313924 219292 313976 219298
rect 313924 219234 313976 219240
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 315500 218074 315528 227530
rect 315672 223032 315724 223038
rect 315672 222974 315724 222980
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 315488 218068 315540 218074
rect 315488 218010 315540 218016
rect 314856 217138 314884 218010
rect 315684 217274 315712 222974
rect 316328 222902 316356 231676
rect 316684 223440 316736 223446
rect 316684 223382 316736 223388
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316500 220380 316552 220386
rect 316500 220322 316552 220328
rect 316512 217274 316540 220322
rect 316696 218618 316724 223382
rect 316972 222766 317000 231676
rect 317616 227186 317644 231676
rect 318260 229906 318288 231676
rect 318248 229900 318300 229906
rect 318248 229842 318300 229848
rect 318064 229764 318116 229770
rect 318064 229706 318116 229712
rect 317604 227180 317656 227186
rect 317604 227122 317656 227128
rect 316960 222760 317012 222766
rect 316960 222702 317012 222708
rect 318076 219434 318104 229706
rect 318904 228682 318932 231676
rect 319088 231662 319562 231690
rect 320206 231662 320404 231690
rect 318892 228676 318944 228682
rect 318892 228618 318944 228624
rect 318248 221876 318300 221882
rect 318248 221818 318300 221824
rect 318260 219434 318288 221818
rect 319088 219842 319116 231662
rect 320088 228404 320140 228410
rect 320088 228346 320140 228352
rect 319812 224936 319864 224942
rect 319812 224878 319864 224884
rect 319076 219836 319128 219842
rect 319076 219778 319128 219784
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218612 316736 218618
rect 316684 218554 316736 218560
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 224878
rect 320100 218074 320128 228346
rect 320376 221474 320404 231662
rect 320836 228546 320864 231676
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 321480 223174 321508 231676
rect 322124 227322 322152 231676
rect 322112 227316 322164 227322
rect 322112 227258 322164 227264
rect 322204 227180 322256 227186
rect 322204 227122 322256 227128
rect 321468 223168 321520 223174
rect 321468 223110 321520 223116
rect 321468 222896 321520 222902
rect 321468 222838 321520 222844
rect 320364 221468 320416 221474
rect 320364 221410 320416 221416
rect 320640 218612 320692 218618
rect 320640 218554 320692 218560
rect 320088 218068 320140 218074
rect 320088 218010 320140 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 218554
rect 321480 217274 321508 222838
rect 322216 219434 322244 227122
rect 322768 226166 322796 231676
rect 323412 229634 323440 231676
rect 323400 229628 323452 229634
rect 323400 229570 323452 229576
rect 322756 226160 322808 226166
rect 322756 226102 322808 226108
rect 324056 224534 324084 231676
rect 324228 229900 324280 229906
rect 324228 229842 324280 229848
rect 324044 224528 324096 224534
rect 324044 224470 324096 224476
rect 322848 224392 322900 224398
rect 322848 224334 322900 224340
rect 322204 219428 322256 219434
rect 322204 219370 322256 219376
rect 322860 218074 322888 224334
rect 323952 223168 324004 223174
rect 323952 223110 324004 223116
rect 323964 218074 323992 223110
rect 324240 219434 324268 229842
rect 324700 219434 324728 231676
rect 325344 227730 325372 231676
rect 325516 228540 325568 228546
rect 325516 228482 325568 228488
rect 325332 227724 325384 227730
rect 325332 227666 325384 227672
rect 324148 219406 324268 219434
rect 324608 219406 324728 219434
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 323952 218068 324004 218074
rect 323952 218010 324004 218016
rect 320606 217110 320680 217138
rect 321434 217246 321508 217274
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 324148 217274 324176 219406
rect 324608 218754 324636 219406
rect 325332 219020 325384 219026
rect 325332 218962 325384 218968
rect 324596 218748 324648 218754
rect 324596 218690 324648 218696
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 324176 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325344 217274 325372 218962
rect 325528 218074 325556 228482
rect 325988 224806 326016 231676
rect 326172 231662 326646 231690
rect 325976 224800 326028 224806
rect 325976 224742 326028 224748
rect 326172 220114 326200 231662
rect 326896 228676 326948 228682
rect 326896 228618 326948 228624
rect 326160 220108 326212 220114
rect 326160 220050 326212 220056
rect 326908 218074 326936 228618
rect 327276 223446 327304 231676
rect 327920 225758 327948 231676
rect 328564 226030 328592 231676
rect 329208 228818 329236 231676
rect 329852 230042 329880 231676
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 330496 228954 330524 231676
rect 331140 229090 331168 231676
rect 331416 231662 331798 231690
rect 331128 229084 331180 229090
rect 331128 229026 331180 229032
rect 330484 228948 330536 228954
rect 330484 228890 330536 228896
rect 329196 228812 329248 228818
rect 329196 228754 329248 228760
rect 331036 227792 331088 227798
rect 331036 227734 331088 227740
rect 328552 226024 328604 226030
rect 328552 225966 328604 225972
rect 327908 225752 327960 225758
rect 327908 225694 327960 225700
rect 329748 225752 329800 225758
rect 329748 225694 329800 225700
rect 327724 225616 327776 225622
rect 327724 225558 327776 225564
rect 327264 223440 327316 223446
rect 327264 223382 327316 223388
rect 327736 219026 327764 225558
rect 328092 220516 328144 220522
rect 328092 220458 328144 220464
rect 327724 219020 327776 219026
rect 327724 218962 327776 218968
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 325516 218068 325568 218074
rect 325516 218010 325568 218016
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 325344 217246 325602 217274
rect 324746 217110 324820 217138
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 220458
rect 328920 220108 328972 220114
rect 328920 220050 328972 220056
rect 328932 217274 328960 220050
rect 329760 217274 329788 225694
rect 330484 219020 330536 219026
rect 330484 218962 330536 218968
rect 330496 218618 330524 218962
rect 330484 218612 330536 218618
rect 330484 218554 330536 218560
rect 331048 218074 331076 227734
rect 331416 224262 331444 231662
rect 332428 227186 332456 231676
rect 332796 231662 333086 231690
rect 333440 231662 333730 231690
rect 334084 231662 334374 231690
rect 332416 227180 332468 227186
rect 332416 227122 332468 227128
rect 331864 224800 331916 224806
rect 331864 224742 331916 224748
rect 331404 224256 331456 224262
rect 331404 224198 331456 224204
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 328886 217246 328960 217274
rect 329714 217246 329788 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328886 216988 328914 217246
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 331876 219162 331904 224742
rect 332796 221746 332824 231662
rect 333440 229094 333468 231662
rect 333256 229066 333468 229094
rect 332784 221740 332836 221746
rect 332784 221682 332836 221688
rect 333256 220658 333284 229066
rect 333888 227180 333940 227186
rect 333888 227122 333940 227128
rect 333428 221468 333480 221474
rect 333428 221410 333480 221416
rect 333244 220652 333296 220658
rect 333244 220594 333296 220600
rect 331864 219156 331916 219162
rect 331864 219098 331916 219104
rect 333060 218204 333112 218210
rect 333060 218146 333112 218152
rect 332232 218068 332284 218074
rect 332232 218010 332284 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332244 217138 332272 218010
rect 333072 217138 333100 218146
rect 333440 218074 333468 221410
rect 333704 219156 333756 219162
rect 333704 219098 333756 219104
rect 333428 218068 333480 218074
rect 333428 218010 333480 218016
rect 333716 217274 333744 219098
rect 333900 218210 333928 227122
rect 334084 221610 334112 231662
rect 335004 230450 335032 231676
rect 334992 230444 335044 230450
rect 334992 230386 335044 230392
rect 334256 230036 334308 230042
rect 334256 229978 334308 229984
rect 334268 227798 334296 229978
rect 334256 227792 334308 227798
rect 334256 227734 334308 227740
rect 335176 226024 335228 226030
rect 335176 225966 335228 225972
rect 334072 221604 334124 221610
rect 334072 221546 334124 221552
rect 333888 218204 333940 218210
rect 333888 218146 333940 218152
rect 335188 218074 335216 225966
rect 335648 223310 335676 231676
rect 336292 226302 336320 231676
rect 336464 228812 336516 228818
rect 336464 228754 336516 228760
rect 336280 226296 336332 226302
rect 336280 226238 336332 226244
rect 335636 223304 335688 223310
rect 335636 223246 335688 223252
rect 336476 219434 336504 228754
rect 336936 227458 336964 231676
rect 336924 227452 336976 227458
rect 336924 227394 336976 227400
rect 337580 224806 337608 231676
rect 337752 227452 337804 227458
rect 337752 227394 337804 227400
rect 337568 224800 337620 224806
rect 337568 224742 337620 224748
rect 336384 219406 336504 219434
rect 335544 218204 335596 218210
rect 335544 218146 335596 218152
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 333716 217246 333882 217274
rect 332198 217110 332272 217138
rect 333026 217110 333100 217138
rect 332198 216988 332226 217110
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218146
rect 336384 217274 336412 219406
rect 337764 218074 337792 227394
rect 338224 227050 338252 231676
rect 338212 227044 338264 227050
rect 338212 226986 338264 226992
rect 338672 227044 338724 227050
rect 338672 226986 338724 226992
rect 337936 223304 337988 223310
rect 337936 223246 337988 223252
rect 337200 218068 337252 218074
rect 337200 218010 337252 218016
rect 337752 218068 337804 218074
rect 337752 218010 337804 218016
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218010
rect 337948 217274 337976 223246
rect 338684 218210 338712 226986
rect 338868 224670 338896 231676
rect 339526 231662 339724 231690
rect 338856 224664 338908 224670
rect 338856 224606 338908 224612
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 338672 218204 338724 218210
rect 338672 218146 338724 218152
rect 339420 218074 339448 224198
rect 339696 220250 339724 231662
rect 340156 230178 340184 231676
rect 340432 231662 340814 231690
rect 340144 230172 340196 230178
rect 340144 230114 340196 230120
rect 340432 222018 340460 231662
rect 341444 227594 341472 231676
rect 341720 231662 342102 231690
rect 342456 231662 342746 231690
rect 343008 231662 343390 231690
rect 343836 231662 344034 231690
rect 341432 227588 341484 227594
rect 341432 227530 341484 227536
rect 340696 227316 340748 227322
rect 340696 227258 340748 227264
rect 340420 222012 340472 222018
rect 340420 221954 340472 221960
rect 340328 220380 340380 220386
rect 340328 220322 340380 220328
rect 339684 220244 339736 220250
rect 339684 220186 339736 220192
rect 340340 218890 340368 220322
rect 340328 218884 340380 218890
rect 340328 218826 340380 218832
rect 340512 218340 340564 218346
rect 340512 218282 340564 218288
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217274 340552 218282
rect 340708 218074 340736 227258
rect 341720 225894 341748 231662
rect 341708 225888 341760 225894
rect 341708 225830 341760 225836
rect 341984 225888 342036 225894
rect 341984 225830 342036 225836
rect 341996 219434 342024 225830
rect 342168 224528 342220 224534
rect 342168 224470 342220 224476
rect 342180 219434 342208 224470
rect 342456 220386 342484 231662
rect 343008 220386 343036 231662
rect 343836 221882 343864 231662
rect 344664 223038 344692 231676
rect 345020 229764 345072 229770
rect 345020 229706 345072 229712
rect 345032 227458 345060 229706
rect 345308 229634 345336 231676
rect 345296 229628 345348 229634
rect 345296 229570 345348 229576
rect 345020 227452 345072 227458
rect 345020 227394 345072 227400
rect 345952 224942 345980 231676
rect 345940 224936 345992 224942
rect 345940 224878 345992 224884
rect 346308 224664 346360 224670
rect 346308 224606 346360 224612
rect 344652 223032 344704 223038
rect 344652 222974 344704 222980
rect 345664 222760 345716 222766
rect 345664 222702 345716 222708
rect 343824 221876 343876 221882
rect 343824 221818 343876 221824
rect 344652 221740 344704 221746
rect 344652 221682 344704 221688
rect 342444 220380 342496 220386
rect 342444 220322 342496 220328
rect 342996 220380 343048 220386
rect 342996 220322 343048 220328
rect 342996 220244 343048 220250
rect 342996 220186 343048 220192
rect 341340 219428 341392 219434
rect 341996 219406 342116 219434
rect 342180 219428 342312 219434
rect 342180 219406 342260 219428
rect 341340 219370 341392 219376
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217246 340552 217274
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217246
rect 341352 217138 341380 219370
rect 342088 217274 342116 219406
rect 342260 219370 342312 219376
rect 343008 217274 343036 220186
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342088 217246 342162 217274
rect 341306 217110 341380 217138
rect 341306 216988 341334 217110
rect 342134 216988 342162 217246
rect 342962 217246 343036 217274
rect 342962 216988 342990 217246
rect 343836 217138 343864 219370
rect 344664 217274 344692 221682
rect 345676 218890 345704 222702
rect 345664 218884 345716 218890
rect 345664 218826 345716 218832
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346320 217274 346348 224606
rect 346596 222902 346624 231676
rect 346872 231662 347254 231690
rect 346872 228410 346900 231662
rect 346860 228404 346912 228410
rect 346860 228346 346912 228352
rect 347044 228404 347096 228410
rect 347044 228346 347096 228352
rect 346584 222896 346636 222902
rect 346584 222838 346636 222844
rect 347056 219434 347084 228346
rect 347228 222896 347280 222902
rect 347228 222838 347280 222844
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347044 218884 347096 218890
rect 347044 218826 347096 218832
rect 345446 217110 345520 217138
rect 346274 217246 346348 217274
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347056 217138 347084 218826
rect 347240 218074 347268 222838
rect 347884 222766 347912 231676
rect 348528 223174 348556 231676
rect 349172 228546 349200 231676
rect 349160 228540 349212 228546
rect 349160 228482 349212 228488
rect 349816 224398 349844 231676
rect 350460 229906 350488 231676
rect 350448 229900 350500 229906
rect 350448 229842 350500 229848
rect 351104 228682 351132 231676
rect 351288 231662 351762 231690
rect 351092 228676 351144 228682
rect 351092 228618 351144 228624
rect 350448 228540 350500 228546
rect 350448 228482 350500 228488
rect 350264 224868 350316 224874
rect 350264 224810 350316 224816
rect 349804 224392 349856 224398
rect 349804 224334 349856 224340
rect 348516 223168 348568 223174
rect 348516 223110 348568 223116
rect 349068 223032 349120 223038
rect 349068 222974 349120 222980
rect 347872 222760 347924 222766
rect 347872 222702 347924 222708
rect 348792 221604 348844 221610
rect 348792 221546 348844 221552
rect 347228 218068 347280 218074
rect 347228 218010 347280 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 347976 217138 348004 218010
rect 348804 217274 348832 221546
rect 349080 218074 349108 222974
rect 350276 219434 350304 224810
rect 350460 219434 350488 228482
rect 351092 227792 351144 227798
rect 351092 227734 351144 227740
rect 349620 219428 349672 219434
rect 350276 219406 350396 219434
rect 350460 219428 350592 219434
rect 350460 219406 350540 219428
rect 349620 219370 349672 219376
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 347056 217110 347130 217138
rect 347102 216988 347130 217110
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 219370
rect 350368 217274 350396 219406
rect 350540 219370 350592 219376
rect 351104 218754 351132 227734
rect 351288 220522 351316 231662
rect 352392 225622 352420 231676
rect 353036 227798 353064 231676
rect 353024 227792 353076 227798
rect 353024 227734 353076 227740
rect 352564 227452 352616 227458
rect 352564 227394 352616 227400
rect 352380 225616 352432 225622
rect 352380 225558 352432 225564
rect 351276 220516 351328 220522
rect 351276 220458 351328 220464
rect 351276 220380 351328 220386
rect 351276 220322 351328 220328
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 220322
rect 352576 218346 352604 227394
rect 353680 225758 353708 231676
rect 353956 231662 354338 231690
rect 354784 231662 354982 231690
rect 353668 225752 353720 225758
rect 353668 225694 353720 225700
rect 352932 225616 352984 225622
rect 352932 225558 352984 225564
rect 352564 218340 352616 218346
rect 352564 218282 352616 218288
rect 352104 218068 352156 218074
rect 352104 218010 352156 218016
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 218010
rect 352944 217274 352972 225558
rect 353956 222154 353984 231662
rect 354588 228676 354640 228682
rect 354588 228618 354640 228624
rect 353944 222148 353996 222154
rect 353944 222090 353996 222096
rect 353300 221876 353352 221882
rect 353300 221818 353352 221824
rect 353312 218074 353340 221818
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 353300 218068 353352 218074
rect 353300 218010 353352 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 228618
rect 354784 220114 354812 231662
rect 355612 230042 355640 231676
rect 355600 230036 355652 230042
rect 355600 229978 355652 229984
rect 355784 230036 355836 230042
rect 355784 229978 355836 229984
rect 355232 225004 355284 225010
rect 355232 224946 355284 224952
rect 354772 220108 354824 220114
rect 354772 220050 354824 220056
rect 355244 219230 355272 224946
rect 355796 224874 355824 229978
rect 356256 227186 356284 231676
rect 356244 227180 356296 227186
rect 356244 227122 356296 227128
rect 356900 226030 356928 231676
rect 357256 227180 357308 227186
rect 357256 227122 357308 227128
rect 356888 226024 356940 226030
rect 356888 225966 356940 225972
rect 355784 224868 355836 224874
rect 355784 224810 355836 224816
rect 355416 220108 355468 220114
rect 355416 220050 355468 220056
rect 355232 219224 355284 219230
rect 355232 219166 355284 219172
rect 355428 217274 355456 220050
rect 357072 219020 357124 219026
rect 357072 218962 357124 218968
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 355382 217246 355456 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355382 216988 355410 217246
rect 356256 217138 356284 218010
rect 357084 217138 357112 218962
rect 357268 218074 357296 227122
rect 357544 221474 357572 231676
rect 358188 225010 358216 231676
rect 358832 228818 358860 231676
rect 359200 231662 359490 231690
rect 358820 228812 358872 228818
rect 358820 228754 358872 228760
rect 358176 225004 358228 225010
rect 358176 224946 358228 224952
rect 359200 223310 359228 231662
rect 359924 228812 359976 228818
rect 359924 228754 359976 228760
rect 359464 224392 359516 224398
rect 359464 224334 359516 224340
rect 359188 223304 359240 223310
rect 359188 223246 359240 223252
rect 358544 223168 358596 223174
rect 358544 223110 358596 223116
rect 357532 221468 357584 221474
rect 357532 221410 357584 221416
rect 358556 218074 358584 223110
rect 359476 218210 359504 224334
rect 359936 219434 359964 228754
rect 360120 227050 360148 231676
rect 360764 229770 360792 231676
rect 360752 229764 360804 229770
rect 360752 229706 360804 229712
rect 361212 229764 361264 229770
rect 361212 229706 361264 229712
rect 361224 229094 361252 229706
rect 361040 229066 361252 229094
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359936 219406 360148 219434
rect 358728 218204 358780 218210
rect 358728 218146 358780 218152
rect 359464 218204 359516 218210
rect 359464 218146 359516 218152
rect 357256 218068 357308 218074
rect 357256 218010 357308 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 358544 218068 358596 218074
rect 358544 218010 358596 218016
rect 357912 217138 357940 218010
rect 358740 217138 358768 218146
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227322 361436 231676
rect 361396 227316 361448 227322
rect 361396 227258 361448 227264
rect 361212 226024 361264 226030
rect 361212 225966 361264 225972
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 225966
rect 362052 224534 362080 231676
rect 362328 231662 362710 231690
rect 362040 224528 362092 224534
rect 362040 224470 362092 224476
rect 362328 224262 362356 231662
rect 363340 229094 363368 231676
rect 363524 231662 363998 231690
rect 364536 231662 364642 231690
rect 363524 229094 363552 231662
rect 363248 229066 363368 229094
rect 363432 229066 363552 229094
rect 363248 227458 363276 229066
rect 363236 227452 363288 227458
rect 363236 227394 363288 227400
rect 363432 227338 363460 229066
rect 363340 227310 363460 227338
rect 363604 227316 363656 227322
rect 362776 227044 362828 227050
rect 362776 226986 362828 226992
rect 362316 224256 362368 224262
rect 362316 224198 362368 224204
rect 362040 219156 362092 219162
rect 362040 219098 362092 219104
rect 362052 217274 362080 219098
rect 356210 217110 356284 217138
rect 357038 217110 357112 217138
rect 357866 217110 357940 217138
rect 358694 217110 358768 217138
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362788 217274 362816 226986
rect 363340 220250 363368 227310
rect 363604 227258 363656 227264
rect 363616 220402 363644 227258
rect 364536 221746 364564 231662
rect 365272 225894 365300 231676
rect 365916 228410 365944 231676
rect 365904 228404 365956 228410
rect 365904 228346 365956 228352
rect 365260 225888 365312 225894
rect 365260 225830 365312 225836
rect 365352 225752 365404 225758
rect 365352 225694 365404 225700
rect 364524 221740 364576 221746
rect 364524 221682 364576 221688
rect 364524 220516 364576 220522
rect 364524 220458 364576 220464
rect 363524 220374 363644 220402
rect 363328 220244 363380 220250
rect 363328 220186 363380 220192
rect 363524 218890 363552 220374
rect 363696 220244 363748 220250
rect 363696 220186 363748 220192
rect 363512 218884 363564 218890
rect 363512 218826 363564 218832
rect 363708 217274 363736 220186
rect 364536 217274 364564 220458
rect 365364 217274 365392 225694
rect 366560 224670 366588 231676
rect 366732 229900 366784 229906
rect 366732 229842 366784 229848
rect 366744 229094 366772 229842
rect 366744 229066 366956 229094
rect 366548 224664 366600 224670
rect 366548 224606 366600 224612
rect 366732 224528 366784 224534
rect 366732 224470 366784 224476
rect 366744 219570 366772 224470
rect 366732 219564 366784 219570
rect 366732 219506 366784 219512
rect 366180 219428 366232 219434
rect 366180 219370 366232 219376
rect 362788 217246 362862 217274
rect 356210 216988 356238 217110
rect 357038 216988 357066 217110
rect 357866 216988 357894 217110
rect 358694 216988 358722 217110
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363662 217246 363736 217274
rect 364490 217246 364564 217274
rect 365318 217246 365392 217274
rect 363662 216988 363690 217246
rect 364490 216988 364518 217246
rect 365318 216988 365346 217246
rect 366192 217138 366220 219370
rect 366928 217274 366956 229066
rect 367204 223038 367232 231676
rect 367192 223032 367244 223038
rect 367192 222974 367244 222980
rect 367848 222902 367876 231676
rect 368492 227322 368520 231676
rect 369136 228546 369164 231676
rect 369320 231662 369794 231690
rect 370056 231662 370438 231690
rect 369124 228540 369176 228546
rect 369124 228482 369176 228488
rect 368480 227316 368532 227322
rect 368480 227258 368532 227264
rect 369124 226500 369176 226506
rect 369124 226442 369176 226448
rect 368388 223032 368440 223038
rect 368388 222974 368440 222980
rect 367836 222896 367888 222902
rect 367836 222838 367888 222844
rect 368400 218074 368428 222974
rect 369136 219026 369164 226442
rect 369320 220386 369348 231662
rect 370056 221610 370084 231662
rect 371068 230042 371096 231676
rect 371056 230036 371108 230042
rect 371056 229978 371108 229984
rect 371712 229094 371740 231676
rect 371620 229066 371740 229094
rect 371148 228404 371200 228410
rect 371148 228346 371200 228352
rect 370964 221740 371016 221746
rect 370964 221682 371016 221688
rect 370044 221604 370096 221610
rect 370044 221546 370096 221552
rect 369492 221468 369544 221474
rect 369492 221410 369544 221416
rect 369308 220380 369360 220386
rect 369308 220322 369360 220328
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 368664 218884 368716 218890
rect 368664 218826 368716 218832
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 366146 217110 366220 217138
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218826
rect 369504 217274 369532 221410
rect 370976 219162 371004 221682
rect 370964 219156 371016 219162
rect 370964 219098 371016 219104
rect 370320 219020 370372 219026
rect 370320 218962 370372 218968
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370332 217138 370360 218962
rect 371160 217274 371188 228346
rect 371620 225622 371648 229066
rect 372356 228682 372384 231676
rect 372724 231662 373014 231690
rect 372344 228676 372396 228682
rect 372344 228618 372396 228624
rect 371792 227792 371844 227798
rect 371792 227734 371844 227740
rect 371608 225616 371660 225622
rect 371608 225558 371660 225564
rect 371804 218754 371832 227734
rect 372528 224256 372580 224262
rect 372528 224198 372580 224204
rect 371792 218748 371844 218754
rect 371792 218690 371844 218696
rect 372540 218074 372568 224198
rect 372724 221882 372752 231662
rect 373448 228540 373500 228546
rect 373448 228482 373500 228488
rect 372712 221876 372764 221882
rect 372712 221818 372764 221824
rect 373460 219434 373488 228482
rect 373644 227798 373672 231676
rect 373632 227792 373684 227798
rect 373632 227734 373684 227740
rect 374288 227186 374316 231676
rect 374656 231662 374946 231690
rect 374276 227180 374328 227186
rect 374276 227122 374328 227128
rect 374656 223174 374684 231662
rect 375012 225888 375064 225894
rect 375012 225830 375064 225836
rect 374644 223168 374696 223174
rect 374644 223110 374696 223116
rect 373724 221604 373776 221610
rect 373724 221546 373776 221552
rect 373460 219406 373580 219434
rect 373552 218074 373580 219406
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373540 218068 373592 218074
rect 373540 218010 373592 218016
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373736 217274 373764 221546
rect 375024 218074 375052 225830
rect 375196 222896 375248 222902
rect 375196 222838 375248 222844
rect 374460 218068 374512 218074
rect 374460 218010 374512 218016
rect 375012 218068 375064 218074
rect 375012 218010 375064 218016
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373764 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218010
rect 375208 217274 375236 222838
rect 375576 220114 375604 231676
rect 376220 226506 376248 231676
rect 376864 228818 376892 231676
rect 376852 228812 376904 228818
rect 376852 228754 376904 228760
rect 376668 227180 376720 227186
rect 376668 227122 376720 227128
rect 376208 226500 376260 226506
rect 376208 226442 376260 226448
rect 375564 220108 375616 220114
rect 375564 220050 375616 220056
rect 376680 218074 376708 227122
rect 377508 226030 377536 231676
rect 377772 228676 377824 228682
rect 377772 228618 377824 228624
rect 377496 226024 377548 226030
rect 377496 225966 377548 225972
rect 376944 220380 376996 220386
rect 376944 220322 376996 220328
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 375208 217246 375282 217274
rect 374426 217110 374500 217138
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217274 376984 220322
rect 377784 217274 377812 228618
rect 378152 224398 378180 231676
rect 378796 229770 378824 231676
rect 379072 231662 379454 231690
rect 379716 231662 380098 231690
rect 380360 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 378784 229764 378836 229770
rect 378784 229706 378836 229712
rect 379072 227050 379100 231662
rect 379060 227044 379112 227050
rect 379060 226986 379112 226992
rect 378784 226840 378836 226846
rect 378784 226782 378836 226788
rect 378140 224392 378192 224398
rect 378140 224334 378192 224340
rect 378796 218890 378824 226782
rect 379244 224392 379296 224398
rect 379244 224334 379296 224340
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379256 218074 379284 224334
rect 379716 220522 379744 231662
rect 380360 221882 380388 231662
rect 380348 221876 380400 221882
rect 380348 221818 380400 221824
rect 380072 221740 380124 221746
rect 380072 221682 380124 221688
rect 379704 220516 379756 220522
rect 379704 220458 379756 220464
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217246 376984 217274
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217246
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 219026 380112 221682
rect 381096 220250 381124 231662
rect 381648 224534 381676 231662
rect 382096 227316 382148 227322
rect 382096 227258 382148 227264
rect 381636 224528 381688 224534
rect 381636 224470 381688 224476
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 380256 219020 380308 219026
rect 380256 218962 380308 218968
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 218962
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227258
rect 382660 223038 382688 231676
rect 383304 225758 383332 231676
rect 383948 229906 383976 231676
rect 384132 231662 384606 231690
rect 383936 229900 383988 229906
rect 383936 229842 383988 229848
rect 383292 225752 383344 225758
rect 383292 225694 383344 225700
rect 382924 225616 382976 225622
rect 382924 225558 382976 225564
rect 382648 223032 382700 223038
rect 382648 222974 382700 222980
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225558
rect 383568 223032 383620 223038
rect 383568 222974 383620 222980
rect 383580 218890 383608 222974
rect 384132 221474 384160 231662
rect 384304 229560 384356 229566
rect 384304 229502 384356 229508
rect 384316 221610 384344 229502
rect 385236 228410 385264 231676
rect 385224 228404 385276 228410
rect 385224 228346 385276 228352
rect 385880 226846 385908 231676
rect 386236 228404 386288 228410
rect 386236 228346 386288 228352
rect 385868 226840 385920 226846
rect 385868 226782 385920 226788
rect 386052 226432 386104 226438
rect 386052 226374 386104 226380
rect 384304 221604 384356 221610
rect 384304 221546 384356 221552
rect 384120 221468 384172 221474
rect 384120 221410 384172 221416
rect 384396 221468 384448 221474
rect 384396 221410 384448 221416
rect 383568 218884 383620 218890
rect 383568 218826 383620 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 221410
rect 386064 218074 386092 226374
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 386052 218068 386104 218074
rect 386052 218010 386104 218016
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385236 217138 385264 218010
rect 386248 217274 386276 228346
rect 386524 221746 386552 231676
rect 387168 228546 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228540 387208 228546
rect 387156 228482 387208 228488
rect 387444 224262 387472 230318
rect 387812 225894 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 388444 230240 388496 230246
rect 388444 230182 388496 230188
rect 387800 225888 387852 225894
rect 387800 225830 387852 225836
rect 387708 225752 387760 225758
rect 387708 225694 387760 225700
rect 387432 224256 387484 224262
rect 387432 224198 387484 224204
rect 386512 221740 386564 221746
rect 386512 221682 386564 221688
rect 386880 218884 386932 218890
rect 386880 218826 386932 218832
rect 385190 217110 385264 217138
rect 386018 217246 386276 217274
rect 385190 216988 385218 217110
rect 386018 216988 386046 217246
rect 386892 217138 386920 218826
rect 387720 217274 387748 225694
rect 388456 220386 388484 230182
rect 389100 229566 389128 231676
rect 389088 229560 389140 229566
rect 389088 229502 389140 229508
rect 389744 227186 389772 231676
rect 390388 228682 390416 231676
rect 390376 228676 390428 228682
rect 390376 228618 390428 228624
rect 390468 228540 390520 228546
rect 390468 228482 390520 228488
rect 389732 227180 389784 227186
rect 389732 227122 389784 227128
rect 388628 226296 388680 226302
rect 388628 226238 388680 226244
rect 388444 220380 388496 220386
rect 388444 220322 388496 220328
rect 388444 220244 388496 220250
rect 388444 220186 388496 220192
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388456 217274 388484 220186
rect 388640 219026 388668 226238
rect 390192 224256 390244 224262
rect 390192 224198 390244 224204
rect 388628 219020 388680 219026
rect 388628 218962 388680 218968
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 388456 217246 388530 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 224198
rect 390480 218074 390508 228482
rect 391032 222902 391060 231676
rect 391676 230246 391704 231676
rect 392136 231662 392334 231690
rect 391664 230240 391716 230246
rect 391664 230182 391716 230188
rect 391204 229764 391256 229770
rect 391204 229706 391256 229712
rect 391216 226438 391244 229706
rect 391756 227044 391808 227050
rect 391756 226986 391808 226992
rect 391204 226432 391256 226438
rect 391204 226374 391256 226380
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221604 391072 221610
rect 391020 221546 391072 221552
rect 390468 218068 390520 218074
rect 390468 218010 390520 218016
rect 391032 217274 391060 221546
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 217274 391796 226986
rect 392136 220114 392164 231662
rect 392964 227322 392992 231676
rect 392952 227316 393004 227322
rect 392952 227258 393004 227264
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 393148 218074 393176 227122
rect 393608 224398 393636 231676
rect 394252 226302 394280 231676
rect 394240 226296 394292 226302
rect 394240 226238 394292 226244
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393596 224392 393648 224398
rect 393596 224334 393648 224340
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224392 394568 224398
rect 394516 224334 394568 224340
rect 394528 218074 394556 224334
rect 394896 223038 394924 231676
rect 395172 231662 395554 231690
rect 394884 223032 394936 223038
rect 394884 222974 394936 222980
rect 395172 221474 395200 231662
rect 396184 225622 396212 231676
rect 396368 231662 396842 231690
rect 396172 225616 396224 225622
rect 396172 225558 396224 225564
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221468 395212 221474
rect 395160 221410 395212 221416
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228410 397500 231676
rect 397840 231662 398130 231690
rect 397460 228404 397512 228410
rect 397460 228346 397512 228352
rect 397840 225758 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 225752 397880 225758
rect 397828 225694 397880 225700
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 218890 398144 230318
rect 398760 229770 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 398748 229764 398800 229770
rect 398748 229706 398800 229712
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399864 219434 399892 229706
rect 400048 228546 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 400036 228540 400088 228546
rect 400036 228482 400088 228488
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400416 221610 400444 231662
rect 400404 221604 400456 221610
rect 400404 221546 400456 221552
rect 400968 220250 400996 231662
rect 401980 224262 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 224256 402020 224262
rect 401968 224198 402020 224204
rect 401324 221604 401376 221610
rect 401324 221546 401376 221552
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 218884 398156 218890
rect 398104 218826 398156 218832
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 397656 217274 397684 218010
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 397610 217246 397684 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397610 216988 397638 217246
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400956 218204 401008 218210
rect 400956 218146 401008 218152
rect 400048 217246 400122 217274
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218146
rect 401336 218074 401364 221546
rect 402256 218210 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 401324 218068 401376 218074
rect 401324 218010 401376 218016
rect 401784 218068 401836 218074
rect 401784 218010 401836 218016
rect 401796 217138 401824 218010
rect 402624 217138 402652 218826
rect 402808 218074 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 402796 218068 402848 218074
rect 402796 218010 402848 218016
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224398 404584 231676
rect 404740 231662 405214 231690
rect 404544 224392 404596 224398
rect 404544 224334 404596 224340
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 405568 218074 405596 224198
rect 405844 221610 405872 231676
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405832 221604 405884 221610
rect 405832 221546 405884 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229764 410944 229770
rect 410892 229706 410944 229712
rect 410904 229094 410932 229706
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229770 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229764 417476 229770
rect 417424 229706 417476 229712
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 221808 425020 221814
rect 424968 221750 425020 221756
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 221750
rect 425440 218210 425468 231662
rect 426452 226982 426480 231676
rect 426728 231662 427110 231690
rect 426440 226976 426492 226982
rect 426440 226918 426492 226924
rect 426728 220114 426756 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429212 231662 429686 231690
rect 429856 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 426992 226976 427044 226982
rect 426992 226918 427044 226924
rect 426716 220108 426768 220114
rect 426716 220050 426768 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 226918
rect 427912 224256 427964 224262
rect 427912 224198 427964 224204
rect 427924 218074 427952 224198
rect 428476 218210 428504 229066
rect 428752 224262 428780 231662
rect 428740 224256 428792 224262
rect 428740 224198 428792 224204
rect 429212 221814 429240 231662
rect 429856 229094 429884 231662
rect 429396 229066 429884 229094
rect 429200 221808 429252 221814
rect 429200 221750 429252 221756
rect 429396 218346 429424 229066
rect 429568 220244 429620 220250
rect 429568 220186 429620 220192
rect 429384 218340 429436 218346
rect 429384 218282 429436 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 429108 218204 429160 218210
rect 429108 218146 429160 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 428280 218068 428332 218074
rect 428280 218010 428332 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 218010
rect 429120 217138 429148 218146
rect 429580 218074 429608 220186
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 220250 432092 231662
rect 432052 220244 432104 220250
rect 432052 220186 432104 220192
rect 431960 220108 432012 220114
rect 431960 220050 432012 220056
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429568 218068 429620 218074
rect 429568 218010 429620 218016
rect 429948 217138 429976 218690
rect 430592 218210 430620 219406
rect 430580 218204 430632 218210
rect 430580 218146 430632 218152
rect 430776 217274 430804 219406
rect 431972 218090 432000 220050
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220114 434852 231676
rect 435192 231662 435482 231690
rect 436126 231662 436692 231690
rect 434812 220108 434864 220114
rect 434812 220050 434864 220056
rect 435192 219434 435220 231662
rect 436100 230308 436152 230314
rect 436100 230250 436152 230256
rect 434732 219406 435220 219434
rect 434732 218210 434760 219406
rect 434720 218204 434772 218210
rect 434720 218146 434772 218152
rect 435732 218204 435784 218210
rect 435732 218146 435784 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434904 218068 434956 218074
rect 434904 218010 434956 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218010
rect 435744 217138 435772 218146
rect 436112 217258 436140 230250
rect 436284 220380 436336 220386
rect 436284 220322 436336 220328
rect 436296 218074 436324 220322
rect 436664 218210 436692 231662
rect 436756 230330 436784 231676
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436756 230314 436876 230330
rect 436756 230308 436888 230314
rect 436756 230302 436836 230308
rect 436836 230250 436888 230256
rect 437032 220386 437060 231662
rect 437020 220380 437072 220386
rect 437020 220322 437072 220328
rect 436652 218204 436704 218210
rect 436652 218146 436704 218152
rect 437768 218074 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 224954 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 224954 439360 230318
rect 438872 224926 438992 224954
rect 439056 224926 439360 224954
rect 438872 219434 438900 224926
rect 438216 219428 438268 219434
rect 438216 219370 438268 219376
rect 438860 219428 438912 219434
rect 438860 219370 438912 219376
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437756 218068 437808 218074
rect 437756 218010 437808 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 219370
rect 439056 217274 439084 224926
rect 440344 219434 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 219428 439924 219434
rect 439872 219370 439924 219376
rect 440332 219428 440384 219434
rect 440332 219370 440384 219376
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 219370
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 224954 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 224926 441752 224954
rect 441632 218090 441660 224926
rect 441540 218062 441660 218090
rect 441540 217274 441568 218062
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441494 217246 441568 217274
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230246 443868 231676
rect 444484 230450 444512 231676
rect 444668 231662 445142 231690
rect 444472 230444 444524 230450
rect 444472 230386 444524 230392
rect 444668 230330 444696 231662
rect 444484 230302 444696 230330
rect 443828 230240 443880 230246
rect 443828 230182 443880 230188
rect 443472 229066 443960 229094
rect 443932 217274 443960 229066
rect 444484 224954 444512 230302
rect 444656 230240 444708 230246
rect 444656 230182 444708 230188
rect 444668 224954 444696 230182
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 445772 229066 446444 229094
rect 444484 224926 444604 224954
rect 444668 224926 445616 224954
rect 444576 217274 444604 224926
rect 445588 217274 445616 224926
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447244 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447244 219434 447272 231662
rect 447600 230444 447652 230450
rect 447600 230386 447652 230392
rect 447612 219434 447640 230386
rect 448348 229094 448376 231676
rect 448992 229566 449020 231676
rect 449636 229906 449664 231676
rect 449624 229900 449676 229906
rect 449624 229842 449676 229848
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448796 229424 448848 229430
rect 448796 229366 448848 229372
rect 448808 229094 448836 229366
rect 450280 229294 450308 231676
rect 450544 229900 450596 229906
rect 450544 229842 450596 229848
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 229842
rect 450924 229430 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451372 229560 451424 229566
rect 451372 229502 451424 229508
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 448348 229066 448652 229094
rect 448808 229066 448928 229094
rect 450556 229066 450768 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444576 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441494 216988 441522 217246
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448624 217258 448652 229066
rect 448900 217274 448928 229066
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 451384 224262 451412 229502
rect 451832 229288 451884 229294
rect 451832 229230 451884 229236
rect 451372 224256 451424 224262
rect 451372 224198 451424 224204
rect 451844 219434 451872 229230
rect 452200 224256 452252 224262
rect 452200 224198 452252 224204
rect 451476 219406 451872 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448106 217194 448158 217200
rect 448612 217252 448664 217258
rect 448900 217246 448974 217274
rect 448612 217194 448664 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449762 217252 449814 217258
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 224198
rect 452580 222154 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453500 230246 453528 231676
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 453488 230240 453540 230246
rect 453488 230182 453540 230188
rect 453028 229424 453080 229430
rect 453028 229366 453080 229372
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229366
rect 453316 218074 453344 230182
rect 454144 230110 454172 231676
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 454328 229094 454356 230318
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455788 230240 455840 230246
rect 455788 230182 455840 230188
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220726 455368 230046
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220720 455380 220726
rect 455328 220662 455380 220668
rect 455616 218074 455644 222090
rect 455800 219434 455828 230182
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220862 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220856 456760 220862
rect 456708 220798 456760 220804
rect 457180 219434 457208 230318
rect 457364 230042 457392 231676
rect 457352 230036 457404 230042
rect 457352 229978 457404 229984
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 458824 220720 458876 220726
rect 458824 220662 458876 220668
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220662
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 224942 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224936 460624 224942
rect 460572 224878 460624 224884
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 225762
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 230036 463936 230042
rect 463884 229978 463936 229984
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224936 463200 224942
rect 463148 224878 463200 224884
rect 463160 218074 463188 224878
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229978
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 472176 229362 472204 231676
rect 472834 231662 473216 231690
rect 472164 229356 472216 229362
rect 472164 229298 472216 229304
rect 472992 229356 473044 229362
rect 472992 229298 473044 229304
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471428 220856 471480 220862
rect 471428 220798 471480 220804
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 471440 218074 471468 220798
rect 473004 220386 473032 229298
rect 472992 220380 473044 220386
rect 472992 220322 473044 220328
rect 473188 220250 473216 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220244 473228 220250
rect 473176 220186 473228 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471428 218068 471480 218074
rect 471428 218010 471480 218016
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220794 474044 229842
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475884 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475856 221746 475884 231662
rect 476040 229838 476068 231676
rect 476684 230042 476712 231676
rect 476672 230036 476724 230042
rect 476672 229978 476724 229984
rect 476028 229832 476080 229838
rect 476028 229774 476080 229780
rect 476764 229696 476816 229702
rect 476764 229638 476816 229644
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475844 221740 475896 221746
rect 475844 221682 475896 221688
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229638
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 229832 478656 229838
rect 478604 229774 478656 229780
rect 478616 227186 478644 229774
rect 478800 229094 478828 231662
rect 479260 229906 479288 231676
rect 479248 229900 479300 229906
rect 479248 229842 479300 229848
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 481192 225758 481220 231676
rect 481640 230036 481692 230042
rect 481640 229978 481692 229984
rect 481652 226370 481680 229978
rect 481836 229770 481864 231676
rect 482494 231662 482968 231690
rect 481824 229764 481876 229770
rect 481824 229706 481876 229712
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 481180 225752 481232 225758
rect 481180 225694 481232 225700
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480352 224256 480404 224262
rect 480352 224198 480404 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480364 217274 480392 224198
rect 482756 222630 482784 226442
rect 482744 222624 482796 222630
rect 482744 222566 482796 222572
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222566
rect 482940 220250 482968 231662
rect 483124 223174 483152 231676
rect 483768 224262 483796 231676
rect 484426 231662 484808 231690
rect 484584 228404 484636 228410
rect 484584 228346 484636 228352
rect 483756 224256 483808 224262
rect 483756 224198 483808 224204
rect 483112 223168 483164 223174
rect 483112 223110 483164 223116
rect 484596 222358 484624 228346
rect 484584 222352 484636 222358
rect 484584 222294 484636 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 480364 217246 480438 217274
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 484596 217274 484624 222294
rect 484780 221610 484808 231662
rect 485056 228410 485084 231676
rect 485700 228546 485728 231676
rect 486358 231662 486648 231690
rect 485688 228540 485740 228546
rect 485688 228482 485740 228488
rect 485044 228404 485096 228410
rect 485044 228346 485096 228352
rect 486620 223038 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486608 223032 486660 223038
rect 486608 222974 486660 222980
rect 486148 221740 486200 221746
rect 486148 221682 486200 221688
rect 484768 221604 484820 221610
rect 484768 221546 484820 221552
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485332 217274 485360 218690
rect 486160 217274 486188 221682
rect 486804 219434 486832 227122
rect 486988 227050 487016 231676
rect 487632 230382 487660 231676
rect 487620 230376 487672 230382
rect 487620 230318 487672 230324
rect 488080 229900 488132 229906
rect 488080 229842 488132 229848
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 488092 226370 488120 229842
rect 488276 229362 488304 231676
rect 488934 231662 489408 231690
rect 488448 230376 488500 230382
rect 488448 230318 488500 230324
rect 488264 229356 488316 229362
rect 488264 229298 488316 229304
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 488080 226364 488132 226370
rect 488080 226306 488132 226312
rect 486974 219464 487030 219473
rect 486804 219408 486974 219434
rect 486804 219406 487030 219408
rect 486974 219399 487030 219406
rect 486988 217274 487016 219399
rect 487816 218113 487844 226306
rect 488460 220522 488488 230318
rect 489380 225622 489408 231662
rect 489564 229094 489592 231676
rect 490208 229770 490236 231676
rect 490866 231662 491248 231690
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 490196 229764 490248 229770
rect 490196 229706 490248 229712
rect 489564 229066 489684 229094
rect 488724 225616 488776 225622
rect 488724 225558 488776 225564
rect 489368 225616 489420 225622
rect 489368 225558 489420 225564
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488736 217274 488764 225558
rect 489656 220114 489684 229066
rect 489932 227798 489960 229706
rect 490380 229356 490432 229362
rect 490380 229298 490432 229304
rect 490196 228812 490248 228818
rect 490196 228754 490248 228760
rect 489920 227792 489972 227798
rect 489920 227734 489972 227740
rect 490012 226364 490064 226370
rect 490012 226306 490064 226312
rect 490024 222426 490052 226306
rect 490012 222420 490064 222426
rect 490012 222362 490064 222368
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 489644 220108 489696 220114
rect 489644 220050 489696 220056
rect 485332 217246 485406 217274
rect 486160 217246 486234 217274
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486206 216988 486234 217246
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488764 217274
rect 489472 217274 489500 220050
rect 490024 219434 490052 222362
rect 489932 219406 490052 219434
rect 490208 219434 490236 228754
rect 490392 227186 490420 229298
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229906 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229900 492180 229906
rect 492128 229842 492180 229848
rect 491220 229066 491340 229094
rect 490380 227180 490432 227186
rect 490380 227122 490432 227128
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 492036 222896 492088 222902
rect 492036 222838 492088 222844
rect 490208 219406 490420 219434
rect 489472 217246 489546 217274
rect 489932 217258 489960 219406
rect 490392 218657 490420 219406
rect 490378 218648 490434 218657
rect 490378 218583 490434 218592
rect 490392 217274 490420 218583
rect 492048 218074 492076 222838
rect 492508 221882 492536 230046
rect 492680 225752 492732 225758
rect 492680 225694 492732 225700
rect 492496 221876 492548 221882
rect 492496 221818 492548 221824
rect 492692 218385 492720 225694
rect 492864 224392 492916 224398
rect 492864 224334 492916 224340
rect 492678 218376 492734 218385
rect 492678 218311 492734 218320
rect 492036 218068 492088 218074
rect 492036 218010 492088 218016
rect 488690 217161 488718 217246
rect 488676 217152 488732 217161
rect 488676 217087 488732 217096
rect 488690 216988 488718 217087
rect 489518 216988 489546 217246
rect 489920 217252 489972 217258
rect 489920 217194 489972 217200
rect 490346 217246 490420 217274
rect 491162 217252 491214 217258
rect 490346 216988 490374 217246
rect 491162 217194 491214 217200
rect 491174 216988 491202 217194
rect 492048 217138 492076 218010
rect 492876 217274 492904 224334
rect 493060 223310 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493600 229764 493652 229770
rect 493600 229706 493652 229712
rect 493612 225758 493640 229706
rect 493600 225752 493652 225758
rect 493600 225694 493652 225700
rect 494072 224670 494100 231676
rect 494520 227792 494572 227798
rect 494520 227734 494572 227740
rect 494060 224664 494112 224670
rect 494060 224606 494112 224612
rect 493048 223304 493100 223310
rect 493048 223246 493100 223252
rect 494532 219434 494560 227734
rect 494716 227458 494744 231676
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 494704 227452 494756 227458
rect 494704 227394 494756 227400
rect 496084 223168 496136 223174
rect 496084 223110 496136 223116
rect 495348 220244 495400 220250
rect 495348 220186 495400 220192
rect 494532 219406 494744 219434
rect 494716 218929 494744 219406
rect 494702 218920 494758 218929
rect 494532 218878 494702 218906
rect 493782 218376 493838 218385
rect 493782 218311 493838 218320
rect 493796 217297 493824 218311
rect 492002 217110 492076 217138
rect 492830 217246 492904 217274
rect 493782 217288 493838 217297
rect 492002 216988 492030 217110
rect 492830 216988 492858 217246
rect 494532 217274 494560 218878
rect 494702 218855 494758 218864
rect 495360 217297 495388 220186
rect 493782 217223 493838 217232
rect 494486 217246 494560 217274
rect 495346 217288 495402 217297
rect 493796 217138 493824 217223
rect 493658 217110 493824 217138
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495346 217223 495402 217232
rect 495360 217138 495388 217223
rect 495314 217110 495388 217138
rect 496096 217138 496124 223110
rect 496280 221746 496308 229066
rect 496268 221740 496320 221746
rect 496268 221682 496320 221688
rect 496464 220386 496492 229066
rect 496912 224256 496964 224262
rect 496912 224198 496964 224204
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 496924 218385 496952 224198
rect 497476 220250 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498292 228540 498344 228546
rect 498292 228482 498344 228488
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 498108 221604 498160 221610
rect 498108 221546 498160 221552
rect 498120 220969 498148 221546
rect 497830 220960 497886 220969
rect 497830 220895 497886 220904
rect 498106 220960 498162 220969
rect 498106 220895 498162 220904
rect 497464 220244 497516 220250
rect 497464 220186 497516 220192
rect 496910 218376 496966 218385
rect 496910 218311 496966 218320
rect 496924 217138 496952 218311
rect 497844 217138 497872 220895
rect 498304 217258 498332 228482
rect 498568 228404 498620 228410
rect 498568 228346 498620 228352
rect 498580 224954 498608 228346
rect 498488 224926 498608 224954
rect 498488 217297 498516 224926
rect 499224 224398 499252 231676
rect 499868 228546 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228540 499908 228546
rect 499856 228482 499908 228488
rect 500236 224954 500264 229230
rect 500236 224926 500448 224954
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500040 223032 500092 223038
rect 500040 222974 500092 222980
rect 500052 218210 500080 222974
rect 500224 222488 500276 222494
rect 500224 222430 500276 222436
rect 500236 222222 500264 222430
rect 500224 222216 500276 222222
rect 500224 222158 500276 222164
rect 500420 220658 500448 224926
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500972 224954 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 500972 224926 501092 224954
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500408 220652 500460 220658
rect 500408 220594 500460 220600
rect 501064 219502 501092 224926
rect 501340 221610 501368 231662
rect 502444 228954 502472 231676
rect 503102 231662 503392 231690
rect 502432 228948 502484 228954
rect 502432 228890 502484 228896
rect 503168 227180 503220 227186
rect 503168 227122 503220 227128
rect 502984 225616 503036 225622
rect 502984 225558 503036 225564
rect 501328 221604 501380 221610
rect 501328 221546 501380 221552
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 501052 219496 501104 219502
rect 501052 219438 501104 219444
rect 500040 218204 500092 218210
rect 500040 218146 500092 218152
rect 498474 217288 498530 217297
rect 498292 217252 498344 217258
rect 500052 217274 500080 218146
rect 501064 217274 501092 219438
rect 498474 217223 498530 217232
rect 499442 217252 499494 217258
rect 498292 217194 498344 217200
rect 496096 217110 496170 217138
rect 496924 217110 496998 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217110
rect 496970 216988 496998 217110
rect 497798 217110 497872 217138
rect 498488 217138 498516 217223
rect 500052 217246 500310 217274
rect 501064 217246 501138 217274
rect 499442 217194 499494 217200
rect 498488 217110 498654 217138
rect 497798 216988 497826 217110
rect 498626 216988 498654 217110
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501110 216988 501138 217246
rect 501892 217138 501920 220458
rect 502996 217258 503024 225558
rect 503180 218346 503208 227122
rect 503364 223174 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504376 224126 504404 231676
rect 505020 227186 505048 231676
rect 505192 229764 505244 229770
rect 505192 229706 505244 229712
rect 505008 227180 505060 227186
rect 505008 227122 505060 227128
rect 504364 224120 504416 224126
rect 504364 224062 504416 224068
rect 505204 223786 505232 229706
rect 505664 229294 505692 231676
rect 505652 229288 505704 229294
rect 505652 229230 505704 229236
rect 506308 227050 506336 231676
rect 506296 227044 506348 227050
rect 506296 226986 506348 226992
rect 505376 225752 505428 225758
rect 505376 225694 505428 225700
rect 505192 223780 505244 223786
rect 505192 223722 505244 223728
rect 505388 223650 505416 225694
rect 506952 224806 506980 231676
rect 507124 229900 507176 229906
rect 507124 229842 507176 229848
rect 507136 228410 507164 229842
rect 507596 229770 507624 231676
rect 507584 229764 507636 229770
rect 507584 229706 507636 229712
rect 507124 228404 507176 228410
rect 507124 228346 507176 228352
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 506020 224528 506072 224534
rect 506020 224470 506072 224476
rect 505376 223644 505428 223650
rect 505376 223586 505428 223592
rect 503352 223168 503404 223174
rect 503352 223110 503404 223116
rect 504364 220108 504416 220114
rect 504364 220050 504416 220056
rect 503168 218340 503220 218346
rect 503168 218282 503220 218288
rect 502984 217252 503036 217258
rect 502984 217194 503036 217200
rect 503180 217138 503208 218282
rect 503582 217252 503634 217258
rect 503582 217194 503634 217200
rect 501892 217110 501966 217138
rect 501938 216988 501966 217110
rect 502766 217110 503208 217138
rect 503594 217122 503622 217194
rect 504376 217138 504404 220050
rect 505388 217274 505416 223586
rect 506032 219638 506060 224470
rect 507676 223780 507728 223786
rect 507676 223722 507728 223728
rect 506848 221876 506900 221882
rect 506848 221818 506900 221824
rect 506020 219632 506072 219638
rect 506020 219574 506072 219580
rect 505652 218068 505704 218074
rect 505652 218010 505704 218016
rect 505664 217569 505692 218010
rect 505650 217560 505706 217569
rect 505650 217495 505706 217504
rect 505250 217246 505416 217274
rect 503582 217116 503634 217122
rect 502766 216988 502794 217110
rect 504376 217110 504450 217138
rect 503582 217058 503634 217064
rect 503594 216988 503622 217058
rect 504422 216988 504450 217110
rect 505250 216988 505278 217246
rect 506032 217138 506060 219574
rect 506860 217138 506888 221818
rect 507688 218074 507716 223722
rect 508240 223038 508268 231676
rect 508884 225758 508912 231676
rect 509528 229634 509556 231676
rect 509516 229628 509568 229634
rect 509516 229570 509568 229576
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 508504 223304 508556 223310
rect 508504 223246 508556 223252
rect 508228 223032 508280 223038
rect 508228 222974 508280 222980
rect 507676 218068 507728 218074
rect 507676 218010 507728 218016
rect 507688 217138 507716 218010
rect 508516 217841 508544 223246
rect 509896 220386 509924 229094
rect 510172 225622 510200 231676
rect 510816 229906 510844 231676
rect 511460 230382 511488 231676
rect 511448 230376 511500 230382
rect 511448 230318 511500 230324
rect 510804 229900 510856 229906
rect 510804 229842 510856 229848
rect 511908 229900 511960 229906
rect 511908 229842 511960 229848
rect 510620 229288 510672 229294
rect 510620 229230 510672 229236
rect 510632 227322 510660 229230
rect 511920 229094 511948 229842
rect 511828 229066 511948 229094
rect 511080 227452 511132 227458
rect 511080 227394 511132 227400
rect 510620 227316 510672 227322
rect 510620 227258 510672 227264
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510160 224664 510212 224670
rect 510160 224606 510212 224612
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 509884 220380 509936 220386
rect 509884 220322 509936 220328
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 508516 217138 508544 217767
rect 509344 217274 509372 220322
rect 510172 217841 510200 224606
rect 510158 217832 510214 217841
rect 510158 217767 510214 217776
rect 509344 217246 509418 217274
rect 506032 217110 506106 217138
rect 506860 217110 506934 217138
rect 507688 217110 507762 217138
rect 508516 217110 508590 217138
rect 506078 216988 506106 217110
rect 506906 216988 506934 217110
rect 507734 216988 507762 217110
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510172 217138 510200 217767
rect 511092 217274 511120 227394
rect 511828 220726 511856 229066
rect 512104 228410 512132 231676
rect 512762 231662 513144 231690
rect 512092 228404 512144 228410
rect 512092 228346 512144 228352
rect 512736 228268 512788 228274
rect 512736 228210 512788 228216
rect 511816 220720 511868 220726
rect 511816 220662 511868 220668
rect 511816 220584 511868 220590
rect 511816 220526 511868 220532
rect 511046 217246 511120 217274
rect 511046 217190 511074 217246
rect 511034 217184 511086 217190
rect 510172 217110 510246 217138
rect 511034 217126 511086 217132
rect 511828 217138 511856 220526
rect 512748 218482 512776 228210
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513564 221740 513616 221746
rect 513564 221682 513616 221688
rect 513576 221513 513604 221682
rect 513562 221504 513618 221513
rect 513562 221439 513618 221448
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218476 512788 218482
rect 512736 218418 512788 218424
rect 512748 217274 512776 218418
rect 513576 217274 513604 221439
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 229906 515352 231676
rect 515312 229900 515364 229906
rect 515312 229842 515364 229848
rect 515404 229628 515456 229634
rect 515404 229570 515456 229576
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515416 220250 515444 229570
rect 515772 228676 515824 228682
rect 515772 228618 515824 228624
rect 515784 220862 515812 228618
rect 515968 223922 515996 231676
rect 516612 226030 516640 231676
rect 517256 230042 517284 231676
rect 517520 230376 517572 230382
rect 517520 230318 517572 230324
rect 517244 230036 517296 230042
rect 517244 229978 517296 229984
rect 516784 229764 516836 229770
rect 516784 229706 516836 229712
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 516600 224392 516652 224398
rect 516600 224334 516652 224340
rect 515956 223916 516008 223922
rect 515956 223858 516008 223864
rect 515772 220856 515824 220862
rect 515772 220798 515824 220804
rect 515220 220244 515272 220250
rect 515220 220186 515272 220192
rect 515404 220244 515456 220250
rect 515404 220186 515456 220192
rect 515232 219473 515260 220186
rect 515218 219464 515274 219473
rect 515218 219399 515274 219408
rect 515784 219434 515812 220798
rect 516612 219434 516640 224334
rect 516796 222018 516824 229706
rect 517532 223446 517560 230318
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229158 519216 231676
rect 519360 229288 519412 229294
rect 519360 229230 519412 229236
rect 519176 229152 519228 229158
rect 519176 229094 519228 229100
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 517704 228540 517756 228546
rect 517704 228482 517756 228488
rect 517716 224058 517744 228482
rect 519176 225888 519228 225894
rect 519176 225830 519228 225836
rect 517704 224052 517756 224058
rect 517704 223994 517756 224000
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 516784 222012 516836 222018
rect 516784 221954 516836 221960
rect 517532 220998 517560 222838
rect 517520 220992 517572 220998
rect 517520 220934 517572 220940
rect 517716 219434 517744 223994
rect 518440 220992 518492 220998
rect 518440 220934 518492 220940
rect 515784 219406 515996 219434
rect 516612 219406 516824 219434
rect 515232 217274 515260 219399
rect 514312 217246 514386 217274
rect 510218 216988 510246 217110
rect 511046 216988 511074 217126
rect 511828 217110 511902 217138
rect 511874 216988 511902 217110
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 217246 515260 217274
rect 515968 217274 515996 219406
rect 516796 217274 516824 219406
rect 517624 219406 517744 219434
rect 517624 217274 517652 219406
rect 518452 217274 518480 220934
rect 519188 219434 519216 225830
rect 519372 224942 519400 229230
rect 519360 224936 519412 224942
rect 519360 224878 519412 224884
rect 519832 222902 519860 231676
rect 520476 224670 520504 231676
rect 521120 230178 521148 231676
rect 521108 230172 521160 230178
rect 521108 230114 521160 230120
rect 521016 228948 521068 228954
rect 521016 228890 521068 228896
rect 520464 224664 520516 224670
rect 520464 224606 520516 224612
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 520188 221604 520240 221610
rect 520188 221546 520240 221552
rect 520200 221241 520228 221546
rect 520186 221232 520242 221241
rect 520186 221167 520242 221176
rect 519188 219406 519308 219434
rect 519280 217274 519308 219406
rect 520200 217274 520228 221167
rect 521028 221134 521056 228890
rect 521764 225894 521792 231676
rect 522422 231662 522712 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 521016 221128 521068 221134
rect 521016 221070 521068 221076
rect 521028 217274 521056 221070
rect 515968 217246 516042 217274
rect 516796 217246 516870 217274
rect 517624 217246 517698 217274
rect 518452 217246 518526 217274
rect 519280 217246 519354 217274
rect 515186 216988 515214 217246
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520982 217246 521056 217274
rect 521764 217274 521792 223110
rect 522684 221610 522712 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227186 523724 231676
rect 524248 231662 524354 231690
rect 523040 227180 523092 227186
rect 523040 227122 523092 227128
rect 523684 227180 523736 227186
rect 523684 227122 523736 227128
rect 522672 221604 522724 221610
rect 522672 221546 522724 221552
rect 522580 220380 522632 220386
rect 522580 220322 522632 220328
rect 522592 217841 522620 220322
rect 523052 217870 523080 227122
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 221882 523540 224198
rect 523500 221876 523552 221882
rect 523500 221818 523552 221824
rect 523040 217864 523092 217870
rect 522578 217832 522634 217841
rect 523040 217806 523092 217812
rect 522578 217767 522634 217776
rect 521764 217246 521838 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522592 217138 522620 217767
rect 523512 217274 523540 221818
rect 524248 221746 524276 231662
rect 524984 229158 525012 231676
rect 525536 231662 525642 231690
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 224262 524460 227258
rect 525536 224398 525564 231662
rect 525708 229900 525760 229906
rect 525708 229842 525760 229848
rect 525720 227594 525748 229842
rect 525708 227588 525760 227594
rect 525708 227530 525760 227536
rect 526272 227322 526300 231676
rect 526916 230450 526944 231676
rect 526904 230444 526956 230450
rect 526904 230386 526956 230392
rect 526444 230036 526496 230042
rect 526444 229978 526496 229984
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 526456 226166 526484 229978
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526628 227044 526680 227050
rect 526628 226986 526680 226992
rect 526444 226160 526496 226166
rect 526444 226102 526496 226108
rect 526352 224800 526404 224806
rect 526352 224742 526404 224748
rect 525524 224392 525576 224398
rect 525524 224334 525576 224340
rect 524420 224256 524472 224262
rect 524420 224198 524472 224204
rect 525064 224256 525116 224262
rect 525064 224198 525116 224204
rect 524236 221740 524288 221746
rect 524236 221682 524288 221688
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 523466 217246 523540 217274
rect 522592 217110 522666 217138
rect 522638 216988 522666 217110
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 224198
rect 525984 217728 526036 217734
rect 525984 217670 526036 217676
rect 525996 217274 526024 217670
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526364 217274 526392 224742
rect 526640 219434 526668 226986
rect 527180 223032 527232 223038
rect 527180 222974 527232 222980
rect 527192 221338 527220 222974
rect 527548 222012 527600 222018
rect 527548 221954 527600 221960
rect 527180 221332 527232 221338
rect 527180 221274 527232 221280
rect 527560 219910 527588 221954
rect 528192 221332 528244 221338
rect 528192 221274 528244 221280
rect 527548 219904 527600 219910
rect 527548 219846 527600 219852
rect 526548 219406 526668 219434
rect 526548 217734 526576 219406
rect 526536 217728 526588 217734
rect 526536 217670 526588 217676
rect 526548 217462 526576 217670
rect 526536 217456 526588 217462
rect 526536 217398 526588 217404
rect 527560 217274 527588 219846
rect 528204 219434 528232 221274
rect 528388 220386 528416 231662
rect 528848 230314 528876 231676
rect 528836 230308 528888 230314
rect 528836 230250 528888 230256
rect 529204 230172 529256 230178
rect 529204 230114 529256 230120
rect 529216 229094 529244 230114
rect 529032 229066 529244 229094
rect 529032 220658 529060 229066
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 529020 220652 529072 220658
rect 529020 220594 529072 220600
rect 528376 220380 528428 220386
rect 528376 220322 528428 220328
rect 528204 219406 528416 219434
rect 528388 217274 528416 219406
rect 529216 217274 529244 225694
rect 529492 223174 529520 231676
rect 530136 229634 530164 231676
rect 530124 229628 530176 229634
rect 530124 229570 530176 229576
rect 530780 229498 530808 231676
rect 531136 229628 531188 229634
rect 531136 229570 531188 229576
rect 530768 229492 530820 229498
rect 530768 229434 530820 229440
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 224806 529980 229094
rect 530584 225616 530636 225622
rect 530584 225558 530636 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 529480 223168 529532 223174
rect 529480 223110 529532 223116
rect 530032 220244 530084 220250
rect 530032 220186 530084 220192
rect 530044 219910 530072 220186
rect 530032 219904 530084 219910
rect 530032 219846 530084 219852
rect 530044 217274 530072 219846
rect 530596 217598 530624 225558
rect 531148 220250 531176 229570
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 532068 223038 532096 231676
rect 532712 230178 532740 231676
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 532976 228404 533028 228410
rect 532976 228346 533028 228352
rect 532516 223440 532568 223446
rect 532516 223382 532568 223388
rect 532056 223032 532108 223038
rect 532056 222974 532108 222980
rect 532528 222766 532556 223382
rect 532516 222760 532568 222766
rect 532516 222702 532568 222708
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 531136 220244 531188 220250
rect 531136 220186 531188 220192
rect 530584 217592 530636 217598
rect 530584 217534 530636 217540
rect 530952 217592 531004 217598
rect 530952 217534 531004 217540
rect 526364 217246 526806 217274
rect 527560 217246 527634 217274
rect 528388 217246 528462 217274
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528434 216988 528462 217246
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217534
rect 531700 217274 531728 220458
rect 532528 217274 532556 222702
rect 532988 219434 533016 228346
rect 533356 227050 533384 231676
rect 533344 227044 533396 227050
rect 533344 226986 533396 226992
rect 533528 222760 533580 222766
rect 533528 222702 533580 222708
rect 533540 222494 533568 222702
rect 533344 222488 533396 222494
rect 533344 222430 533396 222436
rect 533528 222488 533580 222494
rect 533528 222430 533580 222436
rect 533356 222222 533384 222430
rect 533344 222216 533396 222222
rect 533344 222158 533396 222164
rect 533160 222080 533212 222086
rect 533160 222022 533212 222028
rect 533172 221474 533200 222022
rect 534000 221950 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534816 229764 534868 229770
rect 534816 229706 534868 229712
rect 534828 223446 534856 229706
rect 535000 224936 535052 224942
rect 535000 224878 535052 224884
rect 534816 223440 534868 223446
rect 534816 223382 534868 223388
rect 533988 221944 534040 221950
rect 533988 221886 534040 221892
rect 533712 221876 533764 221882
rect 533712 221818 533764 221824
rect 533528 221604 533580 221610
rect 533528 221546 533580 221552
rect 533160 221468 533212 221474
rect 533160 221410 533212 221416
rect 533540 221338 533568 221546
rect 533528 221332 533580 221338
rect 533528 221274 533580 221280
rect 533724 221270 533752 221818
rect 533712 221264 533764 221270
rect 533712 221206 533764 221212
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 532988 219406 533476 219434
rect 533448 217734 533476 219406
rect 533436 217728 533488 217734
rect 533436 217670 533488 217676
rect 531700 217246 531774 217274
rect 532528 217246 532602 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532574 216988 532602 217246
rect 533448 217138 533476 217670
rect 534184 217274 534212 220050
rect 535012 217274 535040 224878
rect 535288 224534 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 224528 535328 224534
rect 535276 224470 535328 224476
rect 535460 223304 535512 223310
rect 535460 223246 535512 223252
rect 535472 217870 535500 223246
rect 535748 219434 535776 227394
rect 535932 225758 535960 231676
rect 536104 230444 536156 230450
rect 536104 230386 536156 230392
rect 536116 227458 536144 230386
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 537484 227588 537536 227594
rect 537484 227530 537536 227536
rect 536104 227452 536156 227458
rect 536104 227394 536156 227400
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 535748 219406 535868 219434
rect 535460 217864 535512 217870
rect 535460 217806 535512 217812
rect 535840 217326 535868 219406
rect 537496 218618 537524 227530
rect 538140 220114 538168 231662
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538312 229628 538364 229634
rect 538312 229570 538364 229576
rect 538324 226030 538352 229570
rect 538496 226160 538548 226166
rect 538496 226102 538548 226108
rect 538312 226024 538364 226030
rect 538312 225966 538364 225972
rect 538508 225842 538536 226102
rect 538324 225814 538536 225842
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 538324 219434 538352 225814
rect 538496 223916 538548 223922
rect 538496 223858 538548 223864
rect 538508 219434 538536 223858
rect 538784 222086 538812 231662
rect 539600 230308 539652 230314
rect 539600 230250 539652 230256
rect 539612 228682 539640 230250
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 542452 228948 542504 228954
rect 542452 228890 542504 228896
rect 541624 228812 541676 228818
rect 541624 228754 541676 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540888 228268 540940 228274
rect 540888 228210 540940 228216
rect 539968 226296 540020 226302
rect 539968 226238 540020 226244
rect 539508 223916 539560 223922
rect 539508 223858 539560 223864
rect 539520 222086 539548 223858
rect 539980 223786 540008 226238
rect 539968 223780 540020 223786
rect 539968 223722 540020 223728
rect 538772 222080 538824 222086
rect 538772 222022 538824 222028
rect 539508 222080 539560 222086
rect 539508 222022 539560 222028
rect 538232 219406 538352 219434
rect 538416 219406 538536 219434
rect 537484 218612 537536 218618
rect 537484 218554 537536 218560
rect 536656 217864 536708 217870
rect 536656 217806 536708 217812
rect 536840 217864 536892 217870
rect 536840 217806 536892 217812
rect 535828 217320 535880 217326
rect 534184 217246 534258 217274
rect 535012 217246 535086 217274
rect 535828 217262 535880 217268
rect 533402 217110 533476 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217246
rect 535058 216988 535086 217246
rect 535840 217138 535868 217262
rect 536668 217138 536696 217806
rect 536852 217598 536880 217806
rect 536840 217592 536892 217598
rect 536840 217534 536892 217540
rect 537496 217274 537524 218554
rect 538232 217598 538260 219406
rect 538220 217592 538272 217598
rect 538220 217534 538272 217540
rect 538416 217274 538444 219406
rect 539140 217592 539192 217598
rect 539140 217534 539192 217540
rect 537496 217246 537570 217274
rect 535840 217110 535914 217138
rect 536668 217110 536742 217138
rect 535886 216988 535914 217110
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539152 217138 539180 217534
rect 539980 217274 540008 223722
rect 540900 221785 540928 228210
rect 540886 221776 540942 221785
rect 540886 221711 540942 221720
rect 540612 218748 540664 218754
rect 540612 218690 540664 218696
rect 540624 218482 540652 218690
rect 540612 218476 540664 218482
rect 540612 218418 540664 218424
rect 540900 217274 540928 221711
rect 539980 217246 540054 217274
rect 539152 217110 539226 217138
rect 539198 216988 539226 217110
rect 540026 216988 540054 217246
rect 540854 217246 540928 217274
rect 541636 217274 541664 228754
rect 542464 223922 542492 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 544108 224664 544160 224670
rect 544108 224606 544160 224612
rect 542452 223916 542504 223922
rect 542452 223858 542504 223864
rect 542464 217274 542492 223858
rect 543372 222896 543424 222902
rect 543372 222838 543424 222844
rect 543186 222320 543242 222329
rect 543186 222255 543242 222264
rect 543200 222086 543228 222255
rect 543384 222086 543412 222838
rect 543188 222080 543240 222086
rect 543188 222022 543240 222028
rect 543372 222080 543424 222086
rect 543372 222022 543424 222028
rect 543384 217274 543412 222022
rect 541636 217246 541710 217274
rect 542464 217246 542538 217274
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542510 216988 542538 217246
rect 543338 217246 543412 217274
rect 544120 217274 544148 224606
rect 544936 220652 544988 220658
rect 544936 220594 544988 220600
rect 544948 218890 544976 220594
rect 544936 218884 544988 218890
rect 544936 218826 544988 218832
rect 544948 217274 544976 218826
rect 545776 217598 545804 225830
rect 547156 222086 547184 230114
rect 549260 230036 549312 230042
rect 549260 229978 549312 229984
rect 548156 227180 548208 227186
rect 548156 227122 548208 227128
rect 548168 224210 548196 227122
rect 548340 224800 548392 224806
rect 548340 224742 548392 224748
rect 548352 224398 548380 224742
rect 549272 224670 549300 229978
rect 553216 228540 553268 228546
rect 553216 228482 553268 228488
rect 552480 227452 552532 227458
rect 552480 227394 552532 227400
rect 551560 227316 551612 227322
rect 551560 227258 551612 227264
rect 550824 224800 550876 224806
rect 550824 224742 550876 224748
rect 549076 224664 549128 224670
rect 549076 224606 549128 224612
rect 549260 224664 549312 224670
rect 549260 224606 549312 224612
rect 549088 224482 549116 224606
rect 549088 224454 549300 224482
rect 548340 224392 548392 224398
rect 548340 224334 548392 224340
rect 548524 224392 548576 224398
rect 548524 224334 548576 224340
rect 548168 224182 548380 224210
rect 547512 223440 547564 223446
rect 547512 223382 547564 223388
rect 546960 222080 547012 222086
rect 546958 222048 546960 222057
rect 547144 222080 547196 222086
rect 547012 222048 547014 222057
rect 547144 222022 547196 222028
rect 546958 221983 547014 221992
rect 546774 221776 546830 221785
rect 546774 221711 546830 221720
rect 546788 221474 546816 221711
rect 546592 221468 546644 221474
rect 546592 221410 546644 221416
rect 546776 221468 546828 221474
rect 546776 221410 546828 221416
rect 545764 217592 545816 217598
rect 545764 217534 545816 217540
rect 545776 217274 545804 217534
rect 546604 217274 546632 221410
rect 547524 218754 547552 223382
rect 547694 222320 547750 222329
rect 547694 222255 547750 222264
rect 547708 222170 547736 222255
rect 547708 222142 547920 222170
rect 547892 222086 547920 222142
rect 547696 222080 547748 222086
rect 547696 222022 547748 222028
rect 547880 222080 547932 222086
rect 547880 222022 547932 222028
rect 547708 221898 547736 222022
rect 547708 221870 547920 221898
rect 547892 221814 547920 221870
rect 547880 221808 547932 221814
rect 547694 221776 547750 221785
rect 547880 221750 547932 221756
rect 547694 221711 547696 221720
rect 547748 221711 547750 221720
rect 547696 221682 547748 221688
rect 548352 220522 548380 224182
rect 548536 223922 548564 224334
rect 549272 223922 549300 224454
rect 548524 223916 548576 223922
rect 548524 223858 548576 223864
rect 549260 223916 549312 223922
rect 549260 223858 549312 223864
rect 549904 223916 549956 223922
rect 549904 223858 549956 223864
rect 549074 221776 549130 221785
rect 549074 221711 549130 221720
rect 548340 220516 548392 220522
rect 548340 220458 548392 220464
rect 547512 218748 547564 218754
rect 547512 218690 547564 218696
rect 547524 217274 547552 218690
rect 548352 217274 548380 220458
rect 544120 217246 544194 217274
rect 544948 217246 545022 217274
rect 545776 217246 545850 217274
rect 546604 217246 546678 217274
rect 543338 216988 543366 217246
rect 544166 216988 544194 217246
rect 544994 216988 545022 217246
rect 545822 216988 545850 217246
rect 546650 216988 546678 217246
rect 547478 217246 547552 217274
rect 548306 217246 548380 217274
rect 549088 217274 549116 221711
rect 549916 217274 549944 223858
rect 550836 220658 550864 224742
rect 550824 220652 550876 220658
rect 550824 220594 550876 220600
rect 550836 217274 550864 220594
rect 551192 220516 551244 220522
rect 551192 220458 551244 220464
rect 551204 220153 551232 220458
rect 551190 220144 551246 220153
rect 551190 220079 551246 220088
rect 549088 217246 549162 217274
rect 549916 217246 549990 217274
rect 547478 216988 547506 217246
rect 548306 216988 548334 217246
rect 549134 216988 549162 217246
rect 549962 216988 549990 217246
rect 550790 217246 550864 217274
rect 551572 217274 551600 227258
rect 552296 220244 552348 220250
rect 552296 220186 552348 220192
rect 552308 219201 552336 220186
rect 552492 219434 552520 227394
rect 552664 220244 552716 220250
rect 552664 220186 552716 220192
rect 552676 219910 552704 220186
rect 552846 220144 552902 220153
rect 552846 220079 552902 220088
rect 552860 219910 552888 220079
rect 552664 219904 552716 219910
rect 552664 219846 552716 219852
rect 552848 219904 552900 219910
rect 552848 219846 552900 219852
rect 552492 219406 552704 219434
rect 552294 219192 552350 219201
rect 552676 219162 552704 219406
rect 553228 219366 553256 228482
rect 554056 222902 554084 249047
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 554964 228676 555016 228682
rect 554964 228618 555016 228624
rect 554976 225078 555004 228618
rect 555436 228546 555464 255546
rect 556804 251252 556856 251258
rect 556804 251194 556856 251200
rect 555424 228540 555476 228546
rect 555424 228482 555476 228488
rect 556816 227186 556844 251194
rect 558184 246356 558236 246362
rect 558184 246298 558236 246304
rect 558196 236094 558224 246298
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 556804 227180 556856 227186
rect 556804 227122 556856 227128
rect 556160 226024 556212 226030
rect 556160 225966 556212 225972
rect 554964 225072 555016 225078
rect 554964 225014 555016 225020
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 553858 222048 553914 222057
rect 553858 221983 553914 221992
rect 553872 221882 553900 221983
rect 553860 221876 553912 221882
rect 553860 221818 553912 221824
rect 553492 221808 553544 221814
rect 553490 221776 553492 221785
rect 553544 221776 553546 221785
rect 553490 221711 553546 221720
rect 553952 220380 554004 220386
rect 553952 220322 554004 220328
rect 553216 219360 553268 219366
rect 553216 219302 553268 219308
rect 552294 219127 552350 219136
rect 552664 219156 552716 219162
rect 552664 219098 552716 219104
rect 552480 219020 552532 219026
rect 552480 218962 552532 218968
rect 552492 218618 552520 218962
rect 552480 218612 552532 218618
rect 552480 218554 552532 218560
rect 552676 217274 552704 219098
rect 551572 217246 551646 217274
rect 550790 216988 550818 217246
rect 551618 216988 551646 217246
rect 552446 217246 552704 217274
rect 553228 217274 553256 219302
rect 553964 217274 553992 220322
rect 554976 217274 555004 225014
rect 556172 224806 556200 225966
rect 558184 225616 558236 225622
rect 558184 225558 558236 225564
rect 558196 224954 558224 225558
rect 559104 225072 559156 225078
rect 559104 225014 559156 225020
rect 558012 224926 558224 224954
rect 555792 224800 555844 224806
rect 555792 224742 555844 224748
rect 556160 224800 556212 224806
rect 556160 224742 556212 224748
rect 557356 224800 557408 224806
rect 557356 224742 557408 224748
rect 555804 224505 555832 224742
rect 555790 224496 555846 224505
rect 555790 224431 555846 224440
rect 555700 223168 555752 223174
rect 555700 223110 555752 223116
rect 555712 217841 555740 223110
rect 556526 219192 556582 219201
rect 556526 219127 556582 219136
rect 555976 218884 556028 218890
rect 555976 218826 556028 218832
rect 555988 218618 556016 218826
rect 555976 218612 556028 218618
rect 555976 218554 556028 218560
rect 555698 217832 555754 217841
rect 555698 217767 555754 217776
rect 553228 217246 553302 217274
rect 553964 217246 554130 217274
rect 552446 216988 552474 217246
rect 553274 216988 553302 217246
rect 554102 216988 554130 217246
rect 554930 217246 555004 217274
rect 554930 216988 554958 217246
rect 555712 217138 555740 217767
rect 556540 217138 556568 219127
rect 557368 217274 557396 224742
rect 557816 224664 557868 224670
rect 557816 224606 557868 224612
rect 557828 223922 557856 224606
rect 557816 223916 557868 223922
rect 557816 223858 557868 223864
rect 557540 223168 557592 223174
rect 557540 223110 557592 223116
rect 557552 221785 557580 223110
rect 558012 222465 558040 224926
rect 559116 224806 559144 225014
rect 558828 224800 558880 224806
rect 558828 224742 558880 224748
rect 559104 224800 559156 224806
rect 559104 224742 559156 224748
rect 558840 224398 558868 224742
rect 558184 224392 558236 224398
rect 558184 224334 558236 224340
rect 558828 224392 558880 224398
rect 558828 224334 558880 224340
rect 558196 223922 558224 224334
rect 558184 223916 558236 223922
rect 558184 223858 558236 223864
rect 559012 223032 559064 223038
rect 559012 222974 559064 222980
rect 558184 222760 558236 222766
rect 558184 222702 558236 222708
rect 557998 222456 558054 222465
rect 557998 222391 558054 222400
rect 557538 221776 557594 221785
rect 557538 221711 557594 221720
rect 558012 217274 558040 222391
rect 558196 222222 558224 222702
rect 558184 222216 558236 222222
rect 558184 222158 558236 222164
rect 558184 220380 558236 220386
rect 558184 220322 558236 220328
rect 558196 220114 558224 220322
rect 558184 220108 558236 220114
rect 558184 220050 558236 220056
rect 558368 220040 558420 220046
rect 558368 219982 558420 219988
rect 558380 219774 558408 219982
rect 558368 219768 558420 219774
rect 558368 219710 558420 219716
rect 558552 219768 558604 219774
rect 558552 219710 558604 219716
rect 558564 219366 558592 219710
rect 558552 219360 558604 219366
rect 558552 219302 558604 219308
rect 558184 219156 558236 219162
rect 558184 219098 558236 219104
rect 558196 218754 558224 219098
rect 558184 218748 558236 218754
rect 558184 218690 558236 218696
rect 557368 217246 557442 217274
rect 558012 217246 558270 217274
rect 555712 217110 555786 217138
rect 556540 217110 556614 217138
rect 555758 216988 555786 217110
rect 556586 216988 556614 217110
rect 557414 216988 557442 217246
rect 558242 216988 558270 217246
rect 559024 217138 559052 222974
rect 559378 221776 559434 221785
rect 559576 221746 559604 229842
rect 560760 227044 560812 227050
rect 560760 226986 560812 226992
rect 559932 223168 559984 223174
rect 559932 223110 559984 223116
rect 559378 221711 559380 221720
rect 559432 221711 559434 221720
rect 559564 221740 559616 221746
rect 559380 221682 559432 221688
rect 559564 221682 559616 221688
rect 559944 217138 559972 223110
rect 560772 220522 560800 226986
rect 560956 222154 560984 259422
rect 563704 256760 563756 256766
rect 563704 256702 563756 256708
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 562336 231854 562364 252554
rect 562336 231826 562732 231854
rect 562704 224806 562732 231826
rect 563716 226302 563744 256702
rect 566464 229764 566516 229770
rect 566464 229706 566516 229712
rect 566476 229094 566504 229706
rect 566476 229066 566688 229094
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563704 226296 563756 226302
rect 563704 226238 563756 226244
rect 563060 225752 563112 225758
rect 563060 225694 563112 225700
rect 562692 224800 562744 224806
rect 562692 224742 562744 224748
rect 562140 224664 562192 224670
rect 562192 224612 562364 224618
rect 562140 224606 562364 224612
rect 562152 224590 562364 224606
rect 562336 224534 562364 224590
rect 562140 224528 562192 224534
rect 561678 224496 561734 224505
rect 562140 224470 562192 224476
rect 562324 224528 562376 224534
rect 562324 224470 562376 224476
rect 561678 224431 561734 224440
rect 561692 222193 561720 224431
rect 562152 224369 562180 224470
rect 562138 224360 562194 224369
rect 562138 224295 562194 224304
rect 562876 223168 562928 223174
rect 562876 223110 562928 223116
rect 562888 222222 562916 223110
rect 562876 222216 562928 222222
rect 561678 222184 561734 222193
rect 560944 222148 560996 222154
rect 562690 222184 562746 222193
rect 561678 222119 561734 222128
rect 562508 222148 562560 222154
rect 560944 222090 560996 222096
rect 562876 222158 562928 222164
rect 562690 222119 562746 222128
rect 562508 222090 562560 222096
rect 561494 221776 561550 221785
rect 561494 221711 561550 221720
rect 560760 220516 560812 220522
rect 560760 220458 560812 220464
rect 560772 217274 560800 220458
rect 559024 217110 559098 217138
rect 559070 216988 559098 217110
rect 559898 217110 559972 217138
rect 560726 217246 560800 217274
rect 559898 216988 559926 217110
rect 560726 216988 560754 217246
rect 561508 217138 561536 221711
rect 562520 221626 562548 222090
rect 562704 221746 562732 222119
rect 562692 221740 562744 221746
rect 562692 221682 562744 221688
rect 562876 221740 562928 221746
rect 562876 221682 562928 221688
rect 562888 221626 562916 221682
rect 562520 221598 562916 221626
rect 562874 220688 562930 220697
rect 562874 220623 562930 220632
rect 562888 220522 562916 220623
rect 562876 220516 562928 220522
rect 562876 220458 562928 220464
rect 561864 219292 561916 219298
rect 561864 219234 561916 219240
rect 561876 217190 561904 219234
rect 562322 219192 562378 219201
rect 563072 219162 563100 225694
rect 563242 224360 563298 224369
rect 563242 224295 563298 224304
rect 563256 220658 563284 224295
rect 564806 222184 564862 222193
rect 564806 222119 564862 222128
rect 564820 221785 564848 222119
rect 564806 221776 564862 221785
rect 564806 221711 564862 221720
rect 563244 220652 563296 220658
rect 563244 220594 563296 220600
rect 563256 219434 563284 220594
rect 563256 219406 563376 219434
rect 562322 219127 562378 219136
rect 563060 219156 563112 219162
rect 561864 217184 561916 217190
rect 561508 217110 561582 217138
rect 562336 217172 562364 219127
rect 563060 219098 563112 219104
rect 562520 217926 563008 217954
rect 562336 217144 562410 217172
rect 561864 217126 561916 217132
rect 561554 216988 561582 217110
rect 562382 216988 562410 217144
rect 562520 217122 562548 217926
rect 562980 217841 563008 217926
rect 562690 217832 562746 217841
rect 562690 217767 562746 217776
rect 562966 217832 563022 217841
rect 562966 217767 563022 217776
rect 562704 217172 562732 217767
rect 563348 217274 563376 219406
rect 563980 219156 564032 219162
rect 563980 219098 564032 219104
rect 563210 217246 563376 217274
rect 562876 217184 562928 217190
rect 562704 217144 562876 217172
rect 562876 217126 562928 217132
rect 562508 217116 562560 217122
rect 562508 217058 562560 217064
rect 563210 216988 563238 217246
rect 563992 217138 564020 219098
rect 564820 217274 564848 221711
rect 565648 220425 565676 228346
rect 565634 220416 565690 220425
rect 565634 220351 565690 220360
rect 566464 220380 566516 220386
rect 565084 219292 565136 219298
rect 565084 219234 565136 219240
rect 564820 217246 564894 217274
rect 563992 217110 564066 217138
rect 564038 216988 564066 217110
rect 564866 216988 564894 217246
rect 565096 217190 565124 219234
rect 565648 217274 565676 220351
rect 566464 220322 566516 220328
rect 566476 217274 566504 220322
rect 566660 220318 566688 229066
rect 568120 226296 568172 226302
rect 568120 226238 568172 226244
rect 567014 222456 567070 222465
rect 567014 222391 567070 222400
rect 567028 221898 567056 222391
rect 567028 221870 567240 221898
rect 567212 221746 567240 221870
rect 567016 221740 567068 221746
rect 567016 221682 567068 221688
rect 567200 221740 567252 221746
rect 567200 221682 567252 221688
rect 567028 220726 567056 221682
rect 567212 220782 567700 220810
rect 567212 220726 567240 220782
rect 567016 220720 567068 220726
rect 567016 220662 567068 220668
rect 567200 220720 567252 220726
rect 567200 220662 567252 220668
rect 566832 220652 566884 220658
rect 566832 220594 566884 220600
rect 567384 220652 567436 220658
rect 567384 220594 567436 220600
rect 566648 220312 566700 220318
rect 566648 220254 566700 220260
rect 566844 220153 566872 220594
rect 567396 220425 567424 220594
rect 567672 220425 567700 220782
rect 567382 220416 567438 220425
rect 567382 220351 567438 220360
rect 567658 220416 567714 220425
rect 567658 220351 567714 220360
rect 567844 220380 567896 220386
rect 567844 220322 567896 220328
rect 567154 220312 567206 220318
rect 567206 220260 567240 220266
rect 567154 220254 567240 220260
rect 567166 220238 567240 220254
rect 566830 220144 566886 220153
rect 566830 220079 566886 220088
rect 567212 219434 567240 220238
rect 567856 220153 567884 220322
rect 567842 220144 567898 220153
rect 567842 220079 567898 220088
rect 567212 219406 567332 219434
rect 567304 219162 567332 219406
rect 567292 219156 567344 219162
rect 567292 219098 567344 219104
rect 567304 217274 567332 219098
rect 568132 217274 568160 226238
rect 568396 219292 568448 219298
rect 568396 219234 568448 219240
rect 568408 218482 568436 219234
rect 568592 218482 568620 260850
rect 570616 234598 570644 261462
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 573364 244316 573416 244322
rect 573364 244258 573416 244264
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 571340 228540 571392 228546
rect 571340 228482 571392 228488
rect 570604 227180 570656 227186
rect 570604 227122 570656 227128
rect 569590 221776 569646 221785
rect 569590 221711 569646 221720
rect 568946 220416 569002 220425
rect 568946 220351 569002 220360
rect 568396 218476 568448 218482
rect 568396 218418 568448 218424
rect 568580 218476 568632 218482
rect 568580 218418 568632 218424
rect 568960 217274 568988 220351
rect 569222 219192 569278 219201
rect 569222 219127 569278 219136
rect 569236 218890 569264 219127
rect 569604 219026 569632 221711
rect 569592 219020 569644 219026
rect 569592 218962 569644 218968
rect 569224 218884 569276 218890
rect 569224 218826 569276 218832
rect 569776 218476 569828 218482
rect 569776 218418 569828 218424
rect 565648 217246 565722 217274
rect 566476 217246 566550 217274
rect 567304 217246 567378 217274
rect 568132 217246 568206 217274
rect 568960 217246 569034 217274
rect 565084 217184 565136 217190
rect 565084 217126 565136 217132
rect 565694 216988 565722 217246
rect 566522 216988 566550 217246
rect 567350 216988 567378 217246
rect 568178 216988 568206 217246
rect 569006 216988 569034 217246
rect 569788 217138 569816 218418
rect 570616 217274 570644 227122
rect 571352 218482 571380 228482
rect 571524 224800 571576 224806
rect 571524 224742 571576 224748
rect 571340 218476 571392 218482
rect 571340 218418 571392 218424
rect 571536 217274 571564 224742
rect 573376 220289 573404 244258
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 576766 220688 576822 220697
rect 576766 220623 576822 220632
rect 573362 220280 573418 220289
rect 576780 220250 576808 220623
rect 573362 220215 573418 220224
rect 576768 220244 576820 220250
rect 576768 220186 576820 220192
rect 576584 220176 576636 220182
rect 576584 220118 576636 220124
rect 576596 220017 576624 220118
rect 576780 220102 577176 220130
rect 576780 220046 576808 220102
rect 576768 220040 576820 220046
rect 576582 220008 576638 220017
rect 576768 219982 576820 219988
rect 576952 220040 577004 220046
rect 576952 219982 577004 219988
rect 576582 219943 576638 219952
rect 576768 219632 576820 219638
rect 576964 219586 576992 219982
rect 576820 219580 576992 219586
rect 576768 219574 576992 219580
rect 576780 219558 576992 219574
rect 577148 219452 577176 220102
rect 571628 219422 572484 219450
rect 571628 218770 571656 219422
rect 572456 219366 572484 219422
rect 577136 219446 577188 219452
rect 577136 219388 577188 219394
rect 572444 219360 572496 219366
rect 572444 219302 572496 219308
rect 574652 219360 574704 219366
rect 574652 219302 574704 219308
rect 571984 219292 572036 219298
rect 571984 219234 572036 219240
rect 571628 218754 571748 218770
rect 571996 218754 572024 219234
rect 572626 219192 572682 219201
rect 572626 219127 572682 219136
rect 572640 218890 572668 219127
rect 572444 218884 572496 218890
rect 572444 218826 572496 218832
rect 572628 218884 572680 218890
rect 572628 218826 572680 218832
rect 571628 218748 571760 218754
rect 571628 218742 571708 218748
rect 571708 218690 571760 218696
rect 571984 218748 572036 218754
rect 571984 218690 572036 218696
rect 572456 218482 572484 218826
rect 572260 218476 572312 218482
rect 572260 218418 572312 218424
rect 572444 218476 572496 218482
rect 572444 218418 572496 218424
rect 570616 217246 570690 217274
rect 569788 217110 569862 217138
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571490 217246 571564 217274
rect 571490 216988 571518 217246
rect 572272 217138 572300 218418
rect 574098 217832 574154 217841
rect 574098 217767 574154 217776
rect 572272 217110 572346 217138
rect 572318 216988 572346 217110
rect 574112 216918 574140 217767
rect 574100 216912 574152 216918
rect 574100 216854 574152 216860
rect 574098 216744 574154 216753
rect 574098 216679 574154 216688
rect 574374 216744 574430 216753
rect 574374 216679 574430 216688
rect 574112 213518 574140 216679
rect 574100 213512 574152 213518
rect 574100 213454 574152 213460
rect 574388 213382 574416 216679
rect 574664 214606 574692 219302
rect 575020 218884 575072 218890
rect 575020 218826 575072 218832
rect 574834 217832 574890 217841
rect 574834 217767 574890 217776
rect 574652 214600 574704 214606
rect 574652 214542 574704 214548
rect 574376 213376 574428 213382
rect 574376 213318 574428 213324
rect 574848 213246 574876 217767
rect 575032 214742 575060 218826
rect 575480 218748 575532 218754
rect 575480 218690 575532 218696
rect 575492 214878 575520 218690
rect 575480 214872 575532 214878
rect 575480 214814 575532 214820
rect 575020 214736 575072 214742
rect 575020 214678 575072 214684
rect 574836 213240 574888 213246
rect 574836 213182 574888 213188
rect 577516 99142 577544 240110
rect 596836 231130 596864 245618
rect 648632 242214 648660 278052
rect 650642 256728 650698 256737
rect 650642 256663 650698 256672
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 596824 231124 596876 231130
rect 596824 231066 596876 231072
rect 629956 229094 629984 241470
rect 639604 232552 639656 232558
rect 639604 232494 639656 232500
rect 633624 231124 633676 231130
rect 633624 231066 633676 231072
rect 636844 231124 636896 231130
rect 636844 231066 636896 231072
rect 629956 229066 630076 229094
rect 621020 224936 621072 224942
rect 621020 224878 621072 224884
rect 610992 224800 611044 224806
rect 610992 224742 611044 224748
rect 610624 224664 610676 224670
rect 610624 224606 610676 224612
rect 610636 224058 610664 224606
rect 610808 224528 610860 224534
rect 610808 224470 610860 224476
rect 610624 224052 610676 224058
rect 610624 223994 610676 224000
rect 610820 223922 610848 224470
rect 611004 224058 611032 224742
rect 617064 224664 617116 224670
rect 617064 224606 617116 224612
rect 610992 224052 611044 224058
rect 610992 223994 611044 224000
rect 610624 223916 610676 223922
rect 610624 223858 610676 223864
rect 610808 223916 610860 223922
rect 610808 223858 610860 223864
rect 610636 223650 610664 223858
rect 610624 223644 610676 223650
rect 610624 223586 610676 223592
rect 614948 223508 615000 223514
rect 614948 223450 615000 223456
rect 593972 222624 594024 222630
rect 593972 222566 594024 222572
rect 582470 220280 582526 220289
rect 582470 220215 582526 220224
rect 582484 220114 582512 220215
rect 582472 220108 582524 220114
rect 582472 220050 582524 220056
rect 581644 220040 581696 220046
rect 581828 220040 581880 220046
rect 581644 219982 581696 219988
rect 581826 220008 581828 220017
rect 582334 220040 582386 220046
rect 581880 220008 581882 220017
rect 581656 219638 581684 219982
rect 582386 219988 582696 219994
rect 582334 219982 582696 219988
rect 582346 219966 582696 219982
rect 581826 219943 581882 219952
rect 581644 219632 581696 219638
rect 581644 219574 581696 219580
rect 582334 219632 582386 219638
rect 582334 219574 582386 219580
rect 582472 219632 582524 219638
rect 582472 219574 582524 219580
rect 582346 219178 582374 219574
rect 582484 219366 582512 219574
rect 582668 219366 582696 219966
rect 591580 219496 591632 219502
rect 591632 219444 591988 219450
rect 591580 219438 591988 219444
rect 591592 219422 591988 219438
rect 591960 219366 591988 219422
rect 582472 219360 582524 219366
rect 582472 219302 582524 219308
rect 582656 219360 582708 219366
rect 582656 219302 582708 219308
rect 591948 219360 592000 219366
rect 591948 219302 592000 219308
rect 582346 219150 582420 219178
rect 582392 218890 582420 219150
rect 582380 218884 582432 218890
rect 582380 218826 582432 218832
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578330 211712 578386 211721
rect 578330 211647 578386 211656
rect 578344 211206 578372 211647
rect 578332 211200 578384 211206
rect 578332 211142 578384 211148
rect 578896 208350 578924 213959
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 593984 210202 594012 222566
rect 598572 222080 598624 222086
rect 598572 222022 598624 222028
rect 598584 221354 598612 222022
rect 598756 222012 598808 222018
rect 598756 221954 598808 221960
rect 603080 222012 603132 222018
rect 603080 221954 603132 221960
rect 598768 221610 598796 221954
rect 598940 221876 598992 221882
rect 598940 221818 598992 221824
rect 599124 221876 599176 221882
rect 599124 221818 599176 221824
rect 598952 221610 598980 221818
rect 598756 221604 598808 221610
rect 598756 221546 598808 221552
rect 598940 221604 598992 221610
rect 598940 221546 598992 221552
rect 599136 221474 599164 221818
rect 599490 221504 599546 221513
rect 599124 221468 599176 221474
rect 599490 221439 599546 221448
rect 599124 221410 599176 221416
rect 599308 221400 599360 221406
rect 598584 221348 599308 221354
rect 598584 221342 599360 221348
rect 598584 221326 599348 221342
rect 598388 219904 598440 219910
rect 598388 219846 598440 219852
rect 598572 219904 598624 219910
rect 598572 219846 598624 219852
rect 598400 219450 598428 219846
rect 598584 219638 598612 219846
rect 598572 219632 598624 219638
rect 598572 219574 598624 219580
rect 598940 219496 598992 219502
rect 598400 219444 598940 219450
rect 598400 219438 598992 219444
rect 598400 219422 598980 219438
rect 596824 219360 596876 219366
rect 596824 219302 596876 219308
rect 594798 218648 594854 218657
rect 594798 218583 594854 218592
rect 594812 216782 594840 218583
rect 595166 217560 595222 217569
rect 595166 217495 595222 217504
rect 594800 216776 594852 216782
rect 594800 216718 594852 216724
rect 594800 213512 594852 213518
rect 594800 213454 594852 213460
rect 594812 210202 594840 213454
rect 595180 210202 595208 217495
rect 596362 217288 596418 217297
rect 596362 217223 596418 217232
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596376 210202 596404 217223
rect 596836 210202 596864 219302
rect 597928 218884 597980 218890
rect 597928 218826 597980 218832
rect 597560 216912 597612 216918
rect 597560 216854 597612 216860
rect 597572 210202 597600 216854
rect 597940 210202 597968 218826
rect 598848 218612 598900 218618
rect 598848 218554 598900 218560
rect 598860 217326 598888 218554
rect 598664 217320 598716 217326
rect 598664 217262 598716 217268
rect 598848 217320 598900 217326
rect 598848 217262 598900 217268
rect 598676 216918 598704 217262
rect 599032 217184 599084 217190
rect 599032 217126 599084 217132
rect 598664 216912 598716 216918
rect 598664 216854 598716 216860
rect 598478 215928 598534 215937
rect 598478 215863 598534 215872
rect 598492 210202 598520 215863
rect 599044 210202 599072 217126
rect 599504 210202 599532 221439
rect 601700 221264 601752 221270
rect 601700 221206 601752 221212
rect 601148 221128 601200 221134
rect 601148 221070 601200 221076
rect 600320 220992 600372 220998
rect 600320 220934 600372 220940
rect 600332 219434 600360 220934
rect 600504 220856 600556 220862
rect 600504 220798 600556 220804
rect 600332 219406 600452 219434
rect 600424 212534 600452 219406
rect 600332 212506 600452 212534
rect 600332 211070 600360 212506
rect 600320 211064 600372 211070
rect 600320 211006 600372 211012
rect 600516 210746 600544 220798
rect 600780 217184 600832 217190
rect 600780 217126 600832 217132
rect 600792 216918 600820 217126
rect 600780 216912 600832 216918
rect 600780 216854 600832 216860
rect 600688 211064 600740 211070
rect 600688 211006 600740 211012
rect 600516 210718 600636 210746
rect 600608 210202 600636 210718
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600636 210202
rect 600700 210202 600728 211006
rect 601160 210202 601188 221070
rect 601332 217320 601384 217326
rect 601332 217262 601384 217268
rect 601344 216782 601372 217262
rect 601332 216776 601384 216782
rect 601332 216718 601384 216724
rect 601712 210202 601740 221206
rect 601884 219020 601936 219026
rect 601884 218962 601936 218968
rect 601896 217462 601924 218962
rect 602896 217728 602948 217734
rect 602896 217670 602948 217676
rect 601884 217456 601936 217462
rect 601884 217398 601936 217404
rect 602908 217326 602936 217670
rect 602344 217320 602396 217326
rect 602344 217262 602396 217268
rect 602896 217320 602948 217326
rect 602896 217262 602948 217268
rect 602356 210202 602384 217262
rect 603092 210202 603120 221954
rect 606116 221876 606168 221882
rect 606116 221818 606168 221824
rect 605932 221604 605984 221610
rect 605932 221546 605984 221552
rect 605012 221400 605064 221406
rect 605012 221342 605064 221348
rect 604460 218476 604512 218482
rect 604460 218418 604512 218424
rect 603262 218376 603318 218385
rect 603262 218311 603318 218320
rect 603276 217870 603304 218311
rect 603264 217864 603316 217870
rect 603264 217806 603316 217812
rect 604472 217734 604500 218418
rect 603448 217728 603500 217734
rect 603448 217670 603500 217676
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 603460 210202 603488 217670
rect 604000 217320 604052 217326
rect 604000 217262 604052 217268
rect 604012 210202 604040 217262
rect 604552 217184 604604 217190
rect 604552 217126 604604 217132
rect 604564 210202 604592 217126
rect 605024 210202 605052 221342
rect 605944 214470 605972 221546
rect 605932 214464 605984 214470
rect 605932 214406 605984 214412
rect 606128 210202 606156 221818
rect 609428 221740 609480 221746
rect 609428 221682 609480 221688
rect 607312 220516 607364 220522
rect 607312 220458 607364 220464
rect 606760 217592 606812 217598
rect 606760 217534 606812 217540
rect 606300 214464 606352 214470
rect 606300 214406 606352 214412
rect 600700 210174 601036 210202
rect 601160 210174 601588 210202
rect 601712 210174 602140 210202
rect 602356 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605024 210174 605452 210202
rect 606004 210174 606156 210202
rect 606312 210202 606340 214406
rect 606772 210202 606800 217534
rect 607324 214470 607352 220458
rect 608600 219768 608652 219774
rect 608600 219710 608652 219716
rect 607496 219496 607548 219502
rect 607496 219438 607548 219444
rect 607312 214464 607364 214470
rect 607312 214406 607364 214412
rect 607508 210202 607536 219438
rect 607864 214464 607916 214470
rect 607864 214406 607916 214412
rect 607876 210202 607904 214406
rect 608612 210202 608640 219710
rect 608968 217048 609020 217054
rect 608968 216990 609020 216996
rect 608980 210202 609008 216990
rect 609440 210202 609468 221682
rect 611452 220652 611504 220658
rect 611452 220594 611504 220600
rect 610532 220380 610584 220386
rect 610532 220322 610584 220328
rect 610072 220244 610124 220250
rect 610072 220186 610124 220192
rect 609888 218204 609940 218210
rect 609888 218146 609940 218152
rect 609900 217054 609928 218146
rect 609888 217048 609940 217054
rect 609888 216990 609940 216996
rect 610084 210202 610112 220186
rect 610544 210202 610572 220322
rect 611464 210202 611492 220594
rect 611634 219736 611690 219745
rect 611634 219671 611690 219680
rect 611648 210202 611676 219671
rect 614488 218340 614540 218346
rect 614488 218282 614540 218288
rect 613384 217864 613436 217870
rect 613384 217806 613436 217812
rect 612280 216912 612332 216918
rect 612280 216854 612332 216860
rect 612292 210202 612320 216854
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 217806
rect 614120 217048 614172 217054
rect 614120 216990 614172 216996
rect 614132 210202 614160 216990
rect 614500 210202 614528 218282
rect 614960 210202 614988 223450
rect 615684 218068 615736 218074
rect 615684 218010 615736 218016
rect 615696 210202 615724 218010
rect 616880 217728 616932 217734
rect 616880 217670 616932 217676
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616708 214470 616736 214678
rect 616696 214464 616748 214470
rect 616696 214406 616748 214412
rect 616144 213240 616196 213246
rect 616144 213182 616196 213188
rect 616156 210202 616184 213182
rect 616892 210202 616920 217670
rect 617076 214742 617104 224606
rect 619640 224256 619692 224262
rect 619640 224198 619692 224204
rect 618258 221232 618314 221241
rect 618258 221167 618314 221176
rect 617246 219464 617302 219473
rect 617246 219399 617302 219408
rect 617064 214736 617116 214742
rect 617064 214678 617116 214684
rect 617260 210202 617288 219399
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 221167
rect 618902 215384 618958 215393
rect 618902 215319 618958 215328
rect 618916 210202 618944 215319
rect 619652 210202 619680 224198
rect 620192 224188 620244 224194
rect 620192 224130 620244 224136
rect 620204 223922 620232 224130
rect 620192 223916 620244 223922
rect 620192 223858 620244 223864
rect 620008 219768 620060 219774
rect 620008 219710 620060 219716
rect 619824 219632 619876 219638
rect 619824 219574 619876 219580
rect 619836 214742 619864 219574
rect 619824 214736 619876 214742
rect 619824 214678 619876 214684
rect 620020 210202 620048 219710
rect 621032 214742 621060 224878
rect 626540 224392 626592 224398
rect 626540 224334 626592 224340
rect 625436 224188 625488 224194
rect 625436 224130 625488 224136
rect 625252 223916 625304 223922
rect 625252 223858 625304 223864
rect 622676 223780 622728 223786
rect 622676 223722 622728 223728
rect 622492 223644 622544 223650
rect 622492 223586 622544 223592
rect 621204 222488 621256 222494
rect 621204 222430 621256 222436
rect 620560 214736 620612 214742
rect 620560 214678 620612 214684
rect 621020 214736 621072 214742
rect 621020 214678 621072 214684
rect 620572 210202 620600 214678
rect 621216 210202 621244 222430
rect 622308 214872 622360 214878
rect 622308 214814 622360 214820
rect 621664 214736 621716 214742
rect 621664 214678 621716 214684
rect 621676 210202 621704 214678
rect 622320 214554 622348 214814
rect 622504 214742 622532 223586
rect 622492 214736 622544 214742
rect 622492 214678 622544 214684
rect 622320 214526 622532 214554
rect 622504 210202 622532 214526
rect 622688 210202 622716 223722
rect 623872 216776 623924 216782
rect 623872 216718 623924 216724
rect 623320 214736 623372 214742
rect 623320 214678 623372 214684
rect 623332 210202 623360 214678
rect 623884 210202 623912 216718
rect 625264 214742 625292 223858
rect 625252 214736 625304 214742
rect 625252 214678 625304 214684
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625448 210202 625476 224130
rect 626356 219156 626408 219162
rect 626356 219098 626408 219104
rect 626080 214736 626132 214742
rect 626080 214678 626132 214684
rect 625620 214600 625672 214606
rect 625620 214542 625672 214548
rect 606312 210174 606556 210202
rect 606772 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210174 608764 210202
rect 608980 210174 609316 210202
rect 609440 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611464 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 616892 210174 617044 210202
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621216 210174 621460 210202
rect 621676 210174 622012 210202
rect 622504 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625476 210202
rect 625632 210202 625660 214542
rect 626092 210202 626120 214678
rect 626368 214470 626396 219098
rect 626356 214464 626408 214470
rect 626356 214406 626408 214412
rect 626552 210202 626580 224334
rect 629852 222352 629904 222358
rect 629852 222294 629904 222300
rect 627092 222216 627144 222222
rect 627092 222158 627144 222164
rect 627104 210202 627132 222158
rect 627458 218104 627514 218113
rect 627458 218039 627514 218048
rect 627472 213994 627500 218039
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 627918 216200 627974 216209
rect 627918 216135 627974 216144
rect 627460 213988 627512 213994
rect 627460 213930 627512 213936
rect 627932 210202 627960 216135
rect 628300 210202 628328 217398
rect 628840 214464 628892 214470
rect 628840 214406 628892 214412
rect 628852 210202 628880 214406
rect 629392 213988 629444 213994
rect 629392 213930 629444 213936
rect 629404 210202 629432 213930
rect 629864 210202 629892 222294
rect 630048 214742 630076 229066
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 630680 222624 630732 222630
rect 630680 222566 630732 222572
rect 630036 214736 630088 214742
rect 630036 214678 630088 214684
rect 630692 212430 630720 222566
rect 631322 220960 631378 220969
rect 631322 220895 631378 220904
rect 631138 218376 631194 218385
rect 631138 218311 631194 218320
rect 630680 212424 630732 212430
rect 630680 212366 630732 212372
rect 631152 210202 631180 218311
rect 625632 210174 625876 210202
rect 626092 210174 626428 210202
rect 626552 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630844 210174 631180 210202
rect 631336 210202 631364 220895
rect 632716 212566 632744 222838
rect 633440 220108 633492 220114
rect 633440 220050 633492 220056
rect 633452 219434 633480 220050
rect 633452 219406 633572 219434
rect 632888 214736 632940 214742
rect 632888 214678 632940 214684
rect 632704 212560 632756 212566
rect 632704 212502 632756 212508
rect 631600 212424 631652 212430
rect 631600 212366 631652 212372
rect 631612 210202 631640 212366
rect 632900 210202 632928 214678
rect 633544 212534 633572 219406
rect 633452 212506 633572 212534
rect 633452 211070 633480 212506
rect 633440 211064 633492 211070
rect 633440 211006 633492 211012
rect 633636 210746 633664 231066
rect 634360 212560 634412 212566
rect 634360 212502 634412 212508
rect 633808 211064 633860 211070
rect 633808 211006 633860 211012
rect 633636 210718 633756 210746
rect 633728 210202 633756 210718
rect 631336 210174 631396 210202
rect 631612 210174 631948 210202
rect 632900 210174 633052 210202
rect 633604 210174 633756 210202
rect 633820 210202 633848 211006
rect 634372 210202 634400 212502
rect 636856 210202 636884 231066
rect 639616 229094 639644 232494
rect 650656 231130 650684 256663
rect 650644 231124 650696 231130
rect 650644 231066 650696 231072
rect 639616 229066 639828 229094
rect 639800 210338 639828 229066
rect 652036 227050 652064 288487
rect 652220 233918 652248 291479
rect 652404 283529 652432 295287
rect 652390 283520 652446 283529
rect 652390 283455 652446 283464
rect 652390 282160 652446 282169
rect 652390 282095 652446 282104
rect 652208 233912 652260 233918
rect 652208 233854 652260 233860
rect 652024 227044 652076 227050
rect 652024 226986 652076 226992
rect 652404 226953 652432 282095
rect 652574 280392 652630 280401
rect 652574 280327 652630 280336
rect 652588 229809 652616 280327
rect 654796 232558 654824 300863
rect 656164 297084 656216 297090
rect 656164 297026 656216 297032
rect 656176 271153 656204 297026
rect 656162 271144 656218 271153
rect 656162 271079 656218 271088
rect 654784 232552 654836 232558
rect 654784 232494 654836 232500
rect 652574 229800 652630 229809
rect 652574 229735 652630 229744
rect 652390 226944 652446 226953
rect 652390 226879 652446 226888
rect 654782 226400 654838 226409
rect 654782 226335 654838 226344
rect 652022 225584 652078 225593
rect 652022 225519 652078 225528
rect 651288 224256 651340 224262
rect 651288 224198 651340 224204
rect 650642 222864 650698 222873
rect 650642 222799 650698 222808
rect 649722 221504 649778 221513
rect 649722 221439 649778 221448
rect 644754 220416 644810 220425
rect 644754 220351 644810 220360
rect 642180 217320 642232 217326
rect 642180 217262 642232 217268
rect 638972 210310 639828 210338
rect 638972 210202 639000 210310
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210186 635596 210202
rect 636580 210186 636916 210202
rect 635260 210180 635608 210186
rect 635260 210174 635556 210180
rect 635556 210122 635608 210128
rect 636568 210180 636916 210186
rect 636620 210174 636916 210180
rect 638572 210174 639000 210202
rect 639800 210202 639828 210310
rect 642192 210202 642220 217262
rect 644572 214736 644624 214742
rect 644572 214678 644624 214684
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 643848 210202 643876 213182
rect 639800 210174 640228 210202
rect 641884 210174 642220 210202
rect 643540 210174 643876 210202
rect 644584 210202 644612 214678
rect 644768 210202 644796 220351
rect 648526 218648 648582 218657
rect 648526 218583 648582 218592
rect 646596 218068 646648 218074
rect 646596 218010 646648 218016
rect 646608 210202 646636 218010
rect 648252 216640 648304 216646
rect 648252 216582 648304 216588
rect 647148 213648 647200 213654
rect 647148 213590 647200 213596
rect 647160 210202 647188 213590
rect 648264 210202 648292 216582
rect 648540 210202 648568 218583
rect 649736 213654 649764 221439
rect 649908 213920 649960 213926
rect 649908 213862 649960 213868
rect 649724 213648 649776 213654
rect 649724 213590 649776 213596
rect 649920 210202 649948 213862
rect 650656 213246 650684 222799
rect 651104 213376 651156 213382
rect 651104 213318 651156 213324
rect 650644 213240 650696 213246
rect 650644 213182 650696 213188
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 644584 210174 644644 210202
rect 644768 210174 645196 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647956 210174 648292 210202
rect 648508 210174 648568 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 213318
rect 651300 212770 651328 224198
rect 651470 221776 651526 221785
rect 651470 221711 651526 221720
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 651484 210202 651512 221711
rect 652036 213926 652064 225519
rect 653402 225040 653458 225049
rect 653402 224975 653458 224984
rect 653034 220144 653090 220153
rect 653034 220079 653090 220088
rect 652850 215928 652906 215937
rect 652850 215863 652906 215872
rect 652024 213920 652076 213926
rect 652024 213862 652076 213868
rect 652864 210202 652892 215863
rect 653048 210202 653076 220079
rect 653416 218074 653444 224975
rect 653404 218068 653456 218074
rect 653404 218010 653456 218016
rect 654796 214742 654824 226335
rect 656162 225312 656218 225321
rect 656162 225247 656218 225256
rect 655426 218920 655482 218929
rect 655426 218855 655482 218864
rect 654784 214736 654836 214742
rect 654784 214678 654836 214684
rect 654876 214600 654928 214606
rect 654876 214542 654928 214548
rect 654888 210202 654916 214542
rect 655440 210202 655468 218855
rect 656176 216646 656204 225247
rect 657542 223952 657598 223961
rect 657542 223887 657598 223896
rect 656806 217288 656862 217297
rect 656806 217223 656862 217232
rect 656164 216640 656216 216646
rect 656164 216582 656216 216588
rect 656530 212936 656586 212945
rect 656530 212871 656586 212880
rect 656544 210202 656572 212871
rect 656820 210202 656848 217223
rect 657556 213382 657584 223887
rect 658936 217326 658964 346423
rect 664442 312080 664498 312089
rect 664442 312015 664498 312024
rect 664456 300830 664484 312015
rect 664444 300824 664496 300830
rect 664444 300766 664496 300772
rect 662420 298172 662472 298178
rect 662420 298114 662472 298120
rect 662432 293865 662460 298114
rect 665824 295996 665876 296002
rect 665824 295938 665876 295944
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 662418 293856 662474 293865
rect 662418 293791 662474 293800
rect 663064 292596 663116 292602
rect 663064 292538 663116 292544
rect 660304 289876 660356 289882
rect 660304 289818 660356 289824
rect 660316 232558 660344 289818
rect 661684 288448 661736 288454
rect 661684 288390 661736 288396
rect 661696 234666 661724 288390
rect 661684 234660 661736 234666
rect 661684 234602 661736 234608
rect 660304 232552 660356 232558
rect 660304 232494 660356 232500
rect 663076 231538 663104 292538
rect 664456 248169 664484 293966
rect 665836 268569 665864 295938
rect 667754 295760 667810 295769
rect 667754 295695 667810 295704
rect 667768 293865 667796 295695
rect 667754 293856 667810 293865
rect 667754 293791 667810 293800
rect 667204 282940 667256 282946
rect 667204 282882 667256 282888
rect 665822 268560 665878 268569
rect 665822 268495 665878 268504
rect 664442 248160 664498 248169
rect 664442 248095 664498 248104
rect 665456 231668 665508 231674
rect 665456 231610 665508 231616
rect 663064 231532 663116 231538
rect 663064 231474 663116 231480
rect 662328 231396 662380 231402
rect 662328 231338 662380 231344
rect 660948 229152 661000 229158
rect 660948 229094 661000 229100
rect 660488 227792 660540 227798
rect 660488 227734 660540 227740
rect 659106 222592 659162 222601
rect 659106 222527 659162 222536
rect 658924 217320 658976 217326
rect 658924 217262 658976 217268
rect 658738 214568 658794 214577
rect 658738 214503 658794 214512
rect 657544 213376 657596 213382
rect 657544 213318 657596 213324
rect 658188 212764 658240 212770
rect 658188 212706 658240 212712
rect 658200 210202 658228 212706
rect 658752 210202 658780 214503
rect 659120 212770 659148 222527
rect 659568 213716 659620 213722
rect 659568 213658 659620 213664
rect 659108 212764 659160 212770
rect 659108 212706 659160 212712
rect 659580 210202 659608 213658
rect 660500 210202 660528 227734
rect 660960 210202 660988 229094
rect 662340 219434 662368 231338
rect 664996 231192 665048 231198
rect 664996 231134 665048 231140
rect 663706 229120 663762 229129
rect 665008 229094 665036 231134
rect 665178 229528 665234 229537
rect 665178 229463 665234 229472
rect 665192 229094 665220 229463
rect 665468 229158 665496 231610
rect 665822 230480 665878 230489
rect 665822 230415 665878 230424
rect 665456 229152 665508 229158
rect 665456 229094 665508 229100
rect 665008 229066 665128 229094
rect 665192 229066 665312 229094
rect 663706 229055 663762 229064
rect 663524 228404 663576 228410
rect 663524 228346 663576 228352
rect 662248 219406 662368 219434
rect 662050 217560 662106 217569
rect 662050 217495 662106 217504
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 217495
rect 651116 210174 651268 210202
rect 651484 210174 651820 210202
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654580 210174 654916 210202
rect 655132 210174 655468 210202
rect 656236 210174 656572 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660528 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662248 210202 662276 219406
rect 663156 215348 663208 215354
rect 663156 215290 663208 215296
rect 663168 210202 663196 215290
rect 663536 210202 663564 228346
rect 663720 215354 663748 229055
rect 664442 223680 664498 223689
rect 664442 223615 664498 223624
rect 663708 215348 663760 215354
rect 663708 215290 663760 215296
rect 664456 214606 664484 223615
rect 664444 214600 664496 214606
rect 664444 214542 664496 214548
rect 664812 214396 664864 214402
rect 664812 214338 664864 214344
rect 664260 212764 664312 212770
rect 664260 212706 664312 212712
rect 664272 210202 664300 212706
rect 664824 210202 664852 214338
rect 665100 212770 665128 229066
rect 665284 227798 665312 229066
rect 665272 227792 665324 227798
rect 665272 227734 665324 227740
rect 665546 216200 665602 216209
rect 665546 216135 665602 216144
rect 665560 213722 665588 216135
rect 665836 214402 665864 230415
rect 666468 225072 666520 225078
rect 666468 225014 666520 225020
rect 666480 224262 666508 225014
rect 666468 224256 666520 224262
rect 666468 224198 666520 224204
rect 667018 221096 667074 221105
rect 667018 221031 667074 221040
rect 665824 214396 665876 214402
rect 665824 214338 665876 214344
rect 665548 213716 665600 213722
rect 665548 213658 665600 213664
rect 665088 212764 665140 212770
rect 665088 212706 665140 212712
rect 662248 210174 662308 210202
rect 662860 210174 663196 210202
rect 663412 210174 663564 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 636568 210122 636620 210128
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 579068 124908 579120 124914
rect 579068 124850 579120 124856
rect 578700 124160 578752 124166
rect 578700 124102 578752 124108
rect 578712 123593 578740 124102
rect 578698 123584 578754 123593
rect 578698 123519 578754 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118584 578568 118590
rect 578516 118526 578568 118532
rect 578528 118425 578556 118526
rect 578514 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108996 578384 109002
rect 578332 108938 578384 108944
rect 578344 108361 578372 108938
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 579080 105913 579108 124850
rect 580276 118590 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580264 118584 580316 118590
rect 580264 118526 580316 118532
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110288 579396 110294
rect 579344 110230 579396 110236
rect 579356 110129 579384 110230
rect 579342 110120 579398 110129
rect 579342 110055 579398 110064
rect 580448 109132 580500 109138
rect 580448 109074 580500 109080
rect 580264 106344 580316 106350
rect 580264 106286 580316 106292
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 579344 105664 579396 105670
rect 579344 105606 579396 105612
rect 578516 103420 578568 103426
rect 578516 103362 578568 103368
rect 578528 103193 578556 103362
rect 578514 103184 578570 103193
rect 578514 103119 578570 103128
rect 579160 102128 579212 102134
rect 579160 102070 579212 102076
rect 579172 101697 579200 102070
rect 579158 101688 579214 101697
rect 579158 101623 579214 101632
rect 578608 100020 578660 100026
rect 578608 99962 578660 99968
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578620 97481 578648 99962
rect 578606 97472 578662 97481
rect 578606 97407 578662 97416
rect 578332 95192 578384 95198
rect 578332 95134 578384 95140
rect 578344 95033 578372 95134
rect 578330 95024 578386 95033
rect 578330 94959 578386 94968
rect 579356 93854 579384 105606
rect 579528 99272 579580 99278
rect 579526 99240 579528 99249
rect 579580 99240 579582 99249
rect 579526 99175 579582 99184
rect 579356 93826 579476 93854
rect 579252 93424 579304 93430
rect 579252 93366 579304 93372
rect 579264 93129 579292 93366
rect 579250 93120 579306 93129
rect 579250 93055 579306 93064
rect 577504 91792 577556 91798
rect 577504 91734 577556 91740
rect 576124 58676 576176 58682
rect 576124 58618 576176 58624
rect 574284 56024 574336 56030
rect 574284 55966 574336 55972
rect 460754 53680 460810 53689
rect 460388 53644 460440 53650
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 462594 53680 462650 53689
rect 461674 53615 461730 53624
rect 461952 53644 462004 53650
rect 460388 53586 460440 53592
rect 459468 53508 459520 53514
rect 459468 53450 459520 53456
rect 130384 53372 130436 53378
rect 130384 53314 130436 53320
rect 129188 53236 129240 53242
rect 129188 53178 129240 53184
rect 129004 53100 129056 53106
rect 129004 53042 129056 53048
rect 129016 51074 129044 53042
rect 128832 51046 129044 51074
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 45468 49020 45520 49026
rect 45468 48962 45520 48968
rect 43812 45212 43864 45218
rect 43812 45154 43864 45160
rect 126428 44940 126480 44946
rect 126428 44882 126480 44888
rect 43628 44328 43680 44334
rect 43628 44270 43680 44276
rect 126440 44198 126468 44882
rect 128832 44402 128860 51046
rect 129004 49020 129056 49026
rect 129004 48962 129056 48968
rect 129016 46102 129044 48962
rect 129004 46096 129056 46102
rect 129004 46038 129056 46044
rect 129200 44810 129228 53178
rect 129372 51876 129424 51882
rect 129372 51818 129424 51824
rect 129384 45082 129412 51818
rect 129648 49156 129700 49162
rect 129648 49098 129700 49104
rect 129660 45422 129688 49098
rect 129648 45416 129700 45422
rect 129648 45358 129700 45364
rect 129372 45076 129424 45082
rect 129372 45018 129424 45024
rect 129188 44804 129240 44810
rect 129188 44746 129240 44752
rect 128820 44396 128872 44402
rect 128820 44338 128872 44344
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 126428 44192 126480 44198
rect 126428 44134 126480 44140
rect 130396 44062 130424 53314
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 306024 51746 306052 53108
rect 130568 51740 130620 51746
rect 130568 51682 130620 51688
rect 145380 51740 145432 51746
rect 145380 51682 145432 51688
rect 306012 51740 306064 51746
rect 306012 51682 306064 51688
rect 130580 45966 130608 51682
rect 145392 50810 145420 51682
rect 145084 50782 145420 50810
rect 131028 50380 131080 50386
rect 131028 50322 131080 50328
rect 130568 45960 130620 45966
rect 130568 45902 130620 45908
rect 131040 45370 131068 50322
rect 308048 50289 308076 53108
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53450
rect 459606 52828 459658 52834
rect 459606 52770 459658 52776
rect 459172 52550 459508 52578
rect 459618 52564 459646 52770
rect 460400 52578 460428 53586
rect 460768 52578 460796 53615
rect 461308 53372 461360 53378
rect 461308 53314 461360 53320
rect 461320 52578 461348 53314
rect 461688 52578 461716 53615
rect 461952 53586 462004 53592
rect 462228 53644 462280 53650
rect 462594 53615 462650 53624
rect 463146 53680 463202 53689
rect 473910 53680 473966 53689
rect 463146 53615 463202 53624
rect 464896 53644 464948 53650
rect 462228 53586 462280 53592
rect 461964 53145 461992 53586
rect 461950 53136 462006 53145
rect 461950 53071 462006 53080
rect 462240 52578 462268 53586
rect 462608 52578 462636 53615
rect 463160 52578 463188 53615
rect 464896 53586 464948 53592
rect 465080 53644 465132 53650
rect 465080 53586 465132 53592
rect 465540 53644 465592 53650
rect 465540 53586 465592 53592
rect 465724 53644 465776 53650
rect 465724 53586 465776 53592
rect 469956 53644 470008 53650
rect 469956 53586 470008 53592
rect 472808 53644 472860 53650
rect 564530 53680 564586 53689
rect 473910 53615 473912 53624
rect 472808 53586 472860 53592
rect 473964 53615 473966 53624
rect 476672 53644 476724 53650
rect 473912 53586 473964 53592
rect 476672 53586 476724 53592
rect 478144 53644 478196 53650
rect 564530 53615 564532 53624
rect 478144 53586 478196 53592
rect 564584 53615 564586 53624
rect 564532 53586 564584 53592
rect 464528 53236 464580 53242
rect 464528 53178 464580 53184
rect 463608 52964 463660 52970
rect 463608 52906 463660 52912
rect 463620 52578 463648 52906
rect 463746 52828 463798 52834
rect 463746 52770 463798 52776
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463648 52578
rect 463758 52564 463786 52770
rect 464540 52578 464568 53178
rect 464908 52578 464936 53586
rect 465092 52834 465120 53586
rect 465552 53242 465580 53586
rect 465540 53236 465592 53242
rect 465540 53178 465592 53184
rect 465736 52970 465764 53586
rect 465908 53236 465960 53242
rect 465908 53178 465960 53184
rect 465724 52964 465776 52970
rect 465724 52906 465776 52912
rect 465080 52828 465132 52834
rect 465080 52770 465132 52776
rect 465448 52828 465500 52834
rect 465448 52770 465500 52776
rect 465460 52578 465488 52770
rect 465920 52578 465948 53178
rect 469968 52834 469996 53586
rect 472820 53145 472848 53586
rect 472806 53136 472862 53145
rect 476684 53106 476712 53586
rect 478156 53242 478184 53586
rect 574296 53310 574324 55966
rect 576136 55049 576164 58618
rect 577320 57248 577372 57254
rect 577320 57190 577372 57196
rect 577136 55888 577188 55894
rect 577136 55830 577188 55836
rect 576122 55040 576178 55049
rect 576122 54975 576178 54984
rect 574744 53984 574796 53990
rect 574744 53926 574796 53932
rect 574756 53689 574784 53926
rect 574742 53680 574798 53689
rect 574742 53615 574798 53624
rect 577148 53514 577176 55830
rect 577332 55622 577360 57190
rect 577320 55616 577372 55622
rect 577320 55558 577372 55564
rect 577516 54194 577544 91734
rect 578700 91452 578752 91458
rect 578700 91394 578752 91400
rect 578712 90953 578740 91394
rect 578698 90944 578754 90953
rect 578698 90879 578754 90888
rect 579252 88324 579304 88330
rect 579252 88266 579304 88272
rect 579264 88097 579292 88266
rect 579250 88088 579306 88097
rect 579250 88023 579306 88032
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 579252 84040 579304 84046
rect 579250 84008 579252 84017
rect 579304 84008 579306 84017
rect 579250 83943 579306 83952
rect 578700 82816 578752 82822
rect 578700 82758 578752 82764
rect 578712 82249 578740 82758
rect 578698 82240 578754 82249
rect 578698 82175 578754 82184
rect 579068 82136 579120 82142
rect 579068 82078 579120 82084
rect 578516 78464 578568 78470
rect 578516 78406 578568 78412
rect 578528 77897 578556 78406
rect 578514 77888 578570 77897
rect 578514 77823 578570 77832
rect 579080 75721 579108 82078
rect 579448 80073 579476 93826
rect 579434 80064 579490 80073
rect 579434 79999 579490 80008
rect 580276 78470 580304 106286
rect 580460 86970 580488 109074
rect 580644 109002 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 632152 209568 632204 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 667032 176497 667060 221031
rect 667018 176488 667074 176497
rect 667018 176423 667074 176432
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108996 580684 109002
rect 580632 108938 580684 108944
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 581656 84046 581684 110434
rect 581840 110294 581868 131242
rect 583036 124166 583064 139402
rect 584784 137358 584812 144910
rect 585784 143608 585836 143614
rect 585784 143550 585836 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583392 129192 583444 129198
rect 583392 129134 583444 129140
rect 583024 124160 583076 124166
rect 583024 124102 583076 124108
rect 583208 120760 583260 120766
rect 583208 120702 583260 120708
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110288 581880 110294
rect 581828 110230 581880 110236
rect 582288 107704 582340 107710
rect 582288 107646 582340 107652
rect 582300 105670 582328 107646
rect 582288 105664 582340 105670
rect 582288 105606 582340 105612
rect 581644 84040 581696 84046
rect 581644 83982 581696 83988
rect 583036 82822 583064 113154
rect 583220 99278 583248 120702
rect 583404 116958 583432 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583392 116952 583444 116958
rect 583392 116894 583444 116900
rect 584416 102134 584444 122810
rect 584600 122194 584628 136614
rect 585796 131170 585824 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 132524 586020 132530
rect 585968 132466 586020 132472
rect 585784 131164 585836 131170
rect 585784 131106 585836 131112
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585784 116000 585836 116006
rect 585784 115942 585836 115948
rect 584588 115252 584640 115258
rect 584588 115194 584640 115200
rect 584404 102128 584456 102134
rect 584404 102070 584456 102076
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 99272 583260 99278
rect 583208 99214 583260 99220
rect 583024 82816 583076 82822
rect 583024 82758 583076 82764
rect 583024 79348 583076 79354
rect 583024 79290 583076 79296
rect 580264 78464 580316 78470
rect 580264 78406 580316 78412
rect 580446 77888 580502 77897
rect 580446 77823 580502 77832
rect 579066 75712 579122 75721
rect 579066 75647 579122 75656
rect 578884 75200 578936 75206
rect 578884 75142 578936 75148
rect 578516 71596 578568 71602
rect 578516 71538 578568 71544
rect 578528 71233 578556 71538
rect 578514 71224 578570 71233
rect 578514 71159 578570 71168
rect 578896 60489 578924 75142
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579528 66904 579580 66910
rect 579526 66872 579528 66881
rect 579580 66872 579582 66881
rect 579526 66807 579582 66816
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 579528 62076 579580 62082
rect 579528 62018 579580 62024
rect 579540 61849 579568 62018
rect 579526 61840 579582 61849
rect 579526 61775 579582 61784
rect 578882 60480 578938 60489
rect 578882 60415 578938 60424
rect 578332 60036 578384 60042
rect 578332 59978 578384 59984
rect 577688 58812 577740 58818
rect 577688 58754 577740 58760
rect 577700 54777 577728 58754
rect 578344 56137 578372 59978
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 578330 56128 578386 56137
rect 578330 56063 578386 56072
rect 577686 54768 577742 54777
rect 577686 54703 577742 54712
rect 580460 54670 580488 77823
rect 580448 54664 580500 54670
rect 580448 54606 580500 54612
rect 583036 54398 583064 79290
rect 584416 71602 584444 100098
rect 584600 95198 584628 115194
rect 584588 95192 584640 95198
rect 584588 95134 584640 95140
rect 585796 91458 585824 115942
rect 585980 112878 586008 132466
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588726 129704 588782 129713
rect 588726 129639 588782 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587808 127016 587860 127022
rect 587808 126958 587860 126964
rect 587820 124914 587848 126958
rect 587808 124908 587860 124914
rect 587808 124850 587860 124856
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585968 112872 586020 112878
rect 585968 112814 586020 112820
rect 586152 112464 586204 112470
rect 586152 112406 586204 112412
rect 586164 93430 586192 112406
rect 587164 104916 587216 104922
rect 587164 104858 587216 104864
rect 586152 93424 586204 93430
rect 586152 93366 586204 93372
rect 585784 91452 585836 91458
rect 585784 91394 585836 91400
rect 587176 82142 587204 104858
rect 587360 100026 587388 121450
rect 588542 103592 588598 103601
rect 588542 103527 588598 103536
rect 587348 100020 587400 100026
rect 587348 99962 587400 99968
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 587164 76560 587216 76566
rect 587164 76502 587216 76508
rect 584404 71596 584456 71602
rect 584404 71538 584456 71544
rect 587176 62082 587204 76502
rect 588556 73166 588584 103527
rect 588740 103426 588768 129639
rect 590396 129198 590424 134535
rect 667216 133249 667244 282882
rect 667388 280220 667440 280226
rect 667388 280162 667440 280168
rect 667400 134609 667428 280162
rect 668768 237448 668820 237454
rect 668768 237390 668820 237396
rect 668216 234932 668268 234938
rect 668216 234874 668268 234880
rect 668032 224256 668084 224262
rect 668032 224198 668084 224204
rect 667848 224120 667900 224126
rect 667848 224062 667900 224068
rect 667860 223689 667888 224062
rect 667846 223680 667902 223689
rect 667846 223615 667902 223624
rect 667570 222048 667626 222057
rect 667570 221983 667626 221992
rect 667584 177313 667612 221983
rect 668044 220153 668072 224198
rect 668030 220144 668086 220153
rect 668030 220079 668086 220088
rect 667754 219464 667810 219473
rect 667754 219399 667810 219408
rect 667570 177304 667626 177313
rect 667570 177239 667626 177248
rect 667768 175001 667796 219399
rect 668030 207632 668086 207641
rect 668030 207567 668086 207576
rect 668044 204105 668072 207567
rect 668030 204096 668086 204105
rect 668030 204031 668086 204040
rect 668044 200114 668072 204031
rect 667952 200086 668072 200114
rect 667952 199209 667980 200086
rect 667938 199200 667994 199209
rect 667938 199135 667994 199144
rect 667938 194168 667994 194177
rect 667938 194103 667994 194112
rect 667952 189689 667980 194103
rect 667938 189680 667994 189689
rect 667938 189615 667994 189624
rect 668030 184376 668086 184385
rect 668030 184311 668086 184320
rect 668044 179489 668072 184311
rect 668030 179480 668086 179489
rect 668030 179415 668086 179424
rect 667754 174992 667810 175001
rect 667754 174927 667810 174936
rect 667386 134600 667442 134609
rect 667386 134535 667442 134544
rect 667202 133240 667258 133249
rect 667202 133175 667258 133184
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589922 126440 589978 126449
rect 589922 126375 589978 126384
rect 589370 124808 589426 124817
rect 589370 124743 589426 124752
rect 589384 120766 589412 124743
rect 589554 123176 589610 123185
rect 589554 123111 589610 123120
rect 589568 122874 589596 123111
rect 589556 122868 589608 122874
rect 589556 122810 589608 122816
rect 589936 122058 589964 126375
rect 668044 125361 668072 179415
rect 668228 173097 668256 234874
rect 668400 234524 668452 234530
rect 668400 234466 668452 234472
rect 668214 173088 668270 173097
rect 668214 173023 668270 173032
rect 668412 169697 668440 234466
rect 668584 227180 668636 227186
rect 668584 227122 668636 227128
rect 668596 224210 668624 227122
rect 668596 224182 668716 224210
rect 668398 169688 668454 169697
rect 668398 169623 668454 169632
rect 668216 165232 668268 165238
rect 668216 165174 668268 165180
rect 668228 164937 668256 165174
rect 668214 164928 668270 164937
rect 668214 164863 668270 164872
rect 668216 163328 668268 163334
rect 668214 163296 668216 163305
rect 668268 163296 668270 163305
rect 668214 163231 668270 163240
rect 668688 161474 668716 224182
rect 668596 161446 668716 161474
rect 668216 160064 668268 160070
rect 668214 160032 668216 160041
rect 668268 160032 668270 160041
rect 668214 159967 668270 159976
rect 668596 158409 668624 161446
rect 668582 158400 668638 158409
rect 668582 158335 668638 158344
rect 668308 155168 668360 155174
rect 668306 155136 668308 155145
rect 668360 155136 668362 155145
rect 668306 155071 668362 155080
rect 668216 148776 668268 148782
rect 668216 148718 668268 148724
rect 668228 148617 668256 148718
rect 668214 148608 668270 148617
rect 668214 148543 668270 148552
rect 668216 136264 668268 136270
rect 668216 136206 668268 136212
rect 668228 135561 668256 136206
rect 668214 135552 668270 135561
rect 668214 135487 668270 135496
rect 668780 130665 668808 237390
rect 669044 227792 669096 227798
rect 669044 227734 669096 227740
rect 669056 219434 669084 227734
rect 668964 219406 669084 219434
rect 668964 138825 668992 219406
rect 669240 143721 669268 393751
rect 670606 392592 670662 392601
rect 670606 392527 670662 392536
rect 669962 345672 670018 345681
rect 669962 345607 670018 345616
rect 669596 235340 669648 235346
rect 669596 235282 669648 235288
rect 669412 232960 669464 232966
rect 669412 232902 669464 232908
rect 669424 174729 669452 232902
rect 669410 174720 669466 174729
rect 669410 174655 669466 174664
rect 669410 172000 669466 172009
rect 669410 171935 669466 171944
rect 669424 149025 669452 171935
rect 669608 165238 669636 235282
rect 669778 234424 669834 234433
rect 669778 234359 669834 234368
rect 669596 165232 669648 165238
rect 669596 165174 669648 165180
rect 669792 163334 669820 234359
rect 669780 163328 669832 163334
rect 669780 163270 669832 163276
rect 669410 149016 669466 149025
rect 669410 148951 669466 148960
rect 669226 143712 669282 143721
rect 669226 143647 669282 143656
rect 668950 138816 669006 138825
rect 668950 138751 669006 138760
rect 669976 136270 670004 345607
rect 670422 261352 670478 261361
rect 670422 261287 670478 261296
rect 670238 259720 670294 259729
rect 670238 259655 670294 259664
rect 670252 245721 670280 259655
rect 670436 247081 670464 261287
rect 670422 247072 670478 247081
rect 670422 247007 670478 247016
rect 670238 245712 670294 245721
rect 670238 245647 670294 245656
rect 670148 235952 670200 235958
rect 670148 235894 670200 235900
rect 670160 148782 670188 235894
rect 670332 233096 670384 233102
rect 670332 233038 670384 233044
rect 670344 160070 670372 233038
rect 670620 224954 670648 392527
rect 672000 372609 672028 397151
rect 672722 394768 672778 394777
rect 672722 394703 672778 394712
rect 672736 381041 672764 394703
rect 672722 381032 672778 381041
rect 672722 380967 672778 380976
rect 671986 372600 672042 372609
rect 671986 372535 672042 372544
rect 672538 357096 672594 357105
rect 672538 357031 672594 357040
rect 672354 351384 672410 351393
rect 672354 351319 672410 351328
rect 671986 350160 672042 350169
rect 671986 350095 672042 350104
rect 672000 332353 672028 350095
rect 672368 337249 672396 351319
rect 672354 337240 672410 337249
rect 672354 337175 672410 337184
rect 671986 332344 672042 332353
rect 671986 332279 672042 332288
rect 672552 312497 672580 357031
rect 672920 356833 672948 401231
rect 673196 357513 673224 402047
rect 673366 400616 673422 400625
rect 673366 400551 673422 400560
rect 673182 357504 673238 357513
rect 673182 357439 673238 357448
rect 672906 356824 672962 356833
rect 672906 356759 672962 356768
rect 672722 356280 672778 356289
rect 672722 356215 672778 356224
rect 672538 312488 672594 312497
rect 672538 312423 672594 312432
rect 672736 311894 672764 356215
rect 673380 355881 673408 400551
rect 673918 399800 673974 399809
rect 673918 399735 673974 399744
rect 673734 394088 673790 394097
rect 673734 394023 673790 394032
rect 673748 376689 673776 394023
rect 673734 376680 673790 376689
rect 673734 376615 673790 376624
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673182 355464 673238 355473
rect 673182 355399 673238 355408
rect 672906 348528 672962 348537
rect 672906 348463 672962 348472
rect 672552 311866 672764 311894
rect 672552 311681 672580 311866
rect 672538 311672 672594 311681
rect 672538 311607 672594 311616
rect 672722 311264 672778 311273
rect 672722 311199 672778 311208
rect 672736 310593 672764 311199
rect 672722 310584 672778 310593
rect 672722 310519 672778 310528
rect 672262 305552 672318 305561
rect 672262 305487 672318 305496
rect 672078 304328 672134 304337
rect 672078 304263 672134 304272
rect 671526 302288 671582 302297
rect 671526 302223 671582 302232
rect 671540 263594 671568 302223
rect 672092 287881 672120 304263
rect 672078 287872 672134 287881
rect 672078 287807 672134 287816
rect 672080 285728 672132 285734
rect 672080 285670 672132 285676
rect 672092 281602 672120 285670
rect 672276 285569 672304 305487
rect 672448 287088 672500 287094
rect 672448 287030 672500 287036
rect 672262 285560 672318 285569
rect 672262 285495 672318 285504
rect 672460 282914 672488 287030
rect 672632 284368 672684 284374
rect 672632 284310 672684 284316
rect 672644 282914 672672 284310
rect 672460 282886 672580 282914
rect 672644 282886 672764 282914
rect 672092 281574 672488 281602
rect 671540 263566 671660 263594
rect 671158 262168 671214 262177
rect 671158 262103 671214 262112
rect 670974 250880 671030 250889
rect 670974 250815 671030 250824
rect 670988 248169 671016 250815
rect 670974 248160 671030 248169
rect 670974 248095 671030 248104
rect 670976 235816 671028 235822
rect 670976 235758 671028 235764
rect 670790 232520 670846 232529
rect 670790 232455 670792 232464
rect 670844 232455 670846 232464
rect 670792 232426 670844 232432
rect 670790 231568 670846 231577
rect 670790 231503 670792 231512
rect 670844 231503 670846 231512
rect 670792 231474 670844 231480
rect 670792 226568 670844 226574
rect 670792 226510 670844 226516
rect 670804 226409 670832 226510
rect 670790 226400 670846 226409
rect 670790 226335 670846 226344
rect 670792 226092 670844 226098
rect 670792 226034 670844 226040
rect 670804 225049 670832 226034
rect 670790 225040 670846 225049
rect 670790 224975 670846 224984
rect 670436 224926 670648 224954
rect 670436 215294 670464 224926
rect 670792 224868 670844 224874
rect 670792 224810 670844 224816
rect 670608 224460 670660 224466
rect 670608 224402 670660 224408
rect 670620 216322 670648 224402
rect 670804 223961 670832 224810
rect 670790 223952 670846 223961
rect 670790 223887 670846 223896
rect 670988 223666 671016 235758
rect 671172 234394 671200 262103
rect 671434 258496 671490 258505
rect 671434 258431 671490 258440
rect 671160 234388 671212 234394
rect 671160 234330 671212 234336
rect 671160 234252 671212 234258
rect 671160 234194 671212 234200
rect 671172 225706 671200 234194
rect 671080 225678 671200 225706
rect 671080 224954 671108 225678
rect 671250 225584 671306 225593
rect 671250 225519 671306 225528
rect 671264 225282 671292 225519
rect 671252 225276 671304 225282
rect 671252 225218 671304 225224
rect 671080 224926 671384 224954
rect 670792 223644 670844 223650
rect 670988 223638 671292 223666
rect 670792 223586 670844 223592
rect 670804 223417 670832 223586
rect 670790 223408 670846 223417
rect 670790 223343 670846 223352
rect 671022 223372 671074 223378
rect 671022 223314 671074 223320
rect 671034 223258 671062 223314
rect 671034 223230 671108 223258
rect 670792 223168 670844 223174
rect 670792 223110 670844 223116
rect 670804 222601 670832 223110
rect 670790 222592 670846 222601
rect 670790 222527 670846 222536
rect 670792 222420 670844 222426
rect 670792 222362 670844 222368
rect 670804 218929 670832 222362
rect 670790 218920 670846 218929
rect 670790 218855 670846 218864
rect 671080 217410 671108 223230
rect 670804 217382 671108 217410
rect 670804 217297 670832 217382
rect 670790 217288 670846 217297
rect 670790 217223 670846 217232
rect 670974 216608 671030 216617
rect 670974 216543 671030 216552
rect 670620 216294 670740 216322
rect 670712 215937 670740 216294
rect 670698 215928 670754 215937
rect 670698 215863 670754 215872
rect 670988 215778 671016 216543
rect 670804 215750 671016 215778
rect 670436 215266 670648 215294
rect 670620 169697 670648 215266
rect 670804 202881 670832 215750
rect 671264 215642 671292 223638
rect 670988 215614 671292 215642
rect 670790 202872 670846 202881
rect 670790 202807 670846 202816
rect 670606 169688 670662 169697
rect 670606 169623 670662 169632
rect 670514 169144 670570 169153
rect 670514 169079 670570 169088
rect 670332 160064 670384 160070
rect 670332 160006 670384 160012
rect 670528 150113 670556 169079
rect 670988 157334 671016 215614
rect 671356 215506 671384 224926
rect 671264 215478 671384 215506
rect 671264 215294 671292 215478
rect 671448 215294 671476 258431
rect 671632 237454 671660 263566
rect 671802 260944 671858 260953
rect 671802 260879 671858 260888
rect 671816 246673 671844 260879
rect 671986 256456 672042 256465
rect 671986 256391 672042 256400
rect 671802 246664 671858 246673
rect 671802 246599 671858 246608
rect 671620 237448 671672 237454
rect 671620 237390 671672 237396
rect 671620 236632 671672 236638
rect 671620 236574 671672 236580
rect 671632 224954 671660 236574
rect 671804 236428 671856 236434
rect 671804 236370 671856 236376
rect 671816 234614 671844 236370
rect 671816 234586 671936 234614
rect 671172 215266 671292 215294
rect 671356 215266 671476 215294
rect 671540 224926 671660 224954
rect 671172 177993 671200 215266
rect 671158 177984 671214 177993
rect 671158 177919 671214 177928
rect 670804 157306 671016 157334
rect 670804 155174 670832 157306
rect 670792 155168 670844 155174
rect 670792 155110 670844 155116
rect 670514 150104 670570 150113
rect 670514 150039 670570 150048
rect 670148 148776 670200 148782
rect 670148 148718 670200 148724
rect 671356 138014 671384 215266
rect 671540 145353 671568 224926
rect 671712 224528 671764 224534
rect 671712 224470 671764 224476
rect 671724 221785 671752 224470
rect 671710 221776 671766 221785
rect 671710 221711 671766 221720
rect 671908 215294 671936 234586
rect 671724 215266 671936 215294
rect 671724 150385 671752 215266
rect 672000 210497 672028 256391
rect 672172 236836 672224 236842
rect 672172 236778 672224 236784
rect 672184 235958 672212 236778
rect 672172 235952 672224 235958
rect 672172 235894 672224 235900
rect 672172 233912 672224 233918
rect 672172 233854 672224 233860
rect 672184 233753 672212 233854
rect 672170 233744 672226 233753
rect 672170 233679 672226 233688
rect 672264 233300 672316 233306
rect 672264 233242 672316 233248
rect 672276 230738 672304 233242
rect 672276 230710 672396 230738
rect 672172 230648 672224 230654
rect 672172 230590 672224 230596
rect 672184 228410 672212 230590
rect 672172 228404 672224 228410
rect 672172 228346 672224 228352
rect 672170 226400 672226 226409
rect 672168 226370 672170 226386
rect 672156 226364 672170 226370
rect 672208 226335 672226 226344
rect 672156 226306 672208 226312
rect 672368 225978 672396 230710
rect 672092 225950 672396 225978
rect 672092 225434 672120 225950
rect 672264 225888 672316 225894
rect 672262 225856 672264 225865
rect 672316 225856 672318 225865
rect 672262 225791 672318 225800
rect 672262 225584 672318 225593
rect 672262 225519 672264 225528
rect 672316 225519 672318 225528
rect 672264 225490 672316 225496
rect 672092 225406 672304 225434
rect 672156 225344 672208 225350
rect 672154 225312 672156 225321
rect 672208 225312 672210 225321
rect 672154 225247 672210 225256
rect 672276 225026 672304 225406
rect 672184 224998 672304 225026
rect 672184 215294 672212 224998
rect 672184 215266 672304 215294
rect 671986 210488 672042 210497
rect 671986 210423 672042 210432
rect 671986 209944 672042 209953
rect 671986 209879 672042 209888
rect 672000 193225 672028 209879
rect 672276 203946 672304 215266
rect 672460 208394 672488 281574
rect 672552 277394 672580 282886
rect 672552 277366 672672 277394
rect 672092 203918 672304 203946
rect 672368 208366 672488 208394
rect 672092 198734 672120 203918
rect 672368 203810 672396 208366
rect 672644 208321 672672 277366
rect 672736 208394 672764 282886
rect 672920 244274 672948 348463
rect 673196 311894 673224 355399
rect 673932 355065 673960 399735
rect 674380 396092 674432 396098
rect 674380 396034 674432 396040
rect 674194 393136 674250 393145
rect 674194 393071 674250 393080
rect 674208 379514 674236 393071
rect 674392 382226 674420 396034
rect 674576 395321 674604 403242
rect 676048 402665 676076 410479
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676218 403336 676274 403345
rect 676218 403271 676220 403280
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 676034 402656 676090 402665
rect 676034 402591 676090 402600
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 676048 398886 676076 399327
rect 674840 398880 674892 398886
rect 674840 398822 674892 398828
rect 676036 398880 676088 398886
rect 676036 398822 676088 398828
rect 674562 395312 674618 395321
rect 674562 395247 674618 395256
rect 674656 395140 674708 395146
rect 674656 395082 674708 395088
rect 674380 382220 674432 382226
rect 674380 382162 674432 382168
rect 674208 379486 674420 379514
rect 674392 378146 674420 379486
rect 674380 378140 674432 378146
rect 674380 378082 674432 378088
rect 674668 375238 674696 395082
rect 674852 384810 674880 398822
rect 679622 398440 679678 398449
rect 679622 398375 679678 398384
rect 676218 398032 676274 398041
rect 676218 397967 676274 397976
rect 676232 396234 676260 397967
rect 675024 396228 675076 396234
rect 675024 396170 675076 396176
rect 676220 396228 676272 396234
rect 676220 396170 676272 396176
rect 674840 384804 674892 384810
rect 674840 384746 674892 384752
rect 675036 382582 675064 396170
rect 676034 396128 676090 396137
rect 676034 396063 676036 396072
rect 676088 396063 676090 396072
rect 676036 396034 676088 396040
rect 676218 395584 676274 395593
rect 676218 395519 676274 395528
rect 676232 395146 676260 395519
rect 676220 395140 676272 395146
rect 676220 395082 676272 395088
rect 675206 394496 675262 394505
rect 675206 394431 675262 394440
rect 675220 393145 675248 394431
rect 675206 393136 675262 393145
rect 675206 393071 675262 393080
rect 679636 389162 679664 398375
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 675208 389156 675260 389162
rect 675208 389098 675260 389104
rect 679624 389156 679676 389162
rect 679624 389098 679676 389104
rect 675220 386374 675248 389098
rect 681016 388521 681044 397559
rect 681002 388512 681058 388521
rect 681002 388447 681058 388456
rect 675208 386368 675260 386374
rect 675208 386310 675260 386316
rect 675312 386261 675418 386289
rect 675312 382945 675340 386261
rect 675484 386028 675536 386034
rect 675484 385970 675536 385976
rect 675496 385696 675524 385970
rect 675758 385384 675814 385393
rect 675758 385319 675814 385328
rect 675772 385084 675800 385319
rect 675484 384804 675536 384810
rect 675484 384746 675536 384752
rect 675496 384435 675524 384746
rect 675298 382936 675354 382945
rect 675298 382871 675354 382880
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675116 382220 675168 382226
rect 675758 382191 675814 382200
rect 675116 382162 675168 382168
rect 675128 381426 675156 382162
rect 675772 382024 675800 382191
rect 675128 381398 675418 381426
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377496 675814 377505
rect 675758 377431 675814 377440
rect 675772 377060 675800 377431
rect 675114 376680 675170 376689
rect 675114 376615 675170 376624
rect 675128 376462 675156 376615
rect 675128 376434 675340 376462
rect 675312 376394 675340 376434
rect 675404 376394 675432 376448
rect 675312 376366 675432 376394
rect 674668 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372776 675708 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675574 358320 675630 358329
rect 675574 358255 675630 358264
rect 673918 355056 673974 355065
rect 673918 354991 673974 355000
rect 674102 354648 674158 354657
rect 674102 354583 674158 354592
rect 673734 352608 673790 352617
rect 673734 352543 673790 352552
rect 673366 349752 673422 349761
rect 673366 349687 673422 349696
rect 673380 335617 673408 349687
rect 673550 349344 673606 349353
rect 673550 349279 673606 349288
rect 673366 335608 673422 335617
rect 673366 335543 673422 335552
rect 673564 332761 673592 349279
rect 673748 333985 673776 352543
rect 673918 348936 673974 348945
rect 673918 348871 673974 348880
rect 673734 333976 673790 333985
rect 673734 333911 673790 333920
rect 673550 332752 673606 332761
rect 673550 332687 673606 332696
rect 673932 331265 673960 348871
rect 673918 331256 673974 331265
rect 673918 331191 673974 331200
rect 674116 325694 674144 354583
rect 674746 354240 674802 354249
rect 674746 354175 674802 354184
rect 674286 350976 674342 350985
rect 674286 350911 674342 350920
rect 674300 345014 674328 350911
rect 674562 350568 674618 350577
rect 674562 350503 674618 350512
rect 674576 345014 674604 350503
rect 674300 344986 674420 345014
rect 674576 344986 674696 345014
rect 674392 336598 674420 344986
rect 674380 336592 674432 336598
rect 674380 336534 674432 336540
rect 674668 330049 674696 344986
rect 674760 339402 674788 354175
rect 675588 352889 675616 358255
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356561 675984 357847
rect 675942 356552 675998 356561
rect 675942 356487 675998 356496
rect 675850 353832 675906 353841
rect 675850 353767 675906 353776
rect 675574 352880 675630 352889
rect 675574 352815 675630 352824
rect 675864 351937 675892 353767
rect 675850 351928 675906 351937
rect 675850 351863 675906 351872
rect 676034 351792 676090 351801
rect 676034 351727 676090 351736
rect 676048 347478 676076 351727
rect 683118 347712 683174 347721
rect 683118 347647 683174 347656
rect 676036 347472 676088 347478
rect 676036 347414 676088 347420
rect 676496 347472 676548 347478
rect 676496 347414 676548 347420
rect 676034 347304 676090 347313
rect 676034 347239 676090 347248
rect 676048 345681 676076 347239
rect 676508 346633 676536 347414
rect 676494 346624 676550 346633
rect 676494 346559 676550 346568
rect 683132 346497 683160 347647
rect 683118 346488 683174 346497
rect 683118 346423 683174 346432
rect 676034 345672 676090 345681
rect 676034 345607 676090 345616
rect 675128 341074 675418 341102
rect 674760 339386 674880 339402
rect 674760 339380 674892 339386
rect 674760 339374 674840 339380
rect 674840 339322 674892 339328
rect 675128 338745 675156 341074
rect 675574 340776 675630 340785
rect 675574 340711 675630 340720
rect 675588 340544 675616 340711
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675484 339380 675536 339386
rect 675484 339322 675536 339328
rect 675496 339252 675524 339322
rect 675114 338736 675170 338745
rect 675114 338671 675170 338680
rect 675666 337784 675722 337793
rect 675666 337719 675722 337728
rect 675680 337416 675708 337719
rect 675114 337240 675170 337249
rect 675114 337175 675170 337184
rect 675128 336857 675156 337175
rect 675128 336829 675418 336857
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675114 332344 675170 332353
rect 675114 332279 675170 332288
rect 675128 331889 675156 332279
rect 675128 331861 675418 331889
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 674668 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675128 327542 675418 327570
rect 674116 325666 674512 325694
rect 673366 312080 673422 312089
rect 673366 312015 673422 312024
rect 673104 311866 673224 311894
rect 673104 310865 673132 311866
rect 673090 310856 673146 310865
rect 673090 310791 673146 310800
rect 673182 310584 673238 310593
rect 673182 310519 673238 310528
rect 673196 266665 673224 310519
rect 673380 267481 673408 312015
rect 674484 310049 674512 325666
rect 675128 325281 675156 327542
rect 675312 326454 675432 326482
rect 675312 325553 675340 326454
rect 675404 326332 675432 326454
rect 675298 325544 675354 325553
rect 675298 325479 675354 325488
rect 675114 325272 675170 325281
rect 675114 325207 675170 325216
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313984 676274 313993
rect 676218 313919 676274 313928
rect 674654 310448 674710 310457
rect 674654 310383 674710 310392
rect 674470 310040 674526 310049
rect 674470 309975 674526 309984
rect 674194 309632 674250 309641
rect 674194 309567 674250 309576
rect 674010 303920 674066 303929
rect 674010 303855 674066 303864
rect 674024 286521 674052 303855
rect 674010 286512 674066 286521
rect 674010 286447 674066 286456
rect 673366 267472 673422 267481
rect 673366 267407 673422 267416
rect 673918 267064 673974 267073
rect 673918 266999 673974 267008
rect 673182 266656 673238 266665
rect 673182 266591 673238 266600
rect 673550 266248 673606 266257
rect 673550 266183 673606 266192
rect 673366 260536 673422 260545
rect 673366 260471 673422 260480
rect 673182 258904 673238 258913
rect 673182 258839 673238 258848
rect 672828 244246 672948 244274
rect 672828 227882 672856 244246
rect 673196 241505 673224 258839
rect 673182 241496 673238 241505
rect 673182 241431 673238 241440
rect 673380 240281 673408 260471
rect 673564 241777 673592 266183
rect 673734 265432 673790 265441
rect 673734 265367 673790 265376
rect 673748 242049 673776 265367
rect 673932 244274 673960 266999
rect 674208 265033 674236 309567
rect 674378 305144 674434 305153
rect 674378 305079 674434 305088
rect 674392 287026 674420 305079
rect 674668 304994 674696 310383
rect 675850 309360 675906 309369
rect 676232 309346 676260 313919
rect 675906 309318 676260 309346
rect 675850 309295 675906 309304
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675114 308000 675170 308009
rect 675114 307935 675170 307944
rect 674484 304966 674696 304994
rect 674484 302234 674512 304966
rect 674654 303512 674710 303521
rect 674654 303447 674710 303456
rect 674484 302206 674604 302234
rect 674380 287020 674432 287026
rect 674380 286962 674432 286968
rect 674378 283520 674434 283529
rect 674378 283455 674434 283464
rect 674392 267889 674420 283455
rect 674378 267880 674434 267889
rect 674378 267815 674434 267824
rect 674576 267730 674604 302206
rect 674484 267702 674604 267730
rect 674484 266014 674512 267702
rect 674472 266008 674524 266014
rect 674472 265950 674524 265956
rect 674194 265024 674250 265033
rect 674194 264959 674250 264968
rect 674470 264616 674526 264625
rect 674470 264551 674526 264560
rect 674286 262576 674342 262585
rect 674286 262511 674342 262520
rect 674102 259312 674158 259321
rect 674102 259247 674158 259256
rect 673932 244246 674052 244274
rect 673734 242040 673790 242049
rect 673734 241975 673790 241984
rect 673550 241768 673606 241777
rect 673550 241703 673606 241712
rect 673366 240272 673422 240281
rect 673366 240207 673422 240216
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 672966 236586 672994 236642
rect 672966 236558 673960 236586
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 673196 236178 673224 236234
rect 673196 236150 673500 236178
rect 673276 235952 673328 235958
rect 673276 235894 673328 235900
rect 673000 235748 673052 235754
rect 673000 235690 673052 235696
rect 673012 235634 673040 235690
rect 672920 235606 673040 235634
rect 672920 233186 672948 235606
rect 673092 235544 673144 235550
rect 673092 235486 673144 235492
rect 673104 233306 673132 235486
rect 673288 234433 673316 235894
rect 673274 234424 673330 234433
rect 673274 234359 673330 234368
rect 673092 233300 673144 233306
rect 673092 233242 673144 233248
rect 672920 233158 673040 233186
rect 673012 233102 673040 233158
rect 673000 233096 673052 233102
rect 673000 233038 673052 233044
rect 673472 230602 673500 236150
rect 673642 234832 673698 234841
rect 673642 234767 673644 234776
rect 673696 234767 673698 234776
rect 673644 234738 673696 234744
rect 673472 230574 673684 230602
rect 673458 230480 673514 230489
rect 673458 230415 673460 230424
rect 673512 230415 673514 230424
rect 673460 230386 673512 230392
rect 673184 229424 673236 229430
rect 673184 229366 673236 229372
rect 673196 228585 673224 229366
rect 673368 229152 673420 229158
rect 673368 229094 673420 229100
rect 673182 228576 673238 228585
rect 673182 228511 673238 228520
rect 672828 227854 672948 227882
rect 672920 227798 672948 227854
rect 672908 227792 672960 227798
rect 672908 227734 672960 227740
rect 673380 227089 673408 229094
rect 673656 227202 673684 230574
rect 673932 229786 673960 236558
rect 673564 227186 673684 227202
rect 673552 227180 673684 227186
rect 673604 227174 673684 227180
rect 673748 229758 673960 229786
rect 673552 227122 673604 227128
rect 673366 227080 673422 227089
rect 673366 227015 673422 227024
rect 673552 227044 673604 227050
rect 673552 226986 673604 226992
rect 673564 226817 673592 226986
rect 673550 226808 673606 226817
rect 673550 226743 673606 226752
rect 673000 226568 673052 226574
rect 673000 226510 673052 226516
rect 673012 222873 673040 226510
rect 673458 223408 673514 223417
rect 673458 223343 673514 223352
rect 672998 222864 673054 222873
rect 672998 222799 673054 222808
rect 673472 219434 673500 223343
rect 673000 219428 673052 219434
rect 673000 219370 673052 219376
rect 673460 219428 673512 219434
rect 673460 219370 673512 219376
rect 673012 213625 673040 219370
rect 673182 215792 673238 215801
rect 673182 215727 673238 215736
rect 672998 213616 673054 213625
rect 672998 213551 673054 213560
rect 672906 213344 672962 213353
rect 672906 213279 672962 213288
rect 672736 208366 672856 208394
rect 672630 208312 672686 208321
rect 672630 208247 672686 208256
rect 672828 203833 672856 208366
rect 672920 203946 672948 213279
rect 672920 203918 673040 203946
rect 672184 203782 672396 203810
rect 672814 203824 672870 203833
rect 672184 203266 672212 203782
rect 672814 203759 672870 203768
rect 672722 203416 672778 203425
rect 672722 203351 672778 203360
rect 672736 203266 672764 203351
rect 672184 203238 672488 203266
rect 672092 198706 672304 198734
rect 671986 193216 672042 193225
rect 671986 193151 672042 193160
rect 671986 170368 672042 170377
rect 671986 170303 672042 170312
rect 672000 150385 672028 170303
rect 672276 168201 672304 198706
rect 672460 177721 672488 203238
rect 672552 203238 672764 203266
rect 672552 183554 672580 203238
rect 672814 202600 672870 202609
rect 672814 202535 672870 202544
rect 672828 193066 672856 202535
rect 673012 198734 673040 203918
rect 673196 200841 673224 215727
rect 673550 214976 673606 214985
rect 673550 214911 673606 214920
rect 673366 213752 673422 213761
rect 673366 213687 673422 213696
rect 673182 200832 673238 200841
rect 673182 200767 673238 200776
rect 672920 198706 673040 198734
rect 672920 193214 672948 198706
rect 673380 196081 673408 213687
rect 673564 201113 673592 214911
rect 673550 201104 673606 201113
rect 673550 201039 673606 201048
rect 673366 196072 673422 196081
rect 673366 196007 673422 196016
rect 672920 193186 673132 193214
rect 672828 193050 672948 193066
rect 672828 193044 672960 193050
rect 672828 193038 672908 193044
rect 672908 192986 672960 192992
rect 673104 183554 673132 193186
rect 673368 193044 673420 193050
rect 673368 192986 673420 192992
rect 673380 185609 673408 192986
rect 673366 185600 673422 185609
rect 673366 185535 673422 185544
rect 672552 183526 672764 183554
rect 672446 177712 672502 177721
rect 672446 177647 672502 177656
rect 672262 168192 672318 168201
rect 672262 168127 672318 168136
rect 672262 167920 672318 167929
rect 672318 167878 672580 167906
rect 672262 167855 672318 167864
rect 672354 166288 672410 166297
rect 672354 166223 672410 166232
rect 672170 165608 672226 165617
rect 672170 165543 672226 165552
rect 671710 150376 671766 150385
rect 671710 150311 671766 150320
rect 671986 150376 672042 150385
rect 671986 150311 672042 150320
rect 671526 145344 671582 145353
rect 671526 145279 671582 145288
rect 670804 137986 671384 138014
rect 669964 136264 670016 136270
rect 669964 136206 670016 136212
rect 669226 133784 669282 133793
rect 669226 133719 669282 133728
rect 669240 132977 669268 133719
rect 669226 132968 669282 132977
rect 669226 132903 669282 132912
rect 668950 131200 669006 131209
rect 668950 131135 669006 131144
rect 668766 130656 668822 130665
rect 668766 130591 668822 130600
rect 668584 129192 668636 129198
rect 668584 129134 668636 129140
rect 668596 129033 668624 129134
rect 668582 129024 668638 129033
rect 668582 128959 668638 128968
rect 668582 126984 668638 126993
rect 668582 126919 668638 126928
rect 668030 125352 668086 125361
rect 668030 125287 668086 125296
rect 589924 122052 589976 122058
rect 589924 121994 589976 122000
rect 589554 121544 589610 121553
rect 589554 121479 589556 121488
rect 589608 121479 589610 121488
rect 589556 121450 589608 121456
rect 589372 120760 589424 120766
rect 589372 120702 589424 120708
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589462 110120 589518 110129
rect 589462 110055 589518 110064
rect 589476 109138 589504 110055
rect 589464 109132 589516 109138
rect 589464 109074 589516 109080
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589830 105224 589886 105233
rect 589830 105159 589886 105168
rect 589844 104922 589872 105159
rect 589832 104916 589884 104922
rect 589832 104858 589884 104864
rect 590304 103514 590332 114951
rect 666650 109372 666706 109381
rect 666650 109307 666706 109316
rect 666664 103514 666692 109307
rect 667940 108860 667992 108866
rect 667940 108802 667992 108808
rect 667952 107817 667980 108802
rect 667938 107808 667994 107817
rect 667938 107743 667994 107752
rect 668030 106176 668086 106185
rect 668030 106111 668086 106120
rect 589936 103486 590332 103514
rect 666572 103486 666692 103514
rect 668044 103514 668072 106111
rect 668216 104848 668268 104854
rect 668216 104790 668268 104796
rect 668228 104417 668256 104790
rect 668214 104408 668270 104417
rect 668214 104343 668270 104352
rect 668044 103486 668164 103514
rect 588728 103420 588780 103426
rect 588728 103362 588780 103368
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 88330 589964 103486
rect 592684 100020 592736 100026
rect 592684 99962 592736 99968
rect 595272 100014 595608 100042
rect 596344 100014 596496 100042
rect 592132 97300 592184 97306
rect 592132 97242 592184 97248
rect 591304 96076 591356 96082
rect 591304 96018 591356 96024
rect 590936 94988 590988 94994
rect 590936 94930 590988 94936
rect 590948 91798 590976 94930
rect 590936 91792 590988 91798
rect 590936 91734 590988 91740
rect 589924 88324 589976 88330
rect 589924 88266 589976 88272
rect 588544 73160 588596 73166
rect 588544 73102 588596 73108
rect 587164 62076 587216 62082
rect 587164 62018 587216 62024
rect 591316 54505 591344 96018
rect 592144 94994 592172 97242
rect 592132 94988 592184 94994
rect 592132 94930 592184 94936
rect 592696 64870 592724 99962
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 594064 95940 594116 95946
rect 594064 95882 594116 95888
rect 592684 64864 592736 64870
rect 592684 64806 592736 64812
rect 594076 57934 594104 95882
rect 595272 93854 595300 99078
rect 596180 96960 596232 96966
rect 596180 96902 596232 96908
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 594064 57928 594116 57934
rect 594064 57870 594116 57876
rect 596192 55078 596220 96902
rect 596468 55214 596496 100014
rect 596744 100014 597080 100042
rect 597664 100014 597816 100042
rect 597940 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600332 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602632 100014 602968 100042
rect 603092 100014 603704 100042
rect 596744 96966 596772 100014
rect 596732 96960 596784 96966
rect 596732 96902 596784 96908
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 596180 55072 596232 55078
rect 596180 55014 596232 55020
rect 597664 54942 597692 100014
rect 597652 54936 597704 54942
rect 597652 54878 597704 54884
rect 597940 54806 597968 100014
rect 598952 97306 598980 100014
rect 598940 97300 598992 97306
rect 598940 97242 598992 97248
rect 599504 84194 599532 100014
rect 598952 84166 599532 84194
rect 598952 56030 598980 84166
rect 600332 57254 600360 100014
rect 600884 84194 600912 100014
rect 600516 84166 600912 84194
rect 600516 79354 600544 84166
rect 600504 79348 600556 79354
rect 600504 79290 600556 79296
rect 600320 57248 600372 57254
rect 600320 57190 600372 57196
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 601896 55894 601924 100014
rect 602632 96082 602660 100014
rect 602620 96076 602672 96082
rect 602620 96018 602672 96024
rect 603092 58682 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613884 100042
rect 604426 99742 604500 99770
rect 604472 58818 604500 99742
rect 605484 97442 605512 100014
rect 605472 97436 605524 97442
rect 605472 97378 605524 97384
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 91798 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 91792 606996 91798
rect 606944 91734 606996 91740
rect 607140 75342 607168 96902
rect 607692 94518 607720 100014
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 608520 84182 608548 100014
rect 609164 96762 609192 100014
rect 609152 96756 609204 96762
rect 609152 96698 609204 96704
rect 609704 96756 609756 96762
rect 609704 96698 609756 96704
rect 609716 93158 609744 96698
rect 609704 93152 609756 93158
rect 609704 93094 609756 93100
rect 609900 85406 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 91050 611308 100014
rect 611912 97436 611964 97442
rect 611912 97378 611964 97384
rect 611924 93854 611952 97378
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 91044 611320 91050
rect 611268 90986 611320 90992
rect 609888 85400 609940 85406
rect 609888 85342 609940 85348
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76702 612044 93826
rect 612660 79354 612688 96834
rect 613856 80850 613884 100014
rect 613994 99770 614022 100028
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620140 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613994 99742 614068 99770
rect 613844 80844 613896 80850
rect 613844 80786 613896 80792
rect 614040 79490 614068 99742
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 94994 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 94988 616564 94994
rect 616512 94930 616564 94936
rect 615236 93826 615448 93854
rect 615420 80986 615448 93826
rect 615408 80980 615460 80986
rect 615408 80922 615460 80928
rect 614028 79484 614080 79490
rect 614028 79426 614080 79432
rect 612648 79348 612700 79354
rect 612648 79290 612700 79296
rect 612004 76696 612056 76702
rect 612004 76638 612056 76644
rect 616800 75478 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91186 618208 96834
rect 619560 93838 619588 100014
rect 620112 97170 620140 100014
rect 620284 97436 620336 97442
rect 620284 97378 620336 97384
rect 620100 97164 620152 97170
rect 620100 97106 620152 97112
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618628 93152 618680 93158
rect 618628 93094 618680 93100
rect 618168 91180 618220 91186
rect 618168 91122 618220 91128
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618180 88330 618208 90986
rect 618168 88324 618220 88330
rect 618168 88266 618220 88272
rect 618640 85542 618668 93094
rect 618628 85536 618680 85542
rect 618628 85478 618680 85484
rect 620296 76838 620324 97378
rect 620940 95198 620968 100014
rect 621676 97306 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 623148 97442 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 624620 99074 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 631916 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 624608 99068 624660 99074
rect 624608 99010 624660 99016
rect 625080 98938 625108 99742
rect 625068 98932 625120 98938
rect 625068 98874 625120 98880
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 623136 97436 623188 97442
rect 623136 97378 623188 97384
rect 621664 97300 621716 97306
rect 621664 97242 621716 97248
rect 621664 96076 621716 96082
rect 621664 96018 621716 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620928 94512 620980 94518
rect 620928 94454 620980 94460
rect 620940 89690 620968 94454
rect 620928 89684 620980 89690
rect 620928 89626 620980 89632
rect 621676 86358 621704 96018
rect 625436 95192 625488 95198
rect 625436 95134 625488 95140
rect 624976 94988 625028 94994
rect 624976 94930 625028 94936
rect 622400 91792 622452 91798
rect 622400 91734 622452 91740
rect 622412 88194 622440 91734
rect 624988 88641 625016 94930
rect 625448 94489 625476 95134
rect 625434 94480 625490 94489
rect 625434 94415 625490 94424
rect 625816 92041 625844 97922
rect 626092 96898 626120 100014
rect 626828 97170 626856 100014
rect 627564 97578 627592 100014
rect 628300 97986 628328 100014
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 98326 629800 100014
rect 630508 98598 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98592 630548 98598
rect 630496 98534 630548 98540
rect 629760 98320 629812 98326
rect 629760 98262 629812 98268
rect 628288 97980 628340 97986
rect 628288 97922 628340 97928
rect 627552 97572 627604 97578
rect 627552 97514 627604 97520
rect 629300 97300 629352 97306
rect 629300 97242 629352 97248
rect 626356 97164 626408 97170
rect 626356 97106 626408 97112
rect 626816 97164 626868 97170
rect 626816 97106 626868 97112
rect 626080 96892 626132 96898
rect 626080 96834 626132 96840
rect 626172 93832 626224 93838
rect 626172 93774 626224 93780
rect 626184 92857 626212 93774
rect 626368 93673 626396 97106
rect 629312 95826 629340 97242
rect 630784 95826 630812 99282
rect 631244 97714 631272 100014
rect 631232 97708 631284 97714
rect 631232 97650 631284 97656
rect 631888 97306 631916 100014
rect 632716 97850 632744 100014
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 633268 97442 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 632060 97436 632112 97442
rect 632060 97378 632112 97384
rect 633256 97436 633308 97442
rect 633256 97378 633308 97384
rect 631876 97300 631928 97306
rect 631876 97242 631928 97248
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97378
rect 633452 95826 633480 99146
rect 633624 98184 633676 98190
rect 633624 98126 633676 98132
rect 633636 97578 633664 98126
rect 633624 97572 633676 97578
rect 633624 97514 633676 97520
rect 633808 97572 633860 97578
rect 633808 97514 633860 97520
rect 633820 97170 633848 97514
rect 634188 97170 634216 100014
rect 633808 97164 633860 97170
rect 633808 97106 633860 97112
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 634740 97034 634768 100014
rect 635004 99068 635056 99074
rect 635004 99010 635056 99016
rect 634728 97028 634780 97034
rect 634728 96970 634780 96976
rect 635016 95826 635044 99010
rect 635568 96937 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635554 96928 635610 96937
rect 635554 96863 635610 96872
rect 635752 95985 635780 100014
rect 636292 98932 636344 98938
rect 636292 98874 636344 98880
rect 635738 95976 635794 95985
rect 635738 95911 635794 95920
rect 636304 95826 636332 98874
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96354 637620 99742
rect 637764 96892 637816 96898
rect 637764 96834 637816 96840
rect 637580 96348 637632 96354
rect 637580 96290 637632 96296
rect 637776 95826 637804 96834
rect 638604 96490 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 638592 96484 638644 96490
rect 638592 96426 638644 96432
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639064 95810 639092 99742
rect 639236 97572 639288 97578
rect 639236 97514 639288 97520
rect 639248 95826 639276 97514
rect 640076 96626 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640064 96620 640116 96626
rect 640064 96562 640116 96568
rect 640536 96082 640564 99742
rect 640708 98184 640760 98190
rect 640708 98126 640760 98132
rect 640524 96076 640576 96082
rect 640524 96018 640576 96024
rect 640720 95826 640748 98126
rect 641548 96490 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98048 642232 98054
rect 642180 97990 642232 97996
rect 641994 96520 642050 96529
rect 641352 96484 641404 96490
rect 641352 96426 641404 96432
rect 641536 96484 641588 96490
rect 641994 96455 642050 96464
rect 641536 96426 641588 96432
rect 639052 95804 639104 95810
rect 639248 95798 639584 95826
rect 640720 95798 641056 95826
rect 639052 95746 639104 95752
rect 641364 95470 641392 96426
rect 642192 95826 642220 97990
rect 643020 97578 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97572 643060 97578
rect 643008 97514 643060 97520
rect 642192 95798 642528 95826
rect 643480 95470 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643664 95826 643692 98738
rect 644308 96830 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 96824 644348 96830
rect 644296 96766 644348 96772
rect 644952 96218 644980 99742
rect 645308 98320 645360 98326
rect 645308 98262 645360 98268
rect 645124 96620 645176 96626
rect 645124 96562 645176 96568
rect 644940 96212 644992 96218
rect 644940 96154 644992 96160
rect 643664 95798 644000 95826
rect 645136 95674 645164 96562
rect 645320 95826 645348 98262
rect 645582 96112 645638 96121
rect 645780 96082 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648476 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 646424 96626 646452 99742
rect 647160 98666 647188 99742
rect 647148 98660 647200 98666
rect 647148 98602 647200 98608
rect 646596 98592 646648 98598
rect 646596 98534 646648 98540
rect 646412 96620 646464 96626
rect 646412 96562 646464 96568
rect 645582 96047 645584 96056
rect 645636 96047 645638 96056
rect 645768 96076 645820 96082
rect 645584 96018 645636 96024
rect 645768 96018 645820 96024
rect 646608 95826 646636 98534
rect 647516 97844 647568 97850
rect 647516 97786 647568 97792
rect 647332 97708 647384 97714
rect 647332 97650 647384 97656
rect 647056 97028 647108 97034
rect 647056 96970 647108 96976
rect 645320 95798 645472 95826
rect 646608 95798 646944 95826
rect 645124 95668 645176 95674
rect 645124 95610 645176 95616
rect 641352 95464 641404 95470
rect 641352 95406 641404 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 647068 95198 647096 96970
rect 647056 95192 647108 95198
rect 647056 95134 647108 95140
rect 647344 95033 647372 97650
rect 647330 95024 647386 95033
rect 647330 94959 647386 94968
rect 647528 93770 647556 97786
rect 648066 96520 648122 96529
rect 648066 96455 648068 96464
rect 648120 96455 648122 96464
rect 648068 96426 648120 96432
rect 647884 96212 647936 96218
rect 647884 96154 647936 96160
rect 647896 95849 647924 96154
rect 648068 96076 648120 96082
rect 648068 96018 648120 96024
rect 647882 95840 647938 95849
rect 647882 95775 647938 95784
rect 647884 95464 647936 95470
rect 647884 95406 647936 95412
rect 647700 95328 647752 95334
rect 647700 95270 647752 95276
rect 647516 93764 647568 93770
rect 647516 93706 647568 93712
rect 626354 93664 626410 93673
rect 626354 93599 626410 93608
rect 626170 92848 626226 92857
rect 626170 92783 626226 92792
rect 647712 92478 647740 95270
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 647700 92472 647752 92478
rect 647700 92414 647752 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 625436 89684 625488 89690
rect 625436 89626 625488 89632
rect 625250 89584 625306 89593
rect 625250 89519 625306 89528
rect 625264 88641 625292 89519
rect 625448 88777 625476 89626
rect 625434 88768 625490 88777
rect 625434 88703 625490 88712
rect 624974 88632 625030 88641
rect 624974 88567 625030 88576
rect 625250 88632 625306 88641
rect 625250 88567 625306 88576
rect 625620 88324 625672 88330
rect 625620 88266 625672 88272
rect 622400 88188 622452 88194
rect 622400 88130 622452 88136
rect 625632 87145 625660 88266
rect 626448 88188 626500 88194
rect 626448 88130 626500 88136
rect 626460 87961 626488 88130
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 625618 87136 625674 87145
rect 625618 87071 625674 87080
rect 647896 86630 647924 95406
rect 648080 95402 648108 96018
rect 648068 95396 648120 95402
rect 648068 95338 648120 95344
rect 648252 93764 648304 93770
rect 648252 93706 648304 93712
rect 648264 89593 648292 93706
rect 648250 89584 648306 89593
rect 648250 89519 648306 89528
rect 648448 87038 648476 100014
rect 648620 97300 648672 97306
rect 648620 97242 648672 97248
rect 648632 92041 648660 97242
rect 648908 96490 648936 100014
rect 649080 97164 649132 97170
rect 649080 97106 649132 97112
rect 648896 96484 648948 96490
rect 648896 96426 648948 96432
rect 648802 96112 648858 96121
rect 648802 96047 648804 96056
rect 648856 96047 648858 96056
rect 648804 96018 648856 96024
rect 648804 95804 648856 95810
rect 648804 95746 648856 95752
rect 648618 92032 648674 92041
rect 648618 91967 648674 91976
rect 648816 90846 648844 95746
rect 648804 90840 648856 90846
rect 648804 90782 648856 90788
rect 649092 89714 649120 97106
rect 649262 96520 649318 96529
rect 649262 96455 649318 96464
rect 649276 96218 649304 96455
rect 649264 96212 649316 96218
rect 649264 96154 649316 96160
rect 648632 89686 649120 89714
rect 648436 87032 648488 87038
rect 648436 86974 648488 86980
rect 647884 86624 647936 86630
rect 647884 86566 647936 86572
rect 621664 86352 621716 86358
rect 626448 86352 626500 86358
rect 621664 86294 621716 86300
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 625342 85504 625398 85513
rect 626448 85478 626500 85484
rect 625342 85439 625398 85448
rect 625356 85338 625384 85439
rect 625344 85332 625396 85338
rect 625344 85274 625396 85280
rect 626460 84697 626488 85478
rect 648632 84697 648660 89686
rect 649736 88806 649764 100014
rect 650380 97714 650408 100014
rect 650368 97708 650420 97714
rect 650368 97650 650420 97656
rect 650552 97436 650604 97442
rect 650552 97378 650604 97384
rect 650276 95192 650328 95198
rect 650276 95134 650328 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 626446 84688 626502 84697
rect 626446 84623 626502 84632
rect 648618 84688 648674 84697
rect 648618 84623 648674 84632
rect 625804 84176 625856 84182
rect 625804 84118 625856 84124
rect 625816 83881 625844 84118
rect 625802 83872 625858 83881
rect 625802 83807 625858 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 81122 628788 83263
rect 650288 82249 650316 95134
rect 650564 87145 650592 97378
rect 651300 93634 651328 100014
rect 651852 97442 651880 100014
rect 651840 97436 651892 97442
rect 651840 97378 651892 97384
rect 652024 96620 652076 96626
rect 652024 96562 652076 96568
rect 651288 93628 651340 93634
rect 651288 93570 651340 93576
rect 650550 87136 650606 87145
rect 650550 87071 650606 87080
rect 652036 86494 652064 96562
rect 652588 95810 652616 100014
rect 653324 96626 653352 100014
rect 653968 97850 653996 100014
rect 653956 97844 654008 97850
rect 653956 97786 654008 97792
rect 654796 96966 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655060 97844 655112 97850
rect 655060 97786 655112 97792
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 653312 96620 653364 96626
rect 653312 96562 653364 96568
rect 652576 95804 652628 95810
rect 652576 95746 652628 95752
rect 652208 95668 652260 95674
rect 652208 95610 652260 95616
rect 652220 86766 652248 95610
rect 655072 94217 655100 97786
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655058 94208 655114 94217
rect 655058 94143 655114 94152
rect 655440 93854 655468 96902
rect 655256 93826 655468 93854
rect 654692 93628 654744 93634
rect 654692 93570 654744 93576
rect 654704 93401 654732 93570
rect 654690 93392 654746 93401
rect 654690 93327 654746 93336
rect 655256 88330 655284 93826
rect 655428 92472 655480 92478
rect 655428 92414 655480 92420
rect 655440 91497 655468 92414
rect 655426 91488 655482 91497
rect 655426 91423 655482 91432
rect 655428 90840 655480 90846
rect 655428 90782 655480 90788
rect 655440 90681 655468 90782
rect 655426 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97238 656848 100014
rect 656808 97232 656860 97238
rect 656808 97174 656860 97180
rect 656716 96960 656768 96966
rect 656716 96902 656768 96908
rect 656346 95840 656402 95849
rect 656346 95775 656402 95784
rect 656164 95532 656216 95538
rect 656164 95474 656216 95480
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 656176 88670 656204 95474
rect 656164 88664 656216 88670
rect 656164 88606 656216 88612
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 652208 86760 652260 86766
rect 652208 86702 652260 86708
rect 652024 86488 652076 86494
rect 652024 86430 652076 86436
rect 656360 86358 656388 95775
rect 656728 86902 656756 96902
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658108 99742 658182 99770
rect 658108 97102 658136 99742
rect 658280 97708 658332 97714
rect 658280 97650 658332 97656
rect 658096 97096 658148 97102
rect 658096 97038 658148 97044
rect 658292 95132 658320 97650
rect 659212 97442 659240 100014
rect 659948 97986 659976 100014
rect 660132 100014 660376 100042
rect 659936 97980 659988 97986
rect 659936 97922 659988 97928
rect 659844 97708 659896 97714
rect 659844 97650 659896 97656
rect 659568 97572 659620 97578
rect 659568 97514 659620 97520
rect 659200 97436 659252 97442
rect 659200 97378 659252 97384
rect 658832 96824 658884 96830
rect 658832 96766 658884 96772
rect 658844 95132 658872 96766
rect 659580 95132 659608 97514
rect 659856 95146 659884 97650
rect 660132 96966 660160 100014
rect 661960 98660 662012 98666
rect 661960 98602 662012 98608
rect 661408 97232 661460 97238
rect 661408 97174 661460 97180
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660672 96348 660724 96354
rect 660672 96290 660724 96296
rect 659856 95118 660146 95146
rect 660684 95132 660712 96290
rect 661420 95132 661448 97174
rect 661972 95132 662000 98602
rect 665364 97980 665416 97986
rect 665364 97922 665416 97928
rect 662512 97844 662564 97850
rect 662512 97786 662564 97792
rect 662524 95132 662552 97786
rect 664352 97436 664404 97442
rect 664352 97378 664404 97384
rect 663064 97096 663116 97102
rect 663064 97038 663116 97044
rect 663076 95132 663104 97038
rect 663984 96212 664036 96218
rect 663984 96154 664036 96160
rect 663800 95804 663852 95810
rect 663800 95746 663852 95752
rect 663812 91089 663840 95746
rect 663996 92585 664024 96154
rect 664168 96076 664220 96082
rect 664168 96018 664220 96024
rect 663982 92576 664038 92585
rect 663982 92511 664038 92520
rect 664180 91769 664208 96018
rect 664166 91760 664222 91769
rect 664166 91695 664222 91704
rect 663798 91080 663854 91089
rect 663798 91015 663854 91024
rect 664364 88806 664392 97378
rect 665180 96620 665232 96626
rect 665180 96562 665232 96568
rect 664536 96484 664588 96490
rect 664536 96426 664588 96432
rect 664548 89865 664576 96426
rect 664534 89856 664590 89865
rect 664534 89791 664590 89800
rect 665192 89049 665220 96562
rect 665376 93401 665404 97922
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664352 88800 664404 88806
rect 664352 88742 664404 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 657188 86494 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86766 660160 88196
rect 660120 86760 660172 86766
rect 660120 86702 660172 86708
rect 657176 86488 657228 86494
rect 657176 86430 657228 86436
rect 660684 86358 660712 88196
rect 661420 86630 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86624 661460 86630
rect 661408 86566 661460 86572
rect 656348 86352 656400 86358
rect 656348 86294 656400 86300
rect 660672 86352 660724 86358
rect 660672 86294 660724 86300
rect 650274 82240 650330 82249
rect 650274 82175 650330 82184
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 81116 628800 81122
rect 628748 81058 628800 81064
rect 629220 80034 629248 81631
rect 642456 81116 642508 81122
rect 642456 81058 642508 81064
rect 632808 80974 633144 81002
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77716 628524 77722
rect 628472 77658 628524 77664
rect 628484 77450 628512 77658
rect 624424 77444 624476 77450
rect 624424 77386 624476 77392
rect 628472 77444 628524 77450
rect 628472 77386 628524 77392
rect 623042 77344 623098 77353
rect 623042 77279 623098 77288
rect 620284 76832 620336 76838
rect 620284 76774 620336 76780
rect 616788 75472 616840 75478
rect 616788 75414 616840 75420
rect 607128 75336 607180 75342
rect 607128 75278 607180 75284
rect 604460 58812 604512 58818
rect 604460 58754 604512 58760
rect 603080 58676 603132 58682
rect 603080 58618 603132 58624
rect 601884 55888 601936 55894
rect 601884 55830 601936 55836
rect 597928 54800 597980 54806
rect 597928 54742 597980 54748
rect 591302 54496 591358 54505
rect 591302 54431 591358 54440
rect 583024 54392 583076 54398
rect 583024 54334 583076 54340
rect 577504 54188 577556 54194
rect 577504 54130 577556 54136
rect 623056 53990 623084 77279
rect 624436 60042 624464 77386
rect 625804 77308 625856 77314
rect 625804 77250 625856 77256
rect 624424 60036 624476 60042
rect 624424 59978 624476 59984
rect 625816 54534 625844 77250
rect 628484 75290 628512 77386
rect 631060 77314 631088 77930
rect 632808 77722 632836 80974
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77716 632848 77722
rect 632796 77658 632848 77664
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 77616 639658 77625
rect 639602 77551 639658 77560
rect 639616 75290 639644 77551
rect 642468 75290 642496 81058
rect 643080 80974 643140 81002
rect 643112 77994 643140 80974
rect 646136 80980 646188 80986
rect 646136 80922 646188 80928
rect 645952 79484 646004 79490
rect 645952 79426 646004 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 645964 67130 645992 79426
rect 646148 69193 646176 80922
rect 647332 80844 647384 80850
rect 647332 80786 647384 80792
rect 646504 75472 646556 75478
rect 646504 75414 646556 75420
rect 646320 75336 646372 75342
rect 646320 75278 646372 75284
rect 646332 74225 646360 75278
rect 646318 74216 646374 74225
rect 646318 74151 646374 74160
rect 646516 71777 646544 75414
rect 646502 71768 646558 71777
rect 646502 71703 646558 71712
rect 646134 69184 646190 69193
rect 646134 69119 646190 69128
rect 646134 67144 646190 67153
rect 645964 67102 646134 67130
rect 646134 67079 646190 67088
rect 625988 66904 626040 66910
rect 625988 66846 626040 66852
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 623044 53984 623096 53990
rect 623044 53926 623096 53932
rect 577136 53508 577188 53514
rect 577136 53450 577188 53456
rect 574284 53304 574336 53310
rect 574284 53246 574336 53252
rect 478144 53236 478196 53242
rect 478144 53178 478196 53184
rect 472806 53071 472862 53080
rect 476672 53100 476724 53106
rect 476672 53042 476724 53048
rect 469956 52828 470008 52834
rect 469956 52770 470008 52776
rect 464232 52550 464568 52578
rect 464692 52550 464936 52578
rect 465152 52550 465488 52578
rect 465612 52550 465948 52578
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132408 46096 132460 46102
rect 132408 46038 132460 46044
rect 131040 45354 131436 45370
rect 131040 45348 131448 45354
rect 131040 45342 131396 45348
rect 131396 45290 131448 45296
rect 131132 45218 131436 45234
rect 131120 45212 131448 45218
rect 131172 45206 131396 45212
rect 131120 45154 131172 45160
rect 131396 45154 131448 45160
rect 132420 44470 132448 46038
rect 132592 45960 132644 45966
rect 132592 45902 132644 45908
rect 132408 44464 132460 44470
rect 132604 44422 132632 45902
rect 132960 45348 133012 45354
rect 132960 45290 133012 45296
rect 132408 44406 132460 44412
rect 132592 44416 132644 44422
rect 132592 44358 132644 44364
rect 132972 44310 133000 45290
rect 133144 45212 133196 45218
rect 133144 45154 133196 45160
rect 132960 44304 133012 44310
rect 132960 44246 133012 44252
rect 133156 44198 133184 45154
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 459204 44441 459232 47654
rect 459190 44432 459246 44441
rect 459190 44367 459246 44376
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 133144 44192 133196 44198
rect 133144 44134 133196 44140
rect 255870 44160 255926 44169
rect 255870 44095 255926 44104
rect 130384 44056 130436 44062
rect 130384 43998 130436 44004
rect 255884 42838 255912 44095
rect 307298 43888 307354 43897
rect 307298 43823 307354 43832
rect 440238 43888 440294 43897
rect 440238 43823 440240 43832
rect 187332 42832 187384 42838
rect 187332 42774 187384 42780
rect 255872 42832 255924 42838
rect 255872 42774 255924 42780
rect 187344 42092 187372 42774
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 43823
rect 440292 43823 440294 43832
rect 441066 43888 441122 43897
rect 441066 43823 441068 43832
rect 440240 43794 440292 43800
rect 441120 43823 441122 43832
rect 441068 43794 441120 43800
rect 410892 42900 410944 42906
rect 410892 42842 410944 42848
rect 415584 42900 415636 42906
rect 415584 42842 415636 42848
rect 310428 42764 310480 42770
rect 310428 42706 310480 42712
rect 364524 42764 364576 42770
rect 364524 42706 364576 42712
rect 310440 42106 310468 42706
rect 361764 42492 361816 42498
rect 361764 42434 361816 42440
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 42434
rect 364536 42362 364564 42706
rect 364892 42628 364944 42634
rect 364892 42570 364944 42576
rect 364524 42356 364576 42362
rect 364524 42298 364576 42304
rect 364904 42092 364932 42570
rect 410904 42498 410932 42842
rect 410892 42492 410944 42498
rect 410892 42434 410944 42440
rect 415596 42362 415624 42842
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 453580 42764 453632 42770
rect 453580 42706 453632 42712
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 416594 42392 416650 42401
rect 415584 42356 415636 42362
rect 416594 42327 416650 42336
rect 415584 42298 415636 42304
rect 415766 42120 415822 42129
rect 415426 42078 415766 42106
rect 194322 42055 194378 42064
rect 416608 42092 416636 42327
rect 415766 42055 415822 42064
rect 427096 42022 427124 42570
rect 429108 42492 429160 42498
rect 429108 42434 429160 42440
rect 427084 42016 427136 42022
rect 427084 41958 427136 41964
rect 405646 41848 405702 41857
rect 405582 41806 405646 41834
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 405646 41783 405702 41792
rect 419906 41783 419962 41792
rect 429120 41750 429148 42434
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 441252 42628 441304 42634
rect 441252 42570 441304 42576
rect 446404 42628 446456 42634
rect 446404 42570 446456 42576
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 441264 41886 441292 42570
rect 446218 42256 446274 42265
rect 446218 42191 446274 42200
rect 441252 41880 441304 41886
rect 441252 41822 441304 41828
rect 429108 41744 429160 41750
rect 429108 41686 429160 41692
rect 446232 41585 446260 42191
rect 446416 42022 446444 42570
rect 446404 42016 446456 42022
rect 446404 41958 446456 41964
rect 449176 41750 449204 42706
rect 453592 41750 453620 42706
rect 454684 42628 454736 42634
rect 454684 42570 454736 42576
rect 454500 42492 454552 42498
rect 454500 42434 454552 42440
rect 454512 42022 454540 42434
rect 454500 42016 454552 42022
rect 454500 41958 454552 41964
rect 454696 41886 454724 42570
rect 459940 42106 459968 47654
rect 460124 44169 460152 47654
rect 460110 44160 460166 44169
rect 460110 44095 460166 44104
rect 460860 43489 460888 47654
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461964 44441 461992 47654
rect 462378 47410 462406 47668
rect 462332 47382 462406 47410
rect 462516 47654 462852 47682
rect 462976 47654 463312 47682
rect 461950 44432 462006 44441
rect 461950 44367 462006 44376
rect 462332 43217 462360 47382
rect 462516 44441 462544 47654
rect 462502 44432 462558 44441
rect 462502 44367 462558 44376
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 462976 42634 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464356 47654 464692 47682
rect 462964 42628 463016 42634
rect 462964 42570 463016 42576
rect 463712 42498 463740 47382
rect 463896 44169 463924 47654
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 464356 42770 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 626000 46510 626028 66846
rect 647344 64433 647372 80786
rect 648620 79348 648672 79354
rect 648620 79290 648672 79296
rect 647514 78160 647570 78169
rect 647514 78095 647570 78104
rect 647330 64424 647386 64433
rect 647330 64359 647386 64368
rect 647528 57361 647556 78095
rect 648632 59265 648660 79290
rect 648988 76832 649040 76838
rect 648988 76774 649040 76780
rect 649000 62121 649028 76774
rect 662420 76696 662472 76702
rect 662420 76638 662472 76644
rect 648986 62112 649042 62121
rect 648986 62047 649042 62056
rect 648618 59256 648674 59265
rect 648618 59191 648674 59200
rect 647514 57352 647570 57361
rect 647514 57287 647570 57296
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 625988 46504 626040 46510
rect 625988 46446 626040 46452
rect 661604 45554 661632 48445
rect 661774 47789 661830 47798
rect 661774 47724 661830 47733
rect 661788 46510 661816 47724
rect 662432 47433 662460 76638
rect 666572 75206 666600 103486
rect 667938 102776 667994 102785
rect 667938 102711 667994 102720
rect 667952 100026 667980 102711
rect 667940 100020 667992 100026
rect 667940 99962 667992 99968
rect 668136 95962 668164 103486
rect 668044 95946 668164 95962
rect 668032 95940 668164 95946
rect 668084 95934 668164 95940
rect 668032 95882 668084 95888
rect 668228 76566 668256 104343
rect 668596 102785 668624 126919
rect 668766 122632 668822 122641
rect 668766 122567 668822 122576
rect 668780 115934 668808 122567
rect 668964 119241 668992 131135
rect 669962 130928 670018 130937
rect 669962 130863 670018 130872
rect 669226 119640 669282 119649
rect 669226 119575 669282 119584
rect 668950 119232 669006 119241
rect 668950 119167 669006 119176
rect 668780 115906 668992 115934
rect 668964 112713 668992 115906
rect 669240 114345 669268 119575
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 668950 112704 669006 112713
rect 668950 112639 669006 112648
rect 669976 108866 670004 130863
rect 670804 129198 670832 137986
rect 670792 129192 670844 129198
rect 670792 129134 670844 129140
rect 671342 128344 671398 128353
rect 671342 128279 671398 128288
rect 671356 109034 671384 128279
rect 671526 121408 671582 121417
rect 671526 121343 671582 121352
rect 671540 111081 671568 121343
rect 672184 115841 672212 165543
rect 672368 164234 672396 166223
rect 672368 164206 672488 164234
rect 672460 162330 672488 164206
rect 672276 162302 672488 162330
rect 672276 157334 672304 162302
rect 672276 157306 672396 157334
rect 672368 131209 672396 157306
rect 672354 131200 672410 131209
rect 672354 131135 672410 131144
rect 672354 124808 672410 124817
rect 672354 124743 672410 124752
rect 672170 115832 672226 115841
rect 672170 115767 672226 115776
rect 671526 111072 671582 111081
rect 671526 111007 671582 111016
rect 670804 109006 671384 109034
rect 669964 108860 670016 108866
rect 669964 108802 670016 108808
rect 670804 104854 670832 109006
rect 672368 107001 672396 124743
rect 672552 117609 672580 167878
rect 672736 161401 672764 183526
rect 672920 183526 673132 183554
rect 672722 161392 672778 161401
rect 672722 161327 672778 161336
rect 672722 131744 672778 131753
rect 672722 131679 672778 131688
rect 672538 117600 672594 117609
rect 672538 117535 672594 117544
rect 672354 106992 672410 107001
rect 672354 106927 672410 106936
rect 672736 106185 672764 131679
rect 672920 124137 672948 183526
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 673182 168736 673238 168745
rect 673182 168671 673238 168680
rect 673196 151337 673224 168671
rect 673182 151328 673238 151337
rect 673182 151263 673238 151272
rect 673380 129713 673408 174383
rect 673550 168328 673606 168337
rect 673550 168263 673606 168272
rect 673564 166297 673592 168263
rect 673550 166288 673606 166297
rect 673550 166223 673606 166232
rect 673748 153241 673776 229758
rect 674024 229650 674052 244246
rect 674116 243522 674144 259247
rect 674300 243681 674328 262511
rect 674286 243672 674342 243681
rect 674286 243607 674342 243616
rect 674116 243494 674236 243522
rect 674208 242865 674236 243494
rect 674194 242856 674250 242865
rect 674194 242791 674250 242800
rect 674484 235249 674512 264551
rect 674470 235240 674526 235249
rect 674470 235175 674526 235184
rect 674196 234252 674248 234258
rect 674196 234194 674248 234200
rect 674208 232966 674236 234194
rect 674196 232960 674248 232966
rect 674196 232902 674248 232908
rect 674378 230480 674434 230489
rect 674378 230415 674434 230424
rect 674392 230246 674420 230415
rect 674380 230240 674432 230246
rect 674380 230182 674432 230188
rect 674196 230036 674248 230042
rect 674196 229978 674248 229984
rect 673932 229622 674052 229650
rect 673932 222329 673960 229622
rect 674208 226930 674236 229978
rect 674452 229968 674504 229974
rect 674452 229910 674504 229916
rect 674334 229764 674386 229770
rect 674334 229706 674386 229712
rect 674346 229537 674374 229706
rect 674464 229650 674492 229910
rect 674464 229622 674512 229650
rect 674332 229528 674388 229537
rect 674332 229463 674388 229472
rect 674484 229265 674512 229622
rect 674470 229256 674526 229265
rect 674470 229191 674526 229200
rect 674116 226902 674236 226930
rect 673918 222320 673974 222329
rect 673918 222255 673974 222264
rect 673918 220280 673974 220289
rect 673918 220215 673974 220224
rect 673932 175681 673960 220215
rect 674116 213081 674144 226902
rect 674286 226808 674342 226817
rect 674286 226743 674342 226752
rect 674102 213072 674158 213081
rect 674102 213007 674158 213016
rect 674102 209672 674158 209681
rect 674102 209607 674158 209616
rect 673918 175672 673974 175681
rect 673918 175607 673974 175616
rect 673918 170776 673974 170785
rect 673918 170711 673974 170720
rect 673932 156505 673960 170711
rect 673918 156496 673974 156505
rect 673918 156431 673974 156440
rect 673734 153232 673790 153241
rect 673734 153167 673790 153176
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 673366 126576 673422 126585
rect 673366 126511 673422 126520
rect 672906 124128 672962 124137
rect 672906 124063 672962 124072
rect 673182 123992 673238 124001
rect 673182 123927 673238 123936
rect 673196 106321 673224 123927
rect 673380 123298 673408 126511
rect 673288 123270 673408 123298
rect 673288 118694 673316 123270
rect 673458 123176 673514 123185
rect 673458 123111 673514 123120
rect 673472 119649 673500 123111
rect 673918 122224 673974 122233
rect 673918 122159 673974 122168
rect 673458 119640 673514 119649
rect 673458 119575 673514 119584
rect 673288 118666 673408 118694
rect 673182 106312 673238 106321
rect 673182 106247 673238 106256
rect 672722 106176 672778 106185
rect 672722 106111 672778 106120
rect 670792 104848 670844 104854
rect 670792 104790 670844 104796
rect 668582 102776 668638 102785
rect 668582 102711 668638 102720
rect 673380 101017 673408 118666
rect 673932 102150 673960 122159
rect 674116 120465 674144 209607
rect 674300 178129 674328 226743
rect 674668 223689 674696 303447
rect 675128 302234 675156 307935
rect 676232 307834 676260 308366
rect 676220 307828 676272 307834
rect 676220 307770 676272 307776
rect 676864 307828 676916 307834
rect 676864 307770 676916 307776
rect 676034 307592 676090 307601
rect 676090 307550 676260 307578
rect 676034 307527 676090 307536
rect 676034 305960 676090 305969
rect 676034 305895 676090 305904
rect 675852 304564 675904 304570
rect 675852 304506 675904 304512
rect 675128 302206 675248 302234
rect 674838 302016 674894 302025
rect 674838 301951 674894 301960
rect 674852 288062 674880 301951
rect 675220 297242 675248 302206
rect 675864 302025 675892 304506
rect 675850 302016 675906 302025
rect 675850 301951 675906 301960
rect 676048 300665 676076 305895
rect 676232 304570 676260 307550
rect 676220 304564 676272 304570
rect 676220 304506 676272 304512
rect 676034 300656 676090 300665
rect 676034 300591 676090 300600
rect 676876 298110 676904 307770
rect 679622 306776 679678 306785
rect 679622 306711 679678 306720
rect 677598 306368 677654 306377
rect 677598 306303 677654 306312
rect 676128 298104 676180 298110
rect 676128 298046 676180 298052
rect 676864 298104 676916 298110
rect 676864 298046 676916 298052
rect 675944 297696 675996 297702
rect 675944 297638 675996 297644
rect 675956 297401 675984 297638
rect 675942 297392 675998 297401
rect 675942 297327 675998 297336
rect 675036 297214 675248 297242
rect 675852 297220 675904 297226
rect 675036 292414 675064 297214
rect 675852 297162 675904 297168
rect 675864 296585 675892 297162
rect 676140 296585 676168 298046
rect 677612 297702 677640 306303
rect 677600 297696 677652 297702
rect 677600 297638 677652 297644
rect 679636 297226 679664 306711
rect 683026 302696 683082 302705
rect 683026 302631 683082 302640
rect 683040 299441 683068 302631
rect 683026 299432 683082 299441
rect 683026 299367 683082 299376
rect 679624 297220 679676 297226
rect 679624 297162 679676 297168
rect 675206 296576 675262 296585
rect 675206 296511 675262 296520
rect 675850 296576 675906 296585
rect 675850 296511 675906 296520
rect 676126 296576 676182 296585
rect 676126 296511 676182 296520
rect 675220 295338 675248 296511
rect 675404 295769 675432 296072
rect 675390 295760 675446 295769
rect 675390 295695 675446 295704
rect 675758 295760 675814 295769
rect 675758 295695 675814 295704
rect 675772 295528 675800 295695
rect 675220 295310 675432 295338
rect 675404 294879 675432 295310
rect 675758 294536 675814 294545
rect 675758 294471 675814 294480
rect 675772 294236 675800 294471
rect 675036 292386 675418 292414
rect 675574 292224 675630 292233
rect 675574 292159 675630 292168
rect 675588 291856 675616 292159
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675758 290864 675814 290873
rect 675758 290799 675814 290808
rect 675772 290564 675800 290799
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675116 287020 675168 287026
rect 675116 286962 675168 286968
rect 675128 286906 675156 286962
rect 675128 286878 675340 286906
rect 675312 286770 675340 286878
rect 675404 286770 675432 286892
rect 675312 286742 675432 286770
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675666 283656 675722 283665
rect 675666 283591 675722 283600
rect 675680 283220 675708 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675772 281217 675800 281355
rect 675758 281208 675814 281217
rect 675758 281143 675814 281152
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 683132 268569 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268560 683174 268569
rect 683118 268495 683174 268504
rect 675484 266008 675536 266014
rect 675484 265950 675536 265956
rect 675496 265849 675524 265950
rect 675482 265840 675538 265849
rect 675482 265775 675538 265784
rect 681002 263256 681058 263265
rect 681002 263191 681058 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259622 676260 262783
rect 675852 259616 675904 259622
rect 675852 259558 675904 259564
rect 676220 259616 676272 259622
rect 676220 259558 676272 259564
rect 675864 255377 675892 259558
rect 676218 257136 676274 257145
rect 676218 257071 676274 257080
rect 676232 256465 676260 257071
rect 676218 256456 676274 256465
rect 676218 256391 676274 256400
rect 674838 255368 674894 255377
rect 674838 255303 674894 255312
rect 675850 255368 675906 255377
rect 675850 255303 675906 255312
rect 674852 248130 674880 255303
rect 675852 254720 675904 254726
rect 675852 254662 675904 254668
rect 675864 254266 675892 254662
rect 675128 254238 675892 254266
rect 674840 248124 674892 248130
rect 674840 248066 674892 248072
rect 674838 247888 674894 247897
rect 674838 247823 674894 247832
rect 674852 239970 674880 247823
rect 675128 244274 675156 254238
rect 681016 253910 681044 263191
rect 683026 257544 683082 257553
rect 683026 257479 683082 257488
rect 683040 254726 683068 257479
rect 683028 254720 683080 254726
rect 683028 254662 683080 254668
rect 675852 253904 675904 253910
rect 675852 253846 675904 253852
rect 681004 253904 681056 253910
rect 681004 253846 681056 253852
rect 675864 252226 675892 253846
rect 675220 252198 675892 252226
rect 675220 250730 675248 252198
rect 675496 250889 675524 251056
rect 675482 250880 675538 250889
rect 675482 250815 675538 250824
rect 675220 250702 675432 250730
rect 675404 250512 675432 250702
rect 675758 250200 675814 250209
rect 675758 250135 675814 250144
rect 675772 249900 675800 250135
rect 675482 249520 675538 249529
rect 675482 249455 675538 249464
rect 675496 249220 675524 249455
rect 675300 247988 675352 247994
rect 675300 247930 675352 247936
rect 675312 247398 675340 247930
rect 675312 247370 675418 247398
rect 675298 247072 675354 247081
rect 675298 247007 675354 247016
rect 675312 246854 675340 247007
rect 675312 246826 675418 246854
rect 675298 246664 675354 246673
rect 675298 246599 675354 246608
rect 675312 246213 675340 246599
rect 675312 246185 675418 246213
rect 675298 245712 675354 245721
rect 675298 245647 675354 245656
rect 675312 245562 675340 245647
rect 675312 245534 675418 245562
rect 674944 244246 675156 244274
rect 674944 240122 674972 244246
rect 675114 243672 675170 243681
rect 675114 243607 675170 243616
rect 675128 243085 675156 243607
rect 675128 243057 675418 243085
rect 675114 242856 675170 242865
rect 675114 242791 675170 242800
rect 675128 242533 675156 242791
rect 675128 242505 675418 242533
rect 675758 242312 675814 242321
rect 675758 242247 675814 242256
rect 675772 241876 675800 242247
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675114 240272 675170 240281
rect 675114 240207 675170 240216
rect 674944 240094 675064 240122
rect 674840 239964 674892 239970
rect 674840 239906 674892 239912
rect 675036 239850 675064 240094
rect 675128 240054 675156 240207
rect 675128 240026 675418 240054
rect 675208 239964 675260 239970
rect 675208 239906 675260 239912
rect 675036 239822 675156 239850
rect 675128 237538 675156 239822
rect 675220 238218 675248 239906
rect 675220 238190 675418 238218
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 675128 237510 675340 237538
rect 675404 237524 675432 237646
rect 675128 236354 675418 236382
rect 675128 234122 675156 236354
rect 675850 235240 675906 235249
rect 675850 235175 675906 235184
rect 675390 234832 675446 234841
rect 675390 234767 675446 234776
rect 675116 234116 675168 234122
rect 675116 234058 675168 234064
rect 674932 231668 674984 231674
rect 674932 231610 674984 231616
rect 674944 231146 674972 231610
rect 675116 231396 675168 231402
rect 675116 231338 675168 231344
rect 674944 231118 674996 231146
rect 674968 230858 674996 231118
rect 675128 231062 675156 231338
rect 675116 231056 675168 231062
rect 675116 230998 675168 231004
rect 674956 230852 675008 230858
rect 674956 230794 675008 230800
rect 675022 226400 675078 226409
rect 675022 226335 675078 226344
rect 674838 225856 674894 225865
rect 674838 225791 674894 225800
rect 674654 223680 674710 223689
rect 674654 223615 674710 223624
rect 674852 221513 674880 225791
rect 674838 221504 674894 221513
rect 674838 221439 674894 221448
rect 675036 220561 675064 226335
rect 675206 225312 675262 225321
rect 675206 225247 675262 225256
rect 675022 220552 675078 220561
rect 675022 220487 675078 220496
rect 675220 218657 675248 225247
rect 675206 218648 675262 218657
rect 675206 218583 675262 218592
rect 675022 217832 675078 217841
rect 675022 217767 675078 217776
rect 674654 217016 674710 217025
rect 674654 216951 674710 216960
rect 674668 215294 674696 216951
rect 674838 216200 674894 216209
rect 674838 216135 674894 216144
rect 674668 215266 674788 215294
rect 674470 214160 674526 214169
rect 674470 214095 674526 214104
rect 674484 201385 674512 214095
rect 674470 201376 674526 201385
rect 674470 201311 674526 201320
rect 674760 191162 674788 215266
rect 674852 201634 674880 216135
rect 675036 202209 675064 217767
rect 675404 215294 675432 234767
rect 675864 233986 675892 235175
rect 683396 234048 683448 234054
rect 683396 233990 683448 233996
rect 675852 233980 675904 233986
rect 675852 233922 675904 233928
rect 675852 233776 675904 233782
rect 675850 233744 675852 233753
rect 678244 233776 678296 233782
rect 675904 233744 675906 233753
rect 678244 233718 678296 233724
rect 675850 233679 675906 233688
rect 675852 232552 675904 232558
rect 675850 232520 675852 232529
rect 675904 232520 675906 232529
rect 675850 232455 675906 232464
rect 675850 231568 675906 231577
rect 675850 231503 675852 231512
rect 675904 231503 675906 231512
rect 675852 231474 675904 231480
rect 676586 230480 676642 230489
rect 676586 230415 676642 230424
rect 676034 230208 676090 230217
rect 676034 230143 676090 230152
rect 676048 221513 676076 230143
rect 676218 228576 676274 228585
rect 676218 228511 676274 228520
rect 676034 221504 676090 221513
rect 676034 221439 676090 221448
rect 676034 219056 676090 219065
rect 676034 218991 676036 219000
rect 676088 218991 676090 219000
rect 676036 218962 676088 218968
rect 675852 217592 675904 217598
rect 675574 217560 675630 217569
rect 675630 217540 675852 217546
rect 675630 217534 675904 217540
rect 675630 217518 675892 217534
rect 675574 217495 675630 217504
rect 675944 215552 675996 215558
rect 675942 215520 675944 215529
rect 675996 215520 675998 215529
rect 675942 215455 675998 215464
rect 675312 215266 675432 215294
rect 675312 205889 675340 215266
rect 675942 214704 675998 214713
rect 676232 214690 676260 228511
rect 676600 217598 676628 230415
rect 677046 227080 677102 227089
rect 677046 227015 677102 227024
rect 676864 219020 676916 219026
rect 676864 218962 676916 218968
rect 676588 217592 676640 217598
rect 676588 217534 676640 217540
rect 675998 214662 676260 214690
rect 675942 214639 675998 214648
rect 675850 212120 675906 212129
rect 675850 212055 675906 212064
rect 675864 209681 675892 212055
rect 675850 209672 675906 209681
rect 675850 209607 675906 209616
rect 676876 206961 676904 218962
rect 677060 215558 677088 227015
rect 678256 223825 678284 233718
rect 683212 232552 683264 232558
rect 683212 232494 683264 232500
rect 678242 223816 678298 223825
rect 678242 223751 678298 223760
rect 683224 222737 683252 232494
rect 683210 222728 683266 222737
rect 683210 222663 683266 222672
rect 683408 219881 683436 233990
rect 683580 231532 683632 231538
rect 683580 231474 683632 231480
rect 683592 223145 683620 231474
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683578 223136 683634 223145
rect 683578 223071 683634 223080
rect 683394 219872 683450 219881
rect 683394 219807 683450 219816
rect 683302 218648 683358 218657
rect 683302 218583 683358 218592
rect 677048 215552 677100 215558
rect 677048 215494 677100 215500
rect 683118 212936 683174 212945
rect 683118 212871 683174 212880
rect 678978 211440 679034 211449
rect 678978 211375 679034 211384
rect 678992 207641 679020 211375
rect 683132 211206 683160 212871
rect 680360 211200 680412 211206
rect 680360 211142 680412 211148
rect 683120 211200 683172 211206
rect 683120 211142 683172 211148
rect 680372 210633 680400 211142
rect 680358 210624 680414 210633
rect 680358 210559 680414 210568
rect 683316 210361 683344 218583
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 678978 207632 679034 207641
rect 678978 207567 679034 207576
rect 676862 206952 676918 206961
rect 676862 206887 676918 206896
rect 675312 205861 675418 205889
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675220 204666 675418 204694
rect 675220 202881 675248 204666
rect 675758 204232 675814 204241
rect 675758 204167 675814 204176
rect 675772 204035 675800 204167
rect 675206 202872 675262 202881
rect 675206 202807 675262 202816
rect 675036 202181 675418 202209
rect 675312 201742 675432 201770
rect 675312 201634 675340 201742
rect 674852 201606 675340 201634
rect 675404 201620 675432 201742
rect 675298 201376 675354 201385
rect 675298 201311 675354 201320
rect 675114 201104 675170 201113
rect 675114 201039 675170 201048
rect 675128 196670 675156 201039
rect 675312 197282 675340 201311
rect 675496 200841 675524 201008
rect 675482 200832 675538 200841
rect 675482 200767 675538 200776
rect 675758 200832 675814 200841
rect 675758 200767 675814 200776
rect 675772 200328 675800 200767
rect 675758 198384 675814 198393
rect 675758 198319 675814 198328
rect 675772 197880 675800 198319
rect 675404 197282 675432 197336
rect 675312 197254 675432 197282
rect 675312 196710 675432 196738
rect 675312 196670 675340 196710
rect 675128 196642 675340 196670
rect 675404 196656 675432 196710
rect 675114 196072 675170 196081
rect 675170 196030 675418 196058
rect 675114 196007 675170 196016
rect 675298 195936 675354 195945
rect 675298 195871 675354 195880
rect 675312 194834 675340 195871
rect 675312 194806 675418 194834
rect 675114 193216 675170 193225
rect 675114 193151 675170 193160
rect 675128 192998 675156 193151
rect 675128 192970 675418 192998
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 674760 191134 675418 191162
rect 676862 189680 676918 189689
rect 676862 189615 676918 189624
rect 674286 178120 674342 178129
rect 674286 178055 674342 178064
rect 674286 176896 674342 176905
rect 674286 176831 674342 176840
rect 674300 132161 674328 176831
rect 674470 176080 674526 176089
rect 674470 176015 674526 176024
rect 674286 132152 674342 132161
rect 674286 132087 674342 132096
rect 674484 131345 674512 176015
rect 674654 175264 674710 175273
rect 674654 175199 674710 175208
rect 674470 131336 674526 131345
rect 674470 131271 674526 131280
rect 674668 130529 674696 175199
rect 674930 174040 674986 174049
rect 674930 173975 674986 173984
rect 674944 159497 674972 173975
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 675114 169416 675170 169425
rect 675114 169351 675170 169360
rect 675942 169416 675998 169425
rect 676232 169402 676260 173182
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 675998 169374 676260 169402
rect 675942 169351 675998 169360
rect 675128 164234 675156 169351
rect 676034 167104 676090 167113
rect 676034 167039 676090 167048
rect 676048 165617 676076 167039
rect 676600 166433 676628 169895
rect 676876 166433 676904 189615
rect 683118 185600 683174 185609
rect 683118 185535 683174 185544
rect 683132 178809 683160 185535
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 178800 683174 178809
rect 683118 178735 683174 178744
rect 678242 171592 678298 171601
rect 678242 171527 678298 171536
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676862 166424 676918 166433
rect 676862 166359 676918 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 675036 164206 675156 164234
rect 675036 160358 675064 164206
rect 678256 162858 678284 171527
rect 675852 162852 675904 162858
rect 675852 162794 675904 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675864 162738 675892 162794
rect 675680 162710 675892 162738
rect 675482 161392 675538 161401
rect 675482 161327 675538 161336
rect 675496 160888 675524 161327
rect 675680 161265 675708 162710
rect 675666 161256 675722 161265
rect 675666 161191 675722 161200
rect 675036 160330 675340 160358
rect 675312 160290 675340 160330
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675758 160032 675814 160041
rect 675758 159967 675814 159976
rect 675772 159664 675800 159967
rect 674930 159488 674986 159497
rect 674930 159423 674986 159432
rect 675482 159488 675538 159497
rect 675482 159423 675538 159432
rect 675496 159052 675524 159423
rect 675772 157049 675800 157216
rect 675390 157040 675446 157049
rect 675390 156975 675446 156984
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 675404 156643 675432 156975
rect 675114 156496 675170 156505
rect 675114 156431 675170 156440
rect 675128 156006 675156 156431
rect 675128 155978 675418 156006
rect 675758 155816 675814 155825
rect 675758 155751 675814 155760
rect 675772 155380 675800 155751
rect 675666 153096 675722 153105
rect 675666 153031 675722 153040
rect 675680 152864 675708 153031
rect 674944 152306 675418 152334
rect 674944 150113 674972 152306
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675114 151328 675170 151337
rect 675114 151263 675170 151272
rect 675128 151042 675156 151263
rect 675128 151014 675418 151042
rect 675114 150376 675170 150385
rect 675114 150311 675170 150320
rect 674930 150104 674986 150113
rect 674930 150039 674986 150048
rect 675128 149849 675156 150311
rect 675128 149821 675418 149849
rect 675298 149016 675354 149025
rect 675298 148951 675354 148960
rect 675312 146690 675340 148951
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 676034 134600 676090 134609
rect 676034 134535 676090 134544
rect 676048 132569 676076 134535
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676034 132560 676090 132569
rect 676034 132495 676090 132504
rect 674654 130520 674710 130529
rect 674654 130455 674710 130464
rect 675850 130112 675906 130121
rect 675850 130047 675906 130056
rect 674838 127392 674894 127401
rect 674838 127327 674894 127336
rect 674470 124400 674526 124409
rect 674470 124335 674526 124344
rect 674102 120456 674158 120465
rect 674102 120391 674158 120400
rect 674484 110401 674512 124335
rect 674654 123584 674710 123593
rect 674654 123519 674710 123528
rect 674470 110392 674526 110401
rect 674470 110327 674526 110336
rect 674668 105822 674696 123519
rect 674852 112010 674880 127327
rect 675864 126993 675892 130047
rect 676218 129024 676274 129033
rect 676218 128959 676274 128968
rect 676232 128354 676260 128959
rect 676048 128353 676260 128354
rect 676034 128344 676260 128353
rect 676090 128326 676260 128344
rect 676034 128279 676090 128288
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 675850 126984 675906 126993
rect 675850 126919 675906 126928
rect 676232 125882 676260 127735
rect 682382 126168 682438 126177
rect 682382 126103 682438 126112
rect 675312 125854 676260 125882
rect 675312 125594 675340 125854
rect 676218 125760 676274 125769
rect 676218 125695 676274 125704
rect 675312 125566 675432 125594
rect 675114 116784 675170 116793
rect 675114 116719 675170 116728
rect 675128 114493 675156 116719
rect 675404 115934 675432 125566
rect 675942 122904 675998 122913
rect 676232 122890 676260 125695
rect 678978 125352 679034 125361
rect 678978 125287 679034 125296
rect 675998 122862 676260 122890
rect 675942 122839 675998 122848
rect 678992 121281 679020 125287
rect 678978 121272 679034 121281
rect 678978 121207 679034 121216
rect 682396 117298 682424 126103
rect 683118 125760 683174 125769
rect 683118 125695 683174 125704
rect 683132 121689 683160 125695
rect 683302 124944 683358 124953
rect 683302 124879 683358 124888
rect 683118 121680 683174 121689
rect 683118 121615 683174 121624
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 682384 117292 682436 117298
rect 682384 117234 682436 117240
rect 675864 116793 675892 117234
rect 675850 116784 675906 116793
rect 675850 116719 675906 116728
rect 683316 116521 683344 124879
rect 683302 116512 683358 116521
rect 683302 116447 683358 116456
rect 675312 115906 675432 115934
rect 675312 115410 675340 115906
rect 675482 115832 675538 115841
rect 675482 115767 675538 115776
rect 675496 115668 675524 115767
rect 675312 115382 675432 115410
rect 675404 115124 675432 115382
rect 675128 114465 675418 114493
rect 675758 114200 675814 114209
rect 675758 114135 675814 114144
rect 675772 113832 675800 114135
rect 674852 111982 675418 112010
rect 675758 111752 675814 111761
rect 675758 111687 675814 111696
rect 675772 111452 675800 111687
rect 675666 111344 675722 111353
rect 675666 111279 675722 111288
rect 675680 110772 675708 111279
rect 675114 110392 675170 110401
rect 675114 110327 675170 110336
rect 675128 110174 675156 110327
rect 675128 110146 675418 110174
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675390 106992 675446 107001
rect 675390 106927 675446 106936
rect 675404 106488 675432 106927
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 675666 104816 675722 104825
rect 675666 104751 675722 104760
rect 675680 104652 675708 104751
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 673932 102122 675418 102150
rect 673366 101008 673422 101017
rect 673366 100943 673422 100952
rect 675114 101008 675170 101017
rect 675170 100966 675340 100994
rect 675114 100943 675170 100952
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 668216 76560 668268 76566
rect 668216 76502 668268 76508
rect 666560 75200 666612 75206
rect 666560 75142 666612 75148
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661776 46504 661828 46510
rect 661776 46446 661828 46452
rect 661420 45526 661632 45554
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464344 42764 464396 42770
rect 464344 42706 464396 42712
rect 463700 42492 463752 42498
rect 463988 42486 464050 42514
rect 463700 42434 463752 42440
rect 461122 42256 461178 42265
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 461122 42191 461178 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 454684 41880 454736 41886
rect 454684 41822 454736 41828
rect 449164 41744 449216 41750
rect 449164 41686 449216 41692
rect 453580 41744 453632 41750
rect 453580 41686 453632 41692
rect 446218 41576 446274 41585
rect 446218 41511 446274 41520
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 675850 896688 675906 896744
rect 676034 896280 676090 896336
rect 652022 867584 652078 867640
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 651470 862280 651526 862336
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35438 816856 35494 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814408 35862 814464
rect 41326 813592 41382 813648
rect 40958 812776 41014 812832
rect 39302 811552 39358 811608
rect 33046 811144 33102 811200
rect 31022 809920 31078 809976
rect 31758 806676 31814 806712
rect 31758 806656 31760 806676
rect 31760 806656 31812 806676
rect 31812 806656 31814 806676
rect 33782 809512 33838 809568
rect 41142 812368 41198 812424
rect 42154 810736 42210 810792
rect 41970 810328 42026 810384
rect 41786 809240 41842 809296
rect 40682 809104 40738 809160
rect 41786 808696 41842 808752
rect 40958 808288 41014 808344
rect 41142 807880 41198 807936
rect 41326 806248 41382 806304
rect 41970 805568 42026 805624
rect 41786 805160 41842 805216
rect 42154 804888 42210 804944
rect 40682 801488 40738 801544
rect 39854 801252 39856 801272
rect 39856 801252 39908 801272
rect 39908 801252 39910 801272
rect 39854 801216 39910 801252
rect 40682 800808 40738 800864
rect 39302 800536 39358 800592
rect 42982 807472 43038 807528
rect 42154 797272 42210 797328
rect 42706 796864 42762 796920
rect 41786 796184 41842 796240
rect 42062 794416 42118 794472
rect 41786 793056 41842 793112
rect 41786 790608 41842 790664
rect 42338 790200 42394 790256
rect 42062 789792 42118 789848
rect 41786 788704 41842 788760
rect 42706 789792 42762 789848
rect 42522 789384 42578 789440
rect 42246 788160 42302 788216
rect 42706 789112 42762 789168
rect 35806 774696 35862 774752
rect 41050 774696 41106 774752
rect 35438 773880 35494 773936
rect 35806 773472 35862 773528
rect 41326 773472 41382 773528
rect 42062 773472 42118 773528
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 41694 773064 41750 773120
rect 41786 772792 41842 772848
rect 35622 772656 35678 772712
rect 35346 772248 35402 772304
rect 35530 771860 35586 771896
rect 35530 771840 35532 771860
rect 35532 771840 35584 771860
rect 35584 771840 35586 771860
rect 35806 771840 35862 771896
rect 35806 771024 35862 771080
rect 35622 770616 35678 770672
rect 35806 770208 35862 770264
rect 35346 769392 35402 769448
rect 35530 768984 35586 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 39578 768576 39634 768632
rect 35806 768168 35862 768224
rect 33046 767760 33102 767816
rect 35806 767372 35862 767408
rect 35806 767352 35808 767372
rect 35808 767352 35860 767372
rect 35860 767352 35862 767372
rect 35162 766944 35218 767000
rect 35806 766148 35862 766184
rect 35806 766128 35808 766148
rect 35808 766128 35860 766148
rect 35860 766128 35862 766148
rect 35806 765720 35862 765776
rect 35806 764532 35808 764552
rect 35808 764532 35860 764552
rect 35860 764532 35862 764552
rect 35806 764496 35862 764532
rect 35622 764088 35678 764144
rect 35806 763308 35808 763328
rect 35808 763308 35860 763328
rect 35860 763308 35862 763328
rect 35806 763272 35862 763308
rect 35806 762864 35862 762920
rect 40314 770208 40370 770264
rect 39762 764088 39818 764144
rect 36542 759056 36598 759112
rect 41510 764904 41566 764960
rect 41234 764496 41290 764552
rect 40866 763680 40922 763736
rect 41510 763292 41566 763328
rect 41510 763272 41512 763292
rect 41512 763272 41564 763292
rect 41564 763272 41566 763292
rect 41694 761096 41750 761152
rect 42706 768576 42762 768632
rect 42614 761096 42670 761152
rect 41878 758920 41934 758976
rect 42430 758920 42486 758976
rect 40038 757696 40094 757752
rect 40682 757696 40738 757752
rect 38934 757424 38990 757480
rect 41786 757016 41842 757072
rect 41878 755384 41934 755440
rect 42522 755112 42578 755168
rect 42062 752936 42118 752992
rect 42062 751576 42118 751632
rect 42062 751032 42118 751088
rect 41970 750352 42026 750408
rect 42430 749536 42486 749592
rect 42246 749400 42302 749456
rect 43534 797272 43590 797328
rect 43258 764088 43314 764144
rect 43074 763680 43130 763736
rect 42338 745320 42394 745376
rect 42522 745320 42578 745376
rect 42706 744912 42762 744968
rect 42246 730496 42302 730552
rect 40866 728626 40922 728682
rect 41326 728626 41382 728682
rect 41326 727402 41382 727458
rect 41142 726824 41198 726880
rect 39302 726178 39358 726234
rect 35162 724784 35218 724840
rect 31666 724376 31722 724432
rect 32954 723968 33010 724024
rect 31666 718256 31722 718312
rect 33782 723152 33838 723208
rect 41326 726232 41382 726234
rect 41326 726180 41328 726232
rect 41328 726180 41380 726232
rect 41380 726180 41382 726232
rect 41326 726178 41382 726180
rect 41786 725736 41842 725792
rect 41326 725600 41382 725656
rect 41142 725192 41198 725248
rect 41142 720296 41198 720352
rect 41326 719208 41382 719264
rect 39302 716080 39358 716136
rect 40590 715672 40646 715728
rect 40406 715400 40462 715456
rect 41786 722336 41842 722392
rect 41786 718528 41842 718584
rect 43074 729272 43130 729328
rect 42522 719208 42578 719264
rect 41510 714856 41566 714912
rect 42246 715400 42302 715456
rect 41234 714176 41290 714232
rect 41786 712136 41842 712192
rect 42062 710776 42118 710832
rect 42062 708328 42118 708384
rect 42706 715944 42762 716000
rect 42798 714856 42854 714912
rect 42890 710776 42946 710832
rect 41786 707104 41842 707160
rect 41786 704248 41842 704304
rect 42246 701800 42302 701856
rect 41786 700440 41842 700496
rect 42706 702072 42762 702128
rect 42706 688064 42762 688120
rect 41142 686840 41198 686896
rect 40866 686432 40922 686488
rect 41050 685854 41106 685910
rect 41326 685854 41382 685910
rect 40774 684630 40830 684686
rect 41694 684256 41750 684312
rect 41142 683984 41198 684040
rect 41326 683460 41382 683462
rect 41326 683408 41328 683460
rect 41328 683408 41380 683460
rect 41380 683408 41382 683460
rect 41326 683406 41382 683408
rect 40958 682760 41014 682816
rect 35162 681944 35218 682000
rect 32402 681128 32458 681184
rect 33782 680720 33838 680776
rect 41326 682352 41382 682408
rect 42246 681536 42302 681592
rect 41142 679904 41198 679960
rect 41786 678816 41842 678872
rect 41786 678272 41842 678328
rect 40958 677748 41014 677750
rect 40958 677696 40960 677748
rect 40960 677696 41012 677748
rect 41012 677696 41014 677748
rect 40958 677694 41014 677696
rect 39946 677048 40002 677104
rect 32402 672696 32458 672752
rect 37922 671472 37978 671528
rect 39946 672424 40002 672480
rect 38842 670928 38898 670984
rect 43074 677864 43130 677920
rect 41786 669024 41842 669080
rect 42522 670928 42578 670984
rect 42062 666576 42118 666632
rect 42338 666304 42394 666360
rect 41786 665216 41842 665272
rect 41786 664128 41842 664184
rect 42154 662768 42210 662824
rect 41786 658280 41842 658336
rect 41786 657192 41842 657248
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 39578 644680 39634 644736
rect 38566 644272 38622 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35622 642640 35678 642696
rect 35806 642232 35862 642288
rect 40498 643492 40500 643512
rect 40500 643492 40552 643512
rect 40552 643492 40554 643512
rect 40498 643456 40554 643492
rect 35346 641416 35402 641472
rect 35530 641008 35586 641064
rect 35806 641008 35862 641064
rect 39946 640192 40002 640248
rect 35806 639784 35862 639840
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35622 638560 35678 638616
rect 35162 637744 35218 637800
rect 32034 636928 32090 636984
rect 35806 638152 35862 638208
rect 35530 636540 35586 636576
rect 35530 636520 35532 636540
rect 35532 636520 35584 636540
rect 35584 636520 35586 636540
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35806 634480 35862 634536
rect 35806 633256 35862 633312
rect 35162 629856 35218 629912
rect 37738 629584 37794 629640
rect 39118 636520 39174 636576
rect 39946 633664 40002 633720
rect 39762 632168 39818 632224
rect 41878 633868 41934 633924
rect 41418 631352 41474 631408
rect 40406 630672 40462 630728
rect 39118 630400 39174 630456
rect 37922 627680 37978 627736
rect 42522 636520 42578 636576
rect 42338 629584 42394 629640
rect 42062 627680 42118 627736
rect 41786 627408 41842 627464
rect 41786 627136 41842 627192
rect 42430 624688 42486 624744
rect 42062 624416 42118 624472
rect 42062 623736 42118 623792
rect 42062 623328 42118 623384
rect 42062 622104 42118 622160
rect 41786 620744 41842 620800
rect 42246 619792 42302 619848
rect 42706 620744 42762 620800
rect 42338 616256 42394 616312
rect 42062 615712 42118 615768
rect 42522 615984 42578 616040
rect 42706 615712 42762 615768
rect 42522 615440 42578 615496
rect 42890 613944 42946 614000
rect 43442 757424 43498 757480
rect 43442 752936 43498 752992
rect 43626 751576 43682 751632
rect 43442 731312 43498 731368
rect 43626 723560 43682 723616
rect 43442 687248 43498 687304
rect 43626 680312 43682 680368
rect 43442 676640 43498 676696
rect 43258 612176 43314 612232
rect 44270 774696 44326 774752
rect 44914 772792 44970 772848
rect 44546 770208 44602 770264
rect 44178 728048 44234 728104
rect 44362 727640 44418 727696
rect 62210 790472 62266 790528
rect 62118 789148 62120 789168
rect 62120 789148 62172 789168
rect 62172 789148 62174 789168
rect 62118 789112 62174 789148
rect 62118 787344 62174 787400
rect 62762 787072 62818 787128
rect 61382 786120 61438 786176
rect 62118 784896 62174 784952
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 46202 773064 46258 773120
rect 45098 764904 45154 764960
rect 45282 764496 45338 764552
rect 45558 763272 45614 763328
rect 45098 751032 45154 751088
rect 44914 730088 44970 730144
rect 45190 729680 45246 729736
rect 44454 722744 44510 722800
rect 44638 721520 44694 721576
rect 44454 708328 44510 708384
rect 44822 687656 44878 687712
rect 44270 685208 44326 685264
rect 44454 684256 44510 684312
rect 43994 679496 44050 679552
rect 44638 683848 44694 683904
rect 44454 644680 44510 644736
rect 45006 666576 45062 666632
rect 45006 643456 45062 643512
rect 44362 633664 44418 633720
rect 43994 632168 44050 632224
rect 43718 630400 43774 630456
rect 44178 631352 44234 631408
rect 44086 623328 44142 623384
rect 44362 622104 44418 622160
rect 44086 613944 44142 614000
rect 43764 612196 43820 612232
rect 43764 612176 43766 612196
rect 43766 612176 43818 612196
rect 43818 612176 43820 612196
rect 44086 612060 44142 612096
rect 44086 612040 44088 612060
rect 44088 612040 44140 612060
rect 44140 612040 44142 612060
rect 43994 611788 44050 611824
rect 43994 611768 43996 611788
rect 43996 611768 44048 611788
rect 44048 611768 44050 611788
rect 44086 611532 44088 611552
rect 44088 611532 44140 611552
rect 44140 611532 44142 611552
rect 44086 611496 44142 611532
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 35622 595754 35678 595810
rect 33046 595176 33102 595232
rect 31022 594360 31078 594416
rect 33782 593544 33838 593600
rect 38566 601296 38622 601352
rect 39946 600888 40002 600944
rect 44822 630672 44878 630728
rect 45282 640192 45338 640248
rect 45006 600480 45062 600536
rect 45098 600072 45154 600128
rect 44638 598848 44694 598904
rect 44914 598440 44970 598496
rect 42890 597624 42946 597680
rect 42430 596808 42486 596864
rect 41142 596400 41198 596456
rect 39302 594768 39358 594824
rect 41970 595992 42026 596048
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 41786 594224 41842 594280
rect 41694 592864 41750 592920
rect 41694 591232 41750 591288
rect 41050 590688 41106 590744
rect 39578 585792 39634 585848
rect 39302 585112 39358 585168
rect 41050 585384 41106 585440
rect 40222 584840 40278 584896
rect 39946 584568 40002 584624
rect 41970 586064 42026 586120
rect 42154 585812 42210 585848
rect 42154 585792 42156 585812
rect 42156 585792 42208 585812
rect 42208 585792 42210 585812
rect 42246 585384 42302 585440
rect 41786 584296 41842 584352
rect 41786 583888 41842 583944
rect 42614 581576 42670 581632
rect 42338 581168 42394 581224
rect 42062 580624 42118 580680
rect 41786 580216 41842 580272
rect 42154 578856 42210 578912
rect 42062 578040 42118 578096
rect 41786 577768 41842 577824
rect 42246 575728 42302 575784
rect 41786 574640 41842 574696
rect 42614 572736 42670 572792
rect 41970 572192 42026 572248
rect 42062 571512 42118 571568
rect 42430 571376 42486 571432
rect 41786 570152 41842 570208
rect 43074 596944 43130 597000
rect 44362 593136 44418 593192
rect 44178 591912 44234 591968
rect 43350 591504 43406 591560
rect 43626 590280 43682 590336
rect 42246 558048 42302 558104
rect 40038 553352 40094 553408
rect 40866 553352 40922 553408
rect 34426 551928 34482 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 42982 556416 43038 556472
rect 42798 554784 42854 554840
rect 42246 552608 42302 552664
rect 42982 552336 43038 552392
rect 42798 551112 42854 551168
rect 41786 550568 41842 550624
rect 41878 550296 41934 550352
rect 42062 549888 42118 549944
rect 41878 545672 41934 545728
rect 37830 541320 37886 541376
rect 42062 545400 42118 545456
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42246 540640 42302 540696
rect 42522 539552 42578 539608
rect 42614 538056 42670 538112
rect 43074 549480 43130 549536
rect 42430 537376 42486 537432
rect 41786 536968 41842 537024
rect 42246 536424 42302 536480
rect 42062 535608 42118 535664
rect 42706 532752 42762 532808
rect 42614 530712 42670 530768
rect 42430 529488 42486 529544
rect 41878 528944 41934 529000
rect 42246 528944 42302 529000
rect 42614 527176 42670 527232
rect 35806 430072 35862 430128
rect 41970 427080 42026 427136
rect 41326 425992 41382 426048
rect 41142 425584 41198 425640
rect 40958 425176 41014 425232
rect 32034 424360 32090 424416
rect 41878 424224 41934 424280
rect 41142 418784 41198 418840
rect 42798 423544 42854 423600
rect 42522 419872 42578 419928
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 41970 408040 42026 408096
rect 42430 407768 42486 407824
rect 42246 407496 42302 407552
rect 42062 406680 42118 406736
rect 41786 406272 41842 406328
rect 42246 405592 42302 405648
rect 42430 405592 42486 405648
rect 43258 420688 43314 420744
rect 43074 419464 43130 419520
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 41786 400016 41842 400072
rect 41786 398792 41842 398848
rect 42154 395664 42210 395720
rect 41142 387096 41198 387152
rect 40774 385872 40830 385928
rect 41326 386688 41382 386744
rect 41326 385872 41382 385928
rect 41326 382608 41382 382664
rect 40958 381792 41014 381848
rect 41142 381792 41198 381848
rect 40222 381384 40278 381440
rect 40774 381384 40830 381440
rect 35162 380976 35218 381032
rect 33782 379752 33838 379808
rect 33782 371864 33838 371920
rect 37922 380160 37978 380216
rect 35806 376488 35862 376544
rect 35806 374584 35862 374640
rect 41510 379752 41566 379808
rect 37922 372680 37978 372736
rect 41786 368464 41842 368520
rect 42890 379480 42946 379536
rect 42062 366152 42118 366208
rect 42062 364792 42118 364848
rect 42246 364112 42302 364168
rect 41786 363704 41842 363760
rect 42890 366152 42946 366208
rect 42246 362888 42302 362944
rect 42706 363160 42762 363216
rect 42430 361528 42486 361584
rect 41786 360032 41842 360088
rect 41786 359216 41842 359272
rect 41786 358672 41842 358728
rect 41786 356088 41842 356144
rect 42430 354320 42486 354376
rect 43074 353912 43130 353968
rect 42154 353232 42210 353288
rect 44178 581168 44234 581224
rect 44638 580624 44694 580680
rect 44362 578040 44418 578096
rect 44546 556824 44602 556880
rect 44270 556008 44326 556064
rect 43810 548256 43866 548312
rect 43994 547032 44050 547088
rect 43810 355136 43866 355192
rect 43626 354864 43682 354920
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 62762 747632 62818 747688
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 62394 741784 62450 741840
rect 651470 734168 651526 734224
rect 651470 732944 651526 733000
rect 651470 731720 651526 731776
rect 651470 731040 651526 731096
rect 46202 730904 46258 730960
rect 47214 721112 47270 721168
rect 47030 719888 47086 719944
rect 45742 624416 45798 624472
rect 45558 612040 45614 612096
rect 47030 611768 47086 611824
rect 651470 729816 651526 729872
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 62210 701256 62266 701312
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 62762 700848 62818 700904
rect 61382 699624 61438 699680
rect 62118 698164 62120 698184
rect 62120 698164 62172 698184
rect 62172 698164 62174 698184
rect 62118 698128 62174 698164
rect 651470 689424 651526 689480
rect 651654 688744 651710 688800
rect 651470 687384 651526 687440
rect 651470 686704 651526 686760
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 62118 659540 62120 659560
rect 62120 659540 62172 659560
rect 62172 659540 62174 659560
rect 62118 659504 62174 659540
rect 62118 658280 62174 658336
rect 651470 685208 651526 685264
rect 652574 684392 652630 684448
rect 62762 657600 62818 657656
rect 61382 656512 61438 656568
rect 62118 655288 62174 655344
rect 651470 643184 651526 643240
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 61382 613808 61438 613864
rect 62118 612620 62120 612640
rect 62120 612620 62172 612640
rect 62172 612620 62174 612640
rect 62118 612584 62174 612620
rect 652022 641824 652078 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 62946 618024 63002 618080
rect 62762 612040 62818 612096
rect 47214 611496 47270 611552
rect 45282 598032 45338 598088
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 62946 595720 63002 595776
rect 62762 594088 62818 594144
rect 45558 578856 45614 578912
rect 62118 574776 62174 574832
rect 62118 573552 62174 573608
rect 651470 595448 651526 595504
rect 651654 595176 651710 595232
rect 651470 594088 651526 594144
rect 63130 592864 63186 592920
rect 62946 571104 63002 571160
rect 651470 592728 651526 592784
rect 63130 569880 63186 569936
rect 62762 568520 62818 568576
rect 45098 558728 45154 558784
rect 61382 557504 61438 557560
rect 44914 555600 44970 555656
rect 45650 555192 45706 555248
rect 45190 551520 45246 551576
rect 45006 549072 45062 549128
rect 44730 548664 44786 548720
rect 45006 538056 45062 538112
rect 44730 536832 44786 536888
rect 44730 535608 44786 535664
rect 45374 550704 45430 550760
rect 45374 532752 45430 532808
rect 45190 528944 45246 529000
rect 45098 527176 45154 527232
rect 44546 429664 44602 429720
rect 44638 429256 44694 429312
rect 44270 428848 44326 428904
rect 44270 428440 44326 428496
rect 44454 422320 44510 422376
rect 44454 407496 44510 407552
rect 45834 554376 45890 554432
rect 45650 428032 45706 428088
rect 45650 427624 45706 427680
rect 60002 539552 60058 539608
rect 63406 556688 63462 556744
rect 62946 552608 63002 552664
rect 62302 531140 62358 531176
rect 62302 531120 62304 531140
rect 62304 531120 62356 531140
rect 62356 531120 62358 531140
rect 62118 530576 62174 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 61382 527040 61438 527096
rect 651470 553424 651526 553480
rect 651470 552336 651526 552392
rect 651470 551112 651526 551168
rect 651378 550332 651380 550352
rect 651380 550332 651432 550352
rect 651432 550332 651434 550352
rect 651378 550296 651434 550332
rect 651470 549092 651526 549128
rect 651470 549072 651472 549092
rect 651472 549072 651524 549092
rect 651524 549072 651526 549092
rect 651470 548392 651526 548448
rect 63406 527992 63462 528048
rect 62946 525680 63002 525736
rect 667018 595448 667074 595504
rect 668030 689832 668086 689888
rect 667754 649168 667810 649224
rect 668214 686432 668270 686488
rect 668950 736072 669006 736128
rect 668398 640600 668454 640656
rect 669778 685752 669834 685808
rect 670514 733760 670570 733816
rect 670974 734188 671030 734224
rect 670974 734168 670976 734188
rect 670976 734168 671028 734188
rect 671028 734168 671030 734188
rect 670698 689152 670754 689208
rect 669870 641688 669926 641744
rect 669042 608232 669098 608288
rect 668858 593544 668914 593600
rect 667754 561856 667810 561912
rect 668674 555192 668730 555248
rect 670514 647808 670570 647864
rect 670238 625096 670294 625152
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 675850 893832 675906 893888
rect 676034 893016 676090 893072
rect 672354 695408 672410 695464
rect 671802 690376 671858 690432
rect 670974 643456 671030 643512
rect 670974 638696 671030 638752
rect 670422 552064 670478 552120
rect 671158 622648 671214 622704
rect 671342 607280 671398 607336
rect 670974 548392 671030 548448
rect 672170 685344 672226 685400
rect 671986 652160 672042 652216
rect 671802 620200 671858 620256
rect 671802 600616 671858 600672
rect 671526 534112 671582 534168
rect 670054 455368 670110 455424
rect 676034 892608 676090 892664
rect 679622 891792 679678 891848
rect 675850 891384 675906 891440
rect 675666 890976 675722 891032
rect 675482 886916 675538 886952
rect 675482 886896 675484 886916
rect 675484 886896 675536 886916
rect 675536 886896 675538 886916
rect 676034 890568 676090 890624
rect 676034 890160 676090 890216
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 888548 676090 888584
rect 676034 888528 676036 888548
rect 676036 888528 676088 888548
rect 676088 888528 676090 888548
rect 676034 888140 676090 888176
rect 676034 888120 676036 888140
rect 676036 888120 676088 888140
rect 676088 888120 676090 888140
rect 676034 887440 676090 887496
rect 676678 887304 676734 887360
rect 676034 885692 676090 885728
rect 676034 885672 676036 885692
rect 676036 885672 676088 885692
rect 676088 885672 676090 885692
rect 676678 882544 676734 882600
rect 678242 889752 678298 889808
rect 683302 889344 683358 889400
rect 683026 886080 683082 886136
rect 683026 881864 683082 881920
rect 675942 878464 675998 878520
rect 675666 877784 675722 877840
rect 675482 876424 675538 876480
rect 675022 874112 675078 874168
rect 675482 874112 675538 874168
rect 675574 873432 675630 873488
rect 675758 869760 675814 869816
rect 675758 868672 675814 868728
rect 675114 867176 675170 867232
rect 674838 866224 674894 866280
rect 675390 866224 675446 866280
rect 675114 865680 675170 865736
rect 675758 865408 675814 865464
rect 675390 788024 675446 788080
rect 675482 786664 675538 786720
rect 672722 714040 672778 714096
rect 673274 721520 673330 721576
rect 673090 712816 673146 712872
rect 672906 709144 672962 709200
rect 673274 706288 673330 706344
rect 675482 783808 675538 783864
rect 675758 779864 675814 779920
rect 675390 742464 675446 742520
rect 674838 742192 674894 742248
rect 675206 738112 675262 738168
rect 674930 736344 674986 736400
rect 675114 736344 675170 736400
rect 675482 736072 675538 736128
rect 675298 734984 675354 735040
rect 675482 734168 675538 734224
rect 675482 733760 675538 733816
rect 675758 732944 675814 733000
rect 675758 728320 675814 728376
rect 674838 723152 674894 723208
rect 674102 721792 674158 721848
rect 675942 728048 675998 728104
rect 675022 721656 675078 721712
rect 674010 715708 674012 715728
rect 674012 715708 674064 715728
rect 674064 715708 674066 715728
rect 674010 715672 674066 715708
rect 674010 715300 674012 715320
rect 674012 715300 674064 715320
rect 674064 715300 674066 715320
rect 674010 715264 674066 715300
rect 674010 715012 674066 715048
rect 674010 714992 674012 715012
rect 674012 714992 674064 715012
rect 674064 714992 674066 715012
rect 674010 714484 674012 714504
rect 674012 714484 674064 714504
rect 674064 714484 674066 714504
rect 674010 714448 674066 714484
rect 674010 713668 674012 713688
rect 674012 713668 674064 713688
rect 674064 713668 674066 713688
rect 674010 713632 674066 713668
rect 674010 713244 674066 713280
rect 674010 713224 674012 713244
rect 674012 713224 674064 713244
rect 674064 713224 674066 713244
rect 674010 712428 674066 712464
rect 674010 712408 674012 712428
rect 674012 712408 674064 712428
rect 674064 712408 674066 712428
rect 674010 709996 674012 710016
rect 674012 709996 674064 710016
rect 674064 709996 674066 710016
rect 674010 709960 674066 709996
rect 674010 709588 674012 709608
rect 674012 709588 674064 709608
rect 674064 709588 674066 709608
rect 674010 709552 674066 709588
rect 675666 712000 675722 712056
rect 676034 716508 676090 716544
rect 676034 716488 676036 716508
rect 676036 716488 676088 716508
rect 676088 716488 676090 716508
rect 676034 716080 676090 716136
rect 675850 711184 675906 711240
rect 676034 710776 676090 710832
rect 683302 711592 683358 711648
rect 676034 710368 676090 710424
rect 684130 726416 684186 726472
rect 684130 708736 684186 708792
rect 683486 708328 683542 708384
rect 676034 707548 676036 707568
rect 676036 707548 676088 707568
rect 676088 707548 676090 707568
rect 676034 707512 676090 707548
rect 676034 707140 676036 707160
rect 676036 707140 676088 707160
rect 676088 707140 676090 707160
rect 676034 707104 676090 707140
rect 675850 706696 675906 706752
rect 683118 705472 683174 705528
rect 676034 705064 676090 705120
rect 673182 697176 673238 697232
rect 672906 687792 672962 687848
rect 672722 669432 672778 669488
rect 672722 651344 672778 651400
rect 672354 603744 672410 603800
rect 672538 597352 672594 597408
rect 673182 619384 673238 619440
rect 672906 618160 672962 618216
rect 673090 604152 673146 604208
rect 672722 576544 672778 576600
rect 672906 553288 672962 553344
rect 672722 534964 672724 534984
rect 672724 534964 672776 534984
rect 672776 534964 672778 534984
rect 672722 534928 672778 534964
rect 672722 533432 672778 533488
rect 672722 490048 672778 490104
rect 672630 489640 672686 489696
rect 672446 453908 672448 453928
rect 672448 453908 672500 453928
rect 672500 453908 672502 453928
rect 672446 453872 672502 453908
rect 60002 430616 60058 430672
rect 45834 427352 45890 427408
rect 45558 426808 45614 426864
rect 44914 423136 44970 423192
rect 45098 421504 45154 421560
rect 45282 421096 45338 421152
rect 45282 408040 45338 408096
rect 45098 406680 45154 406736
rect 45282 405592 45338 405648
rect 44914 402872 44970 402928
rect 44638 386416 44694 386472
rect 44270 385600 44326 385656
rect 45098 385192 45154 385248
rect 44362 379072 44418 379128
rect 44178 376216 44234 376272
rect 44546 378664 44602 378720
rect 44362 364112 44418 364168
rect 44730 377848 44786 377904
rect 44914 377440 44970 377496
rect 44730 364792 44786 364848
rect 46018 423952 46074 424008
rect 53838 407768 53894 407824
rect 46018 400152 46074 400208
rect 61382 429256 61438 429312
rect 63130 427080 63186 427136
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400560 62174 400616
rect 657542 403280 657598 403336
rect 652022 400832 652078 400888
rect 63130 400152 63186 400208
rect 62118 399336 62174 399392
rect 61382 398248 61438 398304
rect 51078 395664 51134 395720
rect 61382 386416 61438 386472
rect 45834 384784 45890 384840
rect 46018 384376 46074 384432
rect 45558 383968 45614 384024
rect 45650 383560 45706 383616
rect 45282 381384 45338 381440
rect 44546 361528 44602 361584
rect 44822 355136 44878 355192
rect 44638 354864 44694 354920
rect 43258 353640 43314 353696
rect 42338 352960 42394 353016
rect 35806 344256 35862 344312
rect 35622 343848 35678 343904
rect 35806 343440 35862 343496
rect 40406 343848 40462 343904
rect 35806 341808 35862 341864
rect 39670 341808 39726 341864
rect 39854 341808 39910 341864
rect 35806 341028 35808 341048
rect 35808 341028 35860 341048
rect 35860 341028 35862 341048
rect 35806 340992 35862 341028
rect 40222 342236 40278 342272
rect 40222 342216 40224 342236
rect 40224 342216 40276 342236
rect 40276 342216 40278 342236
rect 45374 362888 45430 362944
rect 45190 343304 45246 343360
rect 45006 342488 45062 342544
rect 45466 342236 45522 342272
rect 45466 342216 45468 342236
rect 45468 342216 45520 342236
rect 45520 342216 45522 342236
rect 42246 341264 42302 341320
rect 40130 341028 40132 341048
rect 40132 341028 40184 341048
rect 40184 341028 40186 341048
rect 40130 340992 40186 341028
rect 45834 353932 45890 353968
rect 45834 353912 45836 353932
rect 45836 353912 45888 353932
rect 45888 353912 45890 353932
rect 45834 353676 45836 353696
rect 45836 353676 45888 353696
rect 45888 353676 45890 353696
rect 45834 353640 45890 353676
rect 47122 383152 47178 383208
rect 46938 382336 46994 382392
rect 46570 363160 46626 363216
rect 47122 354320 47178 354376
rect 63406 385872 63462 385928
rect 62946 381792 63002 381848
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62118 357720 62174 357776
rect 61382 355952 61438 356008
rect 651470 373224 651526 373280
rect 652206 395256 652262 395312
rect 654782 382880 654838 382936
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 673090 528808 673146 528864
rect 672906 482296 672962 482352
rect 673734 696940 673736 696960
rect 673736 696940 673788 696960
rect 673788 696940 673790 696960
rect 673734 696904 673790 696940
rect 673734 690124 673790 690160
rect 673734 690104 673736 690124
rect 673736 690104 673788 690124
rect 673788 690104 673790 690124
rect 673734 688780 673736 688800
rect 673736 688780 673788 688800
rect 673788 688780 673790 688800
rect 673734 688744 673790 688780
rect 673734 688064 673790 688120
rect 673550 687520 673606 687576
rect 673550 671336 673606 671392
rect 673550 670520 673606 670576
rect 673550 668888 673606 668944
rect 673550 667256 673606 667312
rect 673550 666304 673606 666360
rect 673550 625948 673552 625968
rect 673552 625948 673604 625968
rect 673604 625948 673606 625968
rect 673550 625912 673606 625948
rect 675114 697176 675170 697232
rect 675298 696904 675354 696960
rect 675114 696632 675170 696688
rect 675298 695408 675354 695464
rect 674102 689424 674158 689480
rect 673918 671608 673974 671664
rect 673918 670928 673974 670984
rect 673918 670132 673974 670168
rect 673918 670112 673920 670132
rect 673920 670112 673972 670132
rect 673972 670112 673974 670132
rect 673918 669704 673974 669760
rect 673918 668516 673920 668536
rect 673920 668516 673972 668536
rect 673972 668516 673974 668536
rect 673918 668480 673974 668516
rect 673918 668072 673974 668128
rect 673918 667664 673974 667720
rect 673918 666052 673974 666088
rect 673918 666032 673920 666052
rect 673920 666032 673972 666052
rect 673972 666032 673974 666052
rect 673918 665236 673974 665272
rect 673918 665216 673920 665236
rect 673920 665216 673972 665236
rect 673972 665216 673974 665236
rect 673918 664808 673974 664864
rect 673918 664012 673974 664048
rect 673918 663992 673920 664012
rect 673920 663992 673972 664012
rect 673972 663992 673974 664012
rect 673918 661972 673974 662008
rect 673918 661952 673920 661972
rect 673920 661952 673972 661972
rect 673972 661952 673974 661972
rect 673918 661580 673920 661600
rect 673920 661580 673972 661600
rect 673972 661580 673974 661600
rect 673918 661544 673974 661580
rect 673918 661156 673974 661192
rect 673918 661136 673920 661156
rect 673920 661136 673972 661156
rect 673972 661136 673974 661156
rect 673918 660204 673974 660240
rect 673918 660184 673920 660204
rect 673920 660184 673972 660204
rect 673972 660184 673974 660204
rect 673918 659912 673974 659968
rect 673918 655580 673974 655616
rect 673918 655560 673920 655580
rect 673920 655560 673972 655580
rect 673972 655560 673974 655580
rect 674286 688064 674342 688120
rect 675114 690376 675170 690432
rect 674930 690104 674986 690160
rect 675390 689832 675446 689888
rect 675114 689424 675170 689480
rect 675114 689152 675170 689208
rect 674930 688744 674986 688800
rect 674654 687520 674710 687576
rect 675114 687792 675170 687848
rect 675482 686432 675538 686488
rect 674930 686160 674986 686216
rect 675482 685616 675538 685672
rect 675114 685344 675170 685400
rect 674010 648352 674066 648408
rect 673642 620608 673698 620664
rect 673550 617344 673606 617400
rect 674010 647284 674066 647320
rect 674010 647264 674012 647284
rect 674012 647264 674064 647284
rect 674064 647264 674066 647284
rect 674102 644272 674158 644328
rect 674010 643084 674012 643104
rect 674012 643084 674064 643104
rect 674064 643084 674066 643104
rect 674010 643048 674066 643084
rect 674746 671608 674802 671664
rect 681002 678952 681058 679008
rect 675298 666848 675354 666904
rect 681002 665760 681058 665816
rect 674930 664012 674986 664048
rect 674930 663992 674932 664012
rect 674932 663992 674984 664012
rect 674984 663992 674986 664012
rect 676218 663720 676274 663776
rect 674746 663448 674802 663504
rect 683210 662904 683266 662960
rect 674562 660184 674618 660240
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 675114 652160 675170 652216
rect 675114 651344 675170 651400
rect 674746 644816 674802 644872
rect 675390 649168 675446 649224
rect 675390 648352 675446 648408
rect 675390 647808 675446 647864
rect 675114 647264 675170 647320
rect 675298 644272 675354 644328
rect 674010 626320 674066 626376
rect 674010 625504 674066 625560
rect 674010 624708 674066 624744
rect 674010 624688 674012 624708
rect 674012 624688 674064 624708
rect 674064 624688 674066 624708
rect 674010 624316 674012 624336
rect 674012 624316 674064 624336
rect 674064 624316 674066 624336
rect 674010 624280 674066 624316
rect 674010 623892 674066 623928
rect 674010 623872 674012 623892
rect 674012 623872 674064 623892
rect 674064 623872 674066 623892
rect 674010 623500 674012 623520
rect 674012 623500 674064 623520
rect 674064 623500 674066 623520
rect 674010 623464 674066 623500
rect 674010 623076 674066 623112
rect 674010 623056 674012 623076
rect 674012 623056 674064 623076
rect 674064 623056 674066 623076
rect 674010 622260 674066 622296
rect 674010 622240 674012 622260
rect 674012 622240 674064 622260
rect 674064 622240 674066 622260
rect 674010 621424 674066 621480
rect 674010 621052 674012 621072
rect 674012 621052 674064 621072
rect 674064 621052 674066 621072
rect 674010 621016 674066 621052
rect 674010 619792 674066 619848
rect 674010 619012 674012 619032
rect 674012 619012 674064 619032
rect 674064 619012 674066 619032
rect 674010 618976 674066 619012
rect 674194 618568 674250 618624
rect 674010 616956 674066 616992
rect 674010 616936 674012 616956
rect 674012 616936 674064 616956
rect 674064 616936 674066 616956
rect 674010 616564 674012 616584
rect 674012 616564 674064 616584
rect 674064 616564 674066 616584
rect 674010 616528 674066 616564
rect 674010 615476 674012 615496
rect 674012 615476 674064 615496
rect 674064 615476 674066 615496
rect 674010 615440 674066 615476
rect 674010 614916 674066 614952
rect 674010 614896 674012 614916
rect 674012 614896 674064 614916
rect 674064 614896 674066 614916
rect 674010 611380 674066 611416
rect 674010 611360 674012 611380
rect 674012 611360 674064 611380
rect 674064 611360 674066 611380
rect 673826 600364 673882 600400
rect 673826 600344 673828 600364
rect 673828 600344 673880 600364
rect 673880 600344 673882 600364
rect 673642 599800 673698 599856
rect 673826 599428 673828 599448
rect 673828 599428 673880 599448
rect 673880 599428 673882 599448
rect 673826 599392 673882 599428
rect 673826 599120 673882 599176
rect 674194 598576 674250 598632
rect 674010 591368 674066 591424
rect 674010 581052 674066 581088
rect 674010 581032 674012 581052
rect 674012 581032 674064 581052
rect 674064 581032 674066 581052
rect 675114 643048 675170 643104
rect 675482 643456 675538 643512
rect 675298 641688 675354 641744
rect 675390 640600 675446 640656
rect 674930 631352 674986 631408
rect 675298 640328 675354 640384
rect 675482 638696 675538 638752
rect 675022 629720 675078 629776
rect 674930 625912 674986 625968
rect 676494 625676 676496 625696
rect 676496 625676 676548 625696
rect 676548 625676 676550 625696
rect 676494 625640 676550 625676
rect 683946 636792 684002 636848
rect 683946 621968 684002 622024
rect 683302 617888 683358 617944
rect 675114 615476 675116 615496
rect 675116 615476 675168 615496
rect 675168 615476 675170 615496
rect 675114 615440 675170 615476
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 683118 615440 683174 615476
rect 675114 611360 675170 611416
rect 675114 608232 675170 608288
rect 675114 607280 675170 607336
rect 674838 604696 674894 604752
rect 675390 604152 675446 604208
rect 675114 603744 675170 603800
rect 675114 602928 675170 602984
rect 675114 600616 675170 600672
rect 675298 600344 675354 600400
rect 675114 599392 675170 599448
rect 675482 599800 675538 599856
rect 675482 599120 675538 599176
rect 675482 598576 675538 598632
rect 675390 597352 675446 597408
rect 675390 595448 675446 595504
rect 674010 580252 674012 580272
rect 674012 580252 674064 580272
rect 674064 580252 674066 580272
rect 674010 580216 674066 580252
rect 674010 579028 674012 579048
rect 674012 579028 674064 579048
rect 674064 579028 674066 579048
rect 674010 578992 674066 579028
rect 675390 593544 675446 593600
rect 676034 592864 676090 592920
rect 675482 591404 675484 591424
rect 675484 591404 675536 591424
rect 675536 591404 675538 591424
rect 675482 591368 675538 591404
rect 674930 584568 674986 584624
rect 674010 576972 674066 577008
rect 674010 576952 674012 576972
rect 674012 576952 674064 576972
rect 674064 576952 674066 576972
rect 674010 574540 674012 574560
rect 674012 574540 674064 574560
rect 674064 574540 674066 574560
rect 674010 574504 674066 574540
rect 674010 574268 674012 574288
rect 674012 574268 674064 574288
rect 674064 574268 674066 574288
rect 674010 574232 674066 574268
rect 674010 573044 674012 573064
rect 674012 573044 674064 573064
rect 674064 573044 674066 573064
rect 674010 573008 674066 573044
rect 674838 571240 674894 571296
rect 673826 565836 673828 565856
rect 673828 565836 673880 565856
rect 673880 565836 673882 565856
rect 673826 565800 673882 565836
rect 673826 554804 673882 554840
rect 673826 554784 673828 554804
rect 673828 554784 673880 554804
rect 673880 554784 673882 554804
rect 673826 553716 673882 553752
rect 673826 553696 673828 553716
rect 673828 553696 673880 553716
rect 673880 553696 673882 553716
rect 675298 586200 675354 586256
rect 675850 577360 675906 577416
rect 682382 590552 682438 590608
rect 676218 580488 676274 580544
rect 676402 580080 676458 580136
rect 676218 579284 676274 579320
rect 676218 579264 676220 579284
rect 676220 579264 676272 579284
rect 676272 579264 676274 579284
rect 676218 578468 676274 578504
rect 676218 578448 676220 578468
rect 676220 578448 676272 578468
rect 676272 578448 676274 578468
rect 676218 578076 676220 578096
rect 676220 578076 676272 578096
rect 676272 578076 676274 578096
rect 676218 578040 676274 578076
rect 676218 577652 676274 577688
rect 676218 577632 676220 577652
rect 676220 577632 676272 577652
rect 676272 577632 676274 577652
rect 676218 576020 676274 576056
rect 676218 576000 676220 576020
rect 676220 576000 676272 576020
rect 676272 576000 676274 576020
rect 682382 576000 682438 576056
rect 676034 575456 676090 575512
rect 676218 574776 676274 574832
rect 676218 573552 676274 573608
rect 683210 573552 683266 573608
rect 683394 572736 683450 572792
rect 676218 571940 676274 571976
rect 676218 571920 676220 571940
rect 676220 571920 676272 571940
rect 676272 571920 676274 571940
rect 675482 571648 675538 571704
rect 676218 570696 676274 570752
rect 676218 569472 676274 569528
rect 675390 565800 675446 565856
rect 675390 563080 675446 563136
rect 674010 547848 674066 547904
rect 674010 547576 674066 547632
rect 674194 536016 674250 536072
rect 674010 535644 674012 535664
rect 674012 535644 674064 535664
rect 674064 535644 674066 535664
rect 674010 535608 674066 535644
rect 674010 535200 674066 535256
rect 674194 534384 674250 534440
rect 674010 533160 674066 533216
rect 674010 532772 674066 532808
rect 674010 532752 674012 532772
rect 674012 532752 674064 532772
rect 674064 532752 674066 532772
rect 674010 532344 674066 532400
rect 674194 531936 674250 531992
rect 674010 531120 674066 531176
rect 674194 530712 674250 530768
rect 674010 530032 674066 530088
rect 674194 529488 674250 529544
rect 674010 529080 674066 529136
rect 673642 528128 673698 528184
rect 673550 526768 673606 526824
rect 674010 527856 674066 527912
rect 673826 492088 673882 492144
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 673918 489268 673920 489288
rect 673920 489268 673972 489288
rect 673972 489268 673974 489288
rect 673918 489232 673974 489268
rect 673918 488452 673920 488472
rect 673920 488452 673972 488472
rect 673972 488452 673974 488472
rect 673918 488416 673974 488452
rect 673918 485968 673974 486024
rect 674010 485596 674012 485616
rect 674012 485596 674064 485616
rect 674064 485596 674066 485616
rect 674010 485560 674066 485596
rect 674010 485152 674066 485208
rect 674194 484336 674250 484392
rect 674010 483964 674012 483984
rect 674012 483964 674064 483984
rect 674064 483964 674066 483984
rect 674010 483928 674066 483964
rect 675114 561856 675170 561912
rect 675114 559000 675170 559056
rect 675390 555192 675446 555248
rect 675298 554784 675354 554840
rect 675114 553696 675170 553752
rect 675758 553968 675814 554024
rect 675390 553288 675446 553344
rect 675298 552064 675354 552120
rect 675758 550296 675814 550352
rect 675482 548392 675538 548448
rect 675482 547848 675538 547904
rect 675666 547576 675722 547632
rect 678242 547576 678298 547632
rect 675574 545536 675630 545592
rect 674654 483112 674710 483168
rect 674470 482704 674526 482760
rect 683486 547032 683542 547088
rect 682382 546760 682438 546816
rect 678242 531800 678298 531856
rect 682382 530576 682438 530632
rect 684314 527720 684370 527776
rect 683486 527312 683542 527368
rect 683302 526496 683358 526552
rect 683302 525680 683358 525736
rect 683118 525272 683174 525328
rect 677874 524456 677930 524512
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 673090 454960 673146 455016
rect 674286 454996 674288 455016
rect 674288 454996 674340 455016
rect 674340 454996 674342 455016
rect 674286 454960 674342 454996
rect 672906 454708 672962 454744
rect 672906 454688 672908 454708
rect 672908 454688 672960 454708
rect 672960 454688 672962 454708
rect 674286 454724 674288 454744
rect 674288 454724 674340 454744
rect 674340 454724 674342 454744
rect 674286 454688 674342 454724
rect 672814 454436 672870 454472
rect 672814 454416 672816 454436
rect 672816 454416 672868 454436
rect 672868 454416 672870 454436
rect 674286 454452 674288 454472
rect 674288 454452 674340 454472
rect 674340 454452 674342 454472
rect 674286 454416 674342 454452
rect 676034 491700 676090 491736
rect 676034 491680 676036 491700
rect 676036 491680 676088 491700
rect 676088 491680 676090 491700
rect 675850 491272 675906 491328
rect 675850 490456 675906 490512
rect 676034 487600 676090 487656
rect 675666 480664 675722 480720
rect 675298 453872 675354 453928
rect 683578 503648 683634 503704
rect 678242 486784 678298 486840
rect 683578 487192 683634 487248
rect 683210 486376 683266 486432
rect 680358 481888 680414 481944
rect 683118 481072 683174 481128
rect 675942 447752 675998 447808
rect 676034 410488 676090 410544
rect 673182 402056 673238 402112
rect 672630 401648 672686 401704
rect 672906 401240 672962 401296
rect 671986 397160 672042 397216
rect 669226 393760 669282 393816
rect 651470 370640 651526 370696
rect 654782 358536 654838 358592
rect 63406 357312 63462 357368
rect 652022 356632 652078 356688
rect 62946 354456 63002 354512
rect 51722 353232 51778 353288
rect 46938 352960 46994 353016
rect 46018 343848 46074 343904
rect 62946 341672 63002 341728
rect 62762 341400 62818 341456
rect 45650 340720 45706 340776
rect 39670 340176 39726 340232
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 37094 336504 37150 336560
rect 46938 339224 46994 339280
rect 45558 338816 45614 338872
rect 45374 337864 45430 337920
rect 35806 335688 35862 335744
rect 38842 335688 38898 335744
rect 35806 334464 35862 334520
rect 44178 334600 44234 334656
rect 44362 334600 44418 334656
rect 40314 332832 40370 332888
rect 42890 332832 42946 332888
rect 39854 332424 39910 332480
rect 42430 326984 42486 327040
rect 41786 325352 41842 325408
rect 41786 324808 41842 324864
rect 42062 322768 42118 322824
rect 42062 321136 42118 321192
rect 42154 320456 42210 320512
rect 41878 319912 41934 319968
rect 42062 319912 42118 319968
rect 43074 332424 43130 332480
rect 42890 321136 42946 321192
rect 42614 320728 42670 320784
rect 43074 320456 43130 320512
rect 45282 326984 45338 327040
rect 44362 322768 44418 322824
rect 44178 319912 44234 319968
rect 42430 319368 42486 319424
rect 42246 318960 42302 319016
rect 41786 317328 41842 317384
rect 42154 315968 42210 316024
rect 42154 315424 42210 315480
rect 45558 315424 45614 315480
rect 42062 313656 42118 313712
rect 42430 312704 42486 312760
rect 51722 334056 51778 334112
rect 50342 333104 50398 333160
rect 42430 310392 42486 310448
rect 46938 310392 46994 310448
rect 42062 309032 42118 309088
rect 35622 300872 35678 300928
rect 46202 300464 46258 300520
rect 44362 299648 44418 299704
rect 35806 298832 35862 298888
rect 41786 298696 41842 298752
rect 44178 297200 44234 297256
rect 41786 296520 41842 296576
rect 42798 296520 42854 296576
rect 35438 296384 35494 296440
rect 35622 295976 35678 296032
rect 35806 295604 35808 295624
rect 35808 295604 35860 295624
rect 35860 295604 35862 295624
rect 35806 295568 35862 295604
rect 35806 295160 35862 295216
rect 33782 294752 33838 294808
rect 32402 294344 32458 294400
rect 35806 293120 35862 293176
rect 35806 292712 35862 292768
rect 35806 291080 35862 291136
rect 35622 290264 35678 290320
rect 39210 288904 39266 288960
rect 32402 284824 32458 284880
rect 41786 295296 41842 295352
rect 42246 291896 42302 291952
rect 41786 291080 41842 291136
rect 42246 289176 42302 289232
rect 40682 284280 40738 284336
rect 41786 278432 41842 278488
rect 42062 277752 42118 277808
rect 42430 278704 42486 278760
rect 41786 277072 41842 277128
rect 42614 275848 42670 275904
rect 41786 274216 41842 274272
rect 42338 273128 42394 273184
rect 42430 272856 42486 272912
rect 41970 272312 42026 272368
rect 41786 270408 41842 270464
rect 41878 270000 41934 270056
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 42154 266192 42210 266248
rect 43166 295296 43222 295352
rect 42982 291080 43038 291136
rect 43626 288904 43682 288960
rect 35806 255856 35862 255912
rect 39762 255856 39818 255912
rect 42798 255856 42854 255912
rect 35806 253816 35862 253872
rect 35622 253408 35678 253464
rect 43626 277752 43682 277808
rect 44822 298016 44878 298072
rect 44546 293528 44602 293584
rect 44546 273128 44602 273184
rect 44362 256808 44418 256864
rect 44638 256400 44694 256456
rect 44270 254768 44326 254824
rect 44086 254496 44142 254552
rect 35806 253000 35862 253056
rect 39210 253000 39266 253056
rect 42798 253000 42854 253056
rect 35806 252184 35862 252240
rect 40314 252184 40370 252240
rect 35806 250552 35862 250608
rect 35806 249328 35862 249384
rect 39670 249328 39726 249384
rect 35622 247696 35678 247752
rect 41510 247696 41566 247752
rect 35806 246880 35862 246936
rect 39854 245520 39910 245576
rect 42062 240080 42118 240136
rect 42430 237360 42486 237416
rect 41786 236544 41842 236600
rect 42430 235864 42486 235920
rect 42430 234504 42486 234560
rect 42154 233280 42210 233336
rect 42430 232600 42486 232656
rect 42430 231784 42486 231840
rect 41786 230424 41842 230480
rect 41970 228928 42026 228984
rect 42246 226072 42302 226128
rect 42614 225528 42670 225584
rect 42430 224848 42486 224904
rect 42154 223488 42210 223544
rect 35806 217912 35862 217968
rect 35806 214648 35862 214704
rect 35806 214240 35862 214296
rect 35438 212200 35494 212256
rect 42982 252184 43038 252240
rect 43074 249328 43130 249384
rect 35622 211792 35678 211848
rect 39578 211792 39634 211848
rect 42798 211792 42854 211848
rect 35806 211384 35862 211440
rect 35806 210160 35862 210216
rect 35622 208936 35678 208992
rect 35806 208548 35862 208584
rect 35806 208528 35808 208548
rect 35808 208528 35860 208548
rect 35860 208528 35862 208548
rect 40038 208120 40094 208176
rect 35806 207712 35862 207768
rect 35806 206080 35862 206136
rect 40682 206896 40738 206952
rect 41694 207712 41750 207768
rect 42890 206896 42946 206952
rect 41326 206488 41382 206544
rect 41142 206080 41198 206136
rect 40314 205672 40370 205728
rect 35806 204856 35862 204912
rect 35806 204448 35862 204504
rect 28538 203632 28594 203688
rect 41694 204484 41696 204504
rect 41696 204484 41748 204504
rect 41748 204484 41750 204504
rect 41694 204448 41750 204484
rect 41694 204040 41750 204096
rect 40682 203224 40738 203280
rect 28538 199280 28594 199336
rect 42246 199280 42302 199336
rect 42062 196968 42118 197024
rect 41878 195200 41934 195256
rect 42246 194928 42302 194984
rect 41786 193160 41842 193216
rect 42062 191528 42118 191584
rect 42430 190440 42486 190496
rect 43166 206080 43222 206136
rect 43074 203224 43130 203280
rect 42430 186768 42486 186824
rect 41786 186360 41842 186416
rect 41786 185952 41842 186008
rect 41786 184048 41842 184104
rect 42430 180648 42486 180704
rect 42062 179288 42118 179344
rect 43810 247696 43866 247752
rect 43626 245520 43682 245576
rect 43810 234504 43866 234560
rect 44454 251912 44510 251968
rect 44454 233280 44510 233336
rect 45006 293936 45062 293992
rect 48962 289856 49018 289912
rect 45006 272856 45062 272912
rect 46202 258032 46258 258088
rect 45558 255584 45614 255640
rect 44822 255176 44878 255232
rect 44822 252728 44878 252784
rect 45190 251504 45246 251560
rect 45006 249056 45062 249112
rect 45190 240080 45246 240136
rect 45006 231784 45062 231840
rect 44822 226072 44878 226128
rect 44638 213696 44694 213752
rect 45926 251096 45982 251152
rect 45742 248648 45798 248704
rect 45742 232600 45798 232656
rect 46110 248240 46166 248296
rect 47582 246608 47638 246664
rect 46110 235864 46166 235920
rect 45926 224848 45982 224904
rect 45558 212880 45614 212936
rect 44270 212064 44326 212120
rect 46938 209616 46994 209672
rect 44362 208392 44418 208448
rect 44178 207168 44234 207224
rect 43994 204448 44050 204504
rect 43810 204040 43866 204096
rect 43994 191528 44050 191584
rect 44638 205264 44694 205320
rect 44362 196968 44418 197024
rect 44822 204720 44878 204776
rect 44638 190440 44694 190496
rect 44178 186768 44234 186824
rect 46202 203496 46258 203552
rect 46938 180648 46994 180704
rect 47766 214920 47822 214976
rect 47766 213288 47822 213344
rect 47950 210840 48006 210896
rect 48778 206488 48834 206544
rect 48318 194384 48374 194440
rect 48778 192344 48834 192400
rect 47766 190440 47822 190496
rect 49146 247424 49202 247480
rect 49514 207712 49570 207768
rect 49514 196424 49570 196480
rect 50526 290672 50582 290728
rect 50710 179288 50766 179344
rect 53838 320728 53894 320784
rect 53102 319368 53158 319424
rect 62118 317364 62120 317384
rect 62120 317364 62172 317384
rect 62172 317364 62174 317384
rect 62118 317328 62174 317364
rect 62118 315988 62174 316024
rect 62118 315968 62120 315988
rect 62120 315968 62172 315988
rect 62172 315968 62174 315988
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 651378 328072 651434 328128
rect 652390 352552 652446 352608
rect 653402 338680 653458 338736
rect 652390 329704 652446 329760
rect 652022 326848 652078 326904
rect 651378 325644 651434 325680
rect 658922 346432 658978 346488
rect 651378 325624 651380 325644
rect 651380 325624 651432 325644
rect 651432 325624 651434 325644
rect 63130 314064 63186 314120
rect 653402 313248 653458 313304
rect 62946 312976 63002 313032
rect 62762 311752 62818 311808
rect 652298 309848 652354 309904
rect 59910 309032 59966 309088
rect 651378 303320 651434 303376
rect 652298 302096 652354 302152
rect 53102 301280 53158 301336
rect 654782 300872 654838 300928
rect 651470 300600 651526 300656
rect 62762 298696 62818 298752
rect 651470 298696 651526 298752
rect 62118 295452 62174 295488
rect 62118 295432 62120 295452
rect 62120 295432 62172 295452
rect 62172 295432 62174 295452
rect 54482 266192 54538 266248
rect 62118 294092 62174 294128
rect 62118 294072 62120 294092
rect 62120 294072 62172 294092
rect 62172 294072 62174 294092
rect 62302 292712 62358 292768
rect 62118 292460 62174 292496
rect 62118 292440 62120 292460
rect 62120 292440 62172 292460
rect 62172 292440 62174 292460
rect 62118 290944 62174 291000
rect 651470 297472 651526 297528
rect 652666 296792 652722 296848
rect 652390 295296 652446 295352
rect 651470 294208 651526 294264
rect 651470 292984 651526 293040
rect 652206 291488 652262 291544
rect 651470 290400 651526 290456
rect 62762 289720 62818 289776
rect 651470 289176 651526 289232
rect 62118 288516 62174 288552
rect 62118 288496 62120 288516
rect 62120 288496 62172 288516
rect 62172 288496 62174 288516
rect 652022 288496 652078 288552
rect 651470 287408 651526 287464
rect 63130 287136 63186 287192
rect 62118 285912 62174 285968
rect 62118 284436 62174 284472
rect 62118 284416 62120 284436
rect 62120 284416 62172 284436
rect 62172 284416 62174 284436
rect 58622 278704 58678 278760
rect 57242 275848 57298 275904
rect 62762 283192 62818 283248
rect 62118 280880 62174 280936
rect 61382 280336 61438 280392
rect 60002 256672 60058 256728
rect 55862 223488 55918 223544
rect 61290 217912 61346 217968
rect 62946 282104 63002 282160
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 651470 283328 651526 283384
rect 651470 280880 651526 280936
rect 63130 267008 63186 267064
rect 462226 272312 462282 272368
rect 470414 272620 470416 272640
rect 470416 272620 470468 272640
rect 470468 272620 470470 272640
rect 470414 272584 470470 272620
rect 470598 272620 470600 272640
rect 470600 272620 470652 272640
rect 470652 272620 470654 272640
rect 470598 272584 470654 272620
rect 470414 272312 470470 272368
rect 470598 271904 470654 271960
rect 478050 271904 478106 271960
rect 489918 272720 489974 272776
rect 495714 272720 495770 272776
rect 523866 271124 523868 271144
rect 523868 271124 523920 271144
rect 523920 271124 523922 271144
rect 523866 271088 523922 271124
rect 525338 271088 525394 271144
rect 530398 270136 530454 270192
rect 534078 270136 534134 270192
rect 537298 275032 537354 275088
rect 538126 275032 538182 275088
rect 537758 269900 537760 269920
rect 537760 269900 537812 269920
rect 537812 269900 537814 269920
rect 537758 269864 537814 269900
rect 538310 269864 538366 269920
rect 539322 273672 539378 273728
rect 542266 274760 542322 274816
rect 543186 274780 543242 274816
rect 543186 274760 543188 274780
rect 543188 274760 543240 274780
rect 543240 274760 543242 274780
rect 547510 273964 547566 274000
rect 547510 273944 547512 273964
rect 547512 273944 547564 273964
rect 547564 273944 547566 273964
rect 547694 273672 547750 273728
rect 549258 273944 549314 274000
rect 549902 273672 549958 273728
rect 552846 273692 552902 273728
rect 552846 273672 552848 273692
rect 552848 273672 552900 273692
rect 552900 273672 552902 273692
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553490 255604 553546 255640
rect 553490 255584 553492 255604
rect 553492 255584 553544 255604
rect 553544 255584 553546 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553674 242528 553730 242584
rect 62946 225528 63002 225584
rect 140042 229064 140098 229120
rect 139306 228248 139362 228304
rect 141146 226108 141148 226128
rect 141148 226108 141200 226128
rect 141200 226108 141202 226128
rect 141146 226072 141202 226108
rect 142434 230444 142490 230480
rect 142434 230424 142436 230444
rect 142436 230424 142488 230444
rect 142488 230424 142490 230444
rect 142986 228248 143042 228304
rect 140778 220360 140834 220416
rect 142250 220360 142306 220416
rect 141974 219680 142030 219736
rect 144090 230424 144146 230480
rect 143998 229492 144054 229528
rect 143998 229472 144000 229492
rect 144000 229472 144052 229492
rect 144052 229472 144054 229492
rect 145378 229472 145434 229528
rect 146206 229336 146262 229392
rect 145194 226108 145196 226128
rect 145196 226108 145248 226128
rect 145248 226108 145250 226128
rect 145194 226072 145250 226108
rect 145930 222264 145986 222320
rect 144642 220632 144698 220688
rect 144182 219680 144238 219736
rect 147126 229064 147182 229120
rect 147586 229744 147642 229800
rect 147954 229744 148010 229800
rect 147770 229356 147826 229392
rect 147770 229336 147772 229356
rect 147772 229336 147824 229356
rect 147824 229336 147826 229356
rect 147678 223352 147734 223408
rect 147310 222944 147366 223000
rect 147770 222944 147826 223000
rect 147126 222300 147128 222320
rect 147128 222300 147180 222320
rect 147180 222300 147182 222320
rect 147126 222264 147182 222300
rect 150346 229200 150402 229256
rect 149242 220904 149298 220960
rect 150898 220632 150954 220688
rect 152278 223352 152334 223408
rect 152186 222672 152242 222728
rect 155130 222672 155186 222728
rect 156786 229900 156842 229936
rect 156786 229880 156788 229900
rect 156788 229880 156840 229900
rect 156840 229880 156842 229900
rect 157430 229880 157486 229936
rect 156878 228792 156934 228848
rect 156878 227432 156934 227488
rect 157522 228792 157578 228848
rect 156142 220904 156198 220960
rect 157246 223388 157248 223408
rect 157248 223388 157300 223408
rect 157300 223388 157302 223408
rect 157246 223352 157302 223388
rect 157430 223388 157432 223408
rect 157432 223388 157484 223408
rect 157484 223388 157486 223408
rect 157430 223352 157486 223388
rect 158350 221584 158406 221640
rect 159362 229356 159418 229392
rect 159362 229336 159364 229356
rect 159364 229336 159416 229356
rect 159416 229336 159418 229356
rect 160006 228112 160062 228168
rect 160834 220360 160890 220416
rect 164514 221604 164570 221640
rect 164514 221584 164516 221604
rect 164516 221584 164568 221604
rect 164568 221584 164570 221604
rect 166998 229200 167054 229256
rect 166814 228928 166870 228984
rect 166814 228112 166870 228168
rect 166538 227432 166594 227488
rect 167366 229220 167422 229256
rect 167366 229200 167368 229220
rect 167368 229200 167420 229220
rect 167420 229200 167422 229220
rect 167366 228948 167422 228984
rect 167366 228928 167368 228948
rect 167368 228928 167420 228948
rect 167420 228928 167422 228948
rect 169482 227316 169538 227352
rect 169482 227296 169484 227316
rect 169484 227296 169536 227316
rect 169536 227296 169538 227316
rect 166998 220904 167054 220960
rect 166538 220360 166594 220416
rect 166906 220224 166962 220280
rect 167090 220224 167146 220280
rect 169574 218476 169630 218512
rect 169574 218456 169576 218476
rect 169576 218456 169628 218476
rect 169628 218456 169630 218476
rect 171230 227568 171286 227624
rect 172150 227568 172206 227624
rect 171690 227296 171746 227352
rect 173346 228792 173402 228848
rect 174818 228812 174874 228848
rect 174818 228792 174820 228812
rect 174820 228792 174872 228812
rect 174872 228792 174874 228812
rect 172886 218456 172942 218512
rect 175554 220904 175610 220960
rect 176474 221332 176530 221368
rect 176474 221312 176476 221332
rect 176476 221312 176528 221332
rect 176528 221312 176530 221332
rect 177302 221312 177358 221368
rect 176474 220788 176530 220824
rect 176474 220768 176476 220788
rect 176476 220768 176528 220788
rect 176528 220768 176530 220788
rect 179878 220768 179934 220824
rect 180522 220088 180578 220144
rect 184662 221720 184718 221776
rect 185766 221740 185822 221776
rect 185766 221720 185768 221740
rect 185768 221720 185820 221740
rect 185820 221720 185822 221740
rect 185766 220088 185822 220144
rect 195886 219544 195942 219600
rect 196346 219544 196402 219600
rect 202878 229084 202934 229120
rect 202878 229064 202880 229084
rect 202880 229064 202932 229084
rect 202932 229064 202934 229084
rect 202418 219680 202474 219736
rect 203154 219700 203210 219736
rect 203154 219680 203156 219700
rect 203156 219680 203208 219700
rect 203208 219680 203210 219700
rect 205178 229064 205234 229120
rect 219438 227432 219494 227488
rect 220450 227432 220506 227488
rect 486974 219408 487030 219464
rect 487802 218048 487858 218104
rect 490378 218592 490434 218648
rect 492678 218320 492734 218376
rect 488676 217096 488732 217152
rect 493782 218320 493838 218376
rect 493782 217232 493838 217288
rect 494702 218864 494758 218920
rect 495346 217232 495402 217288
rect 497830 220904 497886 220960
rect 498106 220904 498162 220960
rect 496910 218320 496966 218376
rect 498474 217232 498530 217288
rect 505650 217504 505706 217560
rect 508502 217776 508558 217832
rect 510158 217776 510214 217832
rect 513562 221448 513618 221504
rect 515218 219408 515274 219464
rect 520186 221176 520242 221232
rect 522578 217776 522634 217832
rect 540886 221720 540942 221776
rect 543186 222264 543242 222320
rect 546958 222028 546960 222048
rect 546960 222028 547012 222048
rect 547012 222028 547014 222048
rect 546958 221992 547014 222028
rect 546774 221720 546830 221776
rect 547694 222264 547750 222320
rect 547694 221740 547750 221776
rect 547694 221720 547696 221740
rect 547696 221720 547748 221740
rect 547748 221720 547750 221740
rect 549074 221720 549130 221776
rect 551190 220088 551246 220144
rect 552846 220088 552902 220144
rect 552294 219136 552350 219192
rect 554502 244704 554558 244760
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 553858 221992 553914 222048
rect 553490 221756 553492 221776
rect 553492 221756 553544 221776
rect 553544 221756 553546 221776
rect 553490 221720 553546 221756
rect 555790 224440 555846 224496
rect 556526 219136 556582 219192
rect 555698 217776 555754 217832
rect 557998 222400 558054 222456
rect 557538 221720 557594 221776
rect 559378 221740 559434 221776
rect 559378 221720 559380 221740
rect 559380 221720 559432 221740
rect 559432 221720 559434 221740
rect 561678 224440 561734 224496
rect 562138 224304 562194 224360
rect 561678 222128 561734 222184
rect 562690 222128 562746 222184
rect 561494 221720 561550 221776
rect 562874 220632 562930 220688
rect 562322 219136 562378 219192
rect 563242 224304 563298 224360
rect 564806 222128 564862 222184
rect 564806 221720 564862 221776
rect 562690 217776 562746 217832
rect 562966 217776 563022 217832
rect 565634 220360 565690 220416
rect 567014 222400 567070 222456
rect 567382 220360 567438 220416
rect 567658 220360 567714 220416
rect 566830 220088 566886 220144
rect 567842 220088 567898 220144
rect 569590 221720 569646 221776
rect 568946 220360 569002 220416
rect 569222 219136 569278 219192
rect 576766 220632 576822 220688
rect 573362 220224 573418 220280
rect 576582 219952 576638 220008
rect 572626 219136 572682 219192
rect 574098 217776 574154 217832
rect 574098 216688 574154 216744
rect 574374 216688 574430 216744
rect 574834 217776 574890 217832
rect 650642 256672 650698 256728
rect 582470 220224 582526 220280
rect 581826 219988 581828 220008
rect 581828 219988 581880 220008
rect 581880 219988 581882 220008
rect 581826 219952 581882 219988
rect 578882 213968 578938 214024
rect 578330 211656 578386 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 599490 221448 599546 221504
rect 594798 218592 594854 218648
rect 595166 217504 595222 217560
rect 596362 217232 596418 217288
rect 595718 216960 595774 217016
rect 598478 215872 598534 215928
rect 603262 218320 603318 218376
rect 611634 219680 611690 219736
rect 618258 221176 618314 221232
rect 617246 219408 617302 219464
rect 618902 215328 618958 215384
rect 627458 218048 627514 218104
rect 627918 216144 627974 216200
rect 631322 220904 631378 220960
rect 631138 218320 631194 218376
rect 652390 283464 652446 283520
rect 652390 282104 652446 282160
rect 652574 280336 652630 280392
rect 656162 271088 656218 271144
rect 652574 229744 652630 229800
rect 652390 226888 652446 226944
rect 654782 226344 654838 226400
rect 652022 225528 652078 225584
rect 650642 222808 650698 222864
rect 649722 221448 649778 221504
rect 644754 220360 644810 220416
rect 648526 218592 648582 218648
rect 651470 221720 651526 221776
rect 653402 224984 653458 225040
rect 653034 220088 653090 220144
rect 652850 215872 652906 215928
rect 656162 225256 656218 225312
rect 655426 218864 655482 218920
rect 657542 223896 657598 223952
rect 656806 217232 656862 217288
rect 656530 212880 656586 212936
rect 664442 312024 664498 312080
rect 662418 293800 662474 293856
rect 667754 295704 667810 295760
rect 667754 293800 667810 293856
rect 665822 268504 665878 268560
rect 664442 248104 664498 248160
rect 659106 222536 659162 222592
rect 658738 214512 658794 214568
rect 663706 229064 663762 229120
rect 665178 229472 665234 229528
rect 665822 230424 665878 230480
rect 662050 217504 662106 217560
rect 661498 213424 661554 213480
rect 664442 223624 664498 223680
rect 665546 216144 665602 216200
rect 667018 221040 667074 221096
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578698 123528 578754 123584
rect 578882 121352 578938 121408
rect 578514 118360 578570 118416
rect 578330 108296 578386 108352
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110064 579398 110120
rect 579066 105848 579122 105904
rect 578514 103128 578570 103184
rect 579158 101632 579214 101688
rect 578606 97416 578662 97472
rect 578330 94968 578386 95024
rect 579526 99220 579528 99240
rect 579528 99220 579580 99240
rect 579580 99220 579582 99240
rect 579526 99184 579582 99220
rect 579250 93064 579306 93120
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 463146 53624 463202 53680
rect 461950 53080 462006 53136
rect 473910 53644 473966 53680
rect 473910 53624 473912 53644
rect 473912 53624 473964 53644
rect 473964 53624 473966 53644
rect 564530 53644 564586 53680
rect 564530 53624 564532 53644
rect 564532 53624 564584 53644
rect 564584 53624 564586 53644
rect 472806 53080 472862 53136
rect 576122 54984 576178 55040
rect 574742 53624 574798 53680
rect 578698 90888 578754 90944
rect 579250 88032 579306 88088
rect 578330 86400 578386 86456
rect 579250 83988 579252 84008
rect 579252 83988 579304 84008
rect 579304 83988 579306 84008
rect 579250 83952 579306 83988
rect 578698 82184 578754 82240
rect 578514 77832 578570 77888
rect 579434 80008 579490 80064
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 667018 176432 667074 176488
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 580446 77832 580502 77888
rect 579066 75656 579122 75712
rect 578514 71168 578570 71224
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579526 66852 579528 66872
rect 579528 66852 579580 66872
rect 579580 66852 579582 66872
rect 579526 66816 579582 66852
rect 579526 64504 579582 64560
rect 579526 61784 579582 61840
rect 578882 60424 578938 60480
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 578330 56072 578386 56128
rect 577686 54712 577742 54768
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588726 129648 588782 129704
rect 588542 103536 588598 103592
rect 667846 223624 667902 223680
rect 667570 221992 667626 222048
rect 668030 220088 668086 220144
rect 667754 219408 667810 219464
rect 667570 177248 667626 177304
rect 668030 207576 668086 207632
rect 668030 204040 668086 204096
rect 667938 199144 667994 199200
rect 667938 194112 667994 194168
rect 667938 189624 667994 189680
rect 668030 184320 668086 184376
rect 668030 179424 668086 179480
rect 667754 174936 667810 174992
rect 667386 134544 667442 134600
rect 667202 133184 667258 133240
rect 589462 128016 589518 128072
rect 589922 126384 589978 126440
rect 589370 124752 589426 124808
rect 589554 123120 589610 123176
rect 668214 173032 668270 173088
rect 668398 169632 668454 169688
rect 668214 164872 668270 164928
rect 668214 163276 668216 163296
rect 668216 163276 668268 163296
rect 668268 163276 668270 163296
rect 668214 163240 668270 163276
rect 668214 160012 668216 160032
rect 668216 160012 668268 160032
rect 668268 160012 668270 160032
rect 668214 159976 668270 160012
rect 668582 158344 668638 158400
rect 668306 155116 668308 155136
rect 668308 155116 668360 155136
rect 668360 155116 668362 155136
rect 668306 155080 668362 155116
rect 668214 148552 668270 148608
rect 668214 135496 668270 135552
rect 670606 392536 670662 392592
rect 669962 345616 670018 345672
rect 669410 174664 669466 174720
rect 669410 171944 669466 172000
rect 669778 234368 669834 234424
rect 669410 148960 669466 149016
rect 669226 143656 669282 143712
rect 668950 138760 669006 138816
rect 670422 261296 670478 261352
rect 670238 259664 670294 259720
rect 670422 247016 670478 247072
rect 670238 245656 670294 245712
rect 672722 394712 672778 394768
rect 672722 380976 672778 381032
rect 671986 372544 672042 372600
rect 672538 357040 672594 357096
rect 672354 351328 672410 351384
rect 671986 350104 672042 350160
rect 672354 337184 672410 337240
rect 671986 332288 672042 332344
rect 673366 400560 673422 400616
rect 673182 357448 673238 357504
rect 672906 356768 672962 356824
rect 672722 356224 672778 356280
rect 672538 312432 672594 312488
rect 673918 399744 673974 399800
rect 673734 394032 673790 394088
rect 673734 376624 673790 376680
rect 673366 355816 673422 355872
rect 673182 355408 673238 355464
rect 672906 348472 672962 348528
rect 672538 311616 672594 311672
rect 672722 311208 672778 311264
rect 672722 310528 672778 310584
rect 672262 305496 672318 305552
rect 672078 304272 672134 304328
rect 671526 302232 671582 302288
rect 672078 287816 672134 287872
rect 672262 285504 672318 285560
rect 671158 262112 671214 262168
rect 670974 250824 671030 250880
rect 670974 248104 671030 248160
rect 670790 232484 670846 232520
rect 670790 232464 670792 232484
rect 670792 232464 670844 232484
rect 670844 232464 670846 232484
rect 670790 231532 670846 231568
rect 670790 231512 670792 231532
rect 670792 231512 670844 231532
rect 670844 231512 670846 231532
rect 670790 226344 670846 226400
rect 670790 224984 670846 225040
rect 670790 223896 670846 223952
rect 671434 258440 671490 258496
rect 671250 225528 671306 225584
rect 670790 223352 670846 223408
rect 670790 222536 670846 222592
rect 670790 218864 670846 218920
rect 670790 217232 670846 217288
rect 670974 216552 671030 216608
rect 670698 215872 670754 215928
rect 670790 202816 670846 202872
rect 670606 169632 670662 169688
rect 670514 169088 670570 169144
rect 671802 260888 671858 260944
rect 671986 256400 672042 256456
rect 671802 246608 671858 246664
rect 671158 177928 671214 177984
rect 670514 150048 670570 150104
rect 671710 221720 671766 221776
rect 672170 233688 672226 233744
rect 672170 226364 672226 226400
rect 672170 226344 672208 226364
rect 672208 226344 672226 226364
rect 672262 225836 672264 225856
rect 672264 225836 672316 225856
rect 672316 225836 672318 225856
rect 672262 225800 672318 225836
rect 672262 225548 672318 225584
rect 672262 225528 672264 225548
rect 672264 225528 672316 225548
rect 672316 225528 672318 225548
rect 672154 225292 672156 225312
rect 672156 225292 672208 225312
rect 672208 225292 672210 225312
rect 672154 225256 672210 225292
rect 671986 210432 672042 210488
rect 671986 209888 672042 209944
rect 674194 393080 674250 393136
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 676586 402872 676642 402928
rect 676034 402600 676090 402656
rect 676586 400832 676642 400888
rect 676034 399336 676090 399392
rect 674562 395256 674618 395312
rect 679622 398384 679678 398440
rect 676218 397976 676274 398032
rect 676034 396092 676090 396128
rect 676034 396072 676036 396092
rect 676036 396072 676088 396092
rect 676088 396072 676090 396092
rect 676218 395528 676274 395584
rect 675206 394440 675262 394496
rect 675206 393080 675262 393136
rect 681002 397568 681058 397624
rect 681002 388456 681058 388512
rect 675758 385328 675814 385384
rect 675298 382880 675354 382936
rect 675758 382200 675814 382256
rect 675390 380976 675446 381032
rect 675758 378664 675814 378720
rect 675758 377440 675814 377496
rect 675114 376624 675170 376680
rect 675758 373632 675814 373688
rect 675666 372952 675722 373008
rect 675114 372544 675170 372600
rect 675574 358264 675630 358320
rect 673918 355000 673974 355056
rect 674102 354592 674158 354648
rect 673734 352552 673790 352608
rect 673366 349696 673422 349752
rect 673550 349288 673606 349344
rect 673366 335552 673422 335608
rect 673918 348880 673974 348936
rect 673734 333920 673790 333976
rect 673550 332696 673606 332752
rect 673918 331200 673974 331256
rect 674746 354184 674802 354240
rect 674286 350920 674342 350976
rect 674562 350512 674618 350568
rect 675942 357856 675998 357912
rect 675942 356496 675998 356552
rect 675850 353776 675906 353832
rect 675574 352824 675630 352880
rect 675850 351872 675906 351928
rect 676034 351736 676090 351792
rect 683118 347656 683174 347712
rect 676034 347248 676090 347304
rect 676494 346568 676550 346624
rect 683118 346432 683174 346488
rect 676034 345616 676090 345672
rect 675574 340720 675630 340776
rect 675758 340176 675814 340232
rect 675114 338680 675170 338736
rect 675666 337728 675722 337784
rect 675114 337184 675170 337240
rect 675114 335552 675170 335608
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675114 332288 675170 332344
rect 675114 331200 675170 331256
rect 675758 328344 675814 328400
rect 673366 312024 673422 312080
rect 673090 310800 673146 310856
rect 673182 310528 673238 310584
rect 675298 325488 675354 325544
rect 675114 325216 675170 325272
rect 676218 313928 676274 313984
rect 674654 310392 674710 310448
rect 674470 309984 674526 310040
rect 674194 309576 674250 309632
rect 674010 303864 674066 303920
rect 674010 286456 674066 286512
rect 673366 267416 673422 267472
rect 673918 267008 673974 267064
rect 673182 266600 673238 266656
rect 673550 266192 673606 266248
rect 673366 260480 673422 260536
rect 673182 258848 673238 258904
rect 673182 241440 673238 241496
rect 673734 265376 673790 265432
rect 674378 305088 674434 305144
rect 675850 309304 675906 309360
rect 676034 308352 676090 308408
rect 675114 307944 675170 308000
rect 674654 303456 674710 303512
rect 674378 283464 674434 283520
rect 674378 267824 674434 267880
rect 674194 264968 674250 265024
rect 674470 264560 674526 264616
rect 674286 262520 674342 262576
rect 674102 259256 674158 259312
rect 673734 241984 673790 242040
rect 673550 241712 673606 241768
rect 673366 240216 673422 240272
rect 673274 234368 673330 234424
rect 673642 234796 673698 234832
rect 673642 234776 673644 234796
rect 673644 234776 673696 234796
rect 673696 234776 673698 234796
rect 673458 230444 673514 230480
rect 673458 230424 673460 230444
rect 673460 230424 673512 230444
rect 673512 230424 673514 230444
rect 673182 228520 673238 228576
rect 673366 227024 673422 227080
rect 673550 226752 673606 226808
rect 673458 223352 673514 223408
rect 672998 222808 673054 222864
rect 673182 215736 673238 215792
rect 672998 213560 673054 213616
rect 672906 213288 672962 213344
rect 672630 208256 672686 208312
rect 672814 203768 672870 203824
rect 672722 203360 672778 203416
rect 671986 193160 672042 193216
rect 671986 170312 672042 170368
rect 672814 202544 672870 202600
rect 673550 214920 673606 214976
rect 673366 213696 673422 213752
rect 673182 200776 673238 200832
rect 673550 201048 673606 201104
rect 673366 196016 673422 196072
rect 673366 185544 673422 185600
rect 672446 177656 672502 177712
rect 672262 168136 672318 168192
rect 672262 167864 672318 167920
rect 672354 166232 672410 166288
rect 672170 165552 672226 165608
rect 671710 150320 671766 150376
rect 671986 150320 672042 150376
rect 671526 145288 671582 145344
rect 669226 133728 669282 133784
rect 669226 132912 669282 132968
rect 668950 131144 669006 131200
rect 668766 130600 668822 130656
rect 668582 128968 668638 129024
rect 668582 126928 668638 126984
rect 668030 125296 668086 125352
rect 589554 121508 589610 121544
rect 589554 121488 589556 121508
rect 589556 121488 589608 121508
rect 589608 121488 589610 121508
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589462 110064 589518 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589830 105168 589886 105224
rect 666650 109316 666706 109372
rect 667938 107752 667994 107808
rect 668030 106120 668086 106176
rect 668214 104352 668270 104408
rect 589462 101904 589518 101960
rect 625434 94424 625490 94480
rect 635554 96872 635610 96928
rect 635738 95920 635794 95976
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 645582 96076 645638 96112
rect 645582 96056 645584 96076
rect 645584 96056 645636 96076
rect 645636 96056 645638 96076
rect 647330 94968 647386 95024
rect 648066 96484 648122 96520
rect 648066 96464 648068 96484
rect 648068 96464 648120 96484
rect 648120 96464 648122 96484
rect 647882 95784 647938 95840
rect 626354 93608 626410 93664
rect 626170 92792 626226 92848
rect 625802 91976 625858 92032
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 625250 89528 625306 89584
rect 625434 88712 625490 88768
rect 624974 88576 625030 88632
rect 625250 88576 625306 88632
rect 626446 87896 626502 87952
rect 625618 87080 625674 87136
rect 648250 89528 648306 89584
rect 648802 96076 648858 96112
rect 648802 96056 648804 96076
rect 648804 96056 648856 96076
rect 648856 96056 648858 96076
rect 648618 91976 648674 92032
rect 649262 96464 649318 96520
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 625342 85448 625398 85504
rect 626446 84632 626502 84688
rect 648618 84632 648674 84688
rect 625802 83816 625858 83872
rect 628746 83272 628802 83328
rect 650550 87080 650606 87136
rect 655058 94152 655114 94208
rect 654690 93336 654746 93392
rect 655426 91432 655482 91488
rect 655426 90616 655482 90672
rect 656346 95784 656402 95840
rect 655794 89800 655850 89856
rect 663982 92520 664038 92576
rect 664166 91704 664222 91760
rect 663798 91024 663854 91080
rect 664534 89800 664590 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 650274 82184 650330 82240
rect 629206 81640 629262 81696
rect 623042 77288 623098 77344
rect 591302 54440 591358 54496
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 77560 639658 77616
rect 646318 74160 646374 74216
rect 646502 71712 646558 71768
rect 646134 69128 646190 69184
rect 646134 67088 646190 67144
rect 308034 50224 308090 50280
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 458362 46688 458418 46744
rect 459190 44376 459246 44432
rect 142618 44240 142674 44296
rect 255870 44104 255926 44160
rect 307298 43832 307354 43888
rect 440238 43852 440294 43888
rect 440238 43832 440240 43852
rect 440240 43832 440292 43852
rect 440292 43832 440294 43852
rect 194322 42064 194378 42120
rect 441066 43852 441122 43888
rect 441066 43832 441068 43852
rect 441068 43832 441120 43852
rect 441120 43832 441122 43852
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 405646 41792 405702 41848
rect 419906 41792 419962 41848
rect 446218 42200 446274 42256
rect 460110 44104 460166 44160
rect 460846 43424 460902 43480
rect 461950 44376 462006 44432
rect 462502 44376 462558 44432
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463882 44104 463938 44160
rect 463974 42880 464030 42936
rect 549994 48864 550050 48920
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 647514 78104 647570 78160
rect 647330 64368 647386 64424
rect 648986 62056 649042 62112
rect 648618 59200 648674 59256
rect 647514 57296 647570 57352
rect 661590 48454 661646 48510
rect 661774 47733 661830 47789
rect 667938 102720 667994 102776
rect 668766 122576 668822 122632
rect 669962 130872 670018 130928
rect 669226 119584 669282 119640
rect 668950 119176 669006 119232
rect 669226 114280 669282 114336
rect 668950 112648 669006 112704
rect 671342 128288 671398 128344
rect 671526 121352 671582 121408
rect 672354 131144 672410 131200
rect 672354 124752 672410 124808
rect 672170 115776 672226 115832
rect 671526 111016 671582 111072
rect 672722 161336 672778 161392
rect 672722 131688 672778 131744
rect 672538 117544 672594 117600
rect 672354 106936 672410 106992
rect 673366 174392 673422 174448
rect 673182 168680 673238 168736
rect 673182 151272 673238 151328
rect 673550 168272 673606 168328
rect 673550 166232 673606 166288
rect 674286 243616 674342 243672
rect 674194 242800 674250 242856
rect 674470 235184 674526 235240
rect 674378 230424 674434 230480
rect 674332 229472 674388 229528
rect 674470 229200 674526 229256
rect 673918 222264 673974 222320
rect 673918 220224 673974 220280
rect 674286 226752 674342 226808
rect 674102 213016 674158 213072
rect 674102 209616 674158 209672
rect 673918 175616 673974 175672
rect 673918 170720 673974 170776
rect 673918 156440 673974 156496
rect 673734 153176 673790 153232
rect 673366 129648 673422 129704
rect 673366 126520 673422 126576
rect 672906 124072 672962 124128
rect 673182 123936 673238 123992
rect 673458 123120 673514 123176
rect 673918 122168 673974 122224
rect 673458 119584 673514 119640
rect 673182 106256 673238 106312
rect 672722 106120 672778 106176
rect 668582 102720 668638 102776
rect 676034 307536 676090 307592
rect 676034 305904 676090 305960
rect 674838 301960 674894 302016
rect 675850 301960 675906 302016
rect 676034 300600 676090 300656
rect 679622 306720 679678 306776
rect 677598 306312 677654 306368
rect 675942 297336 675998 297392
rect 683026 302640 683082 302696
rect 683026 299376 683082 299432
rect 675206 296520 675262 296576
rect 675850 296520 675906 296576
rect 676126 296520 676182 296576
rect 675390 295704 675446 295760
rect 675758 295704 675814 295760
rect 675758 294480 675814 294536
rect 675574 292168 675630 292224
rect 675758 291488 675814 291544
rect 675758 290808 675814 290864
rect 675114 287816 675170 287872
rect 675390 286456 675446 286512
rect 675114 285504 675170 285560
rect 675666 283600 675722 283656
rect 675666 282784 675722 282840
rect 675758 281152 675814 281208
rect 683118 271088 683174 271144
rect 683118 268504 683174 268560
rect 675482 265784 675538 265840
rect 681002 263200 681058 263256
rect 676218 262792 676274 262848
rect 676218 257080 676274 257136
rect 676218 256400 676274 256456
rect 674838 255312 674894 255368
rect 675850 255312 675906 255368
rect 674838 247832 674894 247888
rect 683026 257488 683082 257544
rect 675482 250824 675538 250880
rect 675758 250144 675814 250200
rect 675482 249464 675538 249520
rect 675298 247016 675354 247072
rect 675298 246608 675354 246664
rect 675298 245656 675354 245712
rect 675114 243616 675170 243672
rect 675114 242800 675170 242856
rect 675758 242256 675814 242312
rect 675114 241440 675170 241496
rect 675114 240216 675170 240272
rect 675850 235184 675906 235240
rect 675390 234776 675446 234832
rect 675022 226344 675078 226400
rect 674838 225800 674894 225856
rect 674654 223624 674710 223680
rect 674838 221448 674894 221504
rect 675206 225256 675262 225312
rect 675022 220496 675078 220552
rect 675206 218592 675262 218648
rect 675022 217776 675078 217832
rect 674654 216960 674710 217016
rect 674838 216144 674894 216200
rect 674470 214104 674526 214160
rect 674470 201320 674526 201376
rect 675850 233724 675852 233744
rect 675852 233724 675904 233744
rect 675904 233724 675906 233744
rect 675850 233688 675906 233724
rect 675850 232500 675852 232520
rect 675852 232500 675904 232520
rect 675904 232500 675906 232520
rect 675850 232464 675906 232500
rect 675850 231532 675906 231568
rect 675850 231512 675852 231532
rect 675852 231512 675904 231532
rect 675904 231512 675906 231532
rect 676586 230424 676642 230480
rect 676034 230152 676090 230208
rect 676218 228520 676274 228576
rect 676034 221448 676090 221504
rect 676034 219020 676090 219056
rect 676034 219000 676036 219020
rect 676036 219000 676088 219020
rect 676088 219000 676090 219020
rect 675574 217504 675630 217560
rect 675942 215500 675944 215520
rect 675944 215500 675996 215520
rect 675996 215500 675998 215520
rect 675942 215464 675998 215500
rect 675942 214648 675998 214704
rect 677046 227024 677102 227080
rect 675850 212064 675906 212120
rect 675850 209616 675906 209672
rect 678242 223760 678298 223816
rect 683210 222672 683266 222728
rect 683578 223080 683634 223136
rect 683394 219816 683450 219872
rect 683302 218592 683358 218648
rect 683118 212880 683174 212936
rect 678978 211384 679034 211440
rect 680358 210568 680414 210624
rect 683302 210296 683358 210352
rect 678978 207576 679034 207632
rect 676862 206896 676918 206952
rect 675758 205536 675814 205592
rect 675758 204176 675814 204232
rect 675206 202816 675262 202872
rect 675298 201320 675354 201376
rect 675114 201048 675170 201104
rect 675482 200776 675538 200832
rect 675758 200776 675814 200832
rect 675758 198328 675814 198384
rect 675114 196016 675170 196072
rect 675298 195880 675354 195936
rect 675114 193160 675170 193216
rect 675666 192752 675722 192808
rect 676862 189624 676918 189680
rect 674286 178064 674342 178120
rect 674286 176840 674342 176896
rect 674470 176024 674526 176080
rect 674286 132096 674342 132152
rect 674654 175208 674710 175264
rect 674470 131280 674526 131336
rect 674930 173984 674986 174040
rect 676034 173168 676090 173224
rect 675114 169360 675170 169416
rect 675942 169360 675998 169416
rect 676586 169904 676642 169960
rect 676034 167048 676090 167104
rect 683118 185544 683174 185600
rect 683118 178744 683174 178800
rect 678242 171536 678298 171592
rect 676586 166368 676642 166424
rect 676862 166368 676918 166424
rect 676034 165552 676090 165608
rect 675482 161336 675538 161392
rect 675666 161200 675722 161256
rect 675758 159976 675814 160032
rect 674930 159432 674986 159488
rect 675482 159432 675538 159488
rect 675390 156984 675446 157040
rect 675758 156984 675814 157040
rect 675114 156440 675170 156496
rect 675758 155760 675814 155816
rect 675666 153040 675722 153096
rect 675758 151408 675814 151464
rect 675114 151272 675170 151328
rect 675114 150320 675170 150376
rect 674930 150048 674986 150104
rect 675298 148960 675354 149016
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 676034 134544 676090 134600
rect 676034 132504 676090 132560
rect 674654 130464 674710 130520
rect 675850 130056 675906 130112
rect 674838 127336 674894 127392
rect 674470 124344 674526 124400
rect 674102 120400 674158 120456
rect 674654 123528 674710 123584
rect 674470 110336 674526 110392
rect 676218 128968 676274 129024
rect 676034 128288 676090 128344
rect 676218 127744 676274 127800
rect 675850 126928 675906 126984
rect 682382 126112 682438 126168
rect 676218 125704 676274 125760
rect 675114 116728 675170 116784
rect 675942 122848 675998 122904
rect 678978 125296 679034 125352
rect 678978 121216 679034 121272
rect 683118 125704 683174 125760
rect 683302 124888 683358 124944
rect 683118 121624 683174 121680
rect 675850 116728 675906 116784
rect 683302 116456 683358 116512
rect 675482 115776 675538 115832
rect 675758 114144 675814 114200
rect 675758 111696 675814 111752
rect 675666 111288 675722 111344
rect 675114 110336 675170 110392
rect 675758 108160 675814 108216
rect 675390 106936 675446 106992
rect 675114 106256 675170 106312
rect 675666 104760 675722 104816
rect 675758 103128 675814 103184
rect 673366 100952 673422 101008
rect 675114 100952 675170 101008
rect 662418 47368 662474 47424
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 446218 41520 446274 41576
rect 141698 40296 141754 40352
<< metal3 >>
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675702 892196 675708 892260
rect 675772 892258 675778 892260
rect 675772 892198 676292 892258
rect 675772 892196 675778 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 675845 891442 675911 891445
rect 675845 891440 676292 891442
rect 675845 891384 675850 891440
rect 675906 891384 676292 891440
rect 675845 891382 676292 891384
rect 675845 891379 675911 891382
rect 675661 891034 675727 891037
rect 675661 891032 676292 891034
rect 675661 890976 675666 891032
rect 675722 890976 676292 891032
rect 675661 890974 676292 890976
rect 675661 890971 675727 890974
rect 676029 890626 676095 890629
rect 676029 890624 676292 890626
rect 676029 890568 676034 890624
rect 676090 890568 676292 890624
rect 676029 890566 676292 890568
rect 676029 890563 676095 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 683297 889402 683363 889405
rect 683284 889400 683363 889402
rect 683284 889344 683302 889400
rect 683358 889344 683363 889400
rect 683284 889342 683363 889344
rect 683297 889339 683363 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 676029 888178 676095 888181
rect 676029 888176 676292 888178
rect 676029 888120 676034 888176
rect 676090 888120 676292 888176
rect 676029 888118 676292 888120
rect 676029 888115 676095 888118
rect 675886 887708 675892 887772
rect 675956 887770 675962 887772
rect 675956 887710 676292 887770
rect 675956 887708 675962 887710
rect 675518 887436 675524 887500
rect 675588 887498 675594 887500
rect 676029 887498 676095 887501
rect 675588 887496 676095 887498
rect 675588 887440 676034 887496
rect 676090 887440 676095 887496
rect 675588 887438 676095 887440
rect 675588 887436 675594 887438
rect 676029 887435 676095 887438
rect 676673 887362 676739 887365
rect 676660 887360 676739 887362
rect 676660 887304 676678 887360
rect 676734 887304 676739 887360
rect 676660 887302 676739 887304
rect 676673 887299 676739 887302
rect 675477 886954 675543 886957
rect 675477 886952 676000 886954
rect 675477 886896 675482 886952
rect 675538 886920 676000 886952
rect 676262 886920 676322 886924
rect 675538 886896 676322 886920
rect 675477 886894 676322 886896
rect 675477 886891 675543 886894
rect 675940 886860 676322 886894
rect 683070 886141 683130 886516
rect 683021 886136 683130 886141
rect 683021 886080 683026 886136
rect 683082 886108 683130 886136
rect 683082 886080 683100 886108
rect 683021 886078 683100 886080
rect 683021 886075 683087 886078
rect 676029 885730 676095 885733
rect 676029 885728 676292 885730
rect 676029 885672 676034 885728
rect 676090 885672 676292 885728
rect 676029 885670 676292 885672
rect 676029 885667 676095 885670
rect 676673 882604 676739 882605
rect 676622 882602 676628 882604
rect 676582 882542 676628 882602
rect 676692 882600 676739 882604
rect 676734 882544 676739 882600
rect 676622 882540 676628 882542
rect 676692 882540 676739 882544
rect 676673 882539 676739 882540
rect 675702 881860 675708 881924
rect 675772 881922 675778 881924
rect 683021 881922 683087 881925
rect 675772 881920 683087 881922
rect 675772 881864 683026 881920
rect 683082 881864 683087 881920
rect 675772 881862 683087 881864
rect 675772 881860 675778 881862
rect 683021 881859 683087 881862
rect 675937 878522 676003 878525
rect 675710 878520 676003 878522
rect 675710 878464 675942 878520
rect 675998 878464 676003 878520
rect 675710 878462 676003 878464
rect 675710 877845 675770 878462
rect 675937 878459 676003 878462
rect 675661 877840 675770 877845
rect 675661 877784 675666 877840
rect 675722 877784 675770 877840
rect 675661 877782 675770 877784
rect 675661 877779 675727 877782
rect 675477 876484 675543 876485
rect 675477 876482 675524 876484
rect 675432 876480 675524 876482
rect 675432 876424 675482 876480
rect 675432 876422 675524 876424
rect 675477 876420 675524 876422
rect 675588 876420 675594 876484
rect 675477 876419 675543 876420
rect 675017 874170 675083 874173
rect 675477 874170 675543 874173
rect 675017 874168 675543 874170
rect 675017 874112 675022 874168
rect 675078 874112 675482 874168
rect 675538 874112 675543 874168
rect 675017 874110 675543 874112
rect 675017 874107 675083 874110
rect 675477 874107 675543 874110
rect 675569 873492 675635 873493
rect 675518 873490 675524 873492
rect 675478 873430 675524 873490
rect 675588 873488 675635 873492
rect 675630 873432 675635 873488
rect 675518 873428 675524 873430
rect 675588 873428 675635 873432
rect 675569 873427 675635 873428
rect 675753 869818 675819 869821
rect 676254 869818 676260 869820
rect 675753 869816 676260 869818
rect 675753 869760 675758 869816
rect 675814 869760 676260 869816
rect 675753 869758 676260 869760
rect 675753 869755 675819 869758
rect 676254 869756 676260 869758
rect 676324 869756 676330 869820
rect 675753 868730 675819 868733
rect 676622 868730 676628 868732
rect 675753 868728 676628 868730
rect 675753 868672 675758 868728
rect 675814 868672 676628 868728
rect 675753 868670 676628 868672
rect 675753 868667 675819 868670
rect 676622 868668 676628 868670
rect 676692 868668 676698 868732
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 652017 867642 652083 867645
rect 649950 867640 652083 867642
rect 649950 867584 652022 867640
rect 652078 867584 652083 867640
rect 649950 867582 652083 867584
rect 649950 867064 650010 867582
rect 652017 867579 652083 867582
rect 675109 867234 675175 867237
rect 675702 867234 675708 867236
rect 675109 867232 675708 867234
rect 675109 867176 675114 867232
rect 675170 867176 675708 867232
rect 675109 867174 675708 867176
rect 675109 867171 675175 867174
rect 675702 867172 675708 867174
rect 675772 867172 675778 867236
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 674833 866282 674899 866285
rect 675385 866282 675451 866285
rect 674833 866280 675451 866282
rect 674833 866224 674838 866280
rect 674894 866224 675390 866280
rect 675446 866224 675451 866280
rect 674833 866222 675451 866224
rect 674833 866219 674899 866222
rect 675385 866219 675451 866222
rect 675109 865738 675175 865741
rect 675886 865738 675892 865740
rect 675109 865736 675892 865738
rect 675109 865680 675114 865736
rect 675170 865680 675892 865736
rect 675109 865678 675892 865680
rect 675109 865675 675175 865678
rect 675886 865676 675892 865678
rect 675956 865676 675962 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35433 816914 35499 816917
rect 35420 816912 35499 816914
rect 35420 816856 35438 816912
rect 35494 816856 35499 816912
rect 35420 816854 35499 816856
rect 35433 816851 35499 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 40953 812834 41019 812837
rect 40940 812832 41019 812834
rect 40940 812776 40958 812832
rect 41014 812776 41019 812832
rect 40940 812774 41019 812776
rect 40953 812771 41019 812774
rect 41137 812426 41203 812429
rect 41124 812424 41203 812426
rect 41124 812368 41142 812424
rect 41198 812368 41203 812424
rect 41124 812366 41203 812368
rect 41137 812363 41203 812366
rect 41822 812018 41828 812020
rect 41492 811958 41828 812018
rect 41822 811956 41828 811958
rect 41892 811956 41898 812020
rect 39297 811610 39363 811613
rect 39284 811608 39363 811610
rect 39284 811552 39302 811608
rect 39358 811552 39363 811608
rect 39284 811550 39363 811552
rect 39297 811547 39363 811550
rect 33041 811202 33107 811205
rect 33028 811200 33107 811202
rect 33028 811144 33046 811200
rect 33102 811144 33107 811200
rect 33028 811142 33107 811144
rect 33041 811139 33107 811142
rect 42149 810794 42215 810797
rect 41492 810792 42215 810794
rect 41492 810736 42154 810792
rect 42210 810736 42215 810792
rect 41492 810734 42215 810736
rect 42149 810731 42215 810734
rect 41965 810386 42031 810389
rect 41492 810384 42031 810386
rect 41492 810328 41970 810384
rect 42026 810328 42031 810384
rect 41492 810326 42031 810328
rect 41965 810323 42031 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 33777 809570 33843 809573
rect 33764 809568 33843 809570
rect 33764 809512 33782 809568
rect 33838 809512 33843 809568
rect 33764 809510 33843 809512
rect 33777 809507 33843 809510
rect 41781 809300 41847 809301
rect 41781 809296 41828 809300
rect 41892 809298 41898 809300
rect 41781 809240 41786 809296
rect 41781 809236 41828 809240
rect 41892 809238 41938 809298
rect 41892 809236 41898 809238
rect 41781 809235 41847 809236
rect 40677 809162 40743 809165
rect 40677 809160 40756 809162
rect 40677 809104 40682 809160
rect 40738 809104 40756 809160
rect 40677 809102 40756 809104
rect 40677 809099 40743 809102
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 40953 808346 41019 808349
rect 40940 808344 41019 808346
rect 40940 808288 40958 808344
rect 41014 808288 41019 808344
rect 40940 808286 41019 808288
rect 40953 808283 41019 808286
rect 41137 807938 41203 807941
rect 41124 807936 41203 807938
rect 41124 807880 41142 807936
rect 41198 807880 41203 807936
rect 41124 807878 41203 807880
rect 41137 807875 41203 807878
rect 42977 807530 43043 807533
rect 41492 807528 43043 807530
rect 41492 807472 42982 807528
rect 43038 807472 43043 807528
rect 41492 807470 43043 807472
rect 42977 807467 43043 807470
rect 31710 806717 31770 807092
rect 31710 806712 31819 806717
rect 31710 806684 31758 806712
rect 31740 806656 31758 806684
rect 31814 806656 31819 806712
rect 31740 806654 31819 806656
rect 31753 806651 31819 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40718 805564 40724 805628
rect 40788 805626 40794 805628
rect 41965 805626 42031 805629
rect 40788 805624 42031 805626
rect 40788 805568 41970 805624
rect 42026 805568 42031 805624
rect 40788 805566 42031 805568
rect 40788 805564 40794 805566
rect 41965 805563 42031 805566
rect 40902 805156 40908 805220
rect 40972 805218 40978 805220
rect 41781 805218 41847 805221
rect 40972 805216 41847 805218
rect 40972 805160 41786 805216
rect 41842 805160 41847 805216
rect 40972 805158 41847 805160
rect 40972 805156 40978 805158
rect 41781 805155 41847 805158
rect 40534 804884 40540 804948
rect 40604 804946 40610 804948
rect 42149 804946 42215 804949
rect 40604 804944 42215 804946
rect 40604 804888 42154 804944
rect 42210 804888 42215 804944
rect 40604 804886 42215 804888
rect 40604 804884 40610 804886
rect 42149 804883 42215 804886
rect 40677 801546 40743 801549
rect 42006 801546 42012 801548
rect 40677 801544 42012 801546
rect 40677 801488 40682 801544
rect 40738 801488 42012 801544
rect 40677 801486 42012 801488
rect 40677 801483 40743 801486
rect 42006 801484 42012 801486
rect 42076 801484 42082 801548
rect 39849 801274 39915 801277
rect 41270 801274 41276 801276
rect 39849 801272 41276 801274
rect 39849 801216 39854 801272
rect 39910 801216 41276 801272
rect 39849 801214 41276 801216
rect 39849 801211 39915 801214
rect 41270 801212 41276 801214
rect 41340 801212 41346 801276
rect 40677 800866 40743 800869
rect 41086 800866 41092 800868
rect 40677 800864 41092 800866
rect 40677 800808 40682 800864
rect 40738 800808 41092 800864
rect 40677 800806 41092 800808
rect 40677 800803 40743 800806
rect 41086 800804 41092 800806
rect 41156 800804 41162 800868
rect 39297 800594 39363 800597
rect 40350 800594 40356 800596
rect 39297 800592 40356 800594
rect 39297 800536 39302 800592
rect 39358 800536 40356 800592
rect 39297 800534 40356 800536
rect 39297 800531 39363 800534
rect 40350 800532 40356 800534
rect 40420 800532 40426 800596
rect 42149 797330 42215 797333
rect 43529 797330 43595 797333
rect 42149 797328 43595 797330
rect 42149 797272 42154 797328
rect 42210 797272 43534 797328
rect 43590 797272 43595 797328
rect 42149 797270 43595 797272
rect 42149 797267 42215 797270
rect 43529 797267 43595 797270
rect 41086 796860 41092 796924
rect 41156 796922 41162 796924
rect 42701 796922 42767 796925
rect 41156 796920 42767 796922
rect 41156 796864 42706 796920
rect 42762 796864 42767 796920
rect 41156 796862 42767 796864
rect 41156 796860 41162 796862
rect 42701 796859 42767 796862
rect 41270 796180 41276 796244
rect 41340 796242 41346 796244
rect 41781 796242 41847 796245
rect 41340 796240 41847 796242
rect 41340 796184 41786 796240
rect 41842 796184 41847 796240
rect 41340 796182 41847 796184
rect 41340 796180 41346 796182
rect 41781 796179 41847 796182
rect 42057 794476 42123 794477
rect 42006 794474 42012 794476
rect 41966 794414 42012 794474
rect 42076 794472 42123 794476
rect 42118 794416 42123 794472
rect 42006 794412 42012 794414
rect 42076 794412 42123 794416
rect 42057 794411 42123 794412
rect 40350 793052 40356 793116
rect 40420 793114 40426 793116
rect 41781 793114 41847 793117
rect 40420 793112 41847 793114
rect 40420 793056 41786 793112
rect 41842 793056 41847 793112
rect 40420 793054 41847 793056
rect 40420 793052 40426 793054
rect 41781 793051 41847 793054
rect 40902 790604 40908 790668
rect 40972 790666 40978 790668
rect 41781 790666 41847 790669
rect 40972 790664 41847 790666
rect 40972 790608 41786 790664
rect 41842 790608 41847 790664
rect 40972 790606 41847 790608
rect 40972 790604 40978 790606
rect 41781 790603 41847 790606
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 41638 790196 41644 790260
rect 41708 790258 41714 790260
rect 42333 790258 42399 790261
rect 41708 790256 42399 790258
rect 41708 790200 42338 790256
rect 42394 790200 42399 790256
rect 41708 790198 42399 790200
rect 41708 790196 41714 790198
rect 42333 790195 42399 790198
rect 42057 789850 42123 789853
rect 42701 789850 42767 789853
rect 42057 789848 42767 789850
rect 42057 789792 42062 789848
rect 42118 789792 42706 789848
rect 42762 789792 42767 789848
rect 42057 789790 42767 789792
rect 42057 789787 42123 789790
rect 42701 789787 42767 789790
rect 40534 789380 40540 789444
rect 40604 789442 40610 789444
rect 42517 789442 42583 789445
rect 40604 789440 42583 789442
rect 40604 789384 42522 789440
rect 42578 789384 42583 789440
rect 40604 789382 42583 789384
rect 40604 789380 40610 789382
rect 42517 789379 42583 789382
rect 41822 789108 41828 789172
rect 41892 789170 41898 789172
rect 42701 789170 42767 789173
rect 41892 789168 42767 789170
rect 41892 789112 42706 789168
rect 42762 789112 42767 789168
rect 41892 789110 42767 789112
rect 41892 789108 41898 789110
rect 42701 789107 42767 789110
rect 62113 789170 62179 789173
rect 62113 789168 64706 789170
rect 62113 789112 62118 789168
rect 62174 789112 64706 789168
rect 62113 789110 64706 789112
rect 62113 789107 62179 789110
rect 40718 788700 40724 788764
rect 40788 788762 40794 788764
rect 41781 788762 41847 788765
rect 40788 788760 41847 788762
rect 40788 788704 41786 788760
rect 41842 788704 41847 788760
rect 40788 788702 41847 788704
rect 40788 788700 40794 788702
rect 41781 788699 41847 788702
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 675385 788084 675451 788085
rect 675334 788082 675340 788084
rect 675294 788022 675340 788082
rect 675404 788080 675451 788084
rect 675446 788024 675451 788080
rect 675334 788020 675340 788022
rect 675404 788020 675451 788024
rect 675385 788019 675451 788020
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62757 787130 62823 787133
rect 62757 787128 64706 787130
rect 62757 787072 62762 787128
rect 62818 787072 64706 787128
rect 62757 787070 64706 787072
rect 62757 787067 62823 787070
rect 64646 786758 64706 787070
rect 675477 786724 675543 786725
rect 675477 786720 675524 786724
rect 675588 786722 675594 786724
rect 675477 786664 675482 786720
rect 675477 786660 675524 786664
rect 675588 786662 675634 786722
rect 675588 786660 675594 786662
rect 675477 786659 675543 786660
rect 61377 786178 61443 786181
rect 61377 786176 64706 786178
rect 61377 786120 61382 786176
rect 61438 786120 64706 786176
rect 61377 786118 64706 786120
rect 61377 786115 61443 786118
rect 64646 785576 64706 786118
rect 62113 784954 62179 784957
rect 62113 784952 64706 784954
rect 62113 784896 62118 784952
rect 62174 784896 64706 784952
rect 62113 784894 64706 784896
rect 62113 784891 62179 784894
rect 64646 784394 64706 784894
rect 674230 783804 674236 783868
rect 674300 783866 674306 783868
rect 675477 783866 675543 783869
rect 674300 783864 675543 783866
rect 674300 783808 675482 783864
rect 675538 783808 675543 783864
rect 674300 783806 675543 783808
rect 674300 783804 674306 783806
rect 675477 783803 675543 783806
rect 675753 779922 675819 779925
rect 676990 779922 676996 779924
rect 675753 779920 676996 779922
rect 675753 779864 675758 779920
rect 675814 779864 676996 779920
rect 675753 779862 676996 779864
rect 675753 779859 675819 779862
rect 676990 779860 676996 779862
rect 677060 779860 677066 779924
rect 649950 778426 650010 778824
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 649950 776114 650010 776460
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 651465 776051 651531 776054
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 41045 774754 41111 774757
rect 44265 774754 44331 774757
rect 41045 774752 44331 774754
rect 41045 774696 41050 774752
rect 41106 774696 44270 774752
rect 44326 774696 44331 774752
rect 41045 774694 44331 774696
rect 41045 774691 41111 774694
rect 44265 774691 44331 774694
rect 35758 774452 35818 774691
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35390 773941 35450 774044
rect 35390 773936 35499 773941
rect 35390 773880 35438 773936
rect 35494 773880 35499 773936
rect 35390 773878 35499 773880
rect 35433 773875 35499 773878
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 41321 773530 41387 773533
rect 42057 773530 42123 773533
rect 41321 773528 42123 773530
rect 41321 773472 41326 773528
rect 41382 773472 42062 773528
rect 42118 773472 42123 773528
rect 41321 773470 42123 773472
rect 41321 773467 41387 773470
rect 42057 773467 42123 773470
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35758 773125 35818 773228
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 41689 773122 41755 773125
rect 46197 773122 46263 773125
rect 41689 773120 46263 773122
rect 41689 773064 41694 773120
rect 41750 773064 46202 773120
rect 46258 773064 46263 773120
rect 41689 773062 46263 773064
rect 41689 773059 41755 773062
rect 46197 773059 46263 773062
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 41781 772850 41847 772853
rect 44909 772850 44975 772853
rect 41781 772848 44975 772850
rect 35574 772717 35634 772820
rect 41781 772792 41786 772848
rect 41842 772792 44914 772848
rect 44970 772792 44975 772848
rect 41781 772790 44975 772792
rect 41781 772787 41847 772790
rect 44909 772787 44975 772790
rect 35574 772712 35683 772717
rect 35574 772656 35622 772712
rect 35678 772656 35683 772712
rect 35574 772654 35683 772656
rect 35617 772651 35683 772654
rect 35390 772309 35450 772412
rect 35341 772304 35450 772309
rect 35341 772248 35346 772304
rect 35402 772248 35450 772304
rect 35341 772246 35450 772248
rect 35341 772243 35407 772246
rect 35574 771901 35634 772004
rect 35525 771896 35634 771901
rect 35801 771898 35867 771901
rect 35525 771840 35530 771896
rect 35586 771840 35634 771896
rect 35525 771838 35634 771840
rect 35758 771896 35867 771898
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35525 771835 35591 771838
rect 35758 771835 35867 771840
rect 35758 771596 35818 771835
rect 35758 771085 35818 771188
rect 35758 771080 35867 771085
rect 35758 771024 35806 771080
rect 35862 771024 35867 771080
rect 35758 771022 35867 771024
rect 35801 771019 35867 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 40309 770266 40375 770269
rect 44541 770266 44607 770269
rect 40309 770264 44607 770266
rect 40309 770208 40314 770264
rect 40370 770208 44546 770264
rect 44602 770208 44607 770264
rect 40309 770206 44607 770208
rect 40309 770203 40375 770206
rect 44541 770203 44607 770206
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 39573 768634 39639 768637
rect 42701 768634 42767 768637
rect 39573 768632 42767 768634
rect 39573 768576 39578 768632
rect 39634 768576 42706 768632
rect 42762 768576 42767 768632
rect 39573 768574 42767 768576
rect 39573 768571 39639 768574
rect 42701 768571 42767 768574
rect 35758 768229 35818 768332
rect 35758 768224 35867 768229
rect 35758 768168 35806 768224
rect 35862 768168 35867 768224
rect 35758 768166 35867 768168
rect 35801 768163 35867 768166
rect 32998 767821 33058 767924
rect 32998 767816 33107 767821
rect 32998 767760 33046 767816
rect 33102 767760 33107 767816
rect 32998 767758 33107 767760
rect 33041 767755 33107 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 40726 766596 40786 766700
rect 40718 766532 40724 766596
rect 40788 766532 40794 766596
rect 35758 766189 35818 766292
rect 35758 766184 35867 766189
rect 35758 766128 35806 766184
rect 35862 766128 35867 766184
rect 35758 766126 35867 766128
rect 35801 766123 35867 766126
rect 35758 765781 35818 765884
rect 35758 765776 35867 765781
rect 35758 765720 35806 765776
rect 35862 765720 35867 765776
rect 35758 765718 35867 765720
rect 35801 765715 35867 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 41505 764962 41571 764965
rect 45093 764962 45159 764965
rect 41505 764960 45159 764962
rect 41505 764904 41510 764960
rect 41566 764904 45098 764960
rect 45154 764904 45159 764960
rect 41505 764902 45159 764904
rect 41505 764899 41571 764902
rect 45093 764899 45159 764902
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 41229 764554 41295 764557
rect 45277 764554 45343 764557
rect 41229 764552 45343 764554
rect 41229 764496 41234 764552
rect 41290 764496 45282 764552
rect 45338 764496 45343 764552
rect 41229 764494 45343 764496
rect 41229 764491 41295 764494
rect 45277 764491 45343 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 39757 764146 39823 764149
rect 43253 764146 43319 764149
rect 39757 764144 43319 764146
rect 39757 764088 39762 764144
rect 39818 764088 43258 764144
rect 43314 764088 43319 764144
rect 39757 764086 43319 764088
rect 39757 764083 39823 764086
rect 43253 764083 43319 764086
rect 35758 763333 35818 763844
rect 40861 763738 40927 763741
rect 43069 763738 43135 763741
rect 40861 763736 43135 763738
rect 40861 763680 40866 763736
rect 40922 763680 43074 763736
rect 43130 763680 43135 763736
rect 40861 763678 43135 763680
rect 40861 763675 40927 763678
rect 43069 763675 43135 763678
rect 35758 763328 35867 763333
rect 35758 763272 35806 763328
rect 35862 763272 35867 763328
rect 35758 763270 35867 763272
rect 35801 763267 35867 763270
rect 41505 763330 41571 763333
rect 45553 763330 45619 763333
rect 41505 763328 45619 763330
rect 41505 763272 41510 763328
rect 41566 763272 45558 763328
rect 45614 763272 45619 763328
rect 41505 763270 45619 763272
rect 41505 763267 41571 763270
rect 45553 763267 45619 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 41689 761154 41755 761157
rect 42609 761154 42675 761157
rect 41689 761152 42675 761154
rect 41689 761096 41694 761152
rect 41750 761096 42614 761152
rect 42670 761096 42675 761152
rect 41689 761094 42675 761096
rect 41689 761091 41755 761094
rect 42609 761091 42675 761094
rect 36537 759114 36603 759117
rect 41638 759114 41644 759116
rect 36537 759112 41644 759114
rect 36537 759056 36542 759112
rect 36598 759056 41644 759112
rect 36537 759054 41644 759056
rect 36537 759051 36603 759054
rect 41638 759052 41644 759054
rect 41708 759052 41714 759116
rect 41873 758978 41939 758981
rect 42425 758978 42491 758981
rect 41873 758976 42491 758978
rect 41873 758920 41878 758976
rect 41934 758920 42430 758976
rect 42486 758920 42491 758976
rect 41873 758918 42491 758920
rect 41873 758915 41939 758918
rect 42425 758915 42491 758918
rect 40033 757754 40099 757757
rect 40350 757754 40356 757756
rect 40033 757752 40356 757754
rect 40033 757696 40038 757752
rect 40094 757696 40356 757752
rect 40033 757694 40356 757696
rect 40033 757691 40099 757694
rect 40350 757692 40356 757694
rect 40420 757692 40426 757756
rect 40677 757754 40743 757757
rect 41822 757754 41828 757756
rect 40677 757752 41828 757754
rect 40677 757696 40682 757752
rect 40738 757696 41828 757752
rect 40677 757694 41828 757696
rect 40677 757691 40743 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 38929 757482 38995 757485
rect 43437 757482 43503 757485
rect 38929 757480 43503 757482
rect 38929 757424 38934 757480
rect 38990 757424 43442 757480
rect 43498 757424 43503 757480
rect 38929 757422 43503 757424
rect 38929 757419 38995 757422
rect 43437 757419 43503 757422
rect 41781 757074 41847 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 41830 755445 41890 757011
rect 41830 755440 41939 755445
rect 41830 755384 41878 755440
rect 41934 755384 41939 755440
rect 41830 755382 41939 755384
rect 41873 755379 41939 755382
rect 40350 755108 40356 755172
rect 40420 755170 40426 755172
rect 42517 755170 42583 755173
rect 40420 755168 42583 755170
rect 40420 755112 42522 755168
rect 42578 755112 42583 755168
rect 40420 755110 42583 755112
rect 40420 755108 40426 755110
rect 42517 755107 42583 755110
rect 40902 754836 40908 754900
rect 40972 754898 40978 754900
rect 42006 754898 42012 754900
rect 40972 754838 42012 754898
rect 40972 754836 40978 754838
rect 42006 754836 42012 754838
rect 42076 754836 42082 754900
rect 42057 752994 42123 752997
rect 43437 752994 43503 752997
rect 42057 752992 43503 752994
rect 42057 752936 42062 752992
rect 42118 752936 43442 752992
rect 43498 752936 43503 752992
rect 42057 752934 43503 752936
rect 42057 752931 42123 752934
rect 43437 752931 43503 752934
rect 40718 752116 40724 752180
rect 40788 752178 40794 752180
rect 42374 752178 42380 752180
rect 40788 752118 42380 752178
rect 40788 752116 40794 752118
rect 42374 752116 42380 752118
rect 42444 752116 42450 752180
rect 42057 751634 42123 751637
rect 43621 751634 43687 751637
rect 42057 751632 43687 751634
rect 42057 751576 42062 751632
rect 42118 751576 43626 751632
rect 43682 751576 43687 751632
rect 42057 751574 43687 751576
rect 42057 751571 42123 751574
rect 43621 751571 43687 751574
rect 42057 751090 42123 751093
rect 45093 751090 45159 751093
rect 42057 751088 45159 751090
rect 42057 751032 42062 751088
rect 42118 751032 45098 751088
rect 45154 751032 45159 751088
rect 42057 751030 45159 751032
rect 42057 751027 42123 751030
rect 45093 751027 45159 751030
rect 41965 750412 42031 750413
rect 41965 750408 42012 750412
rect 42076 750410 42082 750412
rect 41965 750352 41970 750408
rect 41965 750348 42012 750352
rect 42076 750350 42122 750410
rect 42076 750348 42082 750350
rect 41965 750347 42031 750348
rect 42425 749596 42491 749597
rect 42374 749532 42380 749596
rect 42444 749594 42491 749596
rect 42444 749592 42536 749594
rect 42486 749536 42536 749592
rect 42444 749534 42536 749536
rect 42444 749532 42491 749534
rect 42425 749531 42491 749532
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 62757 747690 62823 747693
rect 62757 747688 64706 747690
rect 62757 747632 62762 747688
rect 62818 747632 64706 747688
rect 62757 747630 64706 747632
rect 62757 747627 62823 747630
rect 64646 747082 64706 747630
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 64646 745900 64706 746134
rect 41638 745588 41644 745652
rect 41708 745650 41714 745652
rect 41708 745590 42626 745650
rect 41708 745588 41714 745590
rect 42566 745381 42626 745590
rect 41454 745316 41460 745380
rect 41524 745378 41530 745380
rect 42333 745378 42399 745381
rect 41524 745376 42399 745378
rect 41524 745320 42338 745376
rect 42394 745320 42399 745376
rect 41524 745318 42399 745320
rect 41524 745316 41530 745318
rect 42333 745315 42399 745318
rect 42517 745376 42626 745381
rect 42517 745320 42522 745376
rect 42578 745320 42626 745376
rect 42517 745318 42626 745320
rect 42517 745315 42583 745318
rect 41822 744908 41828 744972
rect 41892 744970 41898 744972
rect 42701 744970 42767 744973
rect 41892 744968 42767 744970
rect 41892 744912 42706 744968
rect 42762 744912 42767 744968
rect 41892 744910 42767 744912
rect 41892 744908 41898 744910
rect 42701 744907 42767 744910
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 674414 742460 674420 742524
rect 674484 742522 674490 742524
rect 675385 742522 675451 742525
rect 674484 742520 675451 742522
rect 674484 742464 675390 742520
rect 675446 742464 675451 742520
rect 674484 742462 675451 742464
rect 674484 742460 674490 742462
rect 675385 742459 675451 742462
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 674833 742252 674899 742253
rect 674782 742188 674788 742252
rect 674852 742250 674899 742252
rect 674852 742248 674944 742250
rect 674894 742192 674944 742248
rect 674852 742190 674944 742192
rect 674852 742188 674899 742190
rect 674833 742187 674899 742188
rect 62389 741842 62455 741845
rect 62389 741840 64706 741842
rect 62389 741784 62394 741840
rect 62450 741784 64706 741840
rect 62389 741782 64706 741784
rect 62389 741779 62455 741782
rect 64646 741172 64706 741782
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675201 738170 675267 738173
rect 674668 738168 675267 738170
rect 674668 738112 675206 738168
rect 675262 738112 675267 738168
rect 674668 738110 675267 738112
rect 674668 738108 674674 738110
rect 675201 738107 675267 738110
rect 674925 736402 674991 736405
rect 675109 736402 675175 736405
rect 674925 736400 675175 736402
rect 674925 736344 674930 736400
rect 674986 736344 675114 736400
rect 675170 736344 675175 736400
rect 674925 736342 675175 736344
rect 674925 736339 674991 736342
rect 675109 736339 675175 736342
rect 668945 736130 669011 736133
rect 675477 736130 675543 736133
rect 668945 736128 675543 736130
rect 668945 736072 668950 736128
rect 669006 736072 675482 736128
rect 675538 736072 675543 736128
rect 668945 736070 675543 736072
rect 668945 736067 669011 736070
rect 675477 736067 675543 736070
rect 674782 734980 674788 735044
rect 674852 735042 674858 735044
rect 675293 735042 675359 735045
rect 674852 735040 675359 735042
rect 674852 734984 675298 735040
rect 675354 734984 675359 735040
rect 674852 734982 675359 734984
rect 674852 734980 674858 734982
rect 675293 734979 675359 734982
rect 649950 734226 650010 734402
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 670969 734226 671035 734229
rect 675477 734226 675543 734229
rect 670969 734224 675543 734226
rect 670969 734168 670974 734224
rect 671030 734168 675482 734224
rect 675538 734168 675543 734224
rect 670969 734166 675543 734168
rect 670969 734163 671035 734166
rect 675477 734163 675543 734166
rect 670509 733818 670575 733821
rect 675477 733818 675543 733821
rect 670509 733816 675543 733818
rect 670509 733760 670514 733816
rect 670570 733760 675482 733816
rect 675538 733760 675543 733816
rect 670509 733758 675543 733760
rect 670509 733755 670575 733758
rect 675477 733755 675543 733758
rect 649950 733002 650010 733220
rect 651465 733002 651531 733005
rect 649950 733000 651531 733002
rect 649950 732944 651470 733000
rect 651526 732944 651531 733000
rect 649950 732942 651531 732944
rect 651465 732939 651531 732942
rect 675753 733002 675819 733005
rect 676806 733002 676812 733004
rect 675753 733000 676812 733002
rect 675753 732944 675758 733000
rect 675814 732944 676812 733000
rect 675753 732942 676812 732944
rect 675753 732939 675819 732942
rect 676806 732940 676812 732942
rect 676876 732940 676882 733004
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 43437 731370 43503 731373
rect 41492 731368 43503 731370
rect 41492 731312 43442 731368
rect 43498 731312 43503 731368
rect 41492 731310 43503 731312
rect 43437 731307 43503 731310
rect 651465 731098 651531 731101
rect 649950 731096 651531 731098
rect 649950 731040 651470 731096
rect 651526 731040 651531 731096
rect 649950 731038 651531 731040
rect 46197 730962 46263 730965
rect 41492 730960 46263 730962
rect 41492 730904 46202 730960
rect 46258 730904 46263 730960
rect 41492 730902 46263 730904
rect 46197 730899 46263 730902
rect 649950 730856 650010 731038
rect 651465 731035 651531 731038
rect 42241 730554 42307 730557
rect 41492 730552 42307 730554
rect 41492 730496 42246 730552
rect 42302 730496 42307 730552
rect 41492 730494 42307 730496
rect 42241 730491 42307 730494
rect 44909 730146 44975 730149
rect 41492 730144 44975 730146
rect 41492 730088 44914 730144
rect 44970 730088 44975 730144
rect 41492 730086 44975 730088
rect 44909 730083 44975 730086
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 45185 729738 45251 729741
rect 41492 729736 45251 729738
rect 41492 729680 45190 729736
rect 45246 729680 45251 729736
rect 41492 729678 45251 729680
rect 45185 729675 45251 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 43069 729330 43135 729333
rect 41492 729328 43135 729330
rect 41492 729272 43074 729328
rect 43130 729272 43135 729328
rect 41492 729270 43135 729272
rect 43069 729267 43135 729270
rect 41278 728687 41338 728892
rect 40861 728684 40927 728687
rect 40861 728682 40970 728684
rect 40861 728626 40866 728682
rect 40922 728626 40970 728682
rect 40861 728621 40970 728626
rect 41278 728682 41387 728687
rect 41278 728626 41326 728682
rect 41382 728626 41387 728682
rect 41278 728624 41387 728626
rect 41321 728621 41387 728624
rect 40910 728484 40970 728621
rect 651465 728514 651531 728517
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 651465 728451 651531 728454
rect 675518 728316 675524 728380
rect 675588 728378 675594 728380
rect 675753 728378 675819 728381
rect 675588 728376 675819 728378
rect 675588 728320 675758 728376
rect 675814 728320 675819 728376
rect 675588 728318 675819 728320
rect 675588 728316 675594 728318
rect 675753 728315 675819 728318
rect 44173 728106 44239 728109
rect 41492 728104 44239 728106
rect 41492 728048 44178 728104
rect 44234 728048 44239 728104
rect 41492 728046 44239 728048
rect 44173 728043 44239 728046
rect 675334 728044 675340 728108
rect 675404 728106 675410 728108
rect 675937 728106 676003 728109
rect 675404 728104 676003 728106
rect 675404 728048 675942 728104
rect 675998 728048 676003 728104
rect 675404 728046 676003 728048
rect 675404 728044 675410 728046
rect 675937 728043 676003 728046
rect 44357 727698 44423 727701
rect 41492 727696 44423 727698
rect 41492 727640 44362 727696
rect 44418 727640 44423 727696
rect 41492 727638 44423 727640
rect 44357 727635 44423 727638
rect 41321 727460 41387 727463
rect 41278 727458 41387 727460
rect 41278 727402 41326 727458
rect 41382 727402 41387 727458
rect 41278 727397 41387 727402
rect 41278 727260 41338 727397
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 41278 726239 41338 726444
rect 674230 726412 674236 726476
rect 674300 726474 674306 726476
rect 684125 726474 684191 726477
rect 674300 726472 684191 726474
rect 674300 726416 684130 726472
rect 684186 726416 684191 726472
rect 674300 726414 684191 726416
rect 674300 726412 674306 726414
rect 684125 726411 684191 726414
rect 39297 726236 39363 726239
rect 39254 726234 39363 726236
rect 39254 726178 39302 726234
rect 39358 726178 39363 726234
rect 39254 726173 39363 726178
rect 41278 726234 41387 726239
rect 41278 726178 41326 726234
rect 41382 726178 41387 726234
rect 41278 726176 41387 726178
rect 41321 726173 41387 726176
rect 39254 726036 39314 726173
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 41137 725250 41203 725253
rect 41124 725248 41203 725250
rect 41124 725192 41142 725248
rect 41198 725192 41203 725248
rect 41124 725190 41203 725192
rect 41137 725187 41203 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 31661 724434 31727 724437
rect 31661 724432 31740 724434
rect 31661 724376 31666 724432
rect 31722 724376 31740 724432
rect 31661 724374 31740 724376
rect 31661 724371 31727 724374
rect 32949 724026 33015 724029
rect 32949 724024 33028 724026
rect 32949 723968 32954 724024
rect 33010 723968 33028 724024
rect 32949 723966 33028 723968
rect 32949 723963 33015 723966
rect 43621 723618 43687 723621
rect 41492 723616 43687 723618
rect 41492 723560 43626 723616
rect 43682 723560 43687 723616
rect 41492 723558 43687 723560
rect 43621 723555 43687 723558
rect 33777 723210 33843 723213
rect 33764 723208 33843 723210
rect 33764 723152 33782 723208
rect 33838 723152 33843 723208
rect 33764 723150 33843 723152
rect 33777 723147 33843 723150
rect 674833 723210 674899 723213
rect 675150 723210 675156 723212
rect 674833 723208 675156 723210
rect 674833 723152 674838 723208
rect 674894 723152 675156 723208
rect 674833 723150 675156 723152
rect 674833 723147 674899 723150
rect 675150 723148 675156 723150
rect 675220 723148 675226 723212
rect 44449 722802 44515 722805
rect 41492 722800 44515 722802
rect 41492 722744 44454 722800
rect 44510 722744 44515 722800
rect 41492 722742 44515 722744
rect 44449 722739 44515 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 40726 721772 40786 721956
rect 674097 721850 674163 721853
rect 673318 721848 674163 721850
rect 673318 721792 674102 721848
rect 674158 721792 674163 721848
rect 673318 721790 674163 721792
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 673318 721581 673378 721790
rect 674097 721787 674163 721790
rect 675017 721716 675083 721717
rect 674966 721652 674972 721716
rect 675036 721714 675083 721716
rect 675036 721712 675128 721714
rect 675078 721656 675128 721712
rect 675036 721654 675128 721656
rect 675036 721652 675083 721654
rect 675017 721651 675083 721652
rect 44633 721578 44699 721581
rect 41492 721576 44699 721578
rect 41492 721520 44638 721576
rect 44694 721520 44699 721576
rect 41492 721518 44699 721520
rect 44633 721515 44699 721518
rect 673269 721576 673378 721581
rect 673269 721520 673274 721576
rect 673330 721520 673378 721576
rect 673269 721518 673378 721520
rect 673269 721515 673335 721518
rect 47209 721170 47275 721173
rect 41492 721168 47275 721170
rect 41492 721112 47214 721168
rect 47270 721112 47275 721168
rect 41492 721110 47275 721112
rect 47209 721107 47275 721110
rect 41094 720357 41154 720732
rect 41094 720352 41203 720357
rect 41094 720324 41142 720352
rect 41124 720296 41142 720324
rect 41198 720296 41203 720352
rect 41124 720294 41203 720296
rect 41137 720291 41203 720294
rect 47025 719946 47091 719949
rect 41492 719944 47091 719946
rect 41492 719888 47030 719944
rect 47086 719888 47091 719944
rect 41492 719886 47091 719888
rect 47025 719883 47091 719886
rect 41321 719266 41387 719269
rect 42517 719266 42583 719269
rect 41321 719264 42583 719266
rect 41321 719208 41326 719264
rect 41382 719208 42522 719264
rect 42578 719208 42583 719264
rect 41321 719206 42583 719208
rect 41321 719203 41387 719206
rect 42517 719203 42583 719206
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 31661 718314 31727 718317
rect 41638 718314 41644 718316
rect 31661 718312 41644 718314
rect 31661 718256 31666 718312
rect 31722 718256 41644 718312
rect 31661 718254 41644 718256
rect 31661 718251 31727 718254
rect 41638 718252 41644 718254
rect 41708 718252 41714 718316
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 39297 716138 39363 716141
rect 41822 716138 41828 716140
rect 39297 716136 41828 716138
rect 39297 716080 39302 716136
rect 39358 716080 41828 716136
rect 39297 716078 41828 716080
rect 39297 716075 39363 716078
rect 41822 716076 41828 716078
rect 41892 716076 41898 716140
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 42701 716002 42767 716005
rect 42014 716000 42767 716002
rect 42014 715944 42706 716000
rect 42762 715944 42767 716000
rect 42014 715942 42767 715944
rect 40585 715730 40651 715733
rect 42014 715730 42074 715942
rect 42701 715939 42767 715942
rect 40585 715728 42074 715730
rect 40585 715672 40590 715728
rect 40646 715672 42074 715728
rect 40585 715670 42074 715672
rect 674005 715730 674071 715733
rect 674005 715728 676292 715730
rect 674005 715672 674010 715728
rect 674066 715672 676292 715728
rect 674005 715670 676292 715672
rect 40585 715667 40651 715670
rect 674005 715667 674071 715670
rect 40401 715458 40467 715461
rect 42241 715458 42307 715461
rect 40401 715456 42307 715458
rect 40401 715400 40406 715456
rect 40462 715400 42246 715456
rect 42302 715400 42307 715456
rect 40401 715398 42307 715400
rect 40401 715395 40467 715398
rect 42241 715395 42307 715398
rect 674005 715322 674071 715325
rect 674005 715320 676292 715322
rect 674005 715264 674010 715320
rect 674066 715264 676292 715320
rect 674005 715262 676292 715264
rect 674005 715259 674071 715262
rect 674005 715050 674071 715053
rect 674005 715048 674482 715050
rect 674005 714992 674010 715048
rect 674066 714992 674482 715048
rect 674005 714990 674482 714992
rect 674005 714987 674071 714990
rect 41505 714914 41571 714917
rect 42793 714914 42859 714917
rect 41505 714912 42859 714914
rect 41505 714856 41510 714912
rect 41566 714856 42798 714912
rect 42854 714856 42859 714912
rect 41505 714854 42859 714856
rect 674422 714914 674482 714990
rect 674422 714854 676292 714914
rect 41505 714851 41571 714854
rect 42793 714851 42859 714854
rect 674005 714506 674071 714509
rect 674005 714504 676292 714506
rect 674005 714448 674010 714504
rect 674066 714448 676292 714504
rect 674005 714446 676292 714448
rect 674005 714443 674071 714446
rect 41229 714236 41295 714237
rect 41229 714234 41276 714236
rect 41184 714232 41276 714234
rect 41184 714176 41234 714232
rect 41184 714174 41276 714176
rect 41229 714172 41276 714174
rect 41340 714172 41346 714236
rect 41229 714171 41295 714172
rect 672717 714098 672783 714101
rect 672717 714096 676292 714098
rect 672717 714040 672722 714096
rect 672778 714040 676292 714096
rect 672717 714038 676292 714040
rect 672717 714035 672783 714038
rect 674005 713690 674071 713693
rect 674005 713688 676292 713690
rect 674005 713632 674010 713688
rect 674066 713632 676292 713688
rect 674005 713630 676292 713632
rect 674005 713627 674071 713630
rect 674005 713282 674071 713285
rect 674005 713280 676292 713282
rect 674005 713224 674010 713280
rect 674066 713224 676292 713280
rect 674005 713222 676292 713224
rect 674005 713219 674071 713222
rect 673085 712874 673151 712877
rect 673085 712872 676292 712874
rect 673085 712816 673090 712872
rect 673146 712816 676292 712872
rect 673085 712814 676292 712816
rect 673085 712811 673151 712814
rect 674005 712466 674071 712469
rect 674005 712464 676292 712466
rect 674005 712408 674010 712464
rect 674066 712408 676292 712464
rect 674005 712406 676292 712408
rect 674005 712403 674071 712406
rect 41270 712132 41276 712196
rect 41340 712194 41346 712196
rect 41781 712194 41847 712197
rect 41340 712192 41847 712194
rect 41340 712136 41786 712192
rect 41842 712136 41847 712192
rect 41340 712134 41847 712136
rect 41340 712132 41346 712134
rect 41781 712131 41847 712134
rect 675661 712058 675727 712061
rect 675661 712056 676292 712058
rect 675661 712000 675666 712056
rect 675722 712000 676292 712056
rect 675661 711998 676292 712000
rect 675661 711995 675727 711998
rect 683297 711650 683363 711653
rect 683284 711648 683363 711650
rect 683284 711592 683302 711648
rect 683358 711592 683363 711648
rect 683284 711590 683363 711592
rect 683297 711587 683363 711590
rect 675845 711242 675911 711245
rect 675845 711240 676292 711242
rect 675845 711184 675850 711240
rect 675906 711184 676292 711240
rect 675845 711182 676292 711184
rect 675845 711179 675911 711182
rect 42057 710834 42123 710837
rect 42885 710834 42951 710837
rect 42057 710832 42951 710834
rect 42057 710776 42062 710832
rect 42118 710776 42890 710832
rect 42946 710776 42951 710832
rect 42057 710774 42951 710776
rect 42057 710771 42123 710774
rect 42885 710771 42951 710774
rect 676029 710834 676095 710837
rect 676029 710832 676292 710834
rect 676029 710776 676034 710832
rect 676090 710776 676292 710832
rect 676029 710774 676292 710776
rect 676029 710771 676095 710774
rect 676029 710426 676095 710429
rect 676029 710424 676292 710426
rect 676029 710368 676034 710424
rect 676090 710368 676292 710424
rect 676029 710366 676292 710368
rect 676029 710363 676095 710366
rect 674005 710018 674071 710021
rect 674005 710016 676292 710018
rect 674005 709960 674010 710016
rect 674066 709960 676292 710016
rect 674005 709958 676292 709960
rect 674005 709955 674071 709958
rect 674005 709610 674071 709613
rect 674005 709608 676292 709610
rect 674005 709552 674010 709608
rect 674066 709552 676292 709608
rect 674005 709550 676292 709552
rect 674005 709547 674071 709550
rect 672901 709202 672967 709205
rect 672901 709200 676292 709202
rect 672901 709144 672906 709200
rect 672962 709144 676292 709200
rect 672901 709142 676292 709144
rect 672901 709139 672967 709142
rect 684125 708794 684191 708797
rect 684125 708792 684204 708794
rect 684125 708736 684130 708792
rect 684186 708736 684204 708792
rect 684125 708734 684204 708736
rect 684125 708731 684191 708734
rect 42057 708386 42123 708389
rect 44449 708386 44515 708389
rect 683481 708386 683547 708389
rect 42057 708384 44515 708386
rect 42057 708328 42062 708384
rect 42118 708328 44454 708384
rect 44510 708328 44515 708384
rect 42057 708326 44515 708328
rect 683468 708384 683547 708386
rect 683468 708328 683486 708384
rect 683542 708328 683547 708384
rect 683468 708326 683547 708328
rect 42057 708323 42123 708326
rect 44449 708323 44515 708326
rect 683481 708323 683547 708326
rect 677174 707950 677180 708014
rect 677244 707950 677250 708014
rect 677182 707948 677242 707950
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 40718 707100 40724 707164
rect 40788 707162 40794 707164
rect 41781 707162 41847 707165
rect 40788 707160 41847 707162
rect 40788 707104 41786 707160
rect 41842 707104 41847 707160
rect 40788 707102 41847 707104
rect 40788 707100 40794 707102
rect 41781 707099 41847 707102
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 675845 706754 675911 706757
rect 675845 706752 676292 706754
rect 675845 706696 675850 706752
rect 675906 706696 676292 706752
rect 675845 706694 676292 706696
rect 675845 706691 675911 706694
rect 673269 706346 673335 706349
rect 673269 706344 676292 706346
rect 673269 706288 673274 706344
rect 673330 706288 676292 706344
rect 673269 706286 676292 706288
rect 673269 706283 673335 706286
rect 677182 705530 677242 705908
rect 683113 705530 683179 705533
rect 677182 705528 683179 705530
rect 677182 705500 683118 705528
rect 677212 705472 683118 705500
rect 683174 705472 683179 705528
rect 677212 705470 683179 705472
rect 683113 705467 683179 705470
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 40534 704244 40540 704308
rect 40604 704306 40610 704308
rect 41781 704306 41847 704309
rect 40604 704304 41847 704306
rect 40604 704248 41786 704304
rect 41842 704248 41847 704304
rect 40604 704246 41847 704248
rect 40604 704244 40610 704246
rect 41781 704243 41847 704246
rect 64646 703860 64706 704382
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 64646 702678 64706 703294
rect 41822 702068 41828 702132
rect 41892 702130 41898 702132
rect 42701 702130 42767 702133
rect 41892 702128 42767 702130
rect 41892 702072 42706 702128
rect 42762 702072 42767 702128
rect 41892 702070 42767 702072
rect 41892 702068 41898 702070
rect 42701 702067 42767 702070
rect 41638 701796 41644 701860
rect 41708 701858 41714 701860
rect 42241 701858 42307 701861
rect 41708 701856 42307 701858
rect 41708 701800 42246 701856
rect 42302 701800 42307 701856
rect 41708 701798 42307 701800
rect 41708 701796 41714 701798
rect 42241 701795 42307 701798
rect 62205 701314 62271 701317
rect 64646 701314 64706 701496
rect 62205 701312 64706 701314
rect 62205 701256 62210 701312
rect 62266 701256 64706 701312
rect 62205 701254 64706 701256
rect 62205 701251 62271 701254
rect 62757 700906 62823 700909
rect 62757 700904 64706 700906
rect 62757 700848 62762 700904
rect 62818 700848 64706 700904
rect 62757 700846 64706 700848
rect 62757 700843 62823 700846
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 64646 700314 64706 700846
rect 61377 699682 61443 699685
rect 61377 699680 64706 699682
rect 61377 699624 61382 699680
rect 61438 699624 64706 699680
rect 61377 699622 64706 699624
rect 61377 699619 61443 699622
rect 64646 699132 64706 699622
rect 62113 698186 62179 698189
rect 62113 698184 64706 698186
rect 62113 698128 62118 698184
rect 62174 698128 64706 698184
rect 62113 698126 64706 698128
rect 62113 698123 62179 698126
rect 64646 697950 64706 698126
rect 673177 697234 673243 697237
rect 675109 697234 675175 697237
rect 673177 697232 675175 697234
rect 673177 697176 673182 697232
rect 673238 697176 675114 697232
rect 675170 697176 675175 697232
rect 673177 697174 675175 697176
rect 673177 697171 673243 697174
rect 675109 697171 675175 697174
rect 673729 696962 673795 696965
rect 675293 696962 675359 696965
rect 673729 696960 675359 696962
rect 673729 696904 673734 696960
rect 673790 696904 675298 696960
rect 675354 696904 675359 696960
rect 673729 696902 675359 696904
rect 673729 696899 673795 696902
rect 675293 696899 675359 696902
rect 674230 696628 674236 696692
rect 674300 696690 674306 696692
rect 675109 696690 675175 696693
rect 674300 696688 675175 696690
rect 674300 696632 675114 696688
rect 675170 696632 675175 696688
rect 674300 696630 675175 696632
rect 674300 696628 674306 696630
rect 675109 696627 675175 696630
rect 672349 695466 672415 695469
rect 675293 695466 675359 695469
rect 672349 695464 675359 695466
rect 672349 695408 672354 695464
rect 672410 695408 675298 695464
rect 675354 695408 675359 695464
rect 672349 695406 675359 695408
rect 672349 695403 672415 695406
rect 675293 695403 675359 695406
rect 671797 690434 671863 690437
rect 675109 690434 675175 690437
rect 671797 690432 675175 690434
rect 671797 690376 671802 690432
rect 671858 690376 675114 690432
rect 675170 690376 675175 690432
rect 671797 690374 675175 690376
rect 671797 690371 671863 690374
rect 675109 690371 675175 690374
rect 673729 690162 673795 690165
rect 674925 690162 674991 690165
rect 673729 690160 674991 690162
rect 673729 690104 673734 690160
rect 673790 690104 674930 690160
rect 674986 690104 674991 690160
rect 673729 690102 674991 690104
rect 673729 690099 673795 690102
rect 674925 690099 674991 690102
rect 649950 689482 650010 689980
rect 668025 689890 668091 689893
rect 675385 689890 675451 689893
rect 668025 689888 675451 689890
rect 668025 689832 668030 689888
rect 668086 689832 675390 689888
rect 675446 689832 675451 689888
rect 668025 689830 675451 689832
rect 668025 689827 668091 689830
rect 675385 689827 675451 689830
rect 651465 689482 651531 689485
rect 649950 689480 651531 689482
rect 649950 689424 651470 689480
rect 651526 689424 651531 689480
rect 649950 689422 651531 689424
rect 651465 689419 651531 689422
rect 674097 689482 674163 689485
rect 675109 689482 675175 689485
rect 674097 689480 675175 689482
rect 674097 689424 674102 689480
rect 674158 689424 675114 689480
rect 675170 689424 675175 689480
rect 674097 689422 675175 689424
rect 674097 689419 674163 689422
rect 675109 689419 675175 689422
rect 670693 689210 670759 689213
rect 675109 689210 675175 689213
rect 670693 689208 675175 689210
rect 670693 689152 670698 689208
rect 670754 689152 675114 689208
rect 675170 689152 675175 689208
rect 670693 689150 675175 689152
rect 670693 689147 670759 689150
rect 675109 689147 675175 689150
rect 649980 688802 650562 688828
rect 651649 688802 651715 688805
rect 649980 688800 651715 688802
rect 649980 688768 651654 688800
rect 650502 688744 651654 688768
rect 651710 688744 651715 688800
rect 650502 688742 651715 688744
rect 651649 688739 651715 688742
rect 673729 688802 673795 688805
rect 674925 688802 674991 688805
rect 673729 688800 674991 688802
rect 673729 688744 673734 688800
rect 673790 688744 674930 688800
rect 674986 688744 674991 688800
rect 673729 688742 674991 688744
rect 673729 688739 673795 688742
rect 674925 688739 674991 688742
rect 42701 688122 42767 688125
rect 41492 688120 42767 688122
rect 41492 688064 42706 688120
rect 42762 688064 42767 688120
rect 41492 688062 42767 688064
rect 42701 688059 42767 688062
rect 673729 688122 673795 688125
rect 674281 688122 674347 688125
rect 673729 688120 674347 688122
rect 673729 688064 673734 688120
rect 673790 688064 674286 688120
rect 674342 688064 674347 688120
rect 673729 688062 674347 688064
rect 673729 688059 673795 688062
rect 674281 688059 674347 688062
rect 672901 687850 672967 687853
rect 675109 687850 675175 687853
rect 672901 687848 675175 687850
rect 672901 687792 672906 687848
rect 672962 687792 675114 687848
rect 675170 687792 675175 687848
rect 672901 687790 675175 687792
rect 672901 687787 672967 687790
rect 675109 687787 675175 687790
rect 44817 687714 44883 687717
rect 41492 687712 44883 687714
rect 41492 687656 44822 687712
rect 44878 687656 44883 687712
rect 41492 687654 44883 687656
rect 44817 687651 44883 687654
rect 649950 687442 650010 687616
rect 673545 687578 673611 687581
rect 674649 687578 674715 687581
rect 673545 687576 674715 687578
rect 673545 687520 673550 687576
rect 673606 687520 674654 687576
rect 674710 687520 674715 687576
rect 673545 687518 674715 687520
rect 673545 687515 673611 687518
rect 674649 687515 674715 687518
rect 651465 687442 651531 687445
rect 649950 687440 651531 687442
rect 649950 687384 651470 687440
rect 651526 687384 651531 687440
rect 649950 687382 651531 687384
rect 651465 687379 651531 687382
rect 43437 687306 43503 687309
rect 41492 687304 43503 687306
rect 41492 687248 43442 687304
rect 43498 687248 43503 687304
rect 41492 687246 43503 687248
rect 43437 687243 43503 687246
rect 41137 686898 41203 686901
rect 41124 686896 41203 686898
rect 41124 686840 41142 686896
rect 41198 686840 41203 686896
rect 41124 686838 41203 686840
rect 41137 686835 41203 686838
rect 651465 686762 651531 686765
rect 649950 686760 651531 686762
rect 649950 686704 651470 686760
rect 651526 686704 651531 686760
rect 649950 686702 651531 686704
rect 40861 686490 40927 686493
rect 40861 686488 40940 686490
rect 40861 686432 40866 686488
rect 40922 686432 40940 686488
rect 649950 686434 650010 686702
rect 651465 686699 651531 686702
rect 668209 686490 668275 686493
rect 675477 686490 675543 686493
rect 668209 686488 675543 686490
rect 40861 686430 40940 686432
rect 668209 686432 668214 686488
rect 668270 686432 675482 686488
rect 675538 686432 675543 686488
rect 668209 686430 675543 686432
rect 40861 686427 40927 686430
rect 668209 686427 668275 686430
rect 675477 686427 675543 686430
rect 674925 686218 674991 686221
rect 675334 686218 675340 686220
rect 674925 686216 675340 686218
rect 674925 686160 674930 686216
rect 674986 686160 675340 686216
rect 674925 686158 675340 686160
rect 674925 686155 674991 686158
rect 675334 686156 675340 686158
rect 675404 686156 675410 686220
rect 41278 685915 41338 686052
rect 41045 685912 41111 685915
rect 41045 685910 41154 685912
rect 41045 685854 41050 685910
rect 41106 685854 41154 685910
rect 41045 685849 41154 685854
rect 41278 685910 41387 685915
rect 41278 685854 41326 685910
rect 41382 685854 41387 685910
rect 41278 685852 41387 685854
rect 41321 685849 41387 685852
rect 41094 685644 41154 685849
rect 669773 685810 669839 685813
rect 669773 685808 673562 685810
rect 669773 685752 669778 685808
rect 669834 685752 673562 685808
rect 669773 685750 673562 685752
rect 669773 685747 669839 685750
rect 673502 685674 673562 685750
rect 675477 685674 675543 685677
rect 673502 685672 675543 685674
rect 673502 685616 675482 685672
rect 675538 685616 675543 685672
rect 673502 685614 675543 685616
rect 675477 685611 675543 685614
rect 672165 685402 672231 685405
rect 675109 685402 675175 685405
rect 672165 685400 675175 685402
rect 672165 685344 672170 685400
rect 672226 685344 675114 685400
rect 675170 685344 675175 685400
rect 672165 685342 675175 685344
rect 672165 685339 672231 685342
rect 675109 685339 675175 685342
rect 44265 685266 44331 685269
rect 651465 685266 651531 685269
rect 41492 685264 44331 685266
rect 41492 685208 44270 685264
rect 44326 685208 44331 685264
rect 41492 685206 44331 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 44265 685203 44331 685206
rect 651465 685203 651531 685206
rect 40769 684688 40835 684691
rect 41462 684690 41522 684828
rect 40726 684686 40835 684688
rect 40726 684630 40774 684686
rect 40830 684630 40835 684686
rect 40726 684625 40835 684630
rect 41454 684626 41460 684690
rect 41524 684626 41530 684690
rect 40726 684420 40786 684625
rect 652569 684450 652635 684453
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 41689 684314 41755 684317
rect 44449 684314 44515 684317
rect 41689 684312 44515 684314
rect 41689 684256 41694 684312
rect 41750 684256 44454 684312
rect 44510 684256 44515 684312
rect 41689 684254 44515 684256
rect 41689 684251 41755 684254
rect 44449 684251 44515 684254
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 41137 684042 41203 684045
rect 41124 684040 41203 684042
rect 41124 683984 41142 684040
rect 41198 683984 41203 684040
rect 41124 683982 41203 683984
rect 41137 683979 41203 683982
rect 41822 683844 41828 683908
rect 41892 683906 41898 683908
rect 44633 683906 44699 683909
rect 41892 683904 44699 683906
rect 41892 683848 44638 683904
rect 44694 683848 44699 683904
rect 41892 683846 44699 683848
rect 41892 683844 41898 683846
rect 44633 683843 44699 683846
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 41321 683464 41387 683467
rect 41278 683462 41387 683464
rect 41278 683406 41326 683462
rect 41382 683406 41387 683462
rect 41278 683401 41387 683406
rect 41278 683196 41338 683401
rect 40953 682818 41019 682821
rect 40940 682816 41019 682818
rect 40940 682760 40958 682816
rect 41014 682760 41019 682816
rect 40940 682758 41019 682760
rect 40953 682755 41019 682758
rect 41321 682410 41387 682413
rect 41308 682408 41387 682410
rect 41308 682352 41326 682408
rect 41382 682352 41387 682408
rect 41308 682350 41387 682352
rect 41321 682347 41387 682350
rect 35157 682002 35223 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 35157 681939 35223 681942
rect 42241 681594 42307 681597
rect 41492 681592 42307 681594
rect 41492 681536 42246 681592
rect 42302 681536 42307 681592
rect 41492 681534 42307 681536
rect 42241 681531 42307 681534
rect 32397 681186 32463 681189
rect 32397 681184 32476 681186
rect 32397 681128 32402 681184
rect 32458 681128 32476 681184
rect 32397 681126 32476 681128
rect 32397 681123 32463 681126
rect 33777 680778 33843 680781
rect 33764 680776 33843 680778
rect 33764 680720 33782 680776
rect 33838 680720 33843 680776
rect 33764 680718 33843 680720
rect 33777 680715 33843 680718
rect 43621 680370 43687 680373
rect 41492 680368 43687 680370
rect 41492 680312 43626 680368
rect 43682 680312 43687 680368
rect 41492 680310 43687 680312
rect 43621 680307 43687 680310
rect 41137 679962 41203 679965
rect 41124 679960 41203 679962
rect 41124 679904 41142 679960
rect 41198 679904 41203 679960
rect 41124 679902 41203 679904
rect 41137 679899 41203 679902
rect 43989 679554 44055 679557
rect 41492 679552 44055 679554
rect 41492 679496 43994 679552
rect 44050 679496 44055 679552
rect 41492 679494 44055 679496
rect 43989 679491 44055 679494
rect 40542 678992 40602 679116
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 676070 678948 676076 679012
rect 676140 679010 676146 679012
rect 680997 679010 681063 679013
rect 676140 679008 681063 679010
rect 676140 678952 681002 679008
rect 681058 678952 681063 679008
rect 676140 678950 681063 678952
rect 676140 678948 676146 678950
rect 680997 678947 681063 678950
rect 40726 678708 40786 678928
rect 41781 678876 41847 678877
rect 41781 678872 41828 678876
rect 41892 678874 41898 678876
rect 41781 678816 41786 678872
rect 41781 678812 41828 678816
rect 41892 678814 41938 678874
rect 41892 678812 41898 678814
rect 41781 678811 41847 678812
rect 41781 678330 41847 678333
rect 41492 678328 41847 678330
rect 41492 678272 41786 678328
rect 41842 678272 41847 678328
rect 41492 678270 41847 678272
rect 41781 678267 41847 678270
rect 43069 677922 43135 677925
rect 41492 677920 43135 677922
rect 41492 677864 43074 677920
rect 43130 677864 43135 677920
rect 41492 677862 43135 677864
rect 43069 677859 43135 677862
rect 40953 677754 41019 677755
rect 40902 677752 40908 677754
rect 40862 677692 40908 677752
rect 40972 677750 41019 677754
rect 41014 677694 41019 677750
rect 40902 677690 40908 677692
rect 40972 677690 41019 677694
rect 40953 677689 41019 677690
rect 39990 677109 40050 677484
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 43437 676698 43503 676701
rect 41492 676696 43503 676698
rect 41492 676640 43442 676696
rect 43498 676640 43503 676696
rect 41492 676638 43503 676640
rect 43437 676635 43503 676638
rect 32397 672754 32463 672757
rect 41822 672754 41828 672756
rect 32397 672752 41828 672754
rect 32397 672696 32402 672752
rect 32458 672696 41828 672752
rect 32397 672694 41828 672696
rect 32397 672691 32463 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 39941 672482 40007 672485
rect 41086 672482 41092 672484
rect 39941 672480 41092 672482
rect 39941 672424 39946 672480
rect 40002 672424 41092 672480
rect 39941 672422 41092 672424
rect 39941 672419 40007 672422
rect 41086 672420 41092 672422
rect 41156 672420 41162 672484
rect 673913 671666 673979 671669
rect 674741 671666 674807 671669
rect 673913 671664 674807 671666
rect 673913 671608 673918 671664
rect 673974 671608 674746 671664
rect 674802 671608 674807 671664
rect 673913 671606 674807 671608
rect 673913 671603 673979 671606
rect 674741 671603 674807 671606
rect 37917 671530 37983 671533
rect 40350 671530 40356 671532
rect 37917 671528 40356 671530
rect 37917 671472 37922 671528
rect 37978 671472 40356 671528
rect 37917 671470 40356 671472
rect 37917 671467 37983 671470
rect 40350 671468 40356 671470
rect 40420 671468 40426 671532
rect 673545 671394 673611 671397
rect 673545 671392 676292 671394
rect 673545 671336 673550 671392
rect 673606 671336 676292 671392
rect 673545 671334 676292 671336
rect 673545 671331 673611 671334
rect 38837 670986 38903 670989
rect 42517 670986 42583 670989
rect 38837 670984 42583 670986
rect 38837 670928 38842 670984
rect 38898 670928 42522 670984
rect 42578 670928 42583 670984
rect 38837 670926 42583 670928
rect 38837 670923 38903 670926
rect 42517 670923 42583 670926
rect 673913 670986 673979 670989
rect 673913 670984 676292 670986
rect 673913 670928 673918 670984
rect 673974 670928 676292 670984
rect 673913 670926 676292 670928
rect 673913 670923 673979 670926
rect 673545 670578 673611 670581
rect 673545 670576 676292 670578
rect 673545 670520 673550 670576
rect 673606 670520 676292 670576
rect 673545 670518 676292 670520
rect 673545 670515 673611 670518
rect 673913 670170 673979 670173
rect 673913 670168 676292 670170
rect 673913 670112 673918 670168
rect 673974 670112 676292 670168
rect 673913 670110 676292 670112
rect 673913 670107 673979 670110
rect 673913 669762 673979 669765
rect 673913 669760 676292 669762
rect 673913 669704 673918 669760
rect 673974 669704 676292 669760
rect 673913 669702 676292 669704
rect 673913 669699 673979 669702
rect 672717 669490 672783 669493
rect 672717 669488 676322 669490
rect 672717 669432 672722 669488
rect 672778 669432 676322 669488
rect 672717 669430 676322 669432
rect 672717 669427 672783 669430
rect 676262 669324 676322 669430
rect 41086 669020 41092 669084
rect 41156 669082 41162 669084
rect 41781 669082 41847 669085
rect 41156 669080 41847 669082
rect 41156 669024 41786 669080
rect 41842 669024 41847 669080
rect 41156 669022 41847 669024
rect 41156 669020 41162 669022
rect 41781 669019 41847 669022
rect 673545 668946 673611 668949
rect 673545 668944 676292 668946
rect 673545 668888 673550 668944
rect 673606 668888 676292 668944
rect 673545 668886 676292 668888
rect 673545 668883 673611 668886
rect 673913 668538 673979 668541
rect 673913 668536 676292 668538
rect 673913 668480 673918 668536
rect 673974 668480 676292 668536
rect 673913 668478 676292 668480
rect 673913 668475 673979 668478
rect 673913 668130 673979 668133
rect 673913 668128 676292 668130
rect 673913 668072 673918 668128
rect 673974 668072 676292 668128
rect 673913 668070 676292 668072
rect 673913 668067 673979 668070
rect 673913 667722 673979 667725
rect 673913 667720 676292 667722
rect 673913 667664 673918 667720
rect 673974 667664 676292 667720
rect 673913 667662 676292 667664
rect 673913 667659 673979 667662
rect 673545 667314 673611 667317
rect 673545 667312 676292 667314
rect 673545 667256 673550 667312
rect 673606 667256 676292 667312
rect 673545 667254 676292 667256
rect 673545 667251 673611 667254
rect 675293 666906 675359 666909
rect 675293 666904 676292 666906
rect 675293 666848 675298 666904
rect 675354 666848 676292 666904
rect 675293 666846 676292 666848
rect 675293 666843 675359 666846
rect 42057 666634 42123 666637
rect 45001 666634 45067 666637
rect 42057 666632 45067 666634
rect 42057 666576 42062 666632
rect 42118 666576 45006 666632
rect 45062 666576 45067 666632
rect 42057 666574 45067 666576
rect 42057 666571 42123 666574
rect 45001 666571 45067 666574
rect 40350 666300 40356 666364
rect 40420 666362 40426 666364
rect 42333 666362 42399 666365
rect 40420 666360 42399 666362
rect 40420 666304 42338 666360
rect 42394 666304 42399 666360
rect 40420 666302 42399 666304
rect 40420 666300 40426 666302
rect 42333 666299 42399 666302
rect 673545 666362 673611 666365
rect 676262 666362 676322 666468
rect 673545 666360 676322 666362
rect 673545 666304 673550 666360
rect 673606 666304 676322 666360
rect 673545 666302 676322 666304
rect 673545 666299 673611 666302
rect 673913 666090 673979 666093
rect 673913 666088 676292 666090
rect 673913 666032 673918 666088
rect 673974 666032 676292 666088
rect 673913 666030 676292 666032
rect 673913 666027 673979 666030
rect 680997 665818 681063 665821
rect 680997 665816 681106 665818
rect 680997 665760 681002 665816
rect 681058 665760 681106 665816
rect 680997 665755 681106 665760
rect 681046 665652 681106 665755
rect 40902 665212 40908 665276
rect 40972 665274 40978 665276
rect 41781 665274 41847 665277
rect 40972 665272 41847 665274
rect 40972 665216 41786 665272
rect 41842 665216 41847 665272
rect 40972 665214 41847 665216
rect 40972 665212 40978 665214
rect 41781 665211 41847 665214
rect 673913 665274 673979 665277
rect 673913 665272 676292 665274
rect 673913 665216 673918 665272
rect 673974 665216 676292 665272
rect 673913 665214 676292 665216
rect 673913 665211 673979 665214
rect 673913 664866 673979 664869
rect 673913 664864 676292 664866
rect 673913 664808 673918 664864
rect 673974 664808 676292 664864
rect 673913 664806 676292 664808
rect 673913 664803 673979 664806
rect 674414 664396 674420 664460
rect 674484 664458 674490 664460
rect 674484 664398 676292 664458
rect 674484 664396 674490 664398
rect 40718 664124 40724 664188
rect 40788 664186 40794 664188
rect 41781 664186 41847 664189
rect 40788 664184 41847 664186
rect 40788 664128 41786 664184
rect 41842 664128 41847 664184
rect 40788 664126 41847 664128
rect 40788 664124 40794 664126
rect 41781 664123 41847 664126
rect 673913 664050 673979 664053
rect 674925 664050 674991 664053
rect 673913 664048 674991 664050
rect 673913 663992 673918 664048
rect 673974 663992 674930 664048
rect 674986 663992 674991 664048
rect 673913 663990 674991 663992
rect 673913 663987 673979 663990
rect 674925 663987 674991 663990
rect 676262 663781 676322 664020
rect 676213 663776 676322 663781
rect 676213 663720 676218 663776
rect 676274 663720 676322 663776
rect 676213 663718 676322 663720
rect 676213 663715 676279 663718
rect 674741 663506 674807 663509
rect 676262 663506 676322 663612
rect 674741 663504 676322 663506
rect 674741 663448 674746 663504
rect 674802 663448 676322 663504
rect 674741 663446 676322 663448
rect 674741 663443 674807 663446
rect 676806 663308 676812 663372
rect 676876 663308 676882 663372
rect 676814 663204 676874 663308
rect 683205 662962 683271 662965
rect 683205 662960 683314 662962
rect 683205 662904 683210 662960
rect 683266 662904 683314 662960
rect 683205 662899 683314 662904
rect 40534 662764 40540 662828
rect 40604 662826 40610 662828
rect 42149 662826 42215 662829
rect 40604 662824 42215 662826
rect 40604 662768 42154 662824
rect 42210 662768 42215 662824
rect 683254 662796 683314 662899
rect 40604 662766 42215 662768
rect 40604 662764 40610 662766
rect 42149 662763 42215 662766
rect 674598 662356 674604 662420
rect 674668 662418 674674 662420
rect 674668 662358 676292 662418
rect 674668 662356 674674 662358
rect 673913 662010 673979 662013
rect 673913 662008 676292 662010
rect 673913 661952 673918 662008
rect 673974 661952 676292 662008
rect 673913 661950 676292 661952
rect 673913 661947 673979 661950
rect 673913 661602 673979 661605
rect 673913 661600 676292 661602
rect 673913 661544 673918 661600
rect 673974 661544 676292 661600
rect 673913 661542 676292 661544
rect 673913 661539 673979 661542
rect 673913 661194 673979 661197
rect 673913 661192 676292 661194
rect 673913 661136 673918 661192
rect 673974 661136 676292 661192
rect 673913 661134 676292 661136
rect 673913 661131 673979 661134
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 673913 660242 673979 660245
rect 674557 660242 674623 660245
rect 673913 660240 674623 660242
rect 673913 660184 673918 660240
rect 673974 660184 674562 660240
rect 674618 660184 674623 660240
rect 673913 660182 674623 660184
rect 673913 660179 673979 660182
rect 674557 660179 674623 660182
rect 683070 660109 683130 660756
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 683113 660043 683179 660046
rect 673913 659970 673979 659973
rect 673913 659968 676292 659970
rect 673913 659912 673918 659968
rect 673974 659912 676292 659968
rect 673913 659910 676292 659912
rect 673913 659907 673979 659910
rect 62113 659562 62179 659565
rect 62113 659560 64706 659562
rect 62113 659504 62118 659560
rect 62174 659504 64706 659560
rect 62113 659502 64706 659504
rect 62113 659499 62179 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 62757 657658 62823 657661
rect 62757 657656 64706 657658
rect 62757 657600 62762 657656
rect 62818 657600 64706 657656
rect 62757 657598 64706 657600
rect 62757 657595 62823 657598
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 64646 657092 64706 657598
rect 61377 656570 61443 656573
rect 61377 656568 64706 656570
rect 61377 656512 61382 656568
rect 61438 656512 64706 656568
rect 61377 656510 64706 656512
rect 61377 656507 61443 656510
rect 64646 655910 64706 656510
rect 673913 655618 673979 655621
rect 675109 655618 675175 655621
rect 673913 655616 675175 655618
rect 673913 655560 673918 655616
rect 673974 655560 675114 655616
rect 675170 655560 675175 655616
rect 673913 655558 675175 655560
rect 673913 655555 673979 655558
rect 675109 655555 675175 655558
rect 62113 655346 62179 655349
rect 62113 655344 64706 655346
rect 62113 655288 62118 655344
rect 62174 655288 64706 655344
rect 62113 655286 64706 655288
rect 62113 655283 62179 655286
rect 64646 654728 64706 655286
rect 671981 652218 672047 652221
rect 675109 652218 675175 652221
rect 671981 652216 675175 652218
rect 671981 652160 671986 652216
rect 672042 652160 675114 652216
rect 675170 652160 675175 652216
rect 671981 652158 675175 652160
rect 671981 652155 672047 652158
rect 675109 652155 675175 652158
rect 672717 651402 672783 651405
rect 675109 651402 675175 651405
rect 672717 651400 675175 651402
rect 672717 651344 672722 651400
rect 672778 651344 675114 651400
rect 675170 651344 675175 651400
rect 672717 651342 675175 651344
rect 672717 651339 672783 651342
rect 675109 651339 675175 651342
rect 667749 649226 667815 649229
rect 675385 649226 675451 649229
rect 667749 649224 675451 649226
rect 667749 649168 667754 649224
rect 667810 649168 675390 649224
rect 675446 649168 675451 649224
rect 667749 649166 675451 649168
rect 667749 649163 667815 649166
rect 675385 649163 675451 649166
rect 674005 648410 674071 648413
rect 675385 648410 675451 648413
rect 674005 648408 675451 648410
rect 674005 648352 674010 648408
rect 674066 648352 675390 648408
rect 675446 648352 675451 648408
rect 674005 648350 675451 648352
rect 674005 648347 674071 648350
rect 675385 648347 675451 648350
rect 670509 647866 670575 647869
rect 675385 647866 675451 647869
rect 670509 647864 675451 647866
rect 670509 647808 670514 647864
rect 670570 647808 675390 647864
rect 675446 647808 675451 647864
rect 670509 647806 675451 647808
rect 670509 647803 670575 647806
rect 675385 647803 675451 647806
rect 674005 647322 674071 647325
rect 675109 647322 675175 647325
rect 674005 647320 675175 647322
rect 674005 647264 674010 647320
rect 674066 647264 675114 647320
rect 675170 647264 675175 647320
rect 674005 647262 675175 647264
rect 674005 647259 674071 647262
rect 675109 647259 675175 647262
rect 35758 644741 35818 644912
rect 674741 644874 674807 644877
rect 675334 644874 675340 644876
rect 674741 644872 675340 644874
rect 674741 644816 674746 644872
rect 674802 644816 675340 644872
rect 674741 644814 675340 644816
rect 674741 644811 674807 644814
rect 675334 644812 675340 644814
rect 675404 644812 675410 644876
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 39573 644738 39639 644741
rect 44449 644738 44515 644741
rect 39573 644736 44515 644738
rect 39573 644680 39578 644736
rect 39634 644680 44454 644736
rect 44510 644680 44515 644736
rect 39573 644678 44515 644680
rect 39573 644675 39639 644678
rect 44449 644675 44515 644678
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 674097 644330 674163 644333
rect 675293 644330 675359 644333
rect 674097 644328 675359 644330
rect 674097 644272 674102 644328
rect 674158 644272 675298 644328
rect 675354 644272 675359 644328
rect 674097 644270 675359 644272
rect 674097 644267 674163 644270
rect 675293 644267 675359 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 35341 643859 35407 643862
rect 35574 643517 35634 643688
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 40493 643514 40559 643517
rect 45001 643514 45067 643517
rect 40493 643512 45067 643514
rect 40493 643456 40498 643512
rect 40554 643456 45006 643512
rect 45062 643456 45067 643512
rect 40493 643454 45067 643456
rect 40493 643451 40559 643454
rect 45001 643451 45067 643454
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 670969 643514 671035 643517
rect 675477 643514 675543 643517
rect 670969 643512 675543 643514
rect 670969 643456 670974 643512
rect 671030 643456 675482 643512
rect 675538 643456 675543 643512
rect 670969 643454 675543 643456
rect 670969 643451 671035 643454
rect 675477 643451 675543 643454
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 674005 643106 674071 643109
rect 675109 643106 675175 643109
rect 674005 643104 675175 643106
rect 674005 643048 674010 643104
rect 674066 643048 675114 643104
rect 675170 643048 675175 643104
rect 674005 643046 675175 643048
rect 674005 643043 674071 643046
rect 675109 643043 675175 643046
rect 35574 642701 35634 642872
rect 35574 642696 35683 642701
rect 35574 642640 35622 642696
rect 35678 642640 35683 642696
rect 35574 642638 35683 642640
rect 35617 642635 35683 642638
rect 35801 642290 35867 642293
rect 35758 642288 35867 642290
rect 35758 642232 35806 642288
rect 35862 642232 35867 642288
rect 35758 642227 35867 642232
rect 41462 642290 41522 642464
rect 44214 642290 44220 642292
rect 41462 642230 44220 642290
rect 44214 642228 44220 642230
rect 44284 642228 44290 642292
rect 35758 642056 35818 642227
rect 649950 641882 650010 642376
rect 652017 641882 652083 641885
rect 649950 641880 652083 641882
rect 649950 641824 652022 641880
rect 652078 641824 652083 641880
rect 649950 641822 652083 641824
rect 652017 641819 652083 641822
rect 669865 641746 669931 641749
rect 675293 641746 675359 641749
rect 669865 641744 675359 641746
rect 669865 641688 669870 641744
rect 669926 641688 675298 641744
rect 675354 641688 675359 641744
rect 669865 641686 675359 641688
rect 669865 641683 669931 641686
rect 675293 641683 675359 641686
rect 35390 641477 35450 641648
rect 35341 641472 35450 641477
rect 35341 641416 35346 641472
rect 35402 641416 35450 641472
rect 35341 641414 35450 641416
rect 35341 641411 35407 641414
rect 35574 641069 35634 641240
rect 35525 641064 35634 641069
rect 35801 641066 35867 641069
rect 35525 641008 35530 641064
rect 35586 641008 35634 641064
rect 35525 641006 35634 641008
rect 35758 641064 35867 641066
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35525 641003 35591 641006
rect 35758 641003 35867 641008
rect 35758 640832 35818 641003
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 668393 640658 668459 640661
rect 675385 640658 675451 640661
rect 668393 640656 675451 640658
rect 668393 640600 668398 640656
rect 668454 640600 675390 640656
rect 675446 640600 675451 640656
rect 668393 640598 675451 640600
rect 41462 640424 41522 640596
rect 668393 640595 668459 640598
rect 675385 640595 675451 640598
rect 675293 640388 675359 640389
rect 675293 640384 675340 640388
rect 675404 640386 675410 640388
rect 675293 640328 675298 640384
rect 675293 640324 675340 640328
rect 675404 640326 675450 640386
rect 675404 640324 675410 640326
rect 675293 640323 675359 640324
rect 39941 640250 40007 640253
rect 45277 640250 45343 640253
rect 39941 640248 45343 640250
rect 39941 640192 39946 640248
rect 40002 640192 45282 640248
rect 45338 640192 45343 640248
rect 39941 640190 45343 640192
rect 39941 640187 40007 640190
rect 45277 640187 45343 640190
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 35758 639845 35818 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 35758 639840 35867 639845
rect 35758 639784 35806 639840
rect 35862 639784 35867 639840
rect 35758 639782 35867 639784
rect 35801 639779 35867 639782
rect 41462 639434 41522 639608
rect 41638 639434 41644 639436
rect 41462 639374 41644 639434
rect 41638 639372 41644 639374
rect 41708 639372 41714 639436
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 670969 638754 671035 638757
rect 675477 638754 675543 638757
rect 670969 638752 675543 638754
rect 670969 638696 670974 638752
rect 671030 638696 675482 638752
rect 675538 638696 675543 638752
rect 670969 638694 675543 638696
rect 670969 638691 671035 638694
rect 675477 638691 675543 638694
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 35206 637805 35266 637976
rect 35157 637800 35266 637805
rect 35157 637744 35162 637800
rect 35218 637744 35266 637800
rect 35157 637742 35266 637744
rect 35157 637739 35223 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 40542 637396 40602 637568
rect 40534 637332 40540 637396
rect 40604 637332 40610 637396
rect 32078 636989 32138 637160
rect 32029 636984 32138 636989
rect 32029 636928 32034 636984
rect 32090 636928 32138 636984
rect 32029 636926 32138 636928
rect 32029 636923 32095 636926
rect 674230 636788 674236 636852
rect 674300 636850 674306 636852
rect 683941 636850 684007 636853
rect 674300 636848 684007 636850
rect 674300 636792 683946 636848
rect 684002 636792 684007 636848
rect 674300 636790 684007 636792
rect 674300 636788 674306 636790
rect 683941 636787 684007 636790
rect 35574 636581 35634 636752
rect 35525 636576 35634 636581
rect 35801 636578 35867 636581
rect 35525 636520 35530 636576
rect 35586 636520 35634 636576
rect 35525 636518 35634 636520
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35525 636515 35591 636518
rect 35758 636515 35867 636520
rect 39113 636578 39179 636581
rect 42517 636578 42583 636581
rect 39113 636576 42583 636578
rect 39113 636520 39118 636576
rect 39174 636520 42522 636576
rect 42578 636520 42583 636576
rect 39113 636518 42583 636520
rect 39113 636515 39179 636518
rect 42517 636515 42583 636518
rect 35758 636344 35818 636515
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 40726 635356 40786 635528
rect 40718 635292 40724 635356
rect 40788 635292 40794 635356
rect 40910 634948 40970 635120
rect 40902 634884 40908 634948
rect 40972 634884 40978 634948
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 41462 633926 41522 634304
rect 41873 633926 41939 633929
rect 41462 633924 41939 633926
rect 41462 633896 41878 633924
rect 41492 633868 41878 633896
rect 41934 633868 41939 633924
rect 41492 633866 41939 633868
rect 41873 633863 41939 633866
rect 39941 633722 40007 633725
rect 44357 633722 44423 633725
rect 39941 633720 44423 633722
rect 39941 633664 39946 633720
rect 40002 633664 44362 633720
rect 44418 633664 44423 633720
rect 39941 633662 44423 633664
rect 39941 633659 40007 633662
rect 44357 633659 44423 633662
rect 35758 633317 35818 633488
rect 35758 633312 35867 633317
rect 35758 633256 35806 633312
rect 35862 633256 35867 633312
rect 35758 633254 35867 633256
rect 35801 633251 35867 633254
rect 39757 632226 39823 632229
rect 43989 632226 44055 632229
rect 39757 632224 44055 632226
rect 39757 632168 39762 632224
rect 39818 632168 43994 632224
rect 44050 632168 44055 632224
rect 39757 632166 44055 632168
rect 39757 632163 39823 632166
rect 43989 632163 44055 632166
rect 41413 631410 41479 631413
rect 44173 631410 44239 631413
rect 41413 631408 44239 631410
rect 41413 631352 41418 631408
rect 41474 631352 44178 631408
rect 44234 631352 44239 631408
rect 41413 631350 44239 631352
rect 41413 631347 41479 631350
rect 44173 631347 44239 631350
rect 674925 631410 674991 631413
rect 675150 631410 675156 631412
rect 674925 631408 675156 631410
rect 674925 631352 674930 631408
rect 674986 631352 675156 631408
rect 674925 631350 675156 631352
rect 674925 631347 674991 631350
rect 675150 631348 675156 631350
rect 675220 631348 675226 631412
rect 40401 630730 40467 630733
rect 44817 630730 44883 630733
rect 40401 630728 44883 630730
rect 40401 630672 40406 630728
rect 40462 630672 44822 630728
rect 44878 630672 44883 630728
rect 40401 630670 44883 630672
rect 40401 630667 40467 630670
rect 44817 630667 44883 630670
rect 39113 630458 39179 630461
rect 43713 630458 43779 630461
rect 39113 630456 43779 630458
rect 39113 630400 39118 630456
rect 39174 630400 43718 630456
rect 43774 630400 43779 630456
rect 39113 630398 43779 630400
rect 39113 630395 39179 630398
rect 43713 630395 43779 630398
rect 35157 629914 35223 629917
rect 41822 629914 41828 629916
rect 35157 629912 41828 629914
rect 35157 629856 35162 629912
rect 35218 629856 41828 629912
rect 35157 629854 41828 629856
rect 35157 629851 35223 629854
rect 41822 629852 41828 629854
rect 41892 629852 41898 629916
rect 675017 629778 675083 629781
rect 676070 629778 676076 629780
rect 675017 629776 676076 629778
rect 675017 629720 675022 629776
rect 675078 629720 676076 629776
rect 675017 629718 676076 629720
rect 675017 629715 675083 629718
rect 676070 629716 676076 629718
rect 676140 629716 676146 629780
rect 37733 629642 37799 629645
rect 42333 629642 42399 629645
rect 37733 629640 42399 629642
rect 37733 629584 37738 629640
rect 37794 629584 42338 629640
rect 42394 629584 42399 629640
rect 37733 629582 42399 629584
rect 37733 629579 37799 629582
rect 42333 629579 42399 629582
rect 37917 627738 37983 627741
rect 42057 627738 42123 627741
rect 37917 627736 42123 627738
rect 37917 627680 37922 627736
rect 37978 627680 42062 627736
rect 42118 627680 42123 627736
rect 37917 627678 42123 627680
rect 37917 627675 37983 627678
rect 42057 627675 42123 627678
rect 41781 627464 41847 627469
rect 41781 627408 41786 627464
rect 41842 627408 41847 627464
rect 41781 627403 41847 627408
rect 41784 627197 41844 627403
rect 41781 627192 41847 627197
rect 41781 627136 41786 627192
rect 41842 627136 41847 627192
rect 41781 627131 41847 627136
rect 674005 626378 674071 626381
rect 674005 626376 676292 626378
rect 674005 626320 674010 626376
rect 674066 626320 676292 626376
rect 674005 626318 676292 626320
rect 674005 626315 674071 626318
rect 673545 625970 673611 625973
rect 674925 625970 674991 625973
rect 673545 625968 674991 625970
rect 673545 625912 673550 625968
rect 673606 625912 674930 625968
rect 674986 625912 674991 625968
rect 673545 625910 674991 625912
rect 673545 625907 673611 625910
rect 674925 625907 674991 625910
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 674054 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 674054 625565 674114 625638
rect 674005 625560 674114 625565
rect 674005 625504 674010 625560
rect 674066 625504 674114 625560
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 674005 625502 674114 625504
rect 674005 625499 674071 625502
rect 670233 625154 670299 625157
rect 670233 625152 676292 625154
rect 670233 625096 670238 625152
rect 670294 625096 676292 625152
rect 670233 625094 676292 625096
rect 670233 625091 670299 625094
rect 42425 624748 42491 624749
rect 42374 624684 42380 624748
rect 42444 624746 42491 624748
rect 674005 624746 674071 624749
rect 42444 624744 42536 624746
rect 42486 624688 42536 624744
rect 42444 624686 42536 624688
rect 674005 624744 676292 624746
rect 674005 624688 674010 624744
rect 674066 624688 676292 624744
rect 674005 624686 676292 624688
rect 42444 624684 42491 624686
rect 42425 624683 42491 624684
rect 674005 624683 674071 624686
rect 42057 624474 42123 624477
rect 45737 624474 45803 624477
rect 42057 624472 45803 624474
rect 42057 624416 42062 624472
rect 42118 624416 45742 624472
rect 45798 624416 45803 624472
rect 42057 624414 45803 624416
rect 42057 624411 42123 624414
rect 45737 624411 45803 624414
rect 674005 624338 674071 624341
rect 674005 624336 676292 624338
rect 674005 624280 674010 624336
rect 674066 624280 676292 624336
rect 674005 624278 676292 624280
rect 674005 624275 674071 624278
rect 674005 623930 674071 623933
rect 674005 623928 676292 623930
rect 674005 623872 674010 623928
rect 674066 623872 676292 623928
rect 674005 623870 676292 623872
rect 674005 623867 674071 623870
rect 40902 623732 40908 623796
rect 40972 623794 40978 623796
rect 42057 623794 42123 623797
rect 40972 623792 42123 623794
rect 40972 623736 42062 623792
rect 42118 623736 42123 623792
rect 40972 623734 42123 623736
rect 40972 623732 40978 623734
rect 42057 623731 42123 623734
rect 674005 623522 674071 623525
rect 674005 623520 676292 623522
rect 674005 623464 674010 623520
rect 674066 623464 676292 623520
rect 674005 623462 676292 623464
rect 674005 623459 674071 623462
rect 42057 623386 42123 623389
rect 44081 623386 44147 623389
rect 42057 623384 44147 623386
rect 42057 623328 42062 623384
rect 42118 623328 44086 623384
rect 44142 623328 44147 623384
rect 42057 623326 44147 623328
rect 42057 623323 42123 623326
rect 44081 623323 44147 623326
rect 674005 623114 674071 623117
rect 674005 623112 676292 623114
rect 674005 623056 674010 623112
rect 674066 623056 676292 623112
rect 674005 623054 676292 623056
rect 674005 623051 674071 623054
rect 671153 622706 671219 622709
rect 671153 622704 676292 622706
rect 671153 622648 671158 622704
rect 671214 622648 676292 622704
rect 671153 622646 676292 622648
rect 671153 622643 671219 622646
rect 674005 622298 674071 622301
rect 674005 622296 676292 622298
rect 674005 622240 674010 622296
rect 674066 622240 676292 622296
rect 674005 622238 676292 622240
rect 674005 622235 674071 622238
rect 42057 622162 42123 622165
rect 44357 622162 44423 622165
rect 42057 622160 44423 622162
rect 42057 622104 42062 622160
rect 42118 622104 44362 622160
rect 44418 622104 44423 622160
rect 42057 622102 44423 622104
rect 42057 622099 42123 622102
rect 44357 622099 44423 622102
rect 683941 622026 684007 622029
rect 683941 622024 684050 622026
rect 683941 621968 683946 622024
rect 684002 621968 684050 622024
rect 683941 621963 684050 621968
rect 683990 621860 684050 621963
rect 674005 621482 674071 621485
rect 674005 621480 676292 621482
rect 674005 621424 674010 621480
rect 674066 621424 676292 621480
rect 674005 621422 676292 621424
rect 674005 621419 674071 621422
rect 674005 621074 674071 621077
rect 674005 621072 676292 621074
rect 674005 621016 674010 621072
rect 674066 621016 676292 621072
rect 674005 621014 676292 621016
rect 674005 621011 674071 621014
rect 40718 620740 40724 620804
rect 40788 620802 40794 620804
rect 41781 620802 41847 620805
rect 40788 620800 41847 620802
rect 40788 620744 41786 620800
rect 41842 620744 41847 620800
rect 40788 620742 41847 620744
rect 40788 620740 40794 620742
rect 41781 620739 41847 620742
rect 42374 620740 42380 620804
rect 42444 620802 42450 620804
rect 42701 620802 42767 620805
rect 42444 620800 42767 620802
rect 42444 620744 42706 620800
rect 42762 620744 42767 620800
rect 42444 620742 42767 620744
rect 42444 620740 42450 620742
rect 42701 620739 42767 620742
rect 673637 620666 673703 620669
rect 673637 620664 676292 620666
rect 673637 620608 673642 620664
rect 673698 620608 676292 620664
rect 673637 620606 676292 620608
rect 673637 620603 673703 620606
rect 671797 620258 671863 620261
rect 671797 620256 676292 620258
rect 671797 620200 671802 620256
rect 671858 620200 676292 620256
rect 671797 620198 676292 620200
rect 671797 620195 671863 620198
rect 40534 619788 40540 619852
rect 40604 619850 40610 619852
rect 42241 619850 42307 619853
rect 40604 619848 42307 619850
rect 40604 619792 42246 619848
rect 42302 619792 42307 619848
rect 40604 619790 42307 619792
rect 40604 619788 40610 619790
rect 42241 619787 42307 619790
rect 674005 619850 674071 619853
rect 674005 619848 676292 619850
rect 674005 619792 674010 619848
rect 674066 619792 676292 619848
rect 674005 619790 676292 619792
rect 674005 619787 674071 619790
rect 673177 619442 673243 619445
rect 673177 619440 676292 619442
rect 673177 619384 673182 619440
rect 673238 619384 676292 619440
rect 673177 619382 676292 619384
rect 673177 619379 673243 619382
rect 674005 619034 674071 619037
rect 674005 619032 676292 619034
rect 674005 618976 674010 619032
rect 674066 618976 676292 619032
rect 674005 618974 676292 618976
rect 674005 618971 674071 618974
rect 674189 618626 674255 618629
rect 674189 618624 676292 618626
rect 674189 618568 674194 618624
rect 674250 618568 676292 618624
rect 674189 618566 676292 618568
rect 674189 618563 674255 618566
rect 672901 618218 672967 618221
rect 672901 618216 676292 618218
rect 672901 618160 672906 618216
rect 672962 618160 676292 618216
rect 672901 618158 676292 618160
rect 672901 618155 672967 618158
rect 62941 618082 63007 618085
rect 62941 618080 64706 618082
rect 62941 618024 62946 618080
rect 63002 618024 64706 618080
rect 62941 618022 64706 618024
rect 62941 618019 63007 618022
rect 64646 617416 64706 618022
rect 683297 617946 683363 617949
rect 683254 617944 683363 617946
rect 683254 617888 683302 617944
rect 683358 617888 683363 617944
rect 683254 617883 683363 617888
rect 683254 617780 683314 617883
rect 673545 617402 673611 617405
rect 673545 617400 676292 617402
rect 673545 617344 673550 617400
rect 673606 617344 676292 617400
rect 673545 617342 676292 617344
rect 673545 617339 673611 617342
rect 674005 616994 674071 616997
rect 674005 616992 676292 616994
rect 674005 616936 674010 616992
rect 674066 616936 676292 616992
rect 674005 616934 676292 616936
rect 674005 616931 674071 616934
rect 62113 616586 62179 616589
rect 674005 616586 674071 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 41454 616252 41460 616316
rect 41524 616314 41530 616316
rect 42333 616314 42399 616317
rect 41524 616312 42399 616314
rect 41524 616256 42338 616312
rect 42394 616256 42399 616312
rect 41524 616254 42399 616256
rect 41524 616252 41530 616254
rect 42333 616251 42399 616254
rect 64646 616234 64706 616526
rect 674005 616584 676292 616586
rect 674005 616528 674010 616584
rect 674066 616528 676292 616584
rect 674005 616526 676292 616528
rect 674005 616523 674071 616526
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 41822 615980 41828 616044
rect 41892 616042 41898 616044
rect 42517 616042 42583 616045
rect 41892 616040 42583 616042
rect 41892 615984 42522 616040
rect 42578 615984 42583 616040
rect 41892 615982 42583 615984
rect 41892 615980 41898 615982
rect 42517 615979 42583 615982
rect 42057 615770 42123 615773
rect 42701 615770 42767 615773
rect 42057 615768 42767 615770
rect 42057 615712 42062 615768
rect 42118 615712 42706 615768
rect 42762 615712 42767 615768
rect 42057 615710 42767 615712
rect 42057 615707 42123 615710
rect 42701 615707 42767 615710
rect 683070 615501 683130 615740
rect 41638 615436 41644 615500
rect 41708 615498 41714 615500
rect 42517 615498 42583 615501
rect 41708 615496 42583 615498
rect 41708 615440 42522 615496
rect 42578 615440 42583 615496
rect 41708 615438 42583 615440
rect 41708 615436 41714 615438
rect 42517 615435 42583 615438
rect 674005 615498 674071 615501
rect 675109 615498 675175 615501
rect 674005 615496 675175 615498
rect 674005 615440 674010 615496
rect 674066 615440 675114 615496
rect 675170 615440 675175 615496
rect 674005 615438 675175 615440
rect 674005 615435 674071 615438
rect 675109 615435 675175 615438
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 674005 614954 674071 614957
rect 674005 614952 676292 614954
rect 674005 614896 674010 614952
rect 674066 614896 676292 614952
rect 674005 614894 676292 614896
rect 674005 614891 674071 614894
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 62113 614619 62179 614622
rect 42885 614002 42951 614005
rect 44081 614002 44147 614005
rect 42885 614000 44147 614002
rect 42885 613944 42890 614000
rect 42946 613944 44086 614000
rect 44142 613944 44147 614000
rect 42885 613942 44147 613944
rect 42885 613939 42951 613942
rect 44081 613939 44147 613942
rect 61377 613866 61443 613869
rect 64646 613866 64706 613870
rect 61377 613864 64706 613866
rect 61377 613808 61382 613864
rect 61438 613808 64706 613864
rect 61377 613806 64706 613808
rect 61377 613803 61443 613806
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 43253 612234 43319 612237
rect 43759 612234 43825 612237
rect 43253 612232 43825 612234
rect 43253 612176 43258 612232
rect 43314 612176 43764 612232
rect 43820 612176 43825 612232
rect 43253 612174 43825 612176
rect 43253 612171 43319 612174
rect 43759 612171 43825 612174
rect 44081 612098 44147 612101
rect 45553 612098 45619 612101
rect 44081 612096 45619 612098
rect 44081 612040 44086 612096
rect 44142 612040 45558 612096
rect 45614 612040 45619 612096
rect 44081 612038 45619 612040
rect 44081 612035 44147 612038
rect 45553 612035 45619 612038
rect 62757 612098 62823 612101
rect 62757 612096 64706 612098
rect 62757 612040 62762 612096
rect 62818 612040 64706 612096
rect 62757 612038 64706 612040
rect 62757 612035 62823 612038
rect 43989 611826 44055 611829
rect 47025 611826 47091 611829
rect 43989 611824 47091 611826
rect 43989 611768 43994 611824
rect 44050 611768 47030 611824
rect 47086 611768 47091 611824
rect 43989 611766 47091 611768
rect 43989 611763 44055 611766
rect 47025 611763 47091 611766
rect 44081 611554 44147 611557
rect 47209 611554 47275 611557
rect 44081 611552 47275 611554
rect 44081 611496 44086 611552
rect 44142 611496 47214 611552
rect 47270 611496 47275 611552
rect 64646 611506 64706 612038
rect 44081 611494 47275 611496
rect 44081 611491 44147 611494
rect 47209 611491 47275 611494
rect 674005 611418 674071 611421
rect 675109 611418 675175 611421
rect 674005 611416 675175 611418
rect 674005 611360 674010 611416
rect 674066 611360 675114 611416
rect 675170 611360 675175 611416
rect 674005 611358 675175 611360
rect 674005 611355 674071 611358
rect 675109 611355 675175 611358
rect 669037 608290 669103 608293
rect 675109 608290 675175 608293
rect 669037 608288 675175 608290
rect 669037 608232 669042 608288
rect 669098 608232 675114 608288
rect 675170 608232 675175 608288
rect 669037 608230 675175 608232
rect 669037 608227 669103 608230
rect 675109 608227 675175 608230
rect 671337 607338 671403 607341
rect 675109 607338 675175 607341
rect 671337 607336 675175 607338
rect 671337 607280 671342 607336
rect 671398 607280 675114 607336
rect 675170 607280 675175 607336
rect 671337 607278 675175 607280
rect 671337 607275 671403 607278
rect 675109 607275 675175 607278
rect 674833 604754 674899 604757
rect 676806 604754 676812 604756
rect 674833 604752 676812 604754
rect 674833 604696 674838 604752
rect 674894 604696 676812 604752
rect 674833 604694 676812 604696
rect 674833 604691 674899 604694
rect 676806 604692 676812 604694
rect 676876 604692 676882 604756
rect 673085 604210 673151 604213
rect 675385 604210 675451 604213
rect 673085 604208 675451 604210
rect 673085 604152 673090 604208
rect 673146 604152 675390 604208
rect 675446 604152 675451 604208
rect 673085 604150 675451 604152
rect 673085 604147 673151 604150
rect 675385 604147 675451 604150
rect 672349 603802 672415 603805
rect 675109 603802 675175 603805
rect 672349 603800 675175 603802
rect 672349 603744 672354 603800
rect 672410 603744 675114 603800
rect 675170 603744 675175 603800
rect 672349 603742 675175 603744
rect 672349 603739 672415 603742
rect 675109 603739 675175 603742
rect 674230 602924 674236 602988
rect 674300 602986 674306 602988
rect 675109 602986 675175 602989
rect 674300 602984 675175 602986
rect 674300 602928 675114 602984
rect 675170 602928 675175 602984
rect 674300 602926 675175 602928
rect 674300 602924 674306 602926
rect 675109 602923 675175 602926
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 38561 601354 38627 601357
rect 38548 601352 38627 601354
rect 38548 601296 38566 601352
rect 38622 601296 38627 601352
rect 38548 601294 38627 601296
rect 38561 601291 38627 601294
rect 39941 600946 40007 600949
rect 39941 600944 40020 600946
rect 39941 600888 39946 600944
rect 40002 600888 40020 600944
rect 39941 600886 40020 600888
rect 39941 600883 40007 600886
rect 671797 600674 671863 600677
rect 675109 600674 675175 600677
rect 671797 600672 675175 600674
rect 671797 600616 671802 600672
rect 671858 600616 675114 600672
rect 675170 600616 675175 600672
rect 671797 600614 675175 600616
rect 671797 600611 671863 600614
rect 675109 600611 675175 600614
rect 45001 600538 45067 600541
rect 41492 600536 45067 600538
rect 41492 600480 45006 600536
rect 45062 600480 45067 600536
rect 41492 600478 45067 600480
rect 45001 600475 45067 600478
rect 673821 600402 673887 600405
rect 675293 600402 675359 600405
rect 673821 600400 675359 600402
rect 673821 600344 673826 600400
rect 673882 600344 675298 600400
rect 675354 600344 675359 600400
rect 673821 600342 675359 600344
rect 673821 600339 673887 600342
rect 675293 600339 675359 600342
rect 45093 600130 45159 600133
rect 41492 600128 45159 600130
rect 41492 600072 45098 600128
rect 45154 600072 45159 600128
rect 41492 600070 45159 600072
rect 45093 600067 45159 600070
rect 673637 599858 673703 599861
rect 675477 599858 675543 599861
rect 673637 599856 675543 599858
rect 673637 599800 673642 599856
rect 673698 599800 675482 599856
rect 675538 599800 675543 599856
rect 673637 599798 675543 599800
rect 673637 599795 673703 599798
rect 675477 599795 675543 599798
rect 44214 599722 44220 599724
rect 41492 599662 44220 599722
rect 44214 599660 44220 599662
rect 44284 599660 44290 599724
rect 673821 599450 673887 599453
rect 675109 599450 675175 599453
rect 673821 599448 675175 599450
rect 673821 599392 673826 599448
rect 673882 599392 675114 599448
rect 675170 599392 675175 599448
rect 673821 599390 675175 599392
rect 673821 599387 673887 599390
rect 675109 599387 675175 599390
rect 43110 599314 43116 599316
rect 41492 599254 43116 599314
rect 43110 599252 43116 599254
rect 43180 599252 43186 599316
rect 673821 599178 673887 599181
rect 675477 599178 675543 599181
rect 673821 599176 675543 599178
rect 673821 599120 673826 599176
rect 673882 599120 675482 599176
rect 675538 599120 675543 599176
rect 673821 599118 675543 599120
rect 673821 599115 673887 599118
rect 675477 599115 675543 599118
rect 44633 598906 44699 598909
rect 41492 598904 44699 598906
rect 41492 598848 44638 598904
rect 44694 598848 44699 598904
rect 41492 598846 44699 598848
rect 44633 598843 44699 598846
rect 674189 598634 674255 598637
rect 675477 598634 675543 598637
rect 674189 598632 675543 598634
rect 674189 598576 674194 598632
rect 674250 598576 675482 598632
rect 675538 598576 675543 598632
rect 674189 598574 675543 598576
rect 674189 598571 674255 598574
rect 675477 598571 675543 598574
rect 44909 598498 44975 598501
rect 41492 598496 44975 598498
rect 41492 598440 44914 598496
rect 44970 598440 44975 598496
rect 41492 598438 44975 598440
rect 44909 598435 44975 598438
rect 45277 598090 45343 598093
rect 41492 598088 45343 598090
rect 41492 598032 45282 598088
rect 45338 598032 45343 598088
rect 41492 598030 45343 598032
rect 45277 598027 45343 598030
rect 649950 597954 650010 598336
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 42885 597682 42951 597685
rect 41492 597680 42951 597682
rect 41492 597624 42890 597680
rect 42946 597624 42951 597680
rect 41492 597622 42951 597624
rect 42885 597619 42951 597622
rect 672533 597410 672599 597413
rect 675385 597410 675451 597413
rect 672533 597408 675451 597410
rect 672533 597352 672538 597408
rect 672594 597352 675390 597408
rect 675446 597352 675451 597408
rect 672533 597350 675451 597352
rect 672533 597347 672599 597350
rect 675385 597347 675451 597350
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 43069 597004 43135 597005
rect 43069 597000 43116 597004
rect 43180 597002 43186 597004
rect 43069 596944 43074 597000
rect 43069 596940 43116 596944
rect 43180 596942 43226 597002
rect 43180 596940 43186 596942
rect 43069 596939 43135 596940
rect 42425 596866 42491 596869
rect 41492 596864 42491 596866
rect 41492 596808 42430 596864
rect 42486 596808 42491 596864
rect 41492 596806 42491 596808
rect 42425 596803 42491 596806
rect 649950 596730 650010 597154
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 41137 596458 41203 596461
rect 41124 596456 41203 596458
rect 41124 596400 41142 596456
rect 41198 596400 41203 596456
rect 41124 596398 41203 596400
rect 41137 596395 41203 596398
rect 41965 596050 42031 596053
rect 41492 596048 42031 596050
rect 41492 595992 41970 596048
rect 42026 595992 42031 596048
rect 41492 595990 42031 595992
rect 41965 595987 42031 595990
rect 35617 595812 35683 595815
rect 35574 595810 35683 595812
rect 35574 595754 35622 595810
rect 35678 595754 35683 595810
rect 35574 595749 35683 595754
rect 41689 595778 41755 595781
rect 62941 595778 63007 595781
rect 41689 595776 63007 595778
rect 35574 595612 35634 595749
rect 41689 595720 41694 595776
rect 41750 595720 62946 595776
rect 63002 595720 63007 595776
rect 41689 595718 63007 595720
rect 41689 595715 41755 595718
rect 62941 595715 63007 595718
rect 649950 595506 650010 595972
rect 651465 595506 651531 595509
rect 649950 595504 651531 595506
rect 649950 595448 651470 595504
rect 651526 595448 651531 595504
rect 649950 595446 651531 595448
rect 651465 595443 651531 595446
rect 667013 595506 667079 595509
rect 675385 595506 675451 595509
rect 667013 595504 675451 595506
rect 667013 595448 667018 595504
rect 667074 595448 675390 595504
rect 675446 595448 675451 595504
rect 667013 595446 675451 595448
rect 667013 595443 667079 595446
rect 675385 595443 675451 595446
rect 33041 595234 33107 595237
rect 651649 595234 651715 595237
rect 33028 595232 33107 595234
rect 33028 595176 33046 595232
rect 33102 595176 33107 595232
rect 33028 595174 33107 595176
rect 33041 595171 33107 595174
rect 649950 595232 651715 595234
rect 649950 595176 651654 595232
rect 651710 595176 651715 595232
rect 649950 595174 651715 595176
rect 39297 594826 39363 594829
rect 39284 594824 39363 594826
rect 39284 594768 39302 594824
rect 39358 594768 39363 594824
rect 649950 594790 650010 595174
rect 651649 595171 651715 595174
rect 39284 594766 39363 594768
rect 39297 594763 39363 594766
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 41781 594282 41847 594285
rect 41781 594280 51090 594282
rect 41781 594224 41786 594280
rect 41842 594224 51090 594280
rect 41781 594222 51090 594224
rect 41781 594219 41847 594222
rect 51030 594146 51090 594222
rect 62757 594146 62823 594149
rect 651465 594146 651531 594149
rect 51030 594144 62823 594146
rect 51030 594088 62762 594144
rect 62818 594088 62823 594144
rect 51030 594086 62823 594088
rect 62757 594083 62823 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 41822 594010 41828 594012
rect 41492 593950 41828 594010
rect 41822 593948 41828 593950
rect 41892 593948 41898 594012
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 33777 593602 33843 593605
rect 33764 593600 33843 593602
rect 33764 593544 33782 593600
rect 33838 593544 33843 593600
rect 33764 593542 33843 593544
rect 33777 593539 33843 593542
rect 668853 593602 668919 593605
rect 675385 593602 675451 593605
rect 668853 593600 675451 593602
rect 668853 593544 668858 593600
rect 668914 593544 675390 593600
rect 675446 593544 675451 593600
rect 668853 593542 675451 593544
rect 668853 593539 668919 593542
rect 675385 593539 675451 593542
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 41689 592922 41755 592925
rect 63125 592922 63191 592925
rect 41689 592920 63191 592922
rect 41689 592864 41694 592920
rect 41750 592864 63130 592920
rect 63186 592864 63191 592920
rect 41689 592862 63191 592864
rect 41689 592859 41755 592862
rect 63125 592859 63191 592862
rect 675150 592860 675156 592924
rect 675220 592922 675226 592924
rect 676029 592922 676095 592925
rect 675220 592920 676095 592922
rect 675220 592864 676034 592920
rect 676090 592864 676095 592920
rect 675220 592862 676095 592864
rect 675220 592860 675226 592862
rect 676029 592859 676095 592862
rect 651465 592786 651531 592789
rect 649950 592784 651531 592786
rect 40726 592550 40786 592756
rect 649950 592728 651470 592784
rect 651526 592728 651531 592784
rect 649950 592726 651531 592728
rect 40718 592486 40724 592550
rect 40788 592486 40794 592550
rect 649950 592426 650010 592726
rect 651465 592723 651531 592726
rect 41822 592378 41828 592380
rect 41492 592318 41828 592378
rect 41822 592316 41828 592318
rect 41892 592316 41898 592380
rect 44173 591970 44239 591973
rect 41492 591968 44239 591970
rect 41492 591912 44178 591968
rect 44234 591912 44239 591968
rect 41492 591910 44239 591912
rect 44173 591907 44239 591910
rect 43345 591562 43411 591565
rect 41492 591560 43411 591562
rect 41492 591504 43350 591560
rect 43406 591504 43411 591560
rect 41492 591502 43411 591504
rect 43345 591499 43411 591502
rect 674005 591426 674071 591429
rect 675477 591426 675543 591429
rect 674005 591424 675543 591426
rect 674005 591368 674010 591424
rect 674066 591368 675482 591424
rect 675538 591368 675543 591424
rect 674005 591366 675543 591368
rect 674005 591363 674071 591366
rect 675477 591363 675543 591366
rect 41689 591290 41755 591293
rect 42190 591290 42196 591292
rect 41689 591288 42196 591290
rect 41689 591232 41694 591288
rect 41750 591232 42196 591288
rect 41689 591230 42196 591232
rect 41689 591227 41755 591230
rect 42190 591228 42196 591230
rect 42260 591228 42266 591292
rect 41094 590749 41154 591124
rect 41045 590744 41154 590749
rect 41045 590688 41050 590744
rect 41106 590716 41154 590744
rect 41106 590688 41124 590716
rect 41045 590686 41124 590688
rect 41045 590683 41111 590686
rect 676070 590548 676076 590612
rect 676140 590610 676146 590612
rect 682377 590610 682443 590613
rect 676140 590608 682443 590610
rect 676140 590552 682382 590608
rect 682438 590552 682443 590608
rect 676140 590550 682443 590552
rect 676140 590548 676146 590550
rect 682377 590547 682443 590550
rect 43621 590338 43687 590341
rect 41492 590336 43687 590338
rect 41492 590280 43626 590336
rect 43682 590280 43687 590336
rect 41492 590278 43687 590280
rect 43621 590275 43687 590278
rect 675293 586258 675359 586261
rect 675886 586258 675892 586260
rect 675293 586256 675892 586258
rect 675293 586200 675298 586256
rect 675354 586200 675892 586256
rect 675293 586198 675892 586200
rect 675293 586195 675359 586198
rect 675886 586196 675892 586198
rect 675956 586196 675962 586260
rect 41965 586124 42031 586125
rect 41965 586122 42012 586124
rect 41920 586120 42012 586122
rect 41920 586064 41970 586120
rect 41920 586062 42012 586064
rect 41965 586060 42012 586062
rect 42076 586060 42082 586124
rect 41965 586059 42031 586060
rect 39573 585850 39639 585853
rect 42149 585850 42215 585853
rect 39573 585848 42215 585850
rect 39573 585792 39578 585848
rect 39634 585792 42154 585848
rect 42210 585792 42215 585848
rect 39573 585790 42215 585792
rect 39573 585787 39639 585790
rect 42149 585787 42215 585790
rect 41045 585442 41111 585445
rect 42241 585442 42307 585445
rect 41045 585440 42307 585442
rect 41045 585384 41050 585440
rect 41106 585384 42246 585440
rect 42302 585384 42307 585440
rect 41045 585382 42307 585384
rect 41045 585379 41111 585382
rect 42241 585379 42307 585382
rect 39297 585170 39363 585173
rect 41822 585170 41828 585172
rect 39297 585168 41828 585170
rect 39297 585112 39302 585168
rect 39358 585112 41828 585168
rect 39297 585110 41828 585112
rect 39297 585107 39363 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 40217 584898 40283 584901
rect 41086 584898 41092 584900
rect 40217 584896 41092 584898
rect 40217 584840 40222 584896
rect 40278 584840 41092 584896
rect 40217 584838 41092 584840
rect 40217 584835 40283 584838
rect 41086 584836 41092 584838
rect 41156 584836 41162 584900
rect 39941 584626 40007 584629
rect 40350 584626 40356 584628
rect 39941 584624 40356 584626
rect 39941 584568 39946 584624
rect 40002 584568 40356 584624
rect 39941 584566 40356 584568
rect 39941 584563 40007 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 674925 584626 674991 584629
rect 676070 584626 676076 584628
rect 674925 584624 676076 584626
rect 674925 584568 674930 584624
rect 674986 584568 676076 584624
rect 674925 584566 676076 584568
rect 674925 584563 674991 584566
rect 676070 584564 676076 584566
rect 676140 584564 676146 584628
rect 41781 584354 41847 584357
rect 41781 584352 41890 584354
rect 41781 584296 41786 584352
rect 41842 584296 41890 584352
rect 41781 584291 41890 584296
rect 41830 583949 41890 584291
rect 41781 583944 41890 583949
rect 41781 583888 41786 583944
rect 41842 583888 41890 583944
rect 41781 583886 41890 583888
rect 41781 583883 41847 583886
rect 40350 581572 40356 581636
rect 40420 581634 40426 581636
rect 42609 581634 42675 581637
rect 40420 581632 42675 581634
rect 40420 581576 42614 581632
rect 42670 581576 42675 581632
rect 40420 581574 42675 581576
rect 40420 581572 40426 581574
rect 42609 581571 42675 581574
rect 42333 581226 42399 581229
rect 44173 581226 44239 581229
rect 42333 581224 44239 581226
rect 42333 581168 42338 581224
rect 42394 581168 44178 581224
rect 44234 581168 44239 581224
rect 42333 581166 44239 581168
rect 42333 581163 42399 581166
rect 44173 581163 44239 581166
rect 674005 581090 674071 581093
rect 674005 581088 676292 581090
rect 674005 581032 674010 581088
rect 674066 581032 676292 581088
rect 674005 581030 676292 581032
rect 674005 581027 674071 581030
rect 42057 580682 42123 580685
rect 44633 580682 44699 580685
rect 42057 580680 44699 580682
rect 42057 580624 42062 580680
rect 42118 580624 44638 580680
rect 44694 580624 44699 580680
rect 42057 580622 44699 580624
rect 42057 580619 42123 580622
rect 44633 580619 44699 580622
rect 676262 580549 676322 580652
rect 676213 580544 676322 580549
rect 676213 580488 676218 580544
rect 676274 580488 676322 580544
rect 676213 580486 676322 580488
rect 676213 580483 676279 580486
rect 41086 580212 41092 580276
rect 41156 580274 41162 580276
rect 41781 580274 41847 580277
rect 41156 580272 41847 580274
rect 41156 580216 41786 580272
rect 41842 580216 41847 580272
rect 41156 580214 41847 580216
rect 41156 580212 41162 580214
rect 41781 580211 41847 580214
rect 674005 580274 674071 580277
rect 674005 580272 676292 580274
rect 674005 580216 674010 580272
rect 674066 580216 676292 580272
rect 674005 580214 676292 580216
rect 674005 580211 674071 580214
rect 676397 580138 676463 580141
rect 676397 580136 676506 580138
rect 676397 580080 676402 580136
rect 676458 580080 676506 580136
rect 676397 580075 676506 580080
rect 676446 579836 676506 580075
rect 676262 579325 676322 579428
rect 676213 579320 676322 579325
rect 676213 579264 676218 579320
rect 676274 579264 676322 579320
rect 676213 579262 676322 579264
rect 676213 579259 676279 579262
rect 674005 579050 674071 579053
rect 674005 579048 676292 579050
rect 674005 578992 674010 579048
rect 674066 578992 676292 579048
rect 674005 578990 676292 578992
rect 674005 578987 674071 578990
rect 42149 578914 42215 578917
rect 45553 578914 45619 578917
rect 42149 578912 45619 578914
rect 42149 578856 42154 578912
rect 42210 578856 45558 578912
rect 45614 578856 45619 578912
rect 42149 578854 45619 578856
rect 42149 578851 42215 578854
rect 45553 578851 45619 578854
rect 676262 578509 676322 578612
rect 676213 578504 676322 578509
rect 676213 578448 676218 578504
rect 676274 578448 676322 578504
rect 676213 578446 676322 578448
rect 676213 578443 676279 578446
rect 676262 578101 676322 578204
rect 42057 578098 42123 578101
rect 44357 578098 44423 578101
rect 42057 578096 44423 578098
rect 42057 578040 42062 578096
rect 42118 578040 44362 578096
rect 44418 578040 44423 578096
rect 42057 578038 44423 578040
rect 42057 578035 42123 578038
rect 44357 578035 44423 578038
rect 676213 578096 676322 578101
rect 676213 578040 676218 578096
rect 676274 578040 676322 578096
rect 676213 578038 676322 578040
rect 676213 578035 676279 578038
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 676262 577693 676322 577796
rect 676213 577688 676322 577693
rect 676213 577632 676218 577688
rect 676274 577632 676322 577688
rect 676213 577630 676322 577632
rect 676213 577627 676279 577630
rect 675845 577418 675911 577421
rect 675845 577416 676292 577418
rect 675845 577360 675850 577416
rect 675906 577360 676292 577416
rect 675845 577358 676292 577360
rect 675845 577355 675911 577358
rect 674005 577010 674071 577013
rect 674005 577008 676292 577010
rect 674005 576952 674010 577008
rect 674066 576952 676292 577008
rect 674005 576950 676292 576952
rect 674005 576947 674071 576950
rect 672717 576602 672783 576605
rect 672717 576600 676292 576602
rect 672717 576544 672722 576600
rect 672778 576544 676292 576600
rect 672717 576542 676292 576544
rect 672717 576539 672783 576542
rect 676262 576061 676322 576164
rect 676213 576056 676322 576061
rect 682377 576058 682443 576061
rect 676213 576000 676218 576056
rect 676274 576000 676322 576056
rect 676213 575998 676322 576000
rect 682334 576056 682443 576058
rect 682334 576000 682382 576056
rect 682438 576000 682443 576056
rect 676213 575995 676279 575998
rect 682334 575995 682443 576000
rect 40534 575724 40540 575788
rect 40604 575786 40610 575788
rect 42241 575786 42307 575789
rect 40604 575784 42307 575786
rect 40604 575728 42246 575784
rect 42302 575728 42307 575784
rect 682334 575756 682394 575995
rect 40604 575726 42307 575728
rect 40604 575724 40610 575726
rect 42241 575723 42307 575726
rect 676029 575514 676095 575517
rect 676029 575512 676322 575514
rect 676029 575456 676034 575512
rect 676090 575456 676322 575512
rect 676029 575454 676322 575456
rect 676029 575451 676095 575454
rect 676262 575348 676322 575454
rect 676262 574837 676322 574940
rect 62113 574834 62179 574837
rect 62113 574832 64706 574834
rect 62113 574776 62118 574832
rect 62174 574776 64706 574832
rect 62113 574774 64706 574776
rect 62113 574771 62179 574774
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 64646 574194 64706 574774
rect 676213 574832 676322 574837
rect 676213 574776 676218 574832
rect 676274 574776 676322 574832
rect 676213 574774 676322 574776
rect 676213 574771 676279 574774
rect 674005 574562 674071 574565
rect 674005 574560 676292 574562
rect 674005 574504 674010 574560
rect 674066 574504 676292 574560
rect 674005 574502 676292 574504
rect 674005 574499 674071 574502
rect 674005 574290 674071 574293
rect 674005 574288 676322 574290
rect 674005 574232 674010 574288
rect 674066 574232 676322 574288
rect 674005 574230 676322 574232
rect 674005 574227 674071 574230
rect 676262 574124 676322 574230
rect 676262 573613 676322 573716
rect 62113 573610 62179 573613
rect 62113 573608 64706 573610
rect 62113 573552 62118 573608
rect 62174 573552 64706 573608
rect 62113 573550 64706 573552
rect 62113 573547 62179 573550
rect 64646 573012 64706 573550
rect 676213 573608 676322 573613
rect 676213 573552 676218 573608
rect 676274 573552 676322 573608
rect 676213 573550 676322 573552
rect 683205 573610 683271 573613
rect 683205 573608 683314 573610
rect 683205 573552 683210 573608
rect 683266 573552 683314 573608
rect 676213 573547 676279 573550
rect 683205 573547 683314 573552
rect 683254 573308 683314 573547
rect 674005 573066 674071 573069
rect 674005 573064 676322 573066
rect 674005 573008 674010 573064
rect 674066 573008 676322 573064
rect 674005 573006 676322 573008
rect 674005 573003 674071 573006
rect 676262 572900 676322 573006
rect 41454 572732 41460 572796
rect 41524 572794 41530 572796
rect 42609 572794 42675 572797
rect 41524 572792 42675 572794
rect 41524 572736 42614 572792
rect 42670 572736 42675 572792
rect 41524 572734 42675 572736
rect 41524 572732 41530 572734
rect 42609 572731 42675 572734
rect 683389 572794 683455 572797
rect 683389 572792 683498 572794
rect 683389 572736 683394 572792
rect 683450 572736 683498 572792
rect 683389 572731 683498 572736
rect 683438 572492 683498 572731
rect 41965 572252 42031 572253
rect 41965 572248 42012 572252
rect 42076 572250 42082 572252
rect 41965 572192 41970 572248
rect 41965 572188 42012 572192
rect 42076 572190 42122 572250
rect 42076 572188 42082 572190
rect 41965 572187 42031 572188
rect 676262 571981 676322 572084
rect 676213 571976 676322 571981
rect 676213 571920 676218 571976
rect 676274 571920 676322 571976
rect 676213 571918 676322 571920
rect 676213 571915 676279 571918
rect 41638 571508 41644 571572
rect 41708 571570 41714 571572
rect 42057 571570 42123 571573
rect 41708 571568 42123 571570
rect 41708 571512 42062 571568
rect 42118 571512 42123 571568
rect 41708 571510 42123 571512
rect 41708 571508 41714 571510
rect 42057 571507 42123 571510
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 675477 571706 675543 571709
rect 675477 571704 676292 571706
rect 675477 571648 675482 571704
rect 675538 571648 676292 571704
rect 675477 571646 676292 571648
rect 675477 571643 675543 571646
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 42425 571371 42491 571374
rect 674833 571298 674899 571301
rect 674833 571296 676292 571298
rect 674833 571240 674838 571296
rect 674894 571240 676292 571296
rect 674833 571238 676292 571240
rect 674833 571235 674899 571238
rect 62941 571162 63007 571165
rect 62941 571160 64706 571162
rect 62941 571104 62946 571160
rect 63002 571104 64706 571160
rect 62941 571102 64706 571104
rect 62941 571099 63007 571102
rect 64646 570648 64706 571102
rect 676262 570757 676322 570860
rect 676213 570752 676322 570757
rect 676213 570696 676218 570752
rect 676274 570696 676322 570752
rect 676213 570694 676322 570696
rect 676213 570691 676279 570694
rect 676806 570692 676812 570756
rect 676876 570692 676882 570756
rect 676814 570482 676874 570692
rect 676476 570452 676874 570482
rect 676446 570422 676844 570452
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 676446 570044 676506 570422
rect 63125 569938 63191 569941
rect 63125 569936 64706 569938
rect 63125 569880 63130 569936
rect 63186 569880 64706 569936
rect 63125 569878 64706 569880
rect 63125 569875 63191 569878
rect 64646 569466 64706 569878
rect 676262 569533 676322 569636
rect 676213 569528 676322 569533
rect 676213 569472 676218 569528
rect 676274 569472 676322 569528
rect 676213 569470 676322 569472
rect 676213 569467 676279 569470
rect 62757 568578 62823 568581
rect 62757 568576 64706 568578
rect 62757 568520 62762 568576
rect 62818 568520 64706 568576
rect 62757 568518 64706 568520
rect 62757 568515 62823 568518
rect 64646 568284 64706 568518
rect 673821 565858 673887 565861
rect 675385 565858 675451 565861
rect 673821 565856 675451 565858
rect 673821 565800 673826 565856
rect 673882 565800 675390 565856
rect 675446 565800 675451 565856
rect 673821 565798 675451 565800
rect 673821 565795 673887 565798
rect 675385 565795 675451 565798
rect 675385 563140 675451 563141
rect 675334 563138 675340 563140
rect 675294 563078 675340 563138
rect 675404 563136 675451 563140
rect 675446 563080 675451 563136
rect 675334 563076 675340 563078
rect 675404 563076 675451 563080
rect 675385 563075 675451 563076
rect 667749 561914 667815 561917
rect 675109 561914 675175 561917
rect 667749 561912 675175 561914
rect 667749 561856 667754 561912
rect 667810 561856 675114 561912
rect 675170 561856 675175 561912
rect 667749 561854 675175 561856
rect 667749 561851 667815 561854
rect 675109 561851 675175 561854
rect 674414 558996 674420 559060
rect 674484 559058 674490 559060
rect 675109 559058 675175 559061
rect 674484 559056 675175 559058
rect 674484 559000 675114 559056
rect 675170 559000 675175 559056
rect 674484 558998 675175 559000
rect 674484 558996 674490 558998
rect 675109 558995 675175 558998
rect 41086 558724 41092 558788
rect 41156 558786 41162 558788
rect 45093 558786 45159 558789
rect 41156 558784 45159 558786
rect 41156 558728 45098 558784
rect 45154 558728 45159 558784
rect 41156 558726 45159 558728
rect 41156 558724 41162 558726
rect 45093 558723 45159 558726
rect 41492 558454 51090 558514
rect 42241 558106 42307 558109
rect 41492 558104 42307 558106
rect 41492 558048 42246 558104
rect 42302 558048 42307 558104
rect 41492 558046 42307 558048
rect 42241 558043 42307 558046
rect 41492 557638 48330 557698
rect 41086 557488 41092 557552
rect 41156 557488 41162 557552
rect 41094 557260 41154 557488
rect 48270 557290 48330 557638
rect 51030 557562 51090 558454
rect 61377 557562 61443 557565
rect 51030 557560 61443 557562
rect 51030 557504 61382 557560
rect 61438 557504 61443 557560
rect 51030 557502 61443 557504
rect 61377 557499 61443 557502
rect 48270 557230 51090 557290
rect 44541 556882 44607 556885
rect 41492 556880 44607 556882
rect 41492 556824 44546 556880
rect 44602 556824 44607 556880
rect 41492 556822 44607 556824
rect 44541 556819 44607 556822
rect 51030 556746 51090 557230
rect 63401 556746 63467 556749
rect 51030 556744 63467 556746
rect 51030 556688 63406 556744
rect 63462 556688 63467 556744
rect 51030 556686 63467 556688
rect 63401 556683 63467 556686
rect 42977 556474 43043 556477
rect 41492 556472 43043 556474
rect 41492 556416 42982 556472
rect 43038 556416 43043 556472
rect 41492 556414 43043 556416
rect 42977 556411 43043 556414
rect 44265 556066 44331 556069
rect 41492 556064 44331 556066
rect 41492 556008 44270 556064
rect 44326 556008 44331 556064
rect 41492 556006 44331 556008
rect 44265 556003 44331 556006
rect 44909 555658 44975 555661
rect 41492 555656 44975 555658
rect 41492 555600 44914 555656
rect 44970 555600 44975 555656
rect 41492 555598 44975 555600
rect 44909 555595 44975 555598
rect 45645 555250 45711 555253
rect 41492 555248 45711 555250
rect 41492 555192 45650 555248
rect 45706 555192 45711 555248
rect 41492 555190 45711 555192
rect 45645 555187 45711 555190
rect 668669 555250 668735 555253
rect 675385 555250 675451 555253
rect 668669 555248 675451 555250
rect 668669 555192 668674 555248
rect 668730 555192 675390 555248
rect 675446 555192 675451 555248
rect 668669 555190 675451 555192
rect 668669 555187 668735 555190
rect 675385 555187 675451 555190
rect 42793 554842 42859 554845
rect 41492 554840 42859 554842
rect 41492 554784 42798 554840
rect 42854 554784 42859 554840
rect 41492 554782 42859 554784
rect 42793 554779 42859 554782
rect 673821 554842 673887 554845
rect 675293 554842 675359 554845
rect 673821 554840 675359 554842
rect 673821 554784 673826 554840
rect 673882 554784 675298 554840
rect 675354 554784 675359 554840
rect 673821 554782 675359 554784
rect 673821 554779 673887 554782
rect 675293 554779 675359 554782
rect 45829 554434 45895 554437
rect 41492 554432 45895 554434
rect 41492 554376 45834 554432
rect 45890 554376 45895 554432
rect 41492 554374 45895 554376
rect 45829 554371 45895 554374
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 675753 554026 675819 554029
rect 676806 554026 676812 554028
rect 675753 554024 676812 554026
rect 675753 553968 675758 554024
rect 675814 553968 676812 554024
rect 675753 553966 676812 553968
rect 675753 553963 675819 553966
rect 676806 553964 676812 553966
rect 676876 553964 676882 554028
rect 39990 553413 40050 553588
rect 649950 553482 650010 553914
rect 673821 553754 673887 553757
rect 675109 553754 675175 553757
rect 673821 553752 675175 553754
rect 673821 553696 673826 553752
rect 673882 553696 675114 553752
rect 675170 553696 675175 553752
rect 673821 553694 675175 553696
rect 673821 553691 673887 553694
rect 675109 553691 675175 553694
rect 651465 553482 651531 553485
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 651465 553419 651531 553422
rect 39990 553408 40099 553413
rect 39990 553352 40038 553408
rect 40094 553352 40099 553408
rect 39990 553350 40099 553352
rect 40033 553347 40099 553350
rect 40861 553410 40927 553413
rect 40861 553408 40970 553410
rect 40861 553352 40866 553408
rect 40922 553352 40970 553408
rect 40861 553347 40970 553352
rect 40910 553180 40970 553347
rect 672901 553346 672967 553349
rect 675385 553346 675451 553349
rect 672901 553344 675451 553346
rect 672901 553288 672906 553344
rect 672962 553288 675390 553344
rect 675446 553288 675451 553344
rect 672901 553286 675451 553288
rect 672901 553283 672967 553286
rect 675385 553283 675451 553286
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 42241 552666 42307 552669
rect 62941 552666 63007 552669
rect 42241 552664 63007 552666
rect 42241 552608 42246 552664
rect 42302 552608 62946 552664
rect 63002 552608 63007 552664
rect 42241 552606 63007 552608
rect 42241 552603 42307 552606
rect 62941 552603 63007 552606
rect 42977 552394 43043 552397
rect 41492 552392 43043 552394
rect 41492 552336 42982 552392
rect 43038 552336 43043 552392
rect 41492 552334 43043 552336
rect 649950 552394 650010 552732
rect 651465 552394 651531 552397
rect 649950 552392 651531 552394
rect 649950 552336 651470 552392
rect 651526 552336 651531 552392
rect 649950 552334 651531 552336
rect 42977 552331 43043 552334
rect 651465 552331 651531 552334
rect 670417 552122 670483 552125
rect 675293 552122 675359 552125
rect 670417 552120 675359 552122
rect 670417 552064 670422 552120
rect 670478 552064 675298 552120
rect 675354 552064 675359 552120
rect 670417 552062 675359 552064
rect 670417 552059 670483 552062
rect 675293 552059 675359 552062
rect 34421 551986 34487 551989
rect 34421 551984 34500 551986
rect 34421 551928 34426 551984
rect 34482 551928 34500 551984
rect 34421 551926 34500 551928
rect 34421 551923 34487 551926
rect 45185 551578 45251 551581
rect 41492 551576 45251 551578
rect 41492 551520 45190 551576
rect 45246 551520 45251 551576
rect 41492 551518 45251 551520
rect 45185 551515 45251 551518
rect 42793 551170 42859 551173
rect 41492 551168 42859 551170
rect 41492 551112 42798 551168
rect 42854 551112 42859 551168
rect 41492 551110 42859 551112
rect 649950 551170 650010 551550
rect 651465 551170 651531 551173
rect 649950 551168 651531 551170
rect 649950 551112 651470 551168
rect 651526 551112 651531 551168
rect 649950 551110 651531 551112
rect 42793 551107 42859 551110
rect 651465 551107 651531 551110
rect 41462 550762 42074 550796
rect 45369 550762 45435 550765
rect 41462 550760 45435 550762
rect 41462 550736 45374 550760
rect 41462 550732 41522 550736
rect 42014 550704 45374 550736
rect 45430 550704 45435 550760
rect 42014 550702 45435 550704
rect 45369 550699 45435 550702
rect 41781 550628 41847 550629
rect 41781 550626 41828 550628
rect 41736 550624 41828 550626
rect 41736 550568 41786 550624
rect 41736 550566 41828 550568
rect 41781 550564 41828 550566
rect 41892 550564 41898 550628
rect 41781 550563 41847 550564
rect 41873 550354 41939 550357
rect 41492 550352 41939 550354
rect 41492 550296 41878 550352
rect 41934 550296 41939 550352
rect 41492 550294 41939 550296
rect 649950 550354 650010 550368
rect 651373 550354 651439 550357
rect 649950 550352 651439 550354
rect 649950 550296 651378 550352
rect 651434 550296 651439 550352
rect 649950 550294 651439 550296
rect 41873 550291 41939 550294
rect 651373 550291 651439 550294
rect 675753 550354 675819 550357
rect 676990 550354 676996 550356
rect 675753 550352 676996 550354
rect 675753 550296 675758 550352
rect 675814 550296 676996 550352
rect 675753 550294 676996 550296
rect 675753 550291 675819 550294
rect 676990 550292 676996 550294
rect 677060 550292 677066 550356
rect 42057 549946 42123 549949
rect 41492 549944 42123 549946
rect 41492 549888 42062 549944
rect 42118 549888 42123 549944
rect 41492 549886 42123 549888
rect 42057 549883 42123 549886
rect 43069 549538 43135 549541
rect 41492 549536 43135 549538
rect 41492 549480 43074 549536
rect 43130 549480 43135 549536
rect 41492 549478 43135 549480
rect 43069 549475 43135 549478
rect 45001 549130 45067 549133
rect 41492 549128 45067 549130
rect 41492 549072 45006 549128
rect 45062 549072 45067 549128
rect 41492 549070 45067 549072
rect 649950 549130 650010 549186
rect 651465 549130 651531 549133
rect 649950 549128 651531 549130
rect 649950 549072 651470 549128
rect 651526 549072 651531 549128
rect 649950 549070 651531 549072
rect 45001 549067 45067 549070
rect 651465 549067 651531 549070
rect 44725 548722 44791 548725
rect 41492 548720 44791 548722
rect 41492 548664 44730 548720
rect 44786 548664 44791 548720
rect 41492 548662 44791 548664
rect 44725 548659 44791 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 43805 548314 43871 548317
rect 41492 548312 43871 548314
rect 41492 548256 43810 548312
rect 43866 548256 43871 548312
rect 41492 548254 43871 548256
rect 43805 548251 43871 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 670969 548450 671035 548453
rect 675477 548450 675543 548453
rect 670969 548448 675543 548450
rect 670969 548392 670974 548448
rect 671030 548392 675482 548448
rect 675538 548392 675543 548448
rect 670969 548390 675543 548392
rect 670969 548387 671035 548390
rect 675477 548387 675543 548390
rect 674005 547906 674071 547909
rect 675477 547906 675543 547909
rect 674005 547904 675543 547906
rect 28766 547498 28826 547890
rect 674005 547848 674010 547904
rect 674066 547848 675482 547904
rect 675538 547848 675543 547904
rect 674005 547846 675543 547848
rect 674005 547843 674071 547846
rect 675477 547843 675543 547846
rect 674005 547634 674071 547637
rect 675661 547634 675727 547637
rect 674005 547632 675727 547634
rect 674005 547576 674010 547632
rect 674066 547576 675666 547632
rect 675722 547576 675727 547632
rect 674005 547574 675727 547576
rect 674005 547571 674071 547574
rect 675661 547571 675727 547574
rect 675886 547572 675892 547636
rect 675956 547634 675962 547636
rect 678237 547634 678303 547637
rect 675956 547632 678303 547634
rect 675956 547576 678242 547632
rect 678298 547576 678303 547632
rect 675956 547574 678303 547576
rect 675956 547572 675962 547574
rect 678237 547571 678303 547574
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 43989 547090 44055 547093
rect 41492 547088 44055 547090
rect 41492 547032 43994 547088
rect 44050 547032 44055 547088
rect 41492 547030 44055 547032
rect 43989 547027 44055 547030
rect 674230 547028 674236 547092
rect 674300 547090 674306 547092
rect 683481 547090 683547 547093
rect 674300 547088 683547 547090
rect 674300 547032 683486 547088
rect 683542 547032 683547 547088
rect 674300 547030 683547 547032
rect 674300 547028 674306 547030
rect 683481 547027 683547 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 682377 546818 682443 546821
rect 676140 546816 682443 546818
rect 676140 546760 682382 546816
rect 682438 546760 682443 546816
rect 676140 546758 682443 546760
rect 676140 546756 676146 546758
rect 682377 546755 682443 546758
rect 40718 545668 40724 545732
rect 40788 545730 40794 545732
rect 41873 545730 41939 545733
rect 40788 545728 41939 545730
rect 40788 545672 41878 545728
rect 41934 545672 41939 545728
rect 40788 545670 41939 545672
rect 40788 545668 40794 545670
rect 41873 545667 41939 545670
rect 675334 545532 675340 545596
rect 675404 545594 675410 545596
rect 675569 545594 675635 545597
rect 675404 545592 675635 545594
rect 675404 545536 675574 545592
rect 675630 545536 675635 545592
rect 675404 545534 675635 545536
rect 675404 545532 675410 545534
rect 675569 545531 675635 545534
rect 40534 545396 40540 545460
rect 40604 545458 40610 545460
rect 42057 545458 42123 545461
rect 40604 545456 42123 545458
rect 40604 545400 42062 545456
rect 42118 545400 42123 545456
rect 40604 545398 42123 545400
rect 40604 545396 40610 545398
rect 42057 545395 42123 545398
rect 37825 541378 37891 541381
rect 37825 541376 40418 541378
rect 37825 541320 37830 541376
rect 37886 541320 40418 541376
rect 37825 541318 40418 541320
rect 37825 541315 37891 541318
rect 40358 540698 40418 541318
rect 41781 541106 41847 541109
rect 41781 541104 42074 541106
rect 41781 541048 41786 541104
rect 41842 541048 42074 541104
rect 41781 541046 42074 541048
rect 41781 541043 41847 541046
rect 41781 540698 41847 540701
rect 40358 540696 41847 540698
rect 40358 540640 41786 540696
rect 41842 540640 41847 540696
rect 40358 540638 41847 540640
rect 42014 540698 42074 541046
rect 42241 540698 42307 540701
rect 42014 540696 42307 540698
rect 42014 540640 42246 540696
rect 42302 540640 42307 540696
rect 42014 540638 42307 540640
rect 41781 540635 41847 540638
rect 42241 540635 42307 540638
rect 42517 539610 42583 539613
rect 59997 539610 60063 539613
rect 42517 539608 60063 539610
rect 42517 539552 42522 539608
rect 42578 539552 60002 539608
rect 60058 539552 60063 539608
rect 42517 539550 60063 539552
rect 42517 539547 42583 539550
rect 59997 539547 60063 539550
rect 42609 538114 42675 538117
rect 45001 538114 45067 538117
rect 42609 538112 45067 538114
rect 42609 538056 42614 538112
rect 42670 538056 45006 538112
rect 45062 538056 45067 538112
rect 42609 538054 45067 538056
rect 42609 538051 42675 538054
rect 45001 538051 45067 538054
rect 40534 537372 40540 537436
rect 40604 537434 40610 537436
rect 42425 537434 42491 537437
rect 40604 537432 42491 537434
rect 40604 537376 42430 537432
rect 42486 537376 42491 537432
rect 40604 537374 42491 537376
rect 40604 537372 40610 537374
rect 42425 537371 42491 537374
rect 40718 536964 40724 537028
rect 40788 537026 40794 537028
rect 41781 537026 41847 537029
rect 40788 537024 41847 537026
rect 40788 536968 41786 537024
rect 41842 536968 41847 537024
rect 40788 536966 41847 536968
rect 40788 536964 40794 536966
rect 41781 536963 41847 536966
rect 44725 536890 44791 536893
rect 42198 536888 44791 536890
rect 42198 536832 44730 536888
rect 44786 536832 44791 536888
rect 42198 536830 44791 536832
rect 42198 536485 42258 536830
rect 44725 536827 44791 536830
rect 42198 536480 42307 536485
rect 42198 536424 42246 536480
rect 42302 536424 42307 536480
rect 42198 536422 42307 536424
rect 42241 536419 42307 536422
rect 674189 536074 674255 536077
rect 676262 536074 676322 536112
rect 674189 536072 676322 536074
rect 674189 536016 674194 536072
rect 674250 536016 676322 536072
rect 674189 536014 676322 536016
rect 674189 536011 674255 536014
rect 42057 535666 42123 535669
rect 44725 535666 44791 535669
rect 42057 535664 44791 535666
rect 42057 535608 42062 535664
rect 42118 535608 44730 535664
rect 44786 535608 44791 535664
rect 42057 535606 44791 535608
rect 42057 535603 42123 535606
rect 44725 535603 44791 535606
rect 674005 535666 674071 535669
rect 676262 535666 676322 535704
rect 674005 535664 676322 535666
rect 674005 535608 674010 535664
rect 674066 535608 676322 535664
rect 674005 535606 676322 535608
rect 674005 535603 674071 535606
rect 674005 535258 674071 535261
rect 676262 535258 676322 535296
rect 674005 535256 676322 535258
rect 674005 535200 674010 535256
rect 674066 535200 676322 535256
rect 674005 535198 676322 535200
rect 674005 535195 674071 535198
rect 672717 534986 672783 534989
rect 672717 534984 676322 534986
rect 672717 534928 672722 534984
rect 672778 534928 676322 534984
rect 672717 534926 676322 534928
rect 672717 534923 672783 534926
rect 676262 534888 676322 534926
rect 674189 534442 674255 534445
rect 676262 534442 676322 534480
rect 674189 534440 676322 534442
rect 674189 534384 674194 534440
rect 674250 534384 676322 534440
rect 674189 534382 676322 534384
rect 674189 534379 674255 534382
rect 671521 534170 671587 534173
rect 671521 534168 676322 534170
rect 671521 534112 671526 534168
rect 671582 534112 676322 534168
rect 671521 534110 676322 534112
rect 671521 534107 671587 534110
rect 676262 534072 676322 534110
rect 672717 533490 672783 533493
rect 676262 533490 676322 533664
rect 672717 533488 676322 533490
rect 672717 533432 672722 533488
rect 672778 533432 676322 533488
rect 672717 533430 676322 533432
rect 672717 533427 672783 533430
rect 674005 533218 674071 533221
rect 676262 533218 676322 533256
rect 674005 533216 676322 533218
rect 674005 533160 674010 533216
rect 674066 533160 676322 533216
rect 674005 533158 676322 533160
rect 674005 533155 674071 533158
rect 42701 532810 42767 532813
rect 45369 532810 45435 532813
rect 42701 532808 45435 532810
rect 42701 532752 42706 532808
rect 42762 532752 45374 532808
rect 45430 532752 45435 532808
rect 42701 532750 45435 532752
rect 42701 532747 42767 532750
rect 45369 532747 45435 532750
rect 674005 532810 674071 532813
rect 676262 532810 676322 532848
rect 674005 532808 676322 532810
rect 674005 532752 674010 532808
rect 674066 532752 676322 532808
rect 674005 532750 676322 532752
rect 674005 532747 674071 532750
rect 674005 532402 674071 532405
rect 676262 532402 676322 532440
rect 674005 532400 676322 532402
rect 674005 532344 674010 532400
rect 674066 532344 676322 532400
rect 674005 532342 676322 532344
rect 674005 532339 674071 532342
rect 674189 531994 674255 531997
rect 676262 531994 676322 532032
rect 674189 531992 676322 531994
rect 674189 531936 674194 531992
rect 674250 531936 676322 531992
rect 674189 531934 676322 531936
rect 674189 531931 674255 531934
rect 678237 531858 678303 531861
rect 678237 531856 678346 531858
rect 678237 531800 678242 531856
rect 678298 531800 678346 531856
rect 678237 531795 678346 531800
rect 678286 531624 678346 531795
rect 62297 531178 62363 531181
rect 674005 531178 674071 531181
rect 676262 531178 676322 531216
rect 62297 531176 64706 531178
rect 62297 531120 62302 531176
rect 62358 531120 64706 531176
rect 62297 531118 64706 531120
rect 674005 531176 676322 531178
rect 674005 531120 674010 531176
rect 674066 531120 676322 531176
rect 674005 531118 676322 531120
rect 62297 531115 62363 531118
rect 674005 531115 674071 531118
rect 41454 530708 41460 530772
rect 41524 530770 41530 530772
rect 42609 530770 42675 530773
rect 41524 530768 42675 530770
rect 41524 530712 42614 530768
rect 42670 530712 42675 530768
rect 41524 530710 42675 530712
rect 41524 530708 41530 530710
rect 42609 530707 42675 530710
rect 674189 530770 674255 530773
rect 676262 530770 676322 530808
rect 674189 530768 676322 530770
rect 674189 530712 674194 530768
rect 674250 530712 676322 530768
rect 674189 530710 676322 530712
rect 674189 530707 674255 530710
rect 62113 530634 62179 530637
rect 682377 530634 682443 530637
rect 62113 530632 64706 530634
rect 62113 530576 62118 530632
rect 62174 530576 64706 530632
rect 62113 530574 64706 530576
rect 62113 530571 62179 530574
rect 64646 529990 64706 530574
rect 682334 530632 682443 530634
rect 682334 530576 682382 530632
rect 682438 530576 682443 530632
rect 682334 530571 682443 530576
rect 682334 530400 682394 530571
rect 674005 530090 674071 530093
rect 674005 530088 676322 530090
rect 674005 530032 674010 530088
rect 674066 530032 676322 530088
rect 674005 530030 676322 530032
rect 674005 530027 674071 530030
rect 676262 529992 676322 530030
rect 41822 529484 41828 529548
rect 41892 529546 41898 529548
rect 42425 529546 42491 529549
rect 41892 529544 42491 529546
rect 41892 529488 42430 529544
rect 42486 529488 42491 529544
rect 41892 529486 42491 529488
rect 41892 529484 41898 529486
rect 42425 529483 42491 529486
rect 674189 529546 674255 529549
rect 676262 529546 676322 529584
rect 674189 529544 676322 529546
rect 674189 529488 674194 529544
rect 674250 529488 676322 529544
rect 674189 529486 676322 529488
rect 674189 529483 674255 529486
rect 41638 529212 41644 529276
rect 41708 529274 41714 529276
rect 41708 529214 41890 529274
rect 41708 529212 41714 529214
rect 41830 529005 41890 529214
rect 674005 529138 674071 529141
rect 676262 529138 676322 529176
rect 674005 529136 676322 529138
rect 674005 529080 674010 529136
rect 674066 529080 676322 529136
rect 674005 529078 676322 529080
rect 674005 529075 674071 529078
rect 41830 529000 41939 529005
rect 41830 528944 41878 529000
rect 41934 528944 41939 529000
rect 41830 528942 41939 528944
rect 41873 528939 41939 528942
rect 42241 529002 42307 529005
rect 45185 529002 45251 529005
rect 42241 529000 45251 529002
rect 42241 528944 42246 529000
rect 42302 528944 45190 529000
rect 45246 528944 45251 529000
rect 42241 528942 45251 528944
rect 42241 528939 42307 528942
rect 45185 528939 45251 528942
rect 673085 528866 673151 528869
rect 673085 528864 676322 528866
rect 673085 528808 673090 528864
rect 673146 528808 676322 528864
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 673085 528806 676322 528808
rect 673085 528803 673151 528806
rect 676262 528768 676322 528806
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 62113 528531 62179 528534
rect 673637 528186 673703 528189
rect 676262 528186 676322 528360
rect 673637 528184 676322 528186
rect 673637 528128 673642 528184
rect 673698 528128 676322 528184
rect 673637 528126 676322 528128
rect 673637 528123 673703 528126
rect 63401 528050 63467 528053
rect 63401 528048 64706 528050
rect 63401 527992 63406 528048
rect 63462 527992 64706 528048
rect 63401 527990 64706 527992
rect 63401 527987 63467 527990
rect 64646 527626 64706 527990
rect 674005 527914 674071 527917
rect 676262 527914 676322 527952
rect 674005 527912 676322 527914
rect 674005 527856 674010 527912
rect 674066 527856 676322 527912
rect 674005 527854 676322 527856
rect 674005 527851 674071 527854
rect 684309 527778 684375 527781
rect 684309 527776 684418 527778
rect 684309 527720 684314 527776
rect 684370 527720 684418 527776
rect 684309 527715 684418 527720
rect 684358 527544 684418 527715
rect 683481 527370 683547 527373
rect 683438 527368 683547 527370
rect 683438 527312 683486 527368
rect 683542 527312 683547 527368
rect 683438 527307 683547 527312
rect 42609 527234 42675 527237
rect 45093 527234 45159 527237
rect 42609 527232 45159 527234
rect 42609 527176 42614 527232
rect 42670 527176 45098 527232
rect 45154 527176 45159 527232
rect 42609 527174 45159 527176
rect 42609 527171 42675 527174
rect 45093 527171 45159 527174
rect 683438 527136 683498 527307
rect 61377 527098 61443 527101
rect 61377 527096 64706 527098
rect 61377 527040 61382 527096
rect 61438 527040 64706 527096
rect 61377 527038 64706 527040
rect 61377 527035 61443 527038
rect 64646 526444 64706 527038
rect 673545 526826 673611 526829
rect 673545 526824 676322 526826
rect 673545 526768 673550 526824
rect 673606 526768 676322 526824
rect 673545 526766 676322 526768
rect 673545 526763 673611 526766
rect 676262 526728 676322 526766
rect 683297 526554 683363 526557
rect 683254 526552 683363 526554
rect 683254 526496 683302 526552
rect 683358 526496 683363 526552
rect 683254 526491 683363 526496
rect 683254 526320 683314 526491
rect 683254 525741 683314 525912
rect 62941 525738 63007 525741
rect 62941 525736 64706 525738
rect 62941 525680 62946 525736
rect 63002 525680 64706 525736
rect 62941 525678 64706 525680
rect 683254 525736 683363 525741
rect 683254 525680 683302 525736
rect 683358 525680 683363 525736
rect 683254 525678 683363 525680
rect 62941 525675 63007 525678
rect 64646 525262 64706 525678
rect 683297 525675 683363 525678
rect 682886 525330 682946 525504
rect 683113 525330 683179 525333
rect 682886 525328 683179 525330
rect 682886 525272 683118 525328
rect 683174 525272 683179 525328
rect 682886 525270 683179 525272
rect 682886 525096 682946 525270
rect 683113 525267 683179 525270
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683573 503706 683639 503709
rect 677060 503704 683639 503706
rect 677060 503648 683578 503704
rect 683634 503648 683639 503704
rect 677060 503646 683639 503648
rect 677060 503644 677066 503646
rect 683573 503643 683639 503646
rect 673821 492146 673887 492149
rect 673821 492144 676292 492146
rect 673821 492088 673826 492144
rect 673882 492088 676292 492144
rect 673821 492086 676292 492088
rect 673821 492083 673887 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 675845 491330 675911 491333
rect 675845 491328 676292 491330
rect 675845 491272 675850 491328
rect 675906 491272 676292 491328
rect 675845 491270 676292 491272
rect 675845 491267 675911 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 675845 490514 675911 490517
rect 675845 490512 676292 490514
rect 675845 490456 675850 490512
rect 675906 490456 676292 490512
rect 675845 490454 676292 490456
rect 675845 490451 675911 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 672625 489698 672691 489701
rect 672625 489696 676292 489698
rect 672625 489640 672630 489696
rect 672686 489640 676292 489696
rect 672625 489638 676292 489640
rect 672625 489635 672691 489638
rect 673913 489290 673979 489293
rect 673913 489288 676292 489290
rect 673913 489232 673918 489288
rect 673974 489232 676292 489288
rect 673913 489230 676292 489232
rect 673913 489227 673979 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 673913 488474 673979 488477
rect 673913 488472 676292 488474
rect 673913 488416 673918 488472
rect 673974 488416 676292 488472
rect 673913 488414 676292 488416
rect 673913 488411 673979 488414
rect 676170 488006 676292 488066
rect 675886 487868 675892 487932
rect 675956 487930 675962 487932
rect 676170 487930 676230 488006
rect 675956 487870 676230 487930
rect 675956 487868 675962 487870
rect 676029 487658 676095 487661
rect 676029 487656 676292 487658
rect 676029 487600 676034 487656
rect 676090 487600 676292 487656
rect 676029 487598 676292 487600
rect 676029 487595 676095 487598
rect 683573 487250 683639 487253
rect 683573 487248 683652 487250
rect 683573 487192 683578 487248
rect 683634 487192 683652 487248
rect 683573 487190 683652 487192
rect 683573 487187 683639 487190
rect 678237 486842 678303 486845
rect 678237 486840 678316 486842
rect 678237 486784 678242 486840
rect 678298 486784 678316 486840
rect 678237 486782 678316 486784
rect 678237 486779 678303 486782
rect 683205 486434 683271 486437
rect 683205 486432 683284 486434
rect 683205 486376 683210 486432
rect 683266 486376 683284 486432
rect 683205 486374 683284 486376
rect 683205 486371 683271 486374
rect 673913 486026 673979 486029
rect 673913 486024 676292 486026
rect 673913 485968 673918 486024
rect 673974 485968 676292 486024
rect 673913 485966 676292 485968
rect 673913 485963 673979 485966
rect 674005 485618 674071 485621
rect 674005 485616 676292 485618
rect 674005 485560 674010 485616
rect 674066 485560 676292 485616
rect 674005 485558 676292 485560
rect 674005 485555 674071 485558
rect 674005 485210 674071 485213
rect 674005 485208 676292 485210
rect 674005 485152 674010 485208
rect 674066 485152 676292 485208
rect 674005 485150 676292 485152
rect 674005 485147 674071 485150
rect 674414 484740 674420 484804
rect 674484 484802 674490 484804
rect 674484 484742 676292 484802
rect 674484 484740 674490 484742
rect 674189 484394 674255 484397
rect 674189 484392 676292 484394
rect 674189 484336 674194 484392
rect 674250 484336 676292 484392
rect 674189 484334 676292 484336
rect 674189 484331 674255 484334
rect 674005 483986 674071 483989
rect 674005 483984 676292 483986
rect 674005 483928 674010 483984
rect 674066 483928 676292 483984
rect 674005 483926 676292 483928
rect 674005 483923 674071 483926
rect 675886 483516 675892 483580
rect 675956 483578 675962 483580
rect 675956 483518 676292 483578
rect 675956 483516 675962 483518
rect 674649 483170 674715 483173
rect 674649 483168 676292 483170
rect 674649 483112 674654 483168
rect 674710 483112 676292 483168
rect 674649 483110 676292 483112
rect 674649 483107 674715 483110
rect 674465 482762 674531 482765
rect 674465 482760 676292 482762
rect 674465 482704 674470 482760
rect 674526 482704 676292 482760
rect 674465 482702 676292 482704
rect 674465 482699 674531 482702
rect 672901 482354 672967 482357
rect 672901 482352 676292 482354
rect 672901 482296 672906 482352
rect 672962 482296 676292 482352
rect 672901 482294 676292 482296
rect 672901 482291 672967 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675661 480722 675727 480725
rect 675661 480720 676292 480722
rect 675661 480664 675666 480720
rect 675722 480664 676292 480720
rect 675661 480662 676292 480664
rect 675661 480659 675727 480662
rect 670049 455426 670115 455429
rect 673269 455426 673335 455429
rect 670049 455424 673335 455426
rect 670049 455368 670054 455424
rect 670110 455368 673274 455424
rect 673330 455368 673335 455424
rect 670049 455366 673335 455368
rect 670049 455363 670115 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 673085 455018 673151 455021
rect 674281 455018 674347 455021
rect 673085 455016 674347 455018
rect 673085 454960 673090 455016
rect 673146 454960 674286 455016
rect 674342 454960 674347 455016
rect 673085 454958 674347 454960
rect 673085 454955 673151 454958
rect 674281 454955 674347 454958
rect 672901 454746 672967 454749
rect 674281 454746 674347 454749
rect 672901 454744 674347 454746
rect 672901 454688 672906 454744
rect 672962 454688 674286 454744
rect 674342 454688 674347 454744
rect 672901 454686 674347 454688
rect 672901 454683 672967 454686
rect 674281 454683 674347 454686
rect 672809 454474 672875 454477
rect 674281 454474 674347 454477
rect 672809 454472 674347 454474
rect 672809 454416 672814 454472
rect 672870 454416 674286 454472
rect 674342 454416 674347 454472
rect 672809 454414 674347 454416
rect 672809 454411 672875 454414
rect 674281 454411 674347 454414
rect 672441 453930 672507 453933
rect 675293 453930 675359 453933
rect 672441 453928 675359 453930
rect 672441 453872 672446 453928
rect 672502 453872 675298 453928
rect 675354 453872 675359 453928
rect 672441 453870 675359 453872
rect 672441 453867 672507 453870
rect 675293 453867 675359 453870
rect 675334 447748 675340 447812
rect 675404 447810 675410 447812
rect 675937 447810 676003 447813
rect 675404 447808 676003 447810
rect 675404 447752 675942 447808
rect 675998 447752 676003 447808
rect 675404 447750 676003 447752
rect 675404 447748 675410 447750
rect 675937 447747 676003 447750
rect 41492 430886 55230 430946
rect 55170 430674 55230 430886
rect 59997 430674 60063 430677
rect 55170 430672 60063 430674
rect 55170 430616 60002 430672
rect 60058 430616 60063 430672
rect 55170 430614 60063 430616
rect 59997 430611 60063 430614
rect 41492 430478 45570 430538
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 44541 429722 44607 429725
rect 41492 429720 44607 429722
rect 41492 429664 44546 429720
rect 44602 429664 44607 429720
rect 41492 429662 44607 429664
rect 44541 429659 44607 429662
rect 44633 429314 44699 429317
rect 41492 429312 44699 429314
rect 41492 429256 44638 429312
rect 44694 429256 44699 429312
rect 41492 429254 44699 429256
rect 45510 429314 45570 430478
rect 61377 429314 61443 429317
rect 45510 429312 61443 429314
rect 45510 429256 61382 429312
rect 61438 429256 61443 429312
rect 45510 429254 61443 429256
rect 44633 429251 44699 429254
rect 61377 429251 61443 429254
rect 44265 428906 44331 428909
rect 41492 428904 44331 428906
rect 41492 428848 44270 428904
rect 44326 428848 44331 428904
rect 41492 428846 44331 428848
rect 44265 428843 44331 428846
rect 44265 428498 44331 428501
rect 41492 428496 44331 428498
rect 41492 428440 44270 428496
rect 44326 428440 44331 428496
rect 41492 428438 44331 428440
rect 44265 428435 44331 428438
rect 45645 428090 45711 428093
rect 41492 428088 45711 428090
rect 41492 428032 45650 428088
rect 45706 428032 45711 428088
rect 41492 428030 45711 428032
rect 45645 428027 45711 428030
rect 45645 427682 45711 427685
rect 41492 427680 45711 427682
rect 41492 427624 45650 427680
rect 45706 427624 45711 427680
rect 41492 427622 45711 427624
rect 45645 427619 45711 427622
rect 45829 427410 45895 427413
rect 41784 427408 45895 427410
rect 41784 427352 45834 427408
rect 45890 427352 45895 427408
rect 41784 427350 45895 427352
rect 41784 427274 41844 427350
rect 45829 427347 45895 427350
rect 41492 427214 41844 427274
rect 41965 427138 42031 427141
rect 63125 427138 63191 427141
rect 41965 427136 63191 427138
rect 41965 427080 41970 427136
rect 42026 427080 63130 427136
rect 63186 427080 63191 427136
rect 41965 427078 63191 427080
rect 41965 427075 42031 427078
rect 63125 427075 63191 427078
rect 45553 426866 45619 426869
rect 41492 426864 45619 426866
rect 41492 426808 45558 426864
rect 45614 426808 45619 426864
rect 41492 426806 45619 426808
rect 45553 426803 45619 426806
rect 41822 426458 41828 426460
rect 41492 426398 41828 426458
rect 41822 426396 41828 426398
rect 41892 426396 41898 426460
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 41137 425642 41203 425645
rect 41124 425640 41203 425642
rect 41124 425584 41142 425640
rect 41198 425584 41203 425640
rect 41124 425582 41203 425584
rect 41137 425579 41203 425582
rect 40953 425234 41019 425237
rect 40940 425232 41019 425234
rect 40940 425176 40958 425232
rect 41014 425176 41019 425232
rect 40940 425174 41019 425176
rect 40953 425171 41019 425174
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 32029 424418 32095 424421
rect 32029 424416 32108 424418
rect 32029 424360 32034 424416
rect 32090 424360 32108 424416
rect 32029 424358 32108 424360
rect 32029 424355 32095 424358
rect 41873 424282 41939 424285
rect 42190 424282 42196 424284
rect 41873 424280 42196 424282
rect 41873 424224 41878 424280
rect 41934 424224 42196 424280
rect 41873 424222 42196 424224
rect 41873 424219 41939 424222
rect 42190 424220 42196 424222
rect 42260 424220 42266 424284
rect 46013 424010 46079 424013
rect 41492 424008 46079 424010
rect 41492 423952 46018 424008
rect 46074 423952 46079 424008
rect 41492 423950 46079 423952
rect 46013 423947 46079 423950
rect 42793 423602 42859 423605
rect 41492 423600 42859 423602
rect 41492 423544 42798 423600
rect 42854 423544 42859 423600
rect 41492 423542 42859 423544
rect 42793 423539 42859 423542
rect 44909 423194 44975 423197
rect 41492 423192 44975 423194
rect 41492 423136 44914 423192
rect 44970 423136 44975 423192
rect 41492 423134 44975 423136
rect 44909 423131 44975 423134
rect 41822 422786 41828 422788
rect 41492 422726 41828 422786
rect 41822 422724 41828 422726
rect 41892 422724 41898 422788
rect 44449 422378 44515 422381
rect 41492 422376 44515 422378
rect 41492 422320 44454 422376
rect 44510 422320 44515 422376
rect 41492 422318 44515 422320
rect 44449 422315 44515 422318
rect 41822 421970 41828 421972
rect 41492 421910 41828 421970
rect 41822 421908 41828 421910
rect 41892 421908 41898 421972
rect 45093 421562 45159 421565
rect 41492 421560 45159 421562
rect 41492 421504 45098 421560
rect 45154 421504 45159 421560
rect 41492 421502 45159 421504
rect 45093 421499 45159 421502
rect 45277 421154 45343 421157
rect 41492 421152 45343 421154
rect 41492 421096 45282 421152
rect 45338 421096 45343 421152
rect 41492 421094 45343 421096
rect 45277 421091 45343 421094
rect 43253 420746 43319 420749
rect 41492 420744 43319 420746
rect 41492 420688 43258 420744
rect 43314 420688 43319 420744
rect 41492 420686 43319 420688
rect 43253 420683 43319 420686
rect 41462 419930 41522 420308
rect 42517 419930 42583 419933
rect 41462 419928 42583 419930
rect 41462 419900 42522 419928
rect 41492 419872 42522 419900
rect 42578 419872 42583 419928
rect 41492 419870 42583 419872
rect 42517 419867 42583 419870
rect 43069 419522 43135 419525
rect 41492 419520 43135 419522
rect 41492 419464 43074 419520
rect 43130 419464 43135 419520
rect 41492 419462 43135 419464
rect 43069 419459 43135 419462
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 41638 413340 41644 413404
rect 41708 413402 41714 413404
rect 42190 413402 42196 413404
rect 41708 413342 42196 413402
rect 41708 413340 41714 413342
rect 42190 413340 42196 413342
rect 42260 413340 42266 413404
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 675334 410484 675340 410548
rect 675404 410546 675410 410548
rect 676029 410546 676095 410549
rect 675404 410544 676095 410546
rect 675404 410488 676034 410544
rect 676090 410488 676095 410544
rect 675404 410486 676095 410488
rect 675404 410484 675410 410486
rect 676029 410483 676095 410486
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 41965 408098 42031 408101
rect 45277 408098 45343 408101
rect 41965 408096 45343 408098
rect 41965 408040 41970 408096
rect 42026 408040 45282 408096
rect 45338 408040 45343 408096
rect 41965 408038 45343 408040
rect 41965 408035 42031 408038
rect 45277 408035 45343 408038
rect 42425 407826 42491 407829
rect 53833 407826 53899 407829
rect 42425 407824 53899 407826
rect 42425 407768 42430 407824
rect 42486 407768 53838 407824
rect 53894 407768 53899 407824
rect 42425 407766 53899 407768
rect 42425 407763 42491 407766
rect 53833 407763 53899 407766
rect 42241 407554 42307 407557
rect 44449 407554 44515 407557
rect 42241 407552 44515 407554
rect 42241 407496 42246 407552
rect 42302 407496 44454 407552
rect 44510 407496 44515 407552
rect 42241 407494 44515 407496
rect 42241 407491 42307 407494
rect 44449 407491 44515 407494
rect 42057 406738 42123 406741
rect 45093 406738 45159 406741
rect 42057 406736 45159 406738
rect 42057 406680 42062 406736
rect 42118 406680 45098 406736
rect 45154 406680 45159 406736
rect 42057 406678 45159 406680
rect 42057 406675 42123 406678
rect 45093 406675 45159 406678
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 40902 405588 40908 405652
rect 40972 405650 40978 405652
rect 42241 405650 42307 405653
rect 40972 405648 42307 405650
rect 40972 405592 42246 405648
rect 42302 405592 42307 405648
rect 40972 405590 42307 405592
rect 40972 405588 40978 405590
rect 42241 405587 42307 405590
rect 42425 405650 42491 405653
rect 45277 405650 45343 405653
rect 42425 405648 45343 405650
rect 42425 405592 42430 405648
rect 42486 405592 45282 405648
rect 45338 405592 45343 405648
rect 42425 405590 45343 405592
rect 42425 405587 42491 405590
rect 45277 405587 45343 405590
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 657537 403338 657603 403341
rect 663750 403338 663810 403686
rect 676262 403341 676322 403444
rect 657537 403336 663810 403338
rect 657537 403280 657542 403336
rect 657598 403280 663810 403336
rect 657537 403278 663810 403280
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 657537 403275 657603 403278
rect 676213 403275 676279 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 44909 402930 44975 402933
rect 42333 402928 44975 402930
rect 42333 402872 42338 402928
rect 42394 402872 44914 402928
rect 44970 402872 44975 402928
rect 42333 402870 44975 402872
rect 42333 402867 42399 402870
rect 44909 402867 44975 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 676029 402658 676095 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 64646 402368 64706 402598
rect 676029 402656 676292 402658
rect 676029 402600 676034 402656
rect 676090 402600 676292 402656
rect 676029 402598 676292 402600
rect 676029 402595 676095 402598
rect 673177 402114 673243 402117
rect 676262 402114 676322 402220
rect 673177 402112 676322 402114
rect 673177 402056 673182 402112
rect 673238 402056 676322 402112
rect 673177 402054 676322 402056
rect 673177 402051 673243 402054
rect 41781 401844 41847 401845
rect 41781 401840 41828 401844
rect 41892 401842 41898 401844
rect 41781 401784 41786 401840
rect 41781 401780 41828 401784
rect 41892 401782 41938 401842
rect 41892 401780 41898 401782
rect 41781 401779 41847 401780
rect 672625 401706 672691 401709
rect 676262 401706 676322 401812
rect 672625 401704 676322 401706
rect 672625 401648 672630 401704
rect 672686 401648 676322 401704
rect 672625 401646 676322 401648
rect 672625 401643 672691 401646
rect 672901 401298 672967 401301
rect 676262 401298 676322 401404
rect 672901 401296 676322 401298
rect 672901 401240 672906 401296
rect 672962 401240 676322 401296
rect 672901 401238 676322 401240
rect 672901 401235 672967 401238
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400618 62179 400621
rect 64646 400618 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400616 64706 400618
rect 62113 400560 62118 400616
rect 62174 400560 64706 400616
rect 62113 400558 64706 400560
rect 673361 400618 673427 400621
rect 673361 400616 676292 400618
rect 673361 400560 673366 400616
rect 673422 400560 676292 400616
rect 673361 400558 676292 400560
rect 62113 400555 62179 400558
rect 673361 400555 673427 400558
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 42425 400210 42491 400213
rect 46013 400210 46079 400213
rect 42425 400208 46079 400210
rect 42425 400152 42430 400208
rect 42486 400152 46018 400208
rect 46074 400152 46079 400208
rect 42425 400150 46079 400152
rect 42425 400147 42491 400150
rect 46013 400147 46079 400150
rect 63125 400210 63191 400213
rect 63125 400208 64706 400210
rect 63125 400152 63130 400208
rect 63186 400152 64706 400208
rect 676814 400180 676874 400420
rect 63125 400150 64706 400152
rect 63125 400147 63191 400150
rect 40534 400012 40540 400076
rect 40604 400074 40610 400076
rect 41781 400074 41847 400077
rect 40604 400072 41847 400074
rect 40604 400016 41786 400072
rect 41842 400016 41847 400072
rect 40604 400014 41847 400016
rect 40604 400012 40610 400014
rect 41781 400011 41847 400014
rect 64646 400004 64706 400150
rect 673913 399802 673979 399805
rect 673913 399800 676292 399802
rect 673913 399744 673918 399800
rect 673974 399744 676292 399800
rect 673913 399742 676292 399744
rect 673913 399739 673979 399742
rect 62113 399394 62179 399397
rect 676029 399394 676095 399397
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 62113 399331 62179 399334
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 679574 398445 679634 398548
rect 679574 398440 679683 398445
rect 679574 398384 679622 398440
rect 679678 398384 679683 398440
rect 679574 398382 679683 398384
rect 679617 398379 679683 398382
rect 61377 398306 61443 398309
rect 61377 398304 64706 398306
rect 61377 398248 61382 398304
rect 61438 398248 64706 398304
rect 61377 398246 64706 398248
rect 61377 398243 61443 398246
rect 64646 397640 64706 398246
rect 676262 398037 676322 398140
rect 676213 398032 676322 398037
rect 676213 397976 676218 398032
rect 676274 397976 676322 398032
rect 676213 397974 676322 397976
rect 676213 397971 676279 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 671981 397218 672047 397221
rect 676262 397218 676322 397324
rect 671981 397216 676322 397218
rect 671981 397160 671986 397216
rect 672042 397160 676322 397216
rect 671981 397158 676322 397160
rect 671981 397155 672047 397158
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 676446 396404 676506 396508
rect 676438 396340 676444 396404
rect 676508 396340 676514 396404
rect 676029 396130 676095 396133
rect 676029 396128 676292 396130
rect 676029 396072 676034 396128
rect 676090 396072 676292 396128
rect 676029 396070 676292 396072
rect 676029 396067 676095 396070
rect 42149 395722 42215 395725
rect 51073 395722 51139 395725
rect 42149 395720 51139 395722
rect 42149 395664 42154 395720
rect 42210 395664 51078 395720
rect 51134 395664 51139 395720
rect 42149 395662 51139 395664
rect 42149 395659 42215 395662
rect 51073 395659 51139 395662
rect 676262 395589 676322 395692
rect 676213 395584 676322 395589
rect 676213 395528 676218 395584
rect 676274 395528 676322 395584
rect 676213 395526 676322 395528
rect 676213 395523 676279 395526
rect 652201 395314 652267 395317
rect 674557 395314 674623 395317
rect 652201 395312 674623 395314
rect 652201 395256 652206 395312
rect 652262 395256 674562 395312
rect 674618 395256 674623 395312
rect 652201 395254 674623 395256
rect 652201 395251 652267 395254
rect 674557 395251 674623 395254
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 672717 394770 672783 394773
rect 676262 394770 676322 394876
rect 672717 394768 676322 394770
rect 672717 394712 672722 394768
rect 672778 394712 676322 394768
rect 672717 394710 676322 394712
rect 672717 394707 672783 394710
rect 675201 394498 675267 394501
rect 675201 394496 676292 394498
rect 675201 394440 675206 394496
rect 675262 394440 676292 394496
rect 675201 394438 676292 394440
rect 675201 394435 675267 394438
rect 673729 394090 673795 394093
rect 673729 394088 676292 394090
rect 673729 394032 673734 394088
rect 673790 394032 676292 394088
rect 673729 394030 676292 394032
rect 673729 394027 673795 394030
rect 669221 393818 669287 393821
rect 669221 393816 676322 393818
rect 669221 393760 669226 393816
rect 669282 393760 676322 393816
rect 669221 393758 676322 393760
rect 669221 393755 669287 393758
rect 676262 393652 676322 393758
rect 674189 393138 674255 393141
rect 675201 393138 675267 393141
rect 674189 393136 675267 393138
rect 674189 393080 674194 393136
rect 674250 393080 675206 393136
rect 675262 393080 675267 393136
rect 674189 393078 675267 393080
rect 674189 393075 674255 393078
rect 675201 393075 675267 393078
rect 675886 392804 675892 392868
rect 675956 392866 675962 392868
rect 676262 392866 676322 393244
rect 675956 392836 676322 392866
rect 675956 392806 676292 392836
rect 675956 392804 675962 392806
rect 670601 392594 670667 392597
rect 670601 392592 676322 392594
rect 670601 392536 670606 392592
rect 670662 392536 676322 392592
rect 670601 392534 676322 392536
rect 670601 392531 670667 392534
rect 676262 392428 676322 392534
rect 675702 388452 675708 388516
rect 675772 388514 675778 388516
rect 680997 388514 681063 388517
rect 675772 388512 681063 388514
rect 675772 388456 681002 388512
rect 681058 388456 681063 388512
rect 675772 388454 681063 388456
rect 675772 388452 675778 388454
rect 680997 388451 681063 388454
rect 41462 387562 41522 387668
rect 41462 387502 51090 387562
rect 41094 387157 41154 387260
rect 41094 387152 41203 387157
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387094 41203 387096
rect 41137 387091 41203 387094
rect 41278 386749 41338 386852
rect 41278 386744 41387 386749
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386686 41387 386688
rect 41321 386683 41387 386686
rect 44633 386474 44699 386477
rect 41492 386472 44699 386474
rect 41492 386416 44638 386472
rect 44694 386416 44699 386472
rect 41492 386414 44699 386416
rect 51030 386474 51090 387502
rect 61377 386474 61443 386477
rect 51030 386472 61443 386474
rect 51030 386416 61382 386472
rect 61438 386416 61443 386472
rect 51030 386414 61443 386416
rect 44633 386411 44699 386414
rect 61377 386411 61443 386414
rect 40726 385933 40786 386036
rect 40726 385928 40835 385933
rect 40726 385872 40774 385928
rect 40830 385872 40835 385928
rect 40726 385870 40835 385872
rect 40769 385867 40835 385870
rect 41321 385930 41387 385933
rect 63401 385930 63467 385933
rect 41321 385928 63467 385930
rect 41321 385872 41326 385928
rect 41382 385872 63406 385928
rect 63462 385872 63467 385928
rect 41321 385870 63467 385872
rect 41321 385867 41387 385870
rect 63401 385867 63467 385870
rect 44265 385658 44331 385661
rect 41492 385656 44331 385658
rect 41492 385600 44270 385656
rect 44326 385600 44331 385656
rect 41492 385598 44331 385600
rect 44265 385595 44331 385598
rect 675753 385386 675819 385389
rect 676622 385386 676628 385388
rect 675753 385384 676628 385386
rect 675753 385328 675758 385384
rect 675814 385328 676628 385384
rect 675753 385326 676628 385328
rect 675753 385323 675819 385326
rect 676622 385324 676628 385326
rect 676692 385324 676698 385388
rect 45093 385250 45159 385253
rect 41492 385248 45159 385250
rect 41492 385192 45098 385248
rect 45154 385192 45159 385248
rect 41492 385190 45159 385192
rect 45093 385187 45159 385190
rect 45829 384842 45895 384845
rect 41492 384840 45895 384842
rect 41492 384784 45834 384840
rect 45890 384784 45895 384840
rect 41492 384782 45895 384784
rect 45829 384779 45895 384782
rect 46013 384434 46079 384437
rect 41492 384432 46079 384434
rect 41492 384376 46018 384432
rect 46074 384376 46079 384432
rect 41492 384374 46079 384376
rect 46013 384371 46079 384374
rect 45553 384026 45619 384029
rect 41492 384024 45619 384026
rect 41492 383968 45558 384024
rect 45614 383968 45619 384024
rect 41492 383966 45619 383968
rect 45553 383963 45619 383966
rect 45645 383618 45711 383621
rect 41492 383616 45711 383618
rect 41492 383560 45650 383616
rect 45706 383560 45711 383616
rect 41492 383558 45711 383560
rect 45645 383555 45711 383558
rect 47117 383210 47183 383213
rect 41492 383208 47183 383210
rect 41492 383152 47122 383208
rect 47178 383152 47183 383208
rect 41492 383150 47183 383152
rect 47117 383147 47183 383150
rect 654777 382938 654843 382941
rect 675293 382938 675359 382941
rect 654777 382936 675359 382938
rect 654777 382880 654782 382936
rect 654838 382880 675298 382936
rect 675354 382880 675359 382936
rect 654777 382878 675359 382880
rect 654777 382875 654843 382878
rect 675293 382875 675359 382878
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 46933 382394 46999 382397
rect 41492 382392 46999 382394
rect 41492 382336 46938 382392
rect 46994 382336 46999 382392
rect 41492 382334 46999 382336
rect 46933 382331 46999 382334
rect 675753 382258 675819 382261
rect 676438 382258 676444 382260
rect 675753 382256 676444 382258
rect 675753 382200 675758 382256
rect 675814 382200 676444 382256
rect 675753 382198 676444 382200
rect 675753 382195 675819 382198
rect 676438 382196 676444 382198
rect 676508 382196 676514 382260
rect 40910 381853 40970 381956
rect 40910 381848 41019 381853
rect 40910 381792 40958 381848
rect 41014 381792 41019 381848
rect 40910 381790 41019 381792
rect 40953 381787 41019 381790
rect 41137 381850 41203 381853
rect 62941 381850 63007 381853
rect 41137 381848 63007 381850
rect 41137 381792 41142 381848
rect 41198 381792 62946 381848
rect 63002 381792 63007 381848
rect 41137 381790 63007 381792
rect 41137 381787 41203 381790
rect 62941 381787 63007 381790
rect 40174 381445 40234 381548
rect 40174 381440 40283 381445
rect 40174 381384 40222 381440
rect 40278 381384 40283 381440
rect 40174 381382 40283 381384
rect 40217 381379 40283 381382
rect 40769 381442 40835 381445
rect 45277 381442 45343 381445
rect 40769 381440 45343 381442
rect 40769 381384 40774 381440
rect 40830 381384 45282 381440
rect 45338 381384 45343 381440
rect 40769 381382 45343 381384
rect 40769 381379 40835 381382
rect 45277 381379 45343 381382
rect 35206 381037 35266 381140
rect 35157 381032 35266 381037
rect 35157 380976 35162 381032
rect 35218 380976 35266 381032
rect 35157 380974 35266 380976
rect 672717 381034 672783 381037
rect 675385 381034 675451 381037
rect 672717 381032 675451 381034
rect 672717 380976 672722 381032
rect 672778 380976 675390 381032
rect 675446 380976 675451 381032
rect 672717 380974 675451 380976
rect 35157 380971 35223 380974
rect 672717 380971 672783 380974
rect 675385 380971 675451 380974
rect 40542 380628 40602 380732
rect 40534 380564 40540 380628
rect 40604 380564 40610 380628
rect 37966 380221 38026 380324
rect 37917 380216 38026 380221
rect 37917 380160 37922 380216
rect 37978 380160 38026 380216
rect 37917 380158 38026 380160
rect 37917 380155 37983 380158
rect 33734 379813 33794 379916
rect 33734 379808 33843 379813
rect 41505 379812 41571 379813
rect 33734 379752 33782 379808
rect 33838 379752 33843 379808
rect 33734 379750 33843 379752
rect 33777 379747 33843 379750
rect 41454 379748 41460 379812
rect 41524 379810 41571 379812
rect 41524 379808 41616 379810
rect 41566 379752 41616 379808
rect 41524 379750 41616 379752
rect 41524 379748 41571 379750
rect 41505 379747 41571 379748
rect 42885 379538 42951 379541
rect 41492 379536 42951 379538
rect 41492 379480 42890 379536
rect 42946 379480 42951 379536
rect 41492 379478 42951 379480
rect 42885 379475 42951 379478
rect 44357 379130 44423 379133
rect 41492 379128 44423 379130
rect 41492 379072 44362 379128
rect 44418 379072 44423 379128
rect 41492 379070 44423 379072
rect 44357 379067 44423 379070
rect 44541 378722 44607 378725
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 41492 378720 44607 378722
rect 41492 378664 44546 378720
rect 44602 378664 44607 378720
rect 41492 378662 44607 378664
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 44541 378659 44607 378662
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 44725 377906 44791 377909
rect 41492 377904 44791 377906
rect 41492 377848 44730 377904
rect 44786 377848 44791 377904
rect 41492 377846 44791 377848
rect 44725 377843 44791 377846
rect 44909 377498 44975 377501
rect 41492 377496 44975 377498
rect 41492 377440 44914 377496
rect 44970 377440 44975 377496
rect 41492 377438 44975 377440
rect 44909 377435 44975 377438
rect 675753 377498 675819 377501
rect 676254 377498 676260 377500
rect 675753 377496 676260 377498
rect 675753 377440 675758 377496
rect 675814 377440 676260 377496
rect 675753 377438 676260 377440
rect 675753 377435 675819 377438
rect 676254 377436 676260 377438
rect 676324 377436 676330 377500
rect 35758 376549 35818 377060
rect 673729 376682 673795 376685
rect 675109 376682 675175 376685
rect 673729 376680 675175 376682
rect 673729 376624 673734 376680
rect 673790 376624 675114 376680
rect 675170 376624 675175 376680
rect 673729 376622 675175 376624
rect 673729 376619 673795 376622
rect 675109 376619 675175 376622
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 44173 376274 44239 376277
rect 41492 376272 44239 376274
rect 41492 376216 44178 376272
rect 44234 376216 44239 376272
rect 41492 376214 44239 376216
rect 44173 376211 44239 376214
rect 35801 374642 35867 374645
rect 41270 374642 41276 374644
rect 35801 374640 41276 374642
rect 35801 374584 35806 374640
rect 35862 374584 41276 374640
rect 35801 374582 41276 374584
rect 35801 374579 35867 374582
rect 41270 374580 41276 374582
rect 41340 374580 41346 374644
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 37917 372738 37983 372741
rect 41638 372738 41644 372740
rect 37917 372736 41644 372738
rect 37917 372680 37922 372736
rect 37978 372680 41644 372736
rect 37917 372678 41644 372680
rect 37917 372675 37983 372678
rect 41638 372676 41644 372678
rect 41708 372676 41714 372740
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675661 373010 675727 373013
rect 675886 373010 675892 373012
rect 675661 373008 675892 373010
rect 675661 372952 675666 373008
rect 675722 372952 675892 373008
rect 675661 372950 675892 372952
rect 675661 372947 675727 372950
rect 675886 372948 675892 372950
rect 675956 372948 675962 373012
rect 671981 372602 672047 372605
rect 675109 372602 675175 372605
rect 671981 372600 675175 372602
rect 671981 372544 671986 372600
rect 672042 372544 675114 372600
rect 675170 372544 675175 372600
rect 671981 372542 675175 372544
rect 671981 372539 672047 372542
rect 675109 372539 675175 372542
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 33777 371922 33843 371925
rect 41822 371922 41828 371924
rect 33777 371920 41828 371922
rect 33777 371864 33782 371920
rect 33838 371864 41828 371920
rect 33777 371862 41828 371864
rect 33777 371859 33843 371862
rect 41822 371860 41828 371862
rect 41892 371860 41898 371924
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 41270 368460 41276 368524
rect 41340 368522 41346 368524
rect 41781 368522 41847 368525
rect 41340 368520 41847 368522
rect 41340 368464 41786 368520
rect 41842 368464 41847 368520
rect 41340 368462 41847 368464
rect 41340 368460 41346 368462
rect 41781 368459 41847 368462
rect 42057 366210 42123 366213
rect 42885 366210 42951 366213
rect 42057 366208 42951 366210
rect 42057 366152 42062 366208
rect 42118 366152 42890 366208
rect 42946 366152 42951 366208
rect 42057 366150 42951 366152
rect 42057 366147 42123 366150
rect 42885 366147 42951 366150
rect 42057 364850 42123 364853
rect 44725 364850 44791 364853
rect 42057 364848 44791 364850
rect 42057 364792 42062 364848
rect 42118 364792 44730 364848
rect 44786 364792 44791 364848
rect 42057 364790 44791 364792
rect 42057 364787 42123 364790
rect 44725 364787 44791 364790
rect 42241 364170 42307 364173
rect 44357 364170 44423 364173
rect 42241 364168 44423 364170
rect 42241 364112 42246 364168
rect 42302 364112 44362 364168
rect 44418 364112 44423 364168
rect 42241 364110 44423 364112
rect 42241 364107 42307 364110
rect 44357 364107 44423 364110
rect 40718 363700 40724 363764
rect 40788 363762 40794 363764
rect 41781 363762 41847 363765
rect 40788 363760 41847 363762
rect 40788 363704 41786 363760
rect 41842 363704 41847 363760
rect 40788 363702 41847 363704
rect 40788 363700 40794 363702
rect 41781 363699 41847 363702
rect 42701 363218 42767 363221
rect 46565 363218 46631 363221
rect 42701 363216 46631 363218
rect 42701 363160 42706 363216
rect 42762 363160 46570 363216
rect 46626 363160 46631 363216
rect 42701 363158 46631 363160
rect 42701 363155 42767 363158
rect 46565 363155 46631 363158
rect 42241 362946 42307 362949
rect 45369 362946 45435 362949
rect 42241 362944 45435 362946
rect 42241 362888 42246 362944
rect 42302 362888 45374 362944
rect 45430 362888 45435 362944
rect 42241 362886 45435 362888
rect 42241 362883 42307 362886
rect 45369 362883 45435 362886
rect 42425 361586 42491 361589
rect 44541 361586 44607 361589
rect 42425 361584 44607 361586
rect 42425 361528 42430 361584
rect 42486 361528 44546 361584
rect 44602 361528 44607 361584
rect 42425 361526 44607 361528
rect 42425 361523 42491 361526
rect 44541 361523 44607 361526
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 41781 360092 41847 360093
rect 41781 360088 41828 360092
rect 41892 360090 41898 360092
rect 41781 360032 41786 360088
rect 41781 360028 41828 360032
rect 41892 360030 41938 360090
rect 41892 360028 41898 360030
rect 41781 360027 41847 360028
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 41638 359484 41644 359548
rect 41708 359546 41714 359548
rect 41708 359486 41890 359546
rect 41708 359484 41714 359486
rect 41830 359277 41890 359486
rect 41781 359272 41890 359277
rect 41781 359216 41786 359272
rect 41842 359216 41890 359272
rect 41781 359214 41890 359216
rect 41781 359211 41847 359214
rect 64646 359146 64706 359758
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 663750 358670 676292 358730
rect 654777 358594 654843 358597
rect 663750 358594 663810 358670
rect 654777 358592 663810 358594
rect 654777 358536 654782 358592
rect 654838 358536 663810 358592
rect 654777 358534 663810 358536
rect 654777 358531 654843 358534
rect 675569 358322 675635 358325
rect 675569 358320 676292 358322
rect 675569 358264 675574 358320
rect 675630 358264 676292 358320
rect 675569 358262 676292 358264
rect 675569 358259 675635 358262
rect 62113 357778 62179 357781
rect 64646 357778 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62113 357776 64706 357778
rect 62113 357720 62118 357776
rect 62174 357720 64706 357776
rect 62113 357718 64706 357720
rect 62113 357715 62179 357718
rect 673177 357506 673243 357509
rect 673177 357504 676292 357506
rect 673177 357448 673182 357504
rect 673238 357448 676292 357504
rect 673177 357446 676292 357448
rect 673177 357443 673243 357446
rect 63401 357370 63467 357373
rect 63401 357368 64706 357370
rect 63401 357312 63406 357368
rect 63462 357312 64706 357368
rect 63401 357310 64706 357312
rect 63401 357307 63467 357310
rect 64646 356782 64706 357310
rect 672533 357098 672599 357101
rect 672533 357096 676292 357098
rect 672533 357040 672538 357096
rect 672594 357040 676292 357096
rect 672533 357038 676292 357040
rect 672533 357035 672599 357038
rect 672901 356826 672967 356829
rect 672901 356824 676230 356826
rect 672901 356768 672906 356824
rect 672962 356768 676230 356824
rect 672901 356766 676230 356768
rect 672901 356763 672967 356766
rect 652017 356690 652083 356693
rect 676170 356690 676230 356766
rect 652017 356688 663810 356690
rect 652017 356632 652022 356688
rect 652078 356632 663810 356688
rect 652017 356630 663810 356632
rect 676170 356630 676292 356690
rect 652017 356627 652083 356630
rect 663750 356554 663810 356630
rect 675937 356554 676003 356557
rect 663750 356552 676003 356554
rect 663750 356496 675942 356552
rect 675998 356496 676003 356552
rect 663750 356494 676003 356496
rect 675937 356491 676003 356494
rect 672717 356282 672783 356285
rect 672717 356280 676292 356282
rect 672717 356224 672722 356280
rect 672778 356224 676292 356280
rect 672717 356222 676292 356224
rect 672717 356219 672783 356222
rect 40534 356084 40540 356148
rect 40604 356146 40610 356148
rect 41781 356146 41847 356149
rect 40604 356144 41847 356146
rect 40604 356088 41786 356144
rect 41842 356088 41847 356144
rect 40604 356086 41847 356088
rect 40604 356084 40610 356086
rect 41781 356083 41847 356086
rect 61377 356010 61443 356013
rect 61377 356008 64706 356010
rect 61377 355952 61382 356008
rect 61438 355952 64706 356008
rect 61377 355950 64706 355952
rect 61377 355947 61443 355950
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 673177 355466 673243 355469
rect 673177 355464 676292 355466
rect 673177 355408 673182 355464
rect 673238 355408 676292 355464
rect 673177 355406 676292 355408
rect 673177 355403 673243 355406
rect 43805 355194 43871 355197
rect 44817 355194 44883 355197
rect 43805 355192 44883 355194
rect 43805 355136 43810 355192
rect 43866 355136 44822 355192
rect 44878 355136 44883 355192
rect 43805 355134 44883 355136
rect 43805 355131 43871 355134
rect 44817 355131 44883 355134
rect 673913 355058 673979 355061
rect 673913 355056 676292 355058
rect 673913 355000 673918 355056
rect 673974 355000 676292 355056
rect 673913 354998 676292 355000
rect 673913 354995 673979 354998
rect 43621 354922 43687 354925
rect 44633 354922 44699 354925
rect 43621 354920 44699 354922
rect 43621 354864 43626 354920
rect 43682 354864 44638 354920
rect 44694 354864 44699 354920
rect 43621 354862 44699 354864
rect 43621 354859 43687 354862
rect 44633 354859 44699 354862
rect 674097 354650 674163 354653
rect 674097 354648 676292 354650
rect 674097 354592 674102 354648
rect 674158 354592 676292 354648
rect 674097 354590 676292 354592
rect 674097 354587 674163 354590
rect 62941 354514 63007 354517
rect 62941 354512 64706 354514
rect 62941 354456 62946 354512
rect 63002 354456 64706 354512
rect 62941 354454 64706 354456
rect 62941 354451 63007 354454
rect 64646 354418 64706 354454
rect 42425 354378 42491 354381
rect 47117 354378 47183 354381
rect 42425 354376 47183 354378
rect 42425 354320 42430 354376
rect 42486 354320 47122 354376
rect 47178 354320 47183 354376
rect 42425 354318 47183 354320
rect 42425 354315 42491 354318
rect 47117 354315 47183 354318
rect 674741 354242 674807 354245
rect 674741 354240 676292 354242
rect 674741 354184 674746 354240
rect 674802 354184 676292 354240
rect 674741 354182 676292 354184
rect 674741 354179 674807 354182
rect 43069 353970 43135 353973
rect 45829 353970 45895 353973
rect 43069 353968 45895 353970
rect 43069 353912 43074 353968
rect 43130 353912 45834 353968
rect 45890 353912 45895 353968
rect 43069 353910 45895 353912
rect 43069 353907 43135 353910
rect 45829 353907 45895 353910
rect 675845 353834 675911 353837
rect 675845 353832 676292 353834
rect 675845 353776 675850 353832
rect 675906 353776 676292 353832
rect 675845 353774 676292 353776
rect 675845 353771 675911 353774
rect 43253 353698 43319 353701
rect 45829 353698 45895 353701
rect 43253 353696 45895 353698
rect 43253 353640 43258 353696
rect 43314 353640 45834 353696
rect 45890 353640 45895 353696
rect 43253 353638 45895 353640
rect 43253 353635 43319 353638
rect 45829 353635 45895 353638
rect 675518 353364 675524 353428
rect 675588 353426 675594 353428
rect 675588 353366 676292 353426
rect 675588 353364 675594 353366
rect 42149 353290 42215 353293
rect 51717 353290 51783 353293
rect 42149 353288 51783 353290
rect 42149 353232 42154 353288
rect 42210 353232 51722 353288
rect 51778 353232 51783 353288
rect 42149 353230 51783 353232
rect 42149 353227 42215 353230
rect 51717 353227 51783 353230
rect 42333 353018 42399 353021
rect 46933 353018 46999 353021
rect 42333 353016 46999 353018
rect 42333 352960 42338 353016
rect 42394 352960 46938 353016
rect 46994 352960 46999 353016
rect 42333 352958 46999 352960
rect 42333 352955 42399 352958
rect 46933 352955 46999 352958
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 675569 352882 675635 352885
rect 669270 352880 675635 352882
rect 669270 352824 675574 352880
rect 675630 352824 675635 352880
rect 669270 352822 675635 352824
rect 652385 352610 652451 352613
rect 669270 352610 669330 352822
rect 675569 352819 675635 352822
rect 652385 352608 669330 352610
rect 652385 352552 652390 352608
rect 652446 352552 669330 352608
rect 652385 352550 669330 352552
rect 673729 352610 673795 352613
rect 673729 352608 676292 352610
rect 673729 352552 673734 352608
rect 673790 352552 676292 352608
rect 673729 352550 676292 352552
rect 652385 352547 652451 352550
rect 673729 352547 673795 352550
rect 675932 352140 675938 352204
rect 676002 352202 676008 352204
rect 676002 352142 676292 352202
rect 676002 352140 676008 352142
rect 675845 351932 675911 351933
rect 675845 351930 675892 351932
rect 675800 351928 675892 351930
rect 675800 351872 675850 351928
rect 675800 351870 675892 351872
rect 675845 351868 675892 351870
rect 675956 351868 675962 351932
rect 675845 351867 675911 351868
rect 676029 351794 676095 351797
rect 676029 351792 676292 351794
rect 676029 351736 676034 351792
rect 676090 351736 676292 351792
rect 676029 351734 676292 351736
rect 676029 351731 676095 351734
rect 672349 351386 672415 351389
rect 672349 351384 676292 351386
rect 672349 351328 672354 351384
rect 672410 351328 676292 351384
rect 672349 351326 676292 351328
rect 672349 351323 672415 351326
rect 674281 350978 674347 350981
rect 674281 350976 676292 350978
rect 674281 350920 674286 350976
rect 674342 350920 676292 350976
rect 674281 350918 676292 350920
rect 674281 350915 674347 350918
rect 674557 350570 674623 350573
rect 674557 350568 676292 350570
rect 674557 350512 674562 350568
rect 674618 350512 676292 350568
rect 674557 350510 676292 350512
rect 674557 350507 674623 350510
rect 671981 350162 672047 350165
rect 671981 350160 676292 350162
rect 671981 350104 671986 350160
rect 672042 350104 676292 350160
rect 671981 350102 676292 350104
rect 671981 350099 672047 350102
rect 673361 349754 673427 349757
rect 673361 349752 676292 349754
rect 673361 349696 673366 349752
rect 673422 349696 676292 349752
rect 673361 349694 676292 349696
rect 673361 349691 673427 349694
rect 673545 349346 673611 349349
rect 673545 349344 676292 349346
rect 673545 349288 673550 349344
rect 673606 349288 676292 349344
rect 673545 349286 676292 349288
rect 673545 349283 673611 349286
rect 673913 348938 673979 348941
rect 673913 348936 676292 348938
rect 673913 348880 673918 348936
rect 673974 348880 676292 348936
rect 673913 348878 676292 348880
rect 673913 348875 673979 348878
rect 672901 348530 672967 348533
rect 672901 348528 676292 348530
rect 672901 348472 672906 348528
rect 672962 348472 676292 348528
rect 672901 348470 676292 348472
rect 672901 348467 672967 348470
rect 683070 347717 683130 348092
rect 683070 347712 683179 347717
rect 683070 347684 683118 347712
rect 683100 347656 683118 347684
rect 683174 347656 683179 347712
rect 683100 347654 683179 347656
rect 683113 347651 683179 347654
rect 676029 347306 676095 347309
rect 676029 347304 676292 347306
rect 676029 347248 676034 347304
rect 676090 347248 676292 347304
rect 676029 347246 676292 347248
rect 676029 347243 676095 347246
rect 658917 346490 658983 346493
rect 676262 346490 676322 346868
rect 676489 346628 676555 346629
rect 676438 346564 676444 346628
rect 676508 346626 676555 346628
rect 676508 346624 676600 346626
rect 676550 346568 676600 346624
rect 676508 346566 676600 346568
rect 676508 346564 676555 346566
rect 676489 346563 676555 346564
rect 683113 346490 683179 346493
rect 658917 346488 676322 346490
rect 658917 346432 658922 346488
rect 658978 346432 676322 346488
rect 658917 346430 676322 346432
rect 676814 346488 683179 346490
rect 676814 346432 683118 346488
rect 683174 346432 683179 346488
rect 676814 346430 683179 346432
rect 658917 346427 658983 346430
rect 676814 346220 676874 346430
rect 683113 346427 683179 346430
rect 676806 346156 676812 346220
rect 676876 346156 676882 346220
rect 669957 345674 670023 345677
rect 676029 345674 676095 345677
rect 669957 345672 676095 345674
rect 669957 345616 669962 345672
rect 670018 345616 676034 345672
rect 676090 345616 676095 345672
rect 669957 345614 676095 345616
rect 669957 345611 670023 345614
rect 676029 345611 676095 345614
rect 35758 344317 35818 344556
rect 35758 344312 35867 344317
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344254 35867 344256
rect 35801 344251 35867 344254
rect 35574 343909 35634 344148
rect 35574 343904 35683 343909
rect 35574 343848 35622 343904
rect 35678 343848 35683 343904
rect 35574 343846 35683 343848
rect 35617 343843 35683 343846
rect 40401 343906 40467 343909
rect 46013 343906 46079 343909
rect 40401 343904 46079 343906
rect 40401 343848 40406 343904
rect 40462 343848 46018 343904
rect 46074 343848 46079 343904
rect 40401 343846 46079 343848
rect 40401 343843 40467 343846
rect 46013 343843 46079 343846
rect 35758 343501 35818 343740
rect 35758 343496 35867 343501
rect 35758 343440 35806 343496
rect 35862 343440 35867 343496
rect 35758 343438 35867 343440
rect 35801 343435 35867 343438
rect 45185 343362 45251 343365
rect 41492 343360 45251 343362
rect 41492 343304 45190 343360
rect 45246 343304 45251 343360
rect 41492 343302 45251 343304
rect 45185 343299 45251 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 45001 342546 45067 342549
rect 41492 342544 45067 342546
rect 41492 342488 45006 342544
rect 45062 342488 45067 342544
rect 41492 342486 45067 342488
rect 45001 342483 45067 342486
rect 40217 342274 40283 342277
rect 45461 342274 45527 342277
rect 40217 342272 45527 342274
rect 40217 342216 40222 342272
rect 40278 342216 45466 342272
rect 45522 342216 45527 342272
rect 40217 342214 45527 342216
rect 40217 342211 40283 342214
rect 45461 342211 45527 342214
rect 39622 341869 39682 342108
rect 35801 341866 35867 341869
rect 35758 341864 35867 341866
rect 35758 341808 35806 341864
rect 35862 341808 35867 341864
rect 35758 341803 35867 341808
rect 39622 341864 39731 341869
rect 39622 341808 39670 341864
rect 39726 341808 39731 341864
rect 39622 341806 39731 341808
rect 39665 341803 39731 341806
rect 39849 341866 39915 341869
rect 39849 341864 45570 341866
rect 39849 341808 39854 341864
rect 39910 341808 45570 341864
rect 39849 341806 45570 341808
rect 39849 341803 39915 341806
rect 35758 341700 35818 341803
rect 45510 341730 45570 341806
rect 62941 341730 63007 341733
rect 45510 341728 63007 341730
rect 45510 341672 62946 341728
rect 63002 341672 63007 341728
rect 45510 341670 63007 341672
rect 62941 341667 63007 341670
rect 44214 341594 44220 341596
rect 42014 341534 44220 341594
rect 42014 341322 42074 341534
rect 44214 341532 44220 341534
rect 44284 341532 44290 341596
rect 62757 341458 62823 341461
rect 45510 341456 62823 341458
rect 45510 341400 62762 341456
rect 62818 341400 62823 341456
rect 45510 341398 62823 341400
rect 41492 341262 42074 341322
rect 42241 341322 42307 341325
rect 45510 341322 45570 341398
rect 62757 341395 62823 341398
rect 42241 341320 45570 341322
rect 42241 341264 42246 341320
rect 42302 341264 45570 341320
rect 42241 341262 45570 341264
rect 42241 341259 42307 341262
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 40125 341050 40191 341053
rect 40125 341048 40418 341050
rect 40125 340992 40130 341048
rect 40186 340992 40418 341048
rect 40125 340990 40418 340992
rect 40125 340987 40191 340990
rect 35758 340884 35818 340987
rect 40358 340778 40418 340990
rect 45645 340778 45711 340781
rect 675569 340780 675635 340781
rect 675518 340778 675524 340780
rect 40358 340776 45711 340778
rect 40358 340720 45650 340776
rect 45706 340720 45711 340776
rect 40358 340718 45711 340720
rect 675478 340718 675524 340778
rect 675588 340776 675635 340780
rect 675630 340720 675635 340776
rect 45645 340715 45711 340718
rect 675518 340716 675524 340718
rect 675588 340716 675635 340720
rect 675569 340715 675635 340716
rect 42742 340506 42748 340508
rect 41492 340446 42748 340506
rect 42742 340444 42748 340446
rect 42812 340444 42818 340508
rect 39665 340234 39731 340237
rect 44582 340234 44588 340236
rect 39665 340232 44588 340234
rect 39665 340176 39670 340232
rect 39726 340176 44588 340232
rect 39665 340174 44588 340176
rect 39665 340171 39731 340174
rect 44582 340172 44588 340174
rect 44652 340172 44658 340236
rect 675753 340234 675819 340237
rect 676438 340234 676444 340236
rect 675753 340232 676444 340234
rect 675753 340176 675758 340232
rect 675814 340176 676444 340232
rect 675753 340174 676444 340176
rect 675753 340171 675819 340174
rect 676438 340172 676444 340174
rect 676508 340172 676514 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 46933 339282 46999 339285
rect 41492 339280 46999 339282
rect 41492 339224 46938 339280
rect 46994 339224 46999 339280
rect 41492 339222 46999 339224
rect 46933 339219 46999 339222
rect 45553 338874 45619 338877
rect 41492 338872 45619 338874
rect 41492 338816 45558 338872
rect 45614 338816 45619 338872
rect 41492 338814 45619 338816
rect 45553 338811 45619 338814
rect 653397 338738 653463 338741
rect 675109 338738 675175 338741
rect 653397 338736 675175 338738
rect 653397 338680 653402 338736
rect 653458 338680 675114 338736
rect 675170 338680 675175 338736
rect 653397 338678 675175 338680
rect 653397 338675 653463 338678
rect 675109 338675 675175 338678
rect 41462 338194 41522 338436
rect 41638 338194 41644 338196
rect 41462 338134 41644 338194
rect 41638 338132 41644 338134
rect 41708 338132 41714 338196
rect 41278 337922 41338 338028
rect 45369 337922 45435 337925
rect 41278 337920 45435 337922
rect 41278 337864 45374 337920
rect 45430 337864 45435 337920
rect 41278 337862 45435 337864
rect 45369 337859 45435 337862
rect 675661 337786 675727 337789
rect 675886 337786 675892 337788
rect 675661 337784 675892 337786
rect 675661 337728 675666 337784
rect 675722 337728 675892 337784
rect 675661 337726 675892 337728
rect 675661 337723 675727 337726
rect 675886 337724 675892 337726
rect 675956 337724 675962 337788
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 43110 337242 43116 337244
rect 41492 337182 43116 337242
rect 43110 337180 43116 337182
rect 43180 337180 43186 337244
rect 672349 337242 672415 337245
rect 675109 337242 675175 337245
rect 672349 337240 675175 337242
rect 672349 337184 672354 337240
rect 672410 337184 675114 337240
rect 675170 337184 675175 337240
rect 672349 337182 675175 337184
rect 672349 337179 672415 337182
rect 675109 337179 675175 337182
rect 40718 336908 40724 336972
rect 40788 336908 40794 336972
rect 40726 336804 40786 336908
rect 37089 336562 37155 336565
rect 42006 336562 42012 336564
rect 37089 336560 42012 336562
rect 37089 336504 37094 336560
rect 37150 336504 42012 336560
rect 37089 336502 42012 336504
rect 37089 336499 37155 336502
rect 42006 336500 42012 336502
rect 42076 336500 42082 336564
rect 41462 336154 41522 336396
rect 41462 336094 44466 336154
rect 35758 335749 35818 335988
rect 35758 335744 35867 335749
rect 35758 335688 35806 335744
rect 35862 335688 35867 335744
rect 35758 335686 35867 335688
rect 35801 335683 35867 335686
rect 38837 335746 38903 335749
rect 41822 335746 41828 335748
rect 38837 335744 41828 335746
rect 38837 335688 38842 335744
rect 38898 335688 41828 335744
rect 38837 335686 41828 335688
rect 38837 335683 38903 335686
rect 41822 335684 41828 335686
rect 41892 335684 41898 335748
rect 40542 335340 40602 335580
rect 40534 335276 40540 335340
rect 40604 335276 40610 335340
rect 41462 334930 41522 335172
rect 41462 334870 41890 334930
rect 35758 334525 35818 334764
rect 41830 334658 41890 334870
rect 44406 334661 44466 336094
rect 673361 335610 673427 335613
rect 675109 335610 675175 335613
rect 673361 335608 675175 335610
rect 673361 335552 673366 335608
rect 673422 335552 675114 335608
rect 675170 335552 675175 335608
rect 673361 335550 675175 335552
rect 673361 335547 673427 335550
rect 675109 335547 675175 335550
rect 44173 334658 44239 334661
rect 41830 334656 44239 334658
rect 41830 334600 44178 334656
rect 44234 334600 44239 334656
rect 41830 334598 44239 334600
rect 44173 334595 44239 334598
rect 44357 334656 44466 334661
rect 44357 334600 44362 334656
rect 44418 334600 44466 334656
rect 44357 334598 44466 334600
rect 44357 334595 44423 334598
rect 35758 334520 35867 334525
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334462 35867 334464
rect 35801 334459 35867 334462
rect 41462 334114 41522 334356
rect 51717 334114 51783 334117
rect 41462 334112 51783 334114
rect 41462 334056 51722 334112
rect 51778 334056 51783 334112
rect 41462 334054 51783 334056
rect 51717 334051 51783 334054
rect 673729 333978 673795 333981
rect 675109 333978 675175 333981
rect 673729 333976 675175 333978
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 673729 333920 673734 333976
rect 673790 333920 675114 333976
rect 675170 333920 675175 333976
rect 673729 333918 675175 333920
rect 673729 333915 673795 333918
rect 675109 333915 675175 333918
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 50337 333162 50403 333165
rect 41492 333160 50403 333162
rect 41492 333104 50342 333160
rect 50398 333104 50403 333160
rect 41492 333102 50403 333104
rect 50337 333099 50403 333102
rect 40309 332890 40375 332893
rect 42885 332890 42951 332893
rect 40309 332888 42951 332890
rect 40309 332832 40314 332888
rect 40370 332832 42890 332888
rect 42946 332832 42951 332888
rect 40309 332830 42951 332832
rect 40309 332827 40375 332830
rect 42885 332827 42951 332830
rect 673545 332754 673611 332757
rect 675109 332754 675175 332757
rect 673545 332752 675175 332754
rect 673545 332696 673550 332752
rect 673606 332696 675114 332752
rect 675170 332696 675175 332752
rect 673545 332694 675175 332696
rect 673545 332691 673611 332694
rect 675109 332691 675175 332694
rect 39849 332482 39915 332485
rect 43069 332482 43135 332485
rect 39849 332480 43135 332482
rect 39849 332424 39854 332480
rect 39910 332424 43074 332480
rect 43130 332424 43135 332480
rect 39849 332422 43135 332424
rect 39849 332419 39915 332422
rect 43069 332419 43135 332422
rect 671981 332346 672047 332349
rect 675109 332346 675175 332349
rect 671981 332344 675175 332346
rect 671981 332288 671986 332344
rect 672042 332288 675114 332344
rect 675170 332288 675175 332344
rect 671981 332286 675175 332288
rect 671981 332283 672047 332286
rect 675109 332283 675175 332286
rect 673913 331258 673979 331261
rect 675109 331258 675175 331261
rect 673913 331256 675175 331258
rect 673913 331200 673918 331256
rect 673974 331200 675114 331256
rect 675170 331200 675175 331256
rect 673913 331198 675175 331200
rect 673913 331195 673979 331198
rect 675109 331195 675175 331198
rect 652385 329762 652451 329765
rect 649950 329760 652451 329762
rect 649950 329704 652390 329760
rect 652446 329704 652451 329760
rect 649950 329702 652451 329704
rect 649950 329234 650010 329702
rect 652385 329699 652451 329702
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 651373 328130 651439 328133
rect 649950 328128 651439 328130
rect 649950 328072 651378 328128
rect 651434 328072 651439 328128
rect 649950 328070 651439 328072
rect 649950 328052 650010 328070
rect 651373 328067 651439 328070
rect 42425 327042 42491 327045
rect 45277 327042 45343 327045
rect 42425 327040 45343 327042
rect 42425 326984 42430 327040
rect 42486 326984 45282 327040
rect 45338 326984 45343 327040
rect 42425 326982 45343 326984
rect 42425 326979 42491 326982
rect 45277 326979 45343 326982
rect 652017 326906 652083 326909
rect 650502 326904 652083 326906
rect 650502 326900 652022 326904
rect 649980 326848 652022 326900
rect 652078 326848 652083 326904
rect 649980 326846 652083 326848
rect 649980 326840 650562 326846
rect 652017 326843 652083 326846
rect 649950 325682 650010 325710
rect 651373 325682 651439 325685
rect 649950 325680 651439 325682
rect 649950 325624 651378 325680
rect 651434 325624 651439 325680
rect 649950 325622 651439 325624
rect 651373 325619 651439 325622
rect 675293 325546 675359 325549
rect 676254 325546 676260 325548
rect 675293 325544 676260 325546
rect 675293 325488 675298 325544
rect 675354 325488 676260 325544
rect 675293 325486 676260 325488
rect 675293 325483 675359 325486
rect 676254 325484 676260 325486
rect 676324 325484 676330 325548
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 675109 325274 675175 325277
rect 676806 325274 676812 325276
rect 675109 325272 676812 325274
rect 675109 325216 675114 325272
rect 675170 325216 676812 325272
rect 675109 325214 676812 325216
rect 675109 325211 675175 325214
rect 676806 325212 676812 325214
rect 676876 325212 676882 325276
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 42057 322826 42123 322829
rect 44357 322826 44423 322829
rect 42057 322824 44423 322826
rect 42057 322768 42062 322824
rect 42118 322768 44362 322824
rect 44418 322768 44423 322824
rect 42057 322766 44423 322768
rect 42057 322763 42123 322766
rect 44357 322763 44423 322766
rect 42057 321194 42123 321197
rect 42885 321194 42951 321197
rect 42057 321192 42951 321194
rect 42057 321136 42062 321192
rect 42118 321136 42890 321192
rect 42946 321136 42951 321192
rect 42057 321134 42951 321136
rect 42057 321131 42123 321134
rect 42885 321131 42951 321134
rect 42609 320786 42675 320789
rect 53833 320786 53899 320789
rect 42609 320784 53899 320786
rect 42609 320728 42614 320784
rect 42670 320728 53838 320784
rect 53894 320728 53899 320784
rect 42609 320726 53899 320728
rect 42609 320723 42675 320726
rect 53833 320723 53899 320726
rect 42149 320514 42215 320517
rect 43069 320514 43135 320517
rect 42149 320512 43135 320514
rect 42149 320456 42154 320512
rect 42210 320456 43074 320512
rect 43130 320456 43135 320512
rect 42149 320454 43135 320456
rect 42149 320451 42215 320454
rect 43069 320451 43135 320454
rect 41873 319972 41939 319973
rect 41822 319970 41828 319972
rect 41782 319910 41828 319970
rect 41892 319968 41939 319972
rect 41934 319912 41939 319968
rect 41822 319908 41828 319910
rect 41892 319908 41939 319912
rect 41873 319907 41939 319908
rect 42057 319970 42123 319973
rect 44173 319970 44239 319973
rect 42057 319968 44239 319970
rect 42057 319912 42062 319968
rect 42118 319912 44178 319968
rect 44234 319912 44239 319968
rect 42057 319910 44239 319912
rect 42057 319907 42123 319910
rect 44173 319907 44239 319910
rect 42425 319426 42491 319429
rect 53097 319426 53163 319429
rect 42425 319424 53163 319426
rect 42425 319368 42430 319424
rect 42486 319368 53102 319424
rect 53158 319368 53163 319424
rect 42425 319366 53163 319368
rect 42425 319363 42491 319366
rect 53097 319363 53163 319366
rect 40718 318956 40724 319020
rect 40788 319018 40794 319020
rect 42241 319018 42307 319021
rect 40788 319016 42307 319018
rect 40788 318960 42246 319016
rect 42302 318960 42307 319016
rect 40788 318958 42307 318960
rect 40788 318956 40794 318958
rect 42241 318955 42307 318958
rect 40534 317324 40540 317388
rect 40604 317386 40610 317388
rect 41781 317386 41847 317389
rect 40604 317384 41847 317386
rect 40604 317328 41786 317384
rect 41842 317328 41847 317384
rect 40604 317326 41847 317328
rect 40604 317324 40610 317326
rect 41781 317323 41847 317326
rect 62113 317386 62179 317389
rect 62113 317384 64706 317386
rect 62113 317328 62118 317384
rect 62174 317328 64706 317384
rect 62113 317326 64706 317328
rect 62113 317323 62179 317326
rect 64646 317106 64706 317326
rect 42149 316026 42215 316029
rect 43110 316026 43116 316028
rect 42149 316024 43116 316026
rect 42149 315968 42154 316024
rect 42210 315968 43116 316024
rect 42149 315966 43116 315968
rect 42149 315963 42215 315966
rect 43110 315964 43116 315966
rect 43180 315964 43186 316028
rect 62113 316026 62179 316029
rect 62113 316024 64706 316026
rect 62113 315968 62118 316024
rect 62174 315968 64706 316024
rect 62113 315966 64706 315968
rect 62113 315963 62179 315966
rect 64646 315924 64706 315966
rect 42149 315482 42215 315485
rect 45553 315482 45619 315485
rect 42149 315480 45619 315482
rect 42149 315424 42154 315480
rect 42210 315424 45558 315480
rect 45614 315424 45619 315480
rect 42149 315422 45619 315424
rect 42149 315419 42215 315422
rect 45553 315419 45619 315422
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 63125 314122 63191 314125
rect 63125 314120 64706 314122
rect 63125 314064 63130 314120
rect 63186 314064 64706 314120
rect 63125 314062 64706 314064
rect 63125 314059 63191 314062
rect 42057 313716 42123 313717
rect 42006 313714 42012 313716
rect 41966 313654 42012 313714
rect 42076 313712 42123 313716
rect 42118 313656 42123 313712
rect 42006 313652 42012 313654
rect 42076 313652 42123 313656
rect 42057 313651 42123 313652
rect 64646 313560 64706 314062
rect 676213 313986 676279 313989
rect 676213 313984 676322 313986
rect 676213 313928 676218 313984
rect 676274 313928 676322 313984
rect 676213 313923 676322 313928
rect 676262 313684 676322 313923
rect 653397 313306 653463 313309
rect 653397 313304 676292 313306
rect 653397 313248 653402 313304
rect 653458 313248 676292 313304
rect 653397 313246 676292 313248
rect 653397 313243 653463 313246
rect 62941 313034 63007 313037
rect 62941 313032 64706 313034
rect 62941 312976 62946 313032
rect 63002 312976 64706 313032
rect 62941 312974 64706 312976
rect 62941 312971 63007 312974
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 64646 312378 64706 312974
rect 669270 312838 676292 312898
rect 664437 312082 664503 312085
rect 669270 312082 669330 312838
rect 672533 312490 672599 312493
rect 672533 312488 676292 312490
rect 672533 312432 672538 312488
rect 672594 312432 676292 312488
rect 672533 312430 676292 312432
rect 672533 312427 672599 312430
rect 664437 312080 669330 312082
rect 664437 312024 664442 312080
rect 664498 312024 669330 312080
rect 664437 312022 669330 312024
rect 673361 312082 673427 312085
rect 673361 312080 676292 312082
rect 673361 312024 673366 312080
rect 673422 312024 676292 312080
rect 673361 312022 676292 312024
rect 664437 312019 664503 312022
rect 673361 312019 673427 312022
rect 62757 311810 62823 311813
rect 62757 311808 64706 311810
rect 62757 311752 62762 311808
rect 62818 311752 64706 311808
rect 62757 311750 64706 311752
rect 62757 311747 62823 311750
rect 64646 311196 64706 311750
rect 672533 311674 672599 311677
rect 672533 311672 676292 311674
rect 672533 311616 672538 311672
rect 672594 311616 676292 311672
rect 672533 311614 676292 311616
rect 672533 311611 672599 311614
rect 672717 311266 672783 311269
rect 672717 311264 676292 311266
rect 672717 311208 672722 311264
rect 672778 311208 676292 311264
rect 672717 311206 676292 311208
rect 672717 311203 672783 311206
rect 673085 310858 673151 310861
rect 673085 310856 676292 310858
rect 673085 310800 673090 310856
rect 673146 310800 676292 310856
rect 673085 310798 676292 310800
rect 673085 310795 673151 310798
rect 672717 310586 672783 310589
rect 673177 310586 673243 310589
rect 672717 310584 673243 310586
rect 672717 310528 672722 310584
rect 672778 310528 673182 310584
rect 673238 310528 673243 310584
rect 672717 310526 673243 310528
rect 672717 310523 672783 310526
rect 673177 310523 673243 310526
rect 42425 310450 42491 310453
rect 46933 310450 46999 310453
rect 42425 310448 46999 310450
rect 42425 310392 42430 310448
rect 42486 310392 46938 310448
rect 46994 310392 46999 310448
rect 42425 310390 46999 310392
rect 42425 310387 42491 310390
rect 46933 310387 46999 310390
rect 674649 310450 674715 310453
rect 674649 310448 676292 310450
rect 674649 310392 674654 310448
rect 674710 310392 676292 310448
rect 674649 310390 676292 310392
rect 674649 310387 674715 310390
rect 674465 310042 674531 310045
rect 674465 310040 676292 310042
rect 674465 309984 674470 310040
rect 674526 309984 676292 310040
rect 674465 309982 676292 309984
rect 674465 309979 674531 309982
rect 652293 309906 652359 309909
rect 652293 309904 663810 309906
rect 652293 309848 652298 309904
rect 652354 309848 663810 309904
rect 652293 309846 663810 309848
rect 652293 309843 652359 309846
rect 663750 309362 663810 309846
rect 674189 309634 674255 309637
rect 674189 309632 676292 309634
rect 674189 309576 674194 309632
rect 674250 309576 676292 309632
rect 674189 309574 676292 309576
rect 674189 309571 674255 309574
rect 675845 309362 675911 309365
rect 663750 309360 675911 309362
rect 663750 309304 675850 309360
rect 675906 309304 675911 309360
rect 663750 309302 675911 309304
rect 675845 309299 675911 309302
rect 676032 309166 676292 309226
rect 42057 309090 42123 309093
rect 59905 309090 59971 309093
rect 42057 309088 59971 309090
rect 42057 309032 42062 309088
rect 42118 309032 59910 309088
rect 59966 309032 59971 309088
rect 42057 309030 59971 309032
rect 42057 309027 42123 309030
rect 59905 309027 59971 309030
rect 675702 309028 675708 309092
rect 675772 309090 675778 309092
rect 676032 309090 676092 309166
rect 675772 309030 676092 309090
rect 675772 309028 675778 309030
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675109 308002 675175 308005
rect 675109 308000 676292 308002
rect 675109 307944 675114 308000
rect 675170 307944 676292 308000
rect 675109 307942 676292 307944
rect 675109 307939 675175 307942
rect 676029 307594 676095 307597
rect 676029 307592 676292 307594
rect 676029 307536 676034 307592
rect 676090 307536 676292 307592
rect 676029 307534 676292 307536
rect 676029 307531 676095 307534
rect 675886 307124 675892 307188
rect 675956 307186 675962 307188
rect 675956 307126 676292 307186
rect 675956 307124 675962 307126
rect 679617 306778 679683 306781
rect 679604 306776 679683 306778
rect 679604 306720 679622 306776
rect 679678 306720 679683 306776
rect 679604 306718 679683 306720
rect 679617 306715 679683 306718
rect 677593 306370 677659 306373
rect 677580 306368 677659 306370
rect 677580 306312 677598 306368
rect 677654 306312 677659 306368
rect 677580 306310 677659 306312
rect 677593 306307 677659 306310
rect 676029 305962 676095 305965
rect 676029 305960 676292 305962
rect 676029 305904 676034 305960
rect 676090 305904 676292 305960
rect 676029 305902 676292 305904
rect 676029 305899 676095 305902
rect 672257 305554 672323 305557
rect 672257 305552 676292 305554
rect 672257 305496 672262 305552
rect 672318 305496 676292 305552
rect 672257 305494 676292 305496
rect 672257 305491 672323 305494
rect 674373 305146 674439 305149
rect 674373 305144 676292 305146
rect 674373 305088 674378 305144
rect 674434 305088 676292 305144
rect 674373 305086 676292 305088
rect 674373 305083 674439 305086
rect 676630 304570 676690 304708
rect 676622 304506 676628 304570
rect 676692 304506 676698 304570
rect 672073 304330 672139 304333
rect 672073 304328 676292 304330
rect 672073 304272 672078 304328
rect 672134 304272 676292 304328
rect 672073 304270 676292 304272
rect 672073 304267 672139 304270
rect 674005 303922 674071 303925
rect 674005 303920 676292 303922
rect 674005 303864 674010 303920
rect 674066 303864 676292 303920
rect 674005 303862 676292 303864
rect 674005 303859 674071 303862
rect 674649 303514 674715 303517
rect 674649 303512 676292 303514
rect 674649 303456 674654 303512
rect 674710 303456 676292 303512
rect 674649 303454 676292 303456
rect 674649 303451 674715 303454
rect 651373 303378 651439 303381
rect 649950 303376 651439 303378
rect 649950 303320 651378 303376
rect 651434 303320 651439 303376
rect 649950 303318 651439 303320
rect 649950 302776 650010 303318
rect 651373 303315 651439 303318
rect 683070 302701 683130 303076
rect 683021 302696 683130 302701
rect 683021 302640 683026 302696
rect 683082 302668 683130 302696
rect 683082 302640 683100 302668
rect 683021 302638 683100 302640
rect 683021 302635 683087 302638
rect 671521 302290 671587 302293
rect 671521 302288 676292 302290
rect 671521 302232 671526 302288
rect 671582 302232 676292 302288
rect 671521 302230 676292 302232
rect 671521 302227 671587 302230
rect 652293 302154 652359 302157
rect 649950 302152 652359 302154
rect 649950 302096 652298 302152
rect 652354 302096 652359 302152
rect 649950 302094 652359 302096
rect 649950 301594 650010 302094
rect 652293 302091 652359 302094
rect 674833 302018 674899 302021
rect 675845 302018 675911 302021
rect 674833 302016 675911 302018
rect 674833 301960 674838 302016
rect 674894 301960 675850 302016
rect 675906 301960 675911 302016
rect 674833 301958 675911 301960
rect 674833 301955 674899 301958
rect 675845 301955 675911 301958
rect 53097 301338 53163 301341
rect 41492 301336 53163 301338
rect 41492 301280 53102 301336
rect 53158 301280 53163 301336
rect 41492 301278 53163 301280
rect 53097 301275 53163 301278
rect 35617 300930 35683 300933
rect 35604 300928 35683 300930
rect 35604 300872 35622 300928
rect 35678 300872 35683 300928
rect 35604 300870 35683 300872
rect 35617 300867 35683 300870
rect 654777 300930 654843 300933
rect 676262 300930 676322 301852
rect 654777 300928 676322 300930
rect 654777 300872 654782 300928
rect 654838 300872 676322 300928
rect 654777 300870 676322 300872
rect 654777 300867 654843 300870
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 46197 300522 46263 300525
rect 41492 300520 46263 300522
rect 41492 300464 46202 300520
rect 46258 300464 46263 300520
rect 41492 300462 46263 300464
rect 46197 300459 46263 300462
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 676029 300658 676095 300661
rect 676438 300658 676444 300660
rect 676029 300656 676444 300658
rect 676029 300600 676034 300656
rect 676090 300600 676444 300656
rect 676029 300598 676444 300600
rect 676029 300595 676095 300598
rect 676438 300596 676444 300598
rect 676508 300596 676514 300660
rect 44398 300114 44404 300116
rect 41492 300054 44404 300114
rect 44398 300052 44404 300054
rect 44468 300052 44474 300116
rect 44357 299706 44423 299709
rect 41492 299704 44423 299706
rect 41492 299648 44362 299704
rect 44418 299648 44423 299704
rect 41492 299646 44423 299648
rect 44357 299643 44423 299646
rect 675702 299372 675708 299436
rect 675772 299434 675778 299436
rect 683021 299434 683087 299437
rect 675772 299432 683087 299434
rect 675772 299376 683026 299432
rect 683082 299376 683087 299432
rect 675772 299374 683087 299376
rect 675772 299372 675778 299374
rect 683021 299371 683087 299374
rect 44582 299298 44588 299300
rect 41492 299238 44588 299298
rect 44582 299236 44588 299238
rect 44652 299236 44658 299300
rect 35801 298890 35867 298893
rect 35788 298888 35867 298890
rect 35788 298832 35806 298888
rect 35862 298832 35867 298888
rect 35788 298830 35867 298832
rect 35801 298827 35867 298830
rect 41781 298754 41847 298757
rect 62757 298754 62823 298757
rect 41781 298752 62823 298754
rect 41781 298696 41786 298752
rect 41842 298696 62762 298752
rect 62818 298696 62823 298752
rect 41781 298694 62823 298696
rect 649950 298754 650010 299230
rect 651465 298754 651531 298757
rect 649950 298752 651531 298754
rect 649950 298696 651470 298752
rect 651526 298696 651531 298752
rect 649950 298694 651531 298696
rect 41781 298691 41847 298694
rect 62757 298691 62823 298694
rect 651465 298691 651531 298694
rect 44214 298482 44220 298484
rect 41492 298422 44220 298482
rect 44214 298420 44220 298422
rect 44284 298420 44290 298484
rect 44817 298074 44883 298077
rect 41492 298072 44883 298074
rect 41492 298016 44822 298072
rect 44878 298016 44883 298072
rect 41492 298014 44883 298016
rect 44817 298011 44883 298014
rect 42742 297666 42748 297668
rect 41492 297606 42748 297666
rect 42742 297604 42748 297606
rect 42812 297604 42818 297668
rect 649950 297530 650010 298048
rect 651465 297530 651531 297533
rect 649950 297528 651531 297530
rect 649950 297472 651470 297528
rect 651526 297472 651531 297528
rect 649950 297470 651531 297472
rect 651465 297467 651531 297470
rect 675518 297332 675524 297396
rect 675588 297394 675594 297396
rect 675937 297394 676003 297397
rect 675588 297392 676003 297394
rect 675588 297336 675942 297392
rect 675998 297336 676003 297392
rect 675588 297334 676003 297336
rect 675588 297332 675594 297334
rect 675937 297331 676003 297334
rect 44173 297258 44239 297261
rect 41492 297256 44239 297258
rect 41492 297200 44178 297256
rect 44234 297200 44239 297256
rect 41492 297198 44239 297200
rect 44173 297195 44239 297198
rect 42006 296850 42012 296852
rect 41492 296790 42012 296850
rect 42006 296788 42012 296790
rect 42076 296788 42082 296852
rect 649950 296850 650010 296866
rect 652661 296850 652727 296853
rect 649950 296848 652727 296850
rect 649950 296792 652666 296848
rect 652722 296792 652727 296848
rect 649950 296790 652727 296792
rect 652661 296787 652727 296790
rect 41781 296578 41847 296581
rect 42793 296578 42859 296581
rect 41781 296576 42859 296578
rect 41781 296520 41786 296576
rect 41842 296520 42798 296576
rect 42854 296520 42859 296576
rect 41781 296518 42859 296520
rect 41781 296515 41847 296518
rect 42793 296515 42859 296518
rect 675201 296578 675267 296581
rect 675845 296578 675911 296581
rect 676121 296578 676187 296581
rect 675201 296576 675911 296578
rect 675201 296520 675206 296576
rect 675262 296520 675850 296576
rect 675906 296520 675911 296576
rect 675201 296518 675911 296520
rect 675201 296515 675267 296518
rect 675845 296515 675911 296518
rect 676078 296576 676187 296578
rect 676078 296520 676126 296576
rect 676182 296520 676187 296576
rect 676078 296515 676187 296520
rect 35433 296442 35499 296445
rect 35420 296440 35499 296442
rect 35420 296384 35438 296440
rect 35494 296384 35499 296440
rect 35420 296382 35499 296384
rect 35433 296379 35499 296382
rect 35617 296034 35683 296037
rect 35604 296032 35683 296034
rect 35604 295976 35622 296032
rect 35678 295976 35683 296032
rect 35604 295974 35683 295976
rect 35617 295971 35683 295974
rect 667749 295762 667815 295765
rect 675385 295762 675451 295765
rect 667749 295760 675451 295762
rect 667749 295704 667754 295760
rect 667810 295704 675390 295760
rect 675446 295704 675451 295760
rect 667749 295702 675451 295704
rect 667749 295699 667815 295702
rect 675385 295699 675451 295702
rect 675753 295762 675819 295765
rect 676078 295762 676138 296515
rect 675753 295760 676138 295762
rect 675753 295704 675758 295760
rect 675814 295704 676138 295760
rect 675753 295702 676138 295704
rect 675753 295699 675819 295702
rect 35801 295626 35867 295629
rect 35788 295624 35867 295626
rect 35788 295568 35806 295624
rect 35862 295568 35867 295624
rect 35788 295566 35867 295568
rect 35801 295563 35867 295566
rect 62113 295490 62179 295493
rect 64646 295490 64706 295684
rect 62113 295488 64706 295490
rect 62113 295432 62118 295488
rect 62174 295432 64706 295488
rect 62113 295430 64706 295432
rect 62113 295427 62179 295430
rect 41781 295354 41847 295357
rect 43161 295354 43227 295357
rect 41781 295352 43227 295354
rect 41781 295296 41786 295352
rect 41842 295296 43166 295352
rect 43222 295296 43227 295352
rect 41781 295294 43227 295296
rect 649950 295354 650010 295684
rect 652385 295354 652451 295357
rect 649950 295352 652451 295354
rect 649950 295296 652390 295352
rect 652446 295296 652451 295352
rect 649950 295294 652451 295296
rect 41781 295291 41847 295294
rect 43161 295291 43227 295294
rect 652385 295291 652451 295294
rect 35801 295218 35867 295221
rect 35788 295216 35867 295218
rect 35788 295160 35806 295216
rect 35862 295160 35867 295216
rect 35788 295158 35867 295160
rect 35801 295155 35867 295158
rect 33777 294810 33843 294813
rect 33764 294808 33843 294810
rect 33764 294752 33782 294808
rect 33838 294752 33843 294808
rect 33764 294750 33843 294752
rect 33777 294747 33843 294750
rect 675753 294538 675819 294541
rect 676254 294538 676260 294540
rect 675753 294536 676260 294538
rect 32397 294402 32463 294405
rect 32397 294400 32476 294402
rect 32397 294344 32402 294400
rect 32458 294344 32476 294400
rect 32397 294342 32476 294344
rect 32397 294339 32463 294342
rect 62113 294130 62179 294133
rect 64646 294130 64706 294502
rect 649950 294266 650010 294502
rect 675753 294480 675758 294536
rect 675814 294480 676260 294536
rect 675753 294478 676260 294480
rect 675753 294475 675819 294478
rect 676254 294476 676260 294478
rect 676324 294476 676330 294540
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 651465 294203 651531 294206
rect 62113 294128 64706 294130
rect 62113 294072 62118 294128
rect 62174 294072 64706 294128
rect 62113 294070 64706 294072
rect 62113 294067 62179 294070
rect 45001 293994 45067 293997
rect 41492 293992 45067 293994
rect 41492 293936 45006 293992
rect 45062 293936 45067 293992
rect 41492 293934 45067 293936
rect 45001 293931 45067 293934
rect 662413 293858 662479 293861
rect 667749 293858 667815 293861
rect 662413 293856 667815 293858
rect 662413 293800 662418 293856
rect 662474 293800 667754 293856
rect 667810 293800 667815 293856
rect 662413 293798 667815 293800
rect 662413 293795 662479 293798
rect 667749 293795 667815 293798
rect 44541 293586 44607 293589
rect 41492 293584 44607 293586
rect 41492 293528 44546 293584
rect 44602 293528 44607 293584
rect 41492 293526 44607 293528
rect 44541 293523 44607 293526
rect 35801 293178 35867 293181
rect 35788 293176 35867 293178
rect 35788 293120 35806 293176
rect 35862 293120 35867 293176
rect 35788 293118 35867 293120
rect 35801 293115 35867 293118
rect 35801 292770 35867 292773
rect 35788 292768 35867 292770
rect 35788 292712 35806 292768
rect 35862 292712 35867 292768
rect 35788 292710 35867 292712
rect 35801 292707 35867 292710
rect 62297 292770 62363 292773
rect 64646 292770 64706 293320
rect 649950 293042 650010 293320
rect 651465 293042 651531 293045
rect 649950 293040 651531 293042
rect 649950 292984 651470 293040
rect 651526 292984 651531 293040
rect 649950 292982 651531 292984
rect 651465 292979 651531 292982
rect 62297 292768 64706 292770
rect 62297 292712 62302 292768
rect 62358 292712 64706 292768
rect 62297 292710 64706 292712
rect 62297 292707 62363 292710
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40542 292332 40602 292528
rect 62113 292498 62179 292501
rect 62113 292496 64706 292498
rect 62113 292440 62118 292496
rect 62174 292440 64706 292496
rect 62113 292438 64706 292440
rect 62113 292435 62179 292438
rect 64646 292138 64706 292438
rect 675569 292228 675635 292229
rect 675518 292164 675524 292228
rect 675588 292226 675635 292228
rect 675588 292224 675680 292226
rect 675630 292168 675680 292224
rect 675588 292166 675680 292168
rect 675588 292164 675635 292166
rect 675569 292163 675635 292164
rect 42241 291954 42307 291957
rect 41492 291952 42307 291954
rect 41492 291896 42246 291952
rect 42302 291896 42307 291952
rect 41492 291894 42307 291896
rect 42241 291891 42307 291894
rect 41822 291546 41828 291548
rect 41492 291486 41828 291546
rect 41822 291484 41828 291486
rect 41892 291484 41898 291548
rect 649950 291546 650010 292138
rect 652201 291546 652267 291549
rect 649950 291544 652267 291546
rect 649950 291488 652206 291544
rect 652262 291488 652267 291544
rect 649950 291486 652267 291488
rect 652201 291483 652267 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 35801 291138 35867 291141
rect 35788 291136 35867 291138
rect 35788 291080 35806 291136
rect 35862 291080 35867 291136
rect 35788 291078 35867 291080
rect 35801 291075 35867 291078
rect 41781 291138 41847 291141
rect 42977 291138 43043 291141
rect 41781 291136 43043 291138
rect 41781 291080 41786 291136
rect 41842 291080 42982 291136
rect 43038 291080 43043 291136
rect 41781 291078 43043 291080
rect 41781 291075 41847 291078
rect 42977 291075 43043 291078
rect 62113 291002 62179 291005
rect 62113 291000 64154 291002
rect 62113 290944 62118 291000
rect 62174 290986 64154 291000
rect 62174 290944 64676 290986
rect 62113 290942 64676 290944
rect 62113 290939 62179 290942
rect 64094 290926 64676 290942
rect 50521 290730 50587 290733
rect 41492 290728 50587 290730
rect 41492 290672 50526 290728
rect 50582 290672 50587 290728
rect 41492 290670 50587 290672
rect 50521 290667 50587 290670
rect 649950 290458 650010 290956
rect 675753 290866 675819 290869
rect 676622 290866 676628 290868
rect 675753 290864 676628 290866
rect 675753 290808 675758 290864
rect 675814 290808 676628 290864
rect 675753 290806 676628 290808
rect 675753 290803 675819 290806
rect 676622 290804 676628 290806
rect 676692 290804 676698 290868
rect 651465 290458 651531 290461
rect 649950 290456 651531 290458
rect 649950 290400 651470 290456
rect 651526 290400 651531 290456
rect 649950 290398 651531 290400
rect 651465 290395 651531 290398
rect 35617 290322 35683 290325
rect 35604 290320 35683 290322
rect 35604 290264 35622 290320
rect 35678 290264 35683 290320
rect 35604 290262 35683 290264
rect 35617 290259 35683 290262
rect 48957 289914 49023 289917
rect 41492 289912 49023 289914
rect 41492 289856 48962 289912
rect 49018 289856 49023 289912
rect 41492 289854 49023 289856
rect 48957 289851 49023 289854
rect 62757 289778 62823 289781
rect 62757 289776 64706 289778
rect 62757 289720 62762 289776
rect 62818 289720 64706 289776
rect 62757 289718 64706 289720
rect 62757 289715 62823 289718
rect 40718 289172 40724 289236
rect 40788 289234 40794 289236
rect 42241 289234 42307 289237
rect 40788 289232 42307 289234
rect 40788 289176 42246 289232
rect 42302 289176 42307 289232
rect 40788 289174 42307 289176
rect 649950 289234 650010 289774
rect 651465 289234 651531 289237
rect 649950 289232 651531 289234
rect 649950 289176 651470 289232
rect 651526 289176 651531 289232
rect 649950 289174 651531 289176
rect 40788 289172 40794 289174
rect 42241 289171 42307 289174
rect 651465 289171 651531 289174
rect 39205 288962 39271 288965
rect 43621 288962 43687 288965
rect 39205 288960 43687 288962
rect 39205 288904 39210 288960
rect 39266 288904 43626 288960
rect 43682 288904 43687 288960
rect 39205 288902 43687 288904
rect 39205 288899 39271 288902
rect 43621 288899 43687 288902
rect 62113 288554 62179 288557
rect 64646 288554 64706 288592
rect 62113 288552 64706 288554
rect 62113 288496 62118 288552
rect 62174 288496 64706 288552
rect 62113 288494 64706 288496
rect 649950 288554 650010 288592
rect 652017 288554 652083 288557
rect 649950 288552 652083 288554
rect 649950 288496 652022 288552
rect 652078 288496 652083 288552
rect 649950 288494 652083 288496
rect 62113 288491 62179 288494
rect 652017 288491 652083 288494
rect 672073 287874 672139 287877
rect 675109 287874 675175 287877
rect 672073 287872 675175 287874
rect 672073 287816 672078 287872
rect 672134 287816 675114 287872
rect 675170 287816 675175 287872
rect 672073 287814 675175 287816
rect 672073 287811 672139 287814
rect 675109 287811 675175 287814
rect 651465 287466 651531 287469
rect 649766 287464 651531 287466
rect 63125 287194 63191 287197
rect 64646 287194 64706 287410
rect 649766 287408 651470 287464
rect 651526 287408 651531 287464
rect 649766 287406 651531 287408
rect 651465 287403 651531 287406
rect 63125 287192 64706 287194
rect 63125 287136 63130 287192
rect 63186 287136 64706 287192
rect 63125 287134 64706 287136
rect 63125 287131 63191 287134
rect 674005 286514 674071 286517
rect 675385 286514 675451 286517
rect 674005 286512 675451 286514
rect 674005 286456 674010 286512
rect 674066 286456 675390 286512
rect 675446 286456 675451 286512
rect 674005 286454 675451 286456
rect 674005 286451 674071 286454
rect 675385 286451 675451 286454
rect 62113 285970 62179 285973
rect 64646 285970 64706 286228
rect 62113 285968 64706 285970
rect 62113 285912 62118 285968
rect 62174 285912 64706 285968
rect 62113 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 62113 285907 62179 285910
rect 651465 285907 651531 285910
rect 672257 285562 672323 285565
rect 675109 285562 675175 285565
rect 672257 285560 675175 285562
rect 672257 285504 672262 285560
rect 672318 285504 675114 285560
rect 675170 285504 675175 285560
rect 672257 285502 675175 285504
rect 672257 285499 672323 285502
rect 675109 285499 675175 285502
rect 32397 284882 32463 284885
rect 41638 284882 41644 284884
rect 32397 284880 41644 284882
rect 32397 284824 32402 284880
rect 32458 284824 41644 284880
rect 32397 284822 41644 284824
rect 32397 284819 32463 284822
rect 41638 284820 41644 284822
rect 41708 284820 41714 284884
rect 62113 284474 62179 284477
rect 64646 284474 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 62113 284472 64706 284474
rect 62113 284416 62118 284472
rect 62174 284416 64706 284472
rect 62113 284414 64706 284416
rect 62113 284411 62179 284414
rect 40677 284338 40743 284341
rect 42006 284338 42012 284340
rect 40677 284336 42012 284338
rect 40677 284280 40682 284336
rect 40738 284280 42012 284336
rect 40677 284278 42012 284280
rect 40677 284275 40743 284278
rect 42006 284276 42012 284278
rect 42076 284276 42082 284340
rect 62757 283250 62823 283253
rect 64646 283250 64706 283864
rect 649950 283386 650010 283864
rect 675661 283658 675727 283661
rect 675886 283658 675892 283660
rect 675661 283656 675892 283658
rect 675661 283600 675666 283656
rect 675722 283600 675892 283656
rect 675661 283598 675892 283600
rect 675661 283595 675727 283598
rect 675886 283596 675892 283598
rect 675956 283596 675962 283660
rect 652385 283522 652451 283525
rect 674373 283522 674439 283525
rect 652385 283520 674439 283522
rect 652385 283464 652390 283520
rect 652446 283464 674378 283520
rect 674434 283464 674439 283520
rect 652385 283462 674439 283464
rect 652385 283459 652451 283462
rect 674373 283459 674439 283462
rect 651465 283386 651531 283389
rect 649950 283384 651531 283386
rect 649950 283328 651470 283384
rect 651526 283328 651531 283384
rect 649950 283326 651531 283328
rect 651465 283323 651531 283326
rect 62757 283248 64706 283250
rect 62757 283192 62762 283248
rect 62818 283192 64706 283248
rect 62757 283190 64706 283192
rect 62757 283187 62823 283190
rect 675661 282844 675727 282845
rect 675661 282840 675708 282844
rect 675772 282842 675778 282844
rect 675661 282784 675666 282840
rect 675661 282780 675708 282784
rect 675772 282782 675818 282842
rect 675772 282780 675778 282782
rect 675661 282779 675727 282780
rect 62941 282162 63007 282165
rect 64646 282162 64706 282682
rect 62941 282160 64706 282162
rect 62941 282104 62946 282160
rect 63002 282104 64706 282160
rect 62941 282102 64706 282104
rect 649950 282162 650010 282682
rect 652385 282162 652451 282165
rect 649950 282160 652451 282162
rect 649950 282104 652390 282160
rect 652446 282104 652451 282160
rect 649950 282102 652451 282104
rect 62941 282099 63007 282102
rect 652385 282099 652451 282102
rect 62113 280938 62179 280941
rect 64646 280938 64706 281500
rect 62113 280936 64706 280938
rect 62113 280880 62118 280936
rect 62174 280880 64706 280936
rect 62113 280878 64706 280880
rect 649950 280938 650010 281500
rect 675753 281210 675819 281213
rect 676070 281210 676076 281212
rect 675753 281208 676076 281210
rect 675753 281152 675758 281208
rect 675814 281152 676076 281208
rect 675753 281150 676076 281152
rect 675753 281147 675819 281150
rect 676070 281148 676076 281150
rect 676140 281148 676146 281212
rect 651465 280938 651531 280941
rect 649950 280936 651531 280938
rect 649950 280880 651470 280936
rect 651526 280880 651531 280936
rect 649950 280878 651531 280880
rect 62113 280875 62179 280878
rect 651465 280875 651531 280878
rect 61377 280394 61443 280397
rect 652569 280394 652635 280397
rect 61377 280392 64706 280394
rect 61377 280336 61382 280392
rect 61438 280336 64706 280392
rect 61377 280334 64706 280336
rect 61377 280331 61443 280334
rect 64646 280318 64706 280334
rect 649950 280392 652635 280394
rect 649950 280336 652574 280392
rect 652630 280336 652635 280392
rect 649950 280334 652635 280336
rect 649950 280318 650010 280334
rect 652569 280331 652635 280334
rect 42425 278762 42491 278765
rect 58617 278762 58683 278765
rect 42425 278760 58683 278762
rect 42425 278704 42430 278760
rect 42486 278704 58622 278760
rect 58678 278704 58683 278760
rect 42425 278702 58683 278704
rect 42425 278699 42491 278702
rect 58617 278699 58683 278702
rect 40902 278428 40908 278492
rect 40972 278490 40978 278492
rect 41781 278490 41847 278493
rect 40972 278488 41847 278490
rect 40972 278432 41786 278488
rect 41842 278432 41847 278488
rect 40972 278430 41847 278432
rect 40972 278428 40978 278430
rect 41781 278427 41847 278430
rect 42057 277810 42123 277813
rect 43621 277810 43687 277813
rect 42057 277808 43687 277810
rect 42057 277752 42062 277808
rect 42118 277752 43626 277808
rect 43682 277752 43687 277808
rect 42057 277750 43687 277752
rect 42057 277747 42123 277750
rect 43621 277747 43687 277750
rect 40718 277068 40724 277132
rect 40788 277130 40794 277132
rect 41781 277130 41847 277133
rect 40788 277128 41847 277130
rect 40788 277072 41786 277128
rect 41842 277072 41847 277128
rect 40788 277070 41847 277072
rect 40788 277068 40794 277070
rect 41781 277067 41847 277070
rect 42609 275906 42675 275909
rect 57237 275906 57303 275909
rect 42609 275904 57303 275906
rect 42609 275848 42614 275904
rect 42670 275848 57242 275904
rect 57298 275848 57303 275904
rect 42609 275846 57303 275848
rect 42609 275843 42675 275846
rect 57237 275843 57303 275846
rect 537293 275090 537359 275093
rect 538121 275090 538187 275093
rect 537293 275088 538187 275090
rect 537293 275032 537298 275088
rect 537354 275032 538126 275088
rect 538182 275032 538187 275088
rect 537293 275030 538187 275032
rect 537293 275027 537359 275030
rect 538121 275027 538187 275030
rect 542261 274818 542327 274821
rect 543181 274818 543247 274821
rect 542261 274816 543247 274818
rect 542261 274760 542266 274816
rect 542322 274760 543186 274816
rect 543242 274760 543247 274816
rect 542261 274758 543247 274760
rect 542261 274755 542327 274758
rect 543181 274755 543247 274758
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 547505 274002 547571 274005
rect 549253 274002 549319 274005
rect 547505 274000 549319 274002
rect 547505 273944 547510 274000
rect 547566 273944 549258 274000
rect 549314 273944 549319 274000
rect 547505 273942 549319 273944
rect 547505 273939 547571 273942
rect 549253 273939 549319 273942
rect 539317 273730 539383 273733
rect 547689 273730 547755 273733
rect 539317 273728 547755 273730
rect 539317 273672 539322 273728
rect 539378 273672 547694 273728
rect 547750 273672 547755 273728
rect 539317 273670 547755 273672
rect 539317 273667 539383 273670
rect 547689 273667 547755 273670
rect 549897 273730 549963 273733
rect 552841 273730 552907 273733
rect 549897 273728 552907 273730
rect 549897 273672 549902 273728
rect 549958 273672 552846 273728
rect 552902 273672 552907 273728
rect 549897 273670 552907 273672
rect 549897 273667 549963 273670
rect 552841 273667 552907 273670
rect 42333 273186 42399 273189
rect 44541 273186 44607 273189
rect 42333 273184 44607 273186
rect 42333 273128 42338 273184
rect 42394 273128 44546 273184
rect 44602 273128 44607 273184
rect 42333 273126 44607 273128
rect 42333 273123 42399 273126
rect 44541 273123 44607 273126
rect 42425 272914 42491 272917
rect 45001 272914 45067 272917
rect 42425 272912 45067 272914
rect 42425 272856 42430 272912
rect 42486 272856 45006 272912
rect 45062 272856 45067 272912
rect 42425 272854 45067 272856
rect 42425 272851 42491 272854
rect 45001 272851 45067 272854
rect 489913 272778 489979 272781
rect 495709 272778 495775 272781
rect 489913 272776 495775 272778
rect 489913 272720 489918 272776
rect 489974 272720 495714 272776
rect 495770 272720 495775 272776
rect 489913 272718 495775 272720
rect 489913 272715 489979 272718
rect 495709 272715 495775 272718
rect 470409 272642 470475 272645
rect 470593 272642 470659 272645
rect 470409 272640 470659 272642
rect 470409 272584 470414 272640
rect 470470 272584 470598 272640
rect 470654 272584 470659 272640
rect 470409 272582 470659 272584
rect 470409 272579 470475 272582
rect 470593 272579 470659 272582
rect 41965 272372 42031 272373
rect 41965 272368 42012 272372
rect 42076 272370 42082 272372
rect 462221 272370 462287 272373
rect 470409 272370 470475 272373
rect 41965 272312 41970 272368
rect 41965 272308 42012 272312
rect 42076 272310 42122 272370
rect 462221 272368 470475 272370
rect 462221 272312 462226 272368
rect 462282 272312 470414 272368
rect 470470 272312 470475 272368
rect 462221 272310 470475 272312
rect 42076 272308 42082 272310
rect 41965 272307 42031 272308
rect 462221 272307 462287 272310
rect 470409 272307 470475 272310
rect 470593 271962 470659 271965
rect 478045 271962 478111 271965
rect 470593 271960 478111 271962
rect 470593 271904 470598 271960
rect 470654 271904 478050 271960
rect 478106 271904 478111 271960
rect 470593 271902 478111 271904
rect 470593 271899 470659 271902
rect 478045 271899 478111 271902
rect 523861 271146 523927 271149
rect 525333 271146 525399 271149
rect 523861 271144 525399 271146
rect 523861 271088 523866 271144
rect 523922 271088 525338 271144
rect 525394 271088 525399 271144
rect 523861 271086 525399 271088
rect 523861 271083 523927 271086
rect 525333 271083 525399 271086
rect 656157 271146 656223 271149
rect 683113 271146 683179 271149
rect 656157 271144 683179 271146
rect 656157 271088 656162 271144
rect 656218 271088 683118 271144
rect 683174 271088 683179 271144
rect 656157 271086 683179 271088
rect 656157 271083 656223 271086
rect 683113 271083 683179 271086
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 530393 270194 530459 270197
rect 534073 270194 534139 270197
rect 530393 270192 534139 270194
rect 530393 270136 530398 270192
rect 530454 270136 534078 270192
rect 534134 270136 534139 270192
rect 530393 270134 534139 270136
rect 530393 270131 530459 270134
rect 534073 270131 534139 270134
rect 41873 270060 41939 270061
rect 41822 270058 41828 270060
rect 41782 269998 41828 270058
rect 41892 270056 41939 270060
rect 41934 270000 41939 270056
rect 41822 269996 41828 269998
rect 41892 269996 41939 270000
rect 41873 269995 41939 269996
rect 537753 269922 537819 269925
rect 538305 269922 538371 269925
rect 537753 269920 538371 269922
rect 537753 269864 537758 269920
rect 537814 269864 538310 269920
rect 538366 269864 538371 269920
rect 537753 269862 538371 269864
rect 537753 269859 537819 269862
rect 538305 269859 538371 269862
rect 665817 268562 665883 268565
rect 676262 268562 676322 268668
rect 683113 268562 683179 268565
rect 665817 268560 676322 268562
rect 665817 268504 665822 268560
rect 665878 268504 676322 268560
rect 665817 268502 676322 268504
rect 683070 268560 683179 268562
rect 683070 268504 683118 268560
rect 683174 268504 683179 268560
rect 665817 268499 665883 268502
rect 683070 268499 683179 268504
rect 683070 268260 683130 268499
rect 674373 267882 674439 267885
rect 674373 267880 676292 267882
rect 674373 267824 674378 267880
rect 674434 267824 676292 267880
rect 674373 267822 676292 267824
rect 674373 267819 674439 267822
rect 673361 267474 673427 267477
rect 673361 267472 676292 267474
rect 673361 267416 673366 267472
rect 673422 267416 676292 267472
rect 673361 267414 676292 267416
rect 673361 267411 673427 267414
rect 40677 267066 40743 267069
rect 63125 267066 63191 267069
rect 40677 267064 63191 267066
rect 40677 267008 40682 267064
rect 40738 267008 63130 267064
rect 63186 267008 63191 267064
rect 40677 267006 63191 267008
rect 40677 267003 40743 267006
rect 63125 267003 63191 267006
rect 673913 267066 673979 267069
rect 673913 267064 676292 267066
rect 673913 267008 673918 267064
rect 673974 267008 676292 267064
rect 673913 267006 676292 267008
rect 673913 267003 673979 267006
rect 673177 266658 673243 266661
rect 673177 266656 676292 266658
rect 673177 266600 673182 266656
rect 673238 266600 676292 266656
rect 673177 266598 676292 266600
rect 673177 266595 673243 266598
rect 42149 266250 42215 266253
rect 54477 266250 54543 266253
rect 42149 266248 54543 266250
rect 42149 266192 42154 266248
rect 42210 266192 54482 266248
rect 54538 266192 54543 266248
rect 42149 266190 54543 266192
rect 42149 266187 42215 266190
rect 54477 266187 54543 266190
rect 673545 266250 673611 266253
rect 673545 266248 676292 266250
rect 673545 266192 673550 266248
rect 673606 266192 676292 266248
rect 673545 266190 676292 266192
rect 673545 266187 673611 266190
rect 675477 265842 675543 265845
rect 675477 265840 676292 265842
rect 675477 265784 675482 265840
rect 675538 265784 676292 265840
rect 675477 265782 676292 265784
rect 675477 265779 675543 265782
rect 673729 265434 673795 265437
rect 673729 265432 676292 265434
rect 673729 265376 673734 265432
rect 673790 265376 676292 265432
rect 673729 265374 676292 265376
rect 673729 265371 673795 265374
rect 674189 265026 674255 265029
rect 674189 265024 676292 265026
rect 674189 264968 674194 265024
rect 674250 264968 676292 265024
rect 674189 264966 676292 264968
rect 674189 264963 674255 264966
rect 674465 264618 674531 264621
rect 674465 264616 676292 264618
rect 674465 264560 674470 264616
rect 674526 264560 676292 264616
rect 674465 264558 676292 264560
rect 674465 264555 674531 264558
rect 674966 264148 674972 264212
rect 675036 264210 675042 264212
rect 675036 264150 676292 264210
rect 675036 264148 675042 264150
rect 676070 263604 676076 263668
rect 676140 263666 676146 263668
rect 676262 263666 676322 263772
rect 676140 263606 676322 263666
rect 676140 263604 676146 263606
rect 681046 263261 681106 263364
rect 680997 263256 681106 263261
rect 680997 263200 681002 263256
rect 681058 263200 681106 263256
rect 680997 263198 681106 263200
rect 680997 263195 681063 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 674281 262578 674347 262581
rect 674281 262576 676292 262578
rect 674281 262520 674286 262576
rect 674342 262520 676292 262576
rect 674281 262518 676292 262520
rect 674281 262515 674347 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671153 262170 671219 262173
rect 671153 262168 676292 262170
rect 671153 262112 671158 262168
rect 671214 262112 676292 262168
rect 671153 262110 676292 262112
rect 671153 262107 671219 262110
rect 676814 261628 676874 261732
rect 676806 261564 676812 261628
rect 676876 261564 676882 261628
rect 670417 261354 670483 261357
rect 670417 261352 676292 261354
rect 670417 261296 670422 261352
rect 670478 261296 676292 261352
rect 670417 261294 676292 261296
rect 670417 261291 670483 261294
rect 671797 260946 671863 260949
rect 671797 260944 676292 260946
rect 671797 260888 671802 260944
rect 671858 260888 676292 260944
rect 671797 260886 676292 260888
rect 671797 260883 671863 260886
rect 673361 260538 673427 260541
rect 673361 260536 676292 260538
rect 673361 260480 673366 260536
rect 673422 260480 676292 260536
rect 673361 260478 676292 260480
rect 673361 260475 673427 260478
rect 554313 259994 554379 259997
rect 676998 259996 677058 260100
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 676990 259932 676996 259996
rect 677060 259932 677066 259996
rect 670233 259722 670299 259725
rect 670233 259720 676292 259722
rect 670233 259664 670238 259720
rect 670294 259664 676292 259720
rect 670233 259662 676292 259664
rect 670233 259659 670299 259662
rect 674097 259314 674163 259317
rect 674097 259312 676292 259314
rect 674097 259256 674102 259312
rect 674158 259256 676292 259312
rect 674097 259254 676292 259256
rect 674097 259251 674163 259254
rect 673177 258906 673243 258909
rect 673177 258904 676292 258906
rect 673177 258848 673182 258904
rect 673238 258848 676292 258904
rect 673177 258846 676292 258848
rect 673177 258843 673243 258846
rect 671429 258498 671495 258501
rect 671429 258496 676292 258498
rect 671429 258440 671434 258496
rect 671490 258440 676292 258496
rect 671429 258438 676292 258440
rect 671429 258435 671495 258438
rect 46197 258090 46263 258093
rect 41492 258088 46263 258090
rect 41492 258032 46202 258088
rect 46258 258032 46263 258088
rect 41492 258030 46263 258032
rect 46197 258027 46263 258030
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 41462 257546 41522 257652
rect 683070 257549 683130 258060
rect 41462 257486 51090 257546
rect 35758 257141 35818 257244
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 44357 256866 44423 256869
rect 41492 256864 44423 256866
rect 41492 256808 44362 256864
rect 44418 256808 44423 256864
rect 41492 256806 44423 256808
rect 44357 256803 44423 256806
rect 51030 256730 51090 257486
rect 683021 257544 683130 257549
rect 683021 257488 683026 257544
rect 683082 257488 683130 257544
rect 683021 257486 683130 257488
rect 683021 257483 683087 257486
rect 676262 257141 676322 257244
rect 676213 257136 676322 257141
rect 676213 257080 676218 257136
rect 676274 257080 676322 257136
rect 676213 257078 676322 257080
rect 676213 257075 676279 257078
rect 59997 256730 60063 256733
rect 51030 256728 60063 256730
rect 51030 256672 60002 256728
rect 60058 256672 60063 256728
rect 51030 256670 60063 256672
rect 59997 256667 60063 256670
rect 650637 256730 650703 256733
rect 676262 256730 676322 256836
rect 650637 256728 676322 256730
rect 650637 256672 650642 256728
rect 650698 256672 676322 256728
rect 650637 256670 676322 256672
rect 650637 256667 650703 256670
rect 44633 256458 44699 256461
rect 41492 256456 44699 256458
rect 41492 256400 44638 256456
rect 44694 256400 44699 256456
rect 41492 256398 44699 256400
rect 44633 256395 44699 256398
rect 671981 256458 672047 256461
rect 676213 256458 676279 256461
rect 671981 256456 676279 256458
rect 671981 256400 671986 256456
rect 672042 256400 676218 256456
rect 676274 256400 676279 256456
rect 671981 256398 676279 256400
rect 671981 256395 672047 256398
rect 676213 256395 676279 256398
rect 35758 255917 35818 256020
rect 35758 255912 35867 255917
rect 35758 255856 35806 255912
rect 35862 255856 35867 255912
rect 35758 255854 35867 255856
rect 35801 255851 35867 255854
rect 39757 255914 39823 255917
rect 42793 255914 42859 255917
rect 39757 255912 42859 255914
rect 39757 255856 39762 255912
rect 39818 255856 42798 255912
rect 42854 255856 42859 255912
rect 39757 255854 42859 255856
rect 39757 255851 39823 255854
rect 42793 255851 42859 255854
rect 45553 255642 45619 255645
rect 553485 255642 553551 255645
rect 41492 255640 45619 255642
rect 41492 255584 45558 255640
rect 45614 255584 45619 255640
rect 41492 255582 45619 255584
rect 552460 255640 553551 255642
rect 552460 255584 553490 255640
rect 553546 255584 553551 255640
rect 552460 255582 553551 255584
rect 45553 255579 45619 255582
rect 553485 255579 553551 255582
rect 674833 255370 674899 255373
rect 675845 255370 675911 255373
rect 674833 255368 675911 255370
rect 674833 255312 674838 255368
rect 674894 255312 675850 255368
rect 675906 255312 675911 255368
rect 674833 255310 675911 255312
rect 674833 255307 674899 255310
rect 675845 255307 675911 255310
rect 44817 255234 44883 255237
rect 41492 255232 44883 255234
rect 41492 255176 44822 255232
rect 44878 255176 44883 255232
rect 41492 255174 44883 255176
rect 44817 255171 44883 255174
rect 44265 254826 44331 254829
rect 41492 254824 44331 254826
rect 41492 254768 44270 254824
rect 44326 254768 44331 254824
rect 41492 254766 44331 254768
rect 44265 254763 44331 254766
rect 44081 254554 44147 254557
rect 41462 254552 44147 254554
rect 41462 254496 44086 254552
rect 44142 254496 44147 254552
rect 41462 254494 44147 254496
rect 41462 254388 41522 254494
rect 44081 254491 44147 254494
rect 35758 253877 35818 253980
rect 35758 253872 35867 253877
rect 35758 253816 35806 253872
rect 35862 253816 35867 253872
rect 35758 253814 35867 253816
rect 35801 253811 35867 253814
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554405 253466 554471 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35617 253403 35683 253406
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 39205 253058 39271 253061
rect 42793 253058 42859 253061
rect 39205 253056 42859 253058
rect 39205 253000 39210 253056
rect 39266 253000 42798 253056
rect 42854 253000 42859 253056
rect 39205 252998 42859 253000
rect 39205 252995 39271 252998
rect 42793 252995 42859 252998
rect 44817 252786 44883 252789
rect 41492 252784 44883 252786
rect 41492 252728 44822 252784
rect 44878 252728 44883 252784
rect 41492 252726 44883 252728
rect 44817 252723 44883 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 40309 252242 40375 252245
rect 42977 252242 43043 252245
rect 40309 252240 43043 252242
rect 40309 252184 40314 252240
rect 40370 252184 42982 252240
rect 43038 252184 43043 252240
rect 40309 252182 43043 252184
rect 40309 252179 40375 252182
rect 42977 252179 43043 252182
rect 44449 251970 44515 251973
rect 41492 251968 44515 251970
rect 41492 251912 44454 251968
rect 44510 251912 44515 251968
rect 41492 251910 44515 251912
rect 44449 251907 44515 251910
rect 45185 251562 45251 251565
rect 41492 251560 45251 251562
rect 41492 251504 45190 251560
rect 45246 251504 45251 251560
rect 41492 251502 45251 251504
rect 45185 251499 45251 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 45921 251154 45987 251157
rect 41492 251152 45987 251154
rect 41492 251096 45926 251152
rect 45982 251096 45987 251152
rect 41492 251094 45987 251096
rect 45921 251091 45987 251094
rect 670969 250882 671035 250885
rect 675477 250882 675543 250885
rect 670969 250880 675543 250882
rect 670969 250824 670974 250880
rect 671030 250824 675482 250880
rect 675538 250824 675543 250880
rect 670969 250822 675543 250824
rect 670969 250819 671035 250822
rect 675477 250819 675543 250822
rect 35758 250613 35818 250716
rect 35758 250608 35867 250613
rect 35758 250552 35806 250608
rect 35862 250552 35867 250608
rect 35758 250550 35867 250552
rect 35801 250547 35867 250550
rect 40542 250204 40602 250308
rect 40534 250140 40540 250204
rect 40604 250140 40610 250204
rect 675753 250202 675819 250205
rect 676806 250202 676812 250204
rect 675753 250200 676812 250202
rect 675753 250144 675758 250200
rect 675814 250144 676812 250200
rect 675753 250142 676812 250144
rect 675753 250139 675819 250142
rect 676806 250140 676812 250142
rect 676876 250140 676882 250204
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 674966 249732 674972 249796
rect 675036 249732 675042 249796
rect 674974 249522 675034 249732
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 675477 249522 675543 249525
rect 674974 249520 675543 249522
rect 35758 249389 35818 249492
rect 674974 249464 675482 249520
rect 675538 249464 675543 249520
rect 674974 249462 675543 249464
rect 675477 249459 675543 249462
rect 35758 249384 35867 249389
rect 35758 249328 35806 249384
rect 35862 249328 35867 249384
rect 35758 249326 35867 249328
rect 35801 249323 35867 249326
rect 39665 249386 39731 249389
rect 43069 249386 43135 249389
rect 39665 249384 43135 249386
rect 39665 249328 39670 249384
rect 39726 249328 43074 249384
rect 43130 249328 43135 249384
rect 39665 249326 43135 249328
rect 39665 249323 39731 249326
rect 43069 249323 43135 249326
rect 45001 249114 45067 249117
rect 554037 249114 554103 249117
rect 41492 249112 45067 249114
rect 41492 249056 45006 249112
rect 45062 249056 45067 249112
rect 41492 249054 45067 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 45001 249051 45067 249054
rect 554037 249051 554103 249054
rect 45737 248706 45803 248709
rect 41492 248704 45803 248706
rect 41492 248648 45742 248704
rect 45798 248648 45803 248704
rect 41492 248646 45803 248648
rect 45737 248643 45803 248646
rect 676078 248434 676138 249596
rect 675526 248374 676138 248434
rect 46105 248298 46171 248301
rect 41492 248296 46171 248298
rect 41492 248240 46110 248296
rect 46166 248240 46171 248296
rect 41492 248238 46171 248240
rect 46105 248235 46171 248238
rect 664437 248162 664503 248165
rect 670969 248162 671035 248165
rect 664437 248160 671035 248162
rect 664437 248104 664442 248160
rect 664498 248104 670974 248160
rect 671030 248104 671035 248160
rect 664437 248102 671035 248104
rect 664437 248099 664503 248102
rect 670969 248099 671035 248102
rect 674833 247890 674899 247893
rect 675526 247890 675586 248374
rect 674833 247888 675586 247890
rect 35574 247757 35634 247860
rect 674833 247832 674838 247888
rect 674894 247832 675586 247888
rect 674833 247830 675586 247832
rect 674833 247827 674899 247830
rect 35574 247752 35683 247757
rect 35574 247696 35622 247752
rect 35678 247696 35683 247752
rect 35574 247694 35683 247696
rect 35617 247691 35683 247694
rect 41505 247754 41571 247757
rect 43805 247754 43871 247757
rect 41505 247752 43871 247754
rect 41505 247696 41510 247752
rect 41566 247696 43810 247752
rect 43866 247696 43871 247752
rect 41505 247694 43871 247696
rect 41505 247691 41571 247694
rect 43805 247691 43871 247694
rect 49141 247482 49207 247485
rect 41492 247480 49207 247482
rect 41492 247424 49146 247480
rect 49202 247424 49207 247480
rect 41492 247422 49207 247424
rect 49141 247419 49207 247422
rect 670417 247074 670483 247077
rect 675293 247074 675359 247077
rect 670417 247072 675359 247074
rect 35758 246941 35818 247044
rect 670417 247016 670422 247072
rect 670478 247016 675298 247072
rect 675354 247016 675359 247072
rect 670417 247014 675359 247016
rect 670417 247011 670483 247014
rect 675293 247011 675359 247014
rect 35758 246936 35867 246941
rect 553853 246938 553919 246941
rect 35758 246880 35806 246936
rect 35862 246880 35867 246936
rect 35758 246878 35867 246880
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 35801 246875 35867 246878
rect 553853 246875 553919 246878
rect 47577 246666 47643 246669
rect 41492 246664 47643 246666
rect 41492 246608 47582 246664
rect 47638 246608 47643 246664
rect 41492 246606 47643 246608
rect 47577 246603 47643 246606
rect 671797 246666 671863 246669
rect 675293 246666 675359 246669
rect 671797 246664 675359 246666
rect 671797 246608 671802 246664
rect 671858 246608 675298 246664
rect 675354 246608 675359 246664
rect 671797 246606 675359 246608
rect 671797 246603 671863 246606
rect 675293 246603 675359 246606
rect 670233 245714 670299 245717
rect 675293 245714 675359 245717
rect 670233 245712 675359 245714
rect 670233 245656 670238 245712
rect 670294 245656 675298 245712
rect 675354 245656 675359 245712
rect 670233 245654 675359 245656
rect 670233 245651 670299 245654
rect 675293 245651 675359 245654
rect 39849 245578 39915 245581
rect 43621 245578 43687 245581
rect 39849 245576 43687 245578
rect 39849 245520 39854 245576
rect 39910 245520 43626 245576
rect 43682 245520 43687 245576
rect 39849 245518 43687 245520
rect 39849 245515 39915 245518
rect 43621 245515 43687 245518
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 674281 243674 674347 243677
rect 675109 243674 675175 243677
rect 674281 243672 675175 243674
rect 674281 243616 674286 243672
rect 674342 243616 675114 243672
rect 675170 243616 675175 243672
rect 674281 243614 675175 243616
rect 674281 243611 674347 243614
rect 675109 243611 675175 243614
rect 674189 242858 674255 242861
rect 675109 242858 675175 242861
rect 674189 242856 675175 242858
rect 674189 242800 674194 242856
rect 674250 242800 675114 242856
rect 675170 242800 675175 242856
rect 674189 242798 675175 242800
rect 674189 242795 674255 242798
rect 675109 242795 675175 242798
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 675753 242314 675819 242317
rect 676990 242314 676996 242316
rect 675753 242312 676996 242314
rect 675753 242256 675758 242312
rect 675814 242256 676996 242312
rect 675753 242254 676996 242256
rect 675753 242251 675819 242254
rect 676990 242252 676996 242254
rect 677060 242252 677066 242316
rect 673729 242042 673795 242045
rect 676806 242042 676812 242044
rect 673729 242040 676812 242042
rect 673729 241984 673734 242040
rect 673790 241984 676812 242040
rect 673729 241982 676812 241984
rect 673729 241979 673795 241982
rect 676806 241980 676812 241982
rect 676876 241980 676882 242044
rect 673545 241770 673611 241773
rect 674966 241770 674972 241772
rect 673545 241768 674972 241770
rect 673545 241712 673550 241768
rect 673606 241712 674972 241768
rect 673545 241710 674972 241712
rect 673545 241707 673611 241710
rect 674966 241708 674972 241710
rect 675036 241708 675042 241772
rect 673177 241498 673243 241501
rect 675109 241498 675175 241501
rect 673177 241496 675175 241498
rect 673177 241440 673182 241496
rect 673238 241440 675114 241496
rect 675170 241440 675175 241496
rect 673177 241438 675175 241440
rect 673177 241435 673243 241438
rect 675109 241435 675175 241438
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 673361 240274 673427 240277
rect 675109 240274 675175 240277
rect 673361 240272 675175 240274
rect 673361 240216 673366 240272
rect 673422 240216 675114 240272
rect 675170 240216 675175 240272
rect 673361 240214 675175 240216
rect 673361 240211 673427 240214
rect 675109 240211 675175 240214
rect 42057 240138 42123 240141
rect 45185 240138 45251 240141
rect 42057 240136 45251 240138
rect 42057 240080 42062 240136
rect 42118 240080 45190 240136
rect 45246 240080 45251 240136
rect 42057 240078 45251 240080
rect 42057 240075 42123 240078
rect 45185 240075 45251 240078
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42425 237418 42491 237421
rect 42076 237416 42491 237418
rect 42076 237360 42430 237416
rect 42486 237360 42491 237416
rect 42076 237358 42491 237360
rect 42076 237356 42082 237358
rect 42425 237355 42491 237358
rect 40718 236540 40724 236604
rect 40788 236602 40794 236604
rect 41781 236602 41847 236605
rect 40788 236600 41847 236602
rect 40788 236544 41786 236600
rect 41842 236544 41847 236600
rect 40788 236542 41847 236544
rect 40788 236540 40794 236542
rect 41781 236539 41847 236542
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 42425 235922 42491 235925
rect 46105 235922 46171 235925
rect 42425 235920 46171 235922
rect 42425 235864 42430 235920
rect 42486 235864 46110 235920
rect 46166 235864 46171 235920
rect 42425 235862 46171 235864
rect 42425 235859 42491 235862
rect 46105 235859 46171 235862
rect 674465 235242 674531 235245
rect 675845 235242 675911 235245
rect 674465 235240 675911 235242
rect 674465 235184 674470 235240
rect 674526 235184 675850 235240
rect 675906 235184 675911 235240
rect 674465 235182 675911 235184
rect 674465 235179 674531 235182
rect 675845 235179 675911 235182
rect 673637 234834 673703 234837
rect 675385 234834 675451 234837
rect 673637 234832 675451 234834
rect 673637 234776 673642 234832
rect 673698 234776 675390 234832
rect 675446 234776 675451 234832
rect 673637 234774 675451 234776
rect 673637 234771 673703 234774
rect 675385 234771 675451 234774
rect 42425 234562 42491 234565
rect 43805 234562 43871 234565
rect 42425 234560 43871 234562
rect 42425 234504 42430 234560
rect 42486 234504 43810 234560
rect 43866 234504 43871 234560
rect 42425 234502 43871 234504
rect 42425 234499 42491 234502
rect 43805 234499 43871 234502
rect 669773 234426 669839 234429
rect 673269 234426 673335 234429
rect 669773 234424 673335 234426
rect 669773 234368 669778 234424
rect 669834 234368 673274 234424
rect 673330 234368 673335 234424
rect 669773 234366 673335 234368
rect 669773 234363 669839 234366
rect 673269 234363 673335 234366
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 672165 233746 672231 233749
rect 675845 233746 675911 233749
rect 672165 233744 675911 233746
rect 672165 233688 672170 233744
rect 672226 233688 675850 233744
rect 675906 233688 675911 233744
rect 672165 233686 675911 233688
rect 672165 233683 672231 233686
rect 675845 233683 675911 233686
rect 42149 233338 42215 233341
rect 44449 233338 44515 233341
rect 42149 233336 44515 233338
rect 42149 233280 42154 233336
rect 42210 233280 44454 233336
rect 44510 233280 44515 233336
rect 42149 233278 44515 233280
rect 42149 233275 42215 233278
rect 44449 233275 44515 233278
rect 42425 232658 42491 232661
rect 45737 232658 45803 232661
rect 42425 232656 45803 232658
rect 42425 232600 42430 232656
rect 42486 232600 45742 232656
rect 45798 232600 45803 232656
rect 42425 232598 45803 232600
rect 42425 232595 42491 232598
rect 45737 232595 45803 232598
rect 670785 232522 670851 232525
rect 675845 232522 675911 232525
rect 670785 232520 675911 232522
rect 670785 232464 670790 232520
rect 670846 232464 675850 232520
rect 675906 232464 675911 232520
rect 670785 232462 675911 232464
rect 670785 232459 670851 232462
rect 675845 232459 675911 232462
rect 42425 231842 42491 231845
rect 45001 231842 45067 231845
rect 42425 231840 45067 231842
rect 42425 231784 42430 231840
rect 42486 231784 45006 231840
rect 45062 231784 45067 231840
rect 42425 231782 45067 231784
rect 42425 231779 42491 231782
rect 45001 231779 45067 231782
rect 670785 231570 670851 231573
rect 675845 231570 675911 231573
rect 670785 231568 675911 231570
rect 670785 231512 670790 231568
rect 670846 231512 675850 231568
rect 675906 231512 675911 231568
rect 670785 231510 675911 231512
rect 670785 231507 670851 231510
rect 675845 231507 675911 231510
rect 40534 230420 40540 230484
rect 40604 230482 40610 230484
rect 41781 230482 41847 230485
rect 40604 230480 41847 230482
rect 40604 230424 41786 230480
rect 41842 230424 41847 230480
rect 40604 230422 41847 230424
rect 40604 230420 40610 230422
rect 41781 230419 41847 230422
rect 142429 230482 142495 230485
rect 144085 230482 144151 230485
rect 142429 230480 144151 230482
rect 142429 230424 142434 230480
rect 142490 230424 144090 230480
rect 144146 230424 144151 230480
rect 142429 230422 144151 230424
rect 142429 230419 142495 230422
rect 144085 230419 144151 230422
rect 665817 230482 665883 230485
rect 673453 230482 673519 230485
rect 665817 230480 673519 230482
rect 665817 230424 665822 230480
rect 665878 230424 673458 230480
rect 673514 230424 673519 230480
rect 665817 230422 673519 230424
rect 665817 230419 665883 230422
rect 673453 230419 673519 230422
rect 674373 230482 674439 230485
rect 676581 230482 676647 230485
rect 674373 230480 676647 230482
rect 674373 230424 674378 230480
rect 674434 230424 676586 230480
rect 676642 230424 676647 230480
rect 674373 230422 676647 230424
rect 674373 230419 674439 230422
rect 676581 230419 676647 230422
rect 674966 230148 674972 230212
rect 675036 230210 675042 230212
rect 676029 230210 676095 230213
rect 675036 230208 676095 230210
rect 675036 230152 676034 230208
rect 676090 230152 676095 230208
rect 675036 230150 676095 230152
rect 675036 230148 675042 230150
rect 676029 230147 676095 230150
rect 156781 229938 156847 229941
rect 157425 229938 157491 229941
rect 156781 229936 157491 229938
rect 156781 229880 156786 229936
rect 156842 229880 157430 229936
rect 157486 229880 157491 229936
rect 156781 229878 157491 229880
rect 156781 229875 156847 229878
rect 157425 229875 157491 229878
rect 147581 229802 147647 229805
rect 147949 229802 148015 229805
rect 147581 229800 148015 229802
rect 147581 229744 147586 229800
rect 147642 229744 147954 229800
rect 148010 229744 148015 229800
rect 147581 229742 148015 229744
rect 147581 229739 147647 229742
rect 147949 229739 148015 229742
rect 652569 229802 652635 229805
rect 674046 229802 674052 229804
rect 652569 229800 674052 229802
rect 652569 229744 652574 229800
rect 652630 229744 674052 229800
rect 652569 229742 674052 229744
rect 652569 229739 652635 229742
rect 674046 229740 674052 229742
rect 674116 229740 674122 229804
rect 143993 229530 144059 229533
rect 145373 229530 145439 229533
rect 143993 229528 145439 229530
rect 143993 229472 143998 229528
rect 144054 229472 145378 229528
rect 145434 229472 145439 229528
rect 143993 229470 145439 229472
rect 143993 229467 144059 229470
rect 145373 229467 145439 229470
rect 665173 229530 665239 229533
rect 674327 229530 674393 229533
rect 665173 229528 674393 229530
rect 665173 229472 665178 229528
rect 665234 229472 674332 229528
rect 674388 229472 674393 229528
rect 665173 229470 674393 229472
rect 665173 229467 665239 229470
rect 674327 229467 674393 229470
rect 146201 229394 146267 229397
rect 147765 229394 147831 229397
rect 159357 229394 159423 229397
rect 146201 229392 147831 229394
rect 146201 229336 146206 229392
rect 146262 229336 147770 229392
rect 147826 229336 147831 229392
rect 146201 229334 147831 229336
rect 146201 229331 146267 229334
rect 147765 229331 147831 229334
rect 154530 229392 159423 229394
rect 154530 229336 159362 229392
rect 159418 229336 159423 229392
rect 154530 229334 159423 229336
rect 150341 229258 150407 229261
rect 154530 229258 154590 229334
rect 159357 229331 159423 229334
rect 150341 229256 154590 229258
rect 150341 229200 150346 229256
rect 150402 229200 154590 229256
rect 150341 229198 154590 229200
rect 166993 229258 167059 229261
rect 167361 229258 167427 229261
rect 674465 229258 674531 229261
rect 166993 229256 167427 229258
rect 166993 229200 166998 229256
rect 167054 229200 167366 229256
rect 167422 229200 167427 229256
rect 166993 229198 167427 229200
rect 150341 229195 150407 229198
rect 166993 229195 167059 229198
rect 167361 229195 167427 229198
rect 663750 229256 674531 229258
rect 663750 229200 674470 229256
rect 674526 229200 674531 229256
rect 663750 229198 674531 229200
rect 663750 229125 663810 229198
rect 674465 229195 674531 229198
rect 140037 229122 140103 229125
rect 147121 229122 147187 229125
rect 140037 229120 147187 229122
rect 140037 229064 140042 229120
rect 140098 229064 147126 229120
rect 147182 229064 147187 229120
rect 140037 229062 147187 229064
rect 140037 229059 140103 229062
rect 147121 229059 147187 229062
rect 202873 229122 202939 229125
rect 205173 229122 205239 229125
rect 202873 229120 205239 229122
rect 202873 229064 202878 229120
rect 202934 229064 205178 229120
rect 205234 229064 205239 229120
rect 202873 229062 205239 229064
rect 202873 229059 202939 229062
rect 205173 229059 205239 229062
rect 663701 229120 663810 229125
rect 663701 229064 663706 229120
rect 663762 229064 663810 229120
rect 663701 229062 663810 229064
rect 663701 229059 663767 229062
rect 41965 228988 42031 228989
rect 41965 228984 42012 228988
rect 42076 228986 42082 228988
rect 166809 228986 166875 228989
rect 167361 228986 167427 228989
rect 41965 228928 41970 228984
rect 41965 228924 42012 228928
rect 42076 228926 42122 228986
rect 166809 228984 167427 228986
rect 166809 228928 166814 228984
rect 166870 228928 167366 228984
rect 167422 228928 167427 228984
rect 166809 228926 167427 228928
rect 42076 228924 42082 228926
rect 41965 228923 42031 228924
rect 166809 228923 166875 228926
rect 167361 228923 167427 228926
rect 156873 228850 156939 228853
rect 157517 228850 157583 228853
rect 156873 228848 157583 228850
rect 156873 228792 156878 228848
rect 156934 228792 157522 228848
rect 157578 228792 157583 228848
rect 156873 228790 157583 228792
rect 156873 228787 156939 228790
rect 157517 228787 157583 228790
rect 173341 228850 173407 228853
rect 174813 228850 174879 228853
rect 173341 228848 174879 228850
rect 173341 228792 173346 228848
rect 173402 228792 174818 228848
rect 174874 228792 174879 228848
rect 173341 228790 174879 228792
rect 173341 228787 173407 228790
rect 174813 228787 174879 228790
rect 673177 228578 673243 228581
rect 676213 228578 676279 228581
rect 673177 228576 676279 228578
rect 673177 228520 673182 228576
rect 673238 228520 676218 228576
rect 676274 228520 676279 228576
rect 673177 228518 676279 228520
rect 673177 228515 673243 228518
rect 676213 228515 676279 228518
rect 139301 228306 139367 228309
rect 142981 228306 143047 228309
rect 139301 228304 143047 228306
rect 139301 228248 139306 228304
rect 139362 228248 142986 228304
rect 143042 228248 143047 228304
rect 139301 228246 143047 228248
rect 139301 228243 139367 228246
rect 142981 228243 143047 228246
rect 160001 228170 160067 228173
rect 166809 228170 166875 228173
rect 160001 228168 166875 228170
rect 160001 228112 160006 228168
rect 160062 228112 166814 228168
rect 166870 228112 166875 228168
rect 160001 228110 166875 228112
rect 160001 228107 160067 228110
rect 166809 228107 166875 228110
rect 171225 227626 171291 227629
rect 172145 227626 172211 227629
rect 171225 227624 172211 227626
rect 171225 227568 171230 227624
rect 171286 227568 172150 227624
rect 172206 227568 172211 227624
rect 171225 227566 172211 227568
rect 171225 227563 171291 227566
rect 172145 227563 172211 227566
rect 156873 227490 156939 227493
rect 166533 227490 166599 227493
rect 156873 227488 166599 227490
rect 156873 227432 156878 227488
rect 156934 227432 166538 227488
rect 166594 227432 166599 227488
rect 156873 227430 166599 227432
rect 156873 227427 156939 227430
rect 166533 227427 166599 227430
rect 219433 227490 219499 227493
rect 220445 227490 220511 227493
rect 219433 227488 220511 227490
rect 219433 227432 219438 227488
rect 219494 227432 220450 227488
rect 220506 227432 220511 227488
rect 219433 227430 220511 227432
rect 219433 227427 219499 227430
rect 220445 227427 220511 227430
rect 169477 227354 169543 227357
rect 171685 227354 171751 227357
rect 169477 227352 171751 227354
rect 169477 227296 169482 227352
rect 169538 227296 171690 227352
rect 171746 227296 171751 227352
rect 169477 227294 171751 227296
rect 169477 227291 169543 227294
rect 171685 227291 171751 227294
rect 672942 227082 672948 227084
rect 663750 227022 672948 227082
rect 652385 226946 652451 226949
rect 663750 226946 663810 227022
rect 672942 227020 672948 227022
rect 673012 227020 673018 227084
rect 673361 227082 673427 227085
rect 677041 227082 677107 227085
rect 673361 227080 677107 227082
rect 673361 227024 673366 227080
rect 673422 227024 677046 227080
rect 677102 227024 677107 227080
rect 673361 227022 677107 227024
rect 673361 227019 673427 227022
rect 677041 227019 677107 227022
rect 652385 226944 663810 226946
rect 652385 226888 652390 226944
rect 652446 226888 663810 226944
rect 652385 226886 663810 226888
rect 652385 226883 652451 226886
rect 673545 226810 673611 226813
rect 674281 226810 674347 226813
rect 673545 226808 674347 226810
rect 673545 226752 673550 226808
rect 673606 226752 674286 226808
rect 674342 226752 674347 226808
rect 673545 226750 674347 226752
rect 673545 226747 673611 226750
rect 674281 226747 674347 226750
rect 654777 226402 654843 226405
rect 670785 226402 670851 226405
rect 654777 226400 670851 226402
rect 654777 226344 654782 226400
rect 654838 226344 670790 226400
rect 670846 226344 670851 226400
rect 654777 226342 670851 226344
rect 654777 226339 654843 226342
rect 670785 226339 670851 226342
rect 672165 226402 672231 226405
rect 675017 226402 675083 226405
rect 672165 226400 675083 226402
rect 672165 226344 672170 226400
rect 672226 226344 675022 226400
rect 675078 226344 675083 226400
rect 672165 226342 675083 226344
rect 672165 226339 672231 226342
rect 675017 226339 675083 226342
rect 42241 226130 42307 226133
rect 44817 226130 44883 226133
rect 42241 226128 44883 226130
rect 42241 226072 42246 226128
rect 42302 226072 44822 226128
rect 44878 226072 44883 226128
rect 42241 226070 44883 226072
rect 42241 226067 42307 226070
rect 44817 226067 44883 226070
rect 141141 226130 141207 226133
rect 145189 226130 145255 226133
rect 141141 226128 145255 226130
rect 141141 226072 141146 226128
rect 141202 226072 145194 226128
rect 145250 226072 145255 226128
rect 141141 226070 145255 226072
rect 141141 226067 141207 226070
rect 145189 226067 145255 226070
rect 672257 225858 672323 225861
rect 674833 225858 674899 225861
rect 672257 225856 674899 225858
rect 672257 225800 672262 225856
rect 672318 225800 674838 225856
rect 674894 225800 674899 225856
rect 672257 225798 674899 225800
rect 672257 225795 672323 225798
rect 674833 225795 674899 225798
rect 42609 225586 42675 225589
rect 62941 225586 63007 225589
rect 42609 225584 63007 225586
rect 42609 225528 42614 225584
rect 42670 225528 62946 225584
rect 63002 225528 63007 225584
rect 42609 225526 63007 225528
rect 42609 225523 42675 225526
rect 62941 225523 63007 225526
rect 652017 225586 652083 225589
rect 671245 225586 671311 225589
rect 672257 225586 672323 225589
rect 652017 225584 671311 225586
rect 652017 225528 652022 225584
rect 652078 225528 671250 225584
rect 671306 225528 671311 225584
rect 652017 225526 671311 225528
rect 652017 225523 652083 225526
rect 671245 225523 671311 225526
rect 671478 225584 672323 225586
rect 671478 225528 672262 225584
rect 672318 225528 672323 225584
rect 671478 225526 672323 225528
rect 656157 225314 656223 225317
rect 671478 225314 671538 225526
rect 672257 225523 672323 225526
rect 656157 225312 671538 225314
rect 656157 225256 656162 225312
rect 656218 225256 671538 225312
rect 656157 225254 671538 225256
rect 672149 225314 672215 225317
rect 675201 225314 675267 225317
rect 672149 225312 675267 225314
rect 672149 225256 672154 225312
rect 672210 225256 675206 225312
rect 675262 225256 675267 225312
rect 672149 225254 675267 225256
rect 656157 225251 656223 225254
rect 672149 225251 672215 225254
rect 675201 225251 675267 225254
rect 653397 225042 653463 225045
rect 670785 225042 670851 225045
rect 653397 225040 670851 225042
rect 653397 224984 653402 225040
rect 653458 224984 670790 225040
rect 670846 224984 670851 225040
rect 653397 224982 670851 224984
rect 653397 224979 653463 224982
rect 670785 224979 670851 224982
rect 42425 224906 42491 224909
rect 45921 224906 45987 224909
rect 42425 224904 45987 224906
rect 42425 224848 42430 224904
rect 42486 224848 45926 224904
rect 45982 224848 45987 224904
rect 42425 224846 45987 224848
rect 42425 224843 42491 224846
rect 45921 224843 45987 224846
rect 555785 224498 555851 224501
rect 561673 224498 561739 224501
rect 555785 224496 561739 224498
rect 555785 224440 555790 224496
rect 555846 224440 561678 224496
rect 561734 224440 561739 224496
rect 555785 224438 561739 224440
rect 555785 224435 555851 224438
rect 561673 224435 561739 224438
rect 562133 224362 562199 224365
rect 563237 224362 563303 224365
rect 562133 224360 563303 224362
rect 562133 224304 562138 224360
rect 562194 224304 563242 224360
rect 563298 224304 563303 224360
rect 562133 224302 563303 224304
rect 562133 224299 562199 224302
rect 563237 224299 563303 224302
rect 657537 223954 657603 223957
rect 670785 223954 670851 223957
rect 657537 223952 670851 223954
rect 657537 223896 657542 223952
rect 657598 223896 670790 223952
rect 670846 223896 670851 223952
rect 657537 223894 670851 223896
rect 657537 223891 657603 223894
rect 670785 223891 670851 223894
rect 678237 223818 678303 223821
rect 678237 223816 678346 223818
rect 678237 223760 678242 223816
rect 678298 223760 678346 223816
rect 678237 223755 678346 223760
rect 664437 223682 664503 223685
rect 667841 223682 667907 223685
rect 664437 223680 667907 223682
rect 664437 223624 664442 223680
rect 664498 223624 667846 223680
rect 667902 223624 667907 223680
rect 664437 223622 667907 223624
rect 664437 223619 664503 223622
rect 667841 223619 667907 223622
rect 673494 223620 673500 223684
rect 673564 223682 673570 223684
rect 674649 223682 674715 223685
rect 673564 223680 674715 223682
rect 673564 223624 674654 223680
rect 674710 223624 674715 223680
rect 673564 223622 674715 223624
rect 673564 223620 673570 223622
rect 674649 223619 674715 223622
rect 42149 223546 42215 223549
rect 55857 223546 55923 223549
rect 42149 223544 55923 223546
rect 42149 223488 42154 223544
rect 42210 223488 55862 223544
rect 55918 223488 55923 223544
rect 678286 223516 678346 223755
rect 42149 223486 55923 223488
rect 42149 223483 42215 223486
rect 55857 223483 55923 223486
rect 147673 223410 147739 223413
rect 152273 223410 152339 223413
rect 147673 223408 152339 223410
rect 147673 223352 147678 223408
rect 147734 223352 152278 223408
rect 152334 223352 152339 223408
rect 147673 223350 152339 223352
rect 147673 223347 147739 223350
rect 152273 223347 152339 223350
rect 157241 223410 157307 223413
rect 157425 223410 157491 223413
rect 157241 223408 157491 223410
rect 157241 223352 157246 223408
rect 157302 223352 157430 223408
rect 157486 223352 157491 223408
rect 157241 223350 157491 223352
rect 157241 223347 157307 223350
rect 157425 223347 157491 223350
rect 670785 223410 670851 223413
rect 673453 223410 673519 223413
rect 670785 223408 673519 223410
rect 670785 223352 670790 223408
rect 670846 223352 673458 223408
rect 673514 223352 673519 223408
rect 670785 223350 673519 223352
rect 670785 223347 670851 223350
rect 673453 223347 673519 223350
rect 683573 223138 683639 223141
rect 683573 223136 683652 223138
rect 683573 223080 683578 223136
rect 683634 223080 683652 223136
rect 683573 223078 683652 223080
rect 683573 223075 683639 223078
rect 147305 223002 147371 223005
rect 147765 223002 147831 223005
rect 147305 223000 147831 223002
rect 147305 222944 147310 223000
rect 147366 222944 147770 223000
rect 147826 222944 147831 223000
rect 147305 222942 147831 222944
rect 147305 222939 147371 222942
rect 147765 222939 147831 222942
rect 650637 222866 650703 222869
rect 672993 222866 673059 222869
rect 650637 222864 673059 222866
rect 650637 222808 650642 222864
rect 650698 222808 672998 222864
rect 673054 222808 673059 222864
rect 650637 222806 673059 222808
rect 650637 222803 650703 222806
rect 672993 222803 673059 222806
rect 152181 222730 152247 222733
rect 155125 222730 155191 222733
rect 152181 222728 155191 222730
rect 152181 222672 152186 222728
rect 152242 222672 155130 222728
rect 155186 222672 155191 222728
rect 152181 222670 155191 222672
rect 152181 222667 152247 222670
rect 155125 222667 155191 222670
rect 683205 222730 683271 222733
rect 683205 222728 683284 222730
rect 683205 222672 683210 222728
rect 683266 222672 683284 222728
rect 683205 222670 683284 222672
rect 683205 222667 683271 222670
rect 659101 222594 659167 222597
rect 670785 222594 670851 222597
rect 659101 222592 670851 222594
rect 659101 222536 659106 222592
rect 659162 222536 670790 222592
rect 670846 222536 670851 222592
rect 659101 222534 670851 222536
rect 659101 222531 659167 222534
rect 670785 222531 670851 222534
rect 557993 222458 558059 222461
rect 567009 222458 567075 222461
rect 557993 222456 567075 222458
rect 557993 222400 557998 222456
rect 558054 222400 567014 222456
rect 567070 222400 567075 222456
rect 557993 222398 567075 222400
rect 557993 222395 558059 222398
rect 567009 222395 567075 222398
rect 145925 222322 145991 222325
rect 147121 222322 147187 222325
rect 145925 222320 147187 222322
rect 145925 222264 145930 222320
rect 145986 222264 147126 222320
rect 147182 222264 147187 222320
rect 145925 222262 147187 222264
rect 145925 222259 145991 222262
rect 147121 222259 147187 222262
rect 543181 222322 543247 222325
rect 547689 222322 547755 222325
rect 543181 222320 547755 222322
rect 543181 222264 543186 222320
rect 543242 222264 547694 222320
rect 547750 222264 547755 222320
rect 543181 222262 547755 222264
rect 543181 222259 543247 222262
rect 547689 222259 547755 222262
rect 673913 222322 673979 222325
rect 673913 222320 676292 222322
rect 673913 222264 673918 222320
rect 673974 222264 676292 222320
rect 673913 222262 676292 222264
rect 673913 222259 673979 222262
rect 561673 222188 561739 222189
rect 561622 222124 561628 222188
rect 561692 222186 561739 222188
rect 562685 222186 562751 222189
rect 564801 222186 564867 222189
rect 561692 222184 561784 222186
rect 561734 222128 561784 222184
rect 561692 222126 561784 222128
rect 562685 222184 564867 222186
rect 562685 222128 562690 222184
rect 562746 222128 564806 222184
rect 564862 222128 564867 222184
rect 562685 222126 564867 222128
rect 561692 222124 561739 222126
rect 561673 222123 561739 222124
rect 562685 222123 562751 222126
rect 564801 222123 564867 222126
rect 546953 222050 547019 222053
rect 553853 222050 553919 222053
rect 546953 222048 553919 222050
rect 546953 221992 546958 222048
rect 547014 221992 553858 222048
rect 553914 221992 553919 222048
rect 546953 221990 553919 221992
rect 546953 221987 547019 221990
rect 553853 221987 553919 221990
rect 667565 222050 667631 222053
rect 667565 222048 672826 222050
rect 667565 221992 667570 222048
rect 667626 221992 672826 222048
rect 667565 221990 672826 221992
rect 667565 221987 667631 221990
rect 672766 221914 672826 221990
rect 672766 221854 676292 221914
rect 184657 221778 184723 221781
rect 185761 221778 185827 221781
rect 184657 221776 185827 221778
rect 184657 221720 184662 221776
rect 184718 221720 185766 221776
rect 185822 221720 185827 221776
rect 184657 221718 185827 221720
rect 184657 221715 184723 221718
rect 185761 221715 185827 221718
rect 540881 221778 540947 221781
rect 546769 221778 546835 221781
rect 540881 221776 546835 221778
rect 540881 221720 540886 221776
rect 540942 221720 546774 221776
rect 546830 221720 546835 221776
rect 540881 221718 546835 221720
rect 540881 221715 540947 221718
rect 546769 221715 546835 221718
rect 547689 221778 547755 221781
rect 549069 221778 549135 221781
rect 547689 221776 549135 221778
rect 547689 221720 547694 221776
rect 547750 221720 549074 221776
rect 549130 221720 549135 221776
rect 547689 221718 549135 221720
rect 547689 221715 547755 221718
rect 549069 221715 549135 221718
rect 553485 221778 553551 221781
rect 557533 221778 557599 221781
rect 553485 221776 557599 221778
rect 553485 221720 553490 221776
rect 553546 221720 557538 221776
rect 557594 221720 557599 221776
rect 553485 221718 557599 221720
rect 553485 221715 553551 221718
rect 557533 221715 557599 221718
rect 559373 221778 559439 221781
rect 561489 221778 561555 221781
rect 559373 221776 561555 221778
rect 559373 221720 559378 221776
rect 559434 221720 561494 221776
rect 561550 221720 561555 221776
rect 559373 221718 561555 221720
rect 559373 221715 559439 221718
rect 561489 221715 561555 221718
rect 564801 221778 564867 221781
rect 569585 221778 569651 221781
rect 564801 221776 569651 221778
rect 564801 221720 564806 221776
rect 564862 221720 569590 221776
rect 569646 221720 569651 221776
rect 564801 221718 569651 221720
rect 564801 221715 564867 221718
rect 569585 221715 569651 221718
rect 651465 221778 651531 221781
rect 671705 221778 671771 221781
rect 651465 221776 671771 221778
rect 651465 221720 651470 221776
rect 651526 221720 671710 221776
rect 671766 221720 671771 221776
rect 651465 221718 671771 221720
rect 651465 221715 651531 221718
rect 671705 221715 671771 221718
rect 158345 221642 158411 221645
rect 164509 221642 164575 221645
rect 158345 221640 164575 221642
rect 158345 221584 158350 221640
rect 158406 221584 164514 221640
rect 164570 221584 164575 221640
rect 158345 221582 164575 221584
rect 158345 221579 158411 221582
rect 164509 221579 164575 221582
rect 513557 221506 513623 221509
rect 599485 221506 599551 221509
rect 513557 221504 599551 221506
rect 513557 221448 513562 221504
rect 513618 221448 599490 221504
rect 599546 221448 599551 221504
rect 513557 221446 599551 221448
rect 513557 221443 513623 221446
rect 599485 221443 599551 221446
rect 649717 221506 649783 221509
rect 674833 221506 674899 221509
rect 649717 221504 674899 221506
rect 649717 221448 649722 221504
rect 649778 221448 674838 221504
rect 674894 221448 674899 221504
rect 649717 221446 674899 221448
rect 649717 221443 649783 221446
rect 674833 221443 674899 221446
rect 676029 221506 676095 221509
rect 676029 221504 676292 221506
rect 676029 221448 676034 221504
rect 676090 221448 676292 221504
rect 676029 221446 676292 221448
rect 676029 221443 676095 221446
rect 176469 221370 176535 221373
rect 177297 221370 177363 221373
rect 176469 221368 177363 221370
rect 176469 221312 176474 221368
rect 176530 221312 177302 221368
rect 177358 221312 177363 221368
rect 176469 221310 177363 221312
rect 176469 221307 176535 221310
rect 177297 221307 177363 221310
rect 520181 221234 520247 221237
rect 618253 221234 618319 221237
rect 520181 221232 618319 221234
rect 520181 221176 520186 221232
rect 520242 221176 618258 221232
rect 618314 221176 618319 221232
rect 520181 221174 618319 221176
rect 520181 221171 520247 221174
rect 618253 221171 618319 221174
rect 667013 221098 667079 221101
rect 667013 221096 676292 221098
rect 667013 221040 667018 221096
rect 667074 221040 676292 221096
rect 667013 221038 676292 221040
rect 667013 221035 667079 221038
rect 149237 220962 149303 220965
rect 156137 220962 156203 220965
rect 149237 220960 156203 220962
rect 149237 220904 149242 220960
rect 149298 220904 156142 220960
rect 156198 220904 156203 220960
rect 149237 220902 156203 220904
rect 149237 220899 149303 220902
rect 156137 220899 156203 220902
rect 166993 220962 167059 220965
rect 175549 220962 175615 220965
rect 166993 220960 175615 220962
rect 166993 220904 166998 220960
rect 167054 220904 175554 220960
rect 175610 220904 175615 220960
rect 166993 220902 175615 220904
rect 166993 220899 167059 220902
rect 175549 220899 175615 220902
rect 497825 220962 497891 220965
rect 498101 220962 498167 220965
rect 631317 220962 631383 220965
rect 497825 220960 631383 220962
rect 497825 220904 497830 220960
rect 497886 220904 498106 220960
rect 498162 220904 631322 220960
rect 631378 220904 631383 220960
rect 497825 220902 631383 220904
rect 497825 220899 497891 220902
rect 498101 220899 498167 220902
rect 631317 220899 631383 220902
rect 176469 220826 176535 220829
rect 179873 220826 179939 220829
rect 176469 220824 179939 220826
rect 176469 220768 176474 220824
rect 176530 220768 179878 220824
rect 179934 220768 179939 220824
rect 176469 220766 179939 220768
rect 176469 220763 176535 220766
rect 179873 220763 179939 220766
rect 144637 220690 144703 220693
rect 150893 220690 150959 220693
rect 144637 220688 150959 220690
rect 144637 220632 144642 220688
rect 144698 220632 150898 220688
rect 150954 220632 150959 220688
rect 144637 220630 150959 220632
rect 144637 220627 144703 220630
rect 150893 220627 150959 220630
rect 562869 220690 562935 220693
rect 576761 220690 576827 220693
rect 562869 220688 576827 220690
rect 562869 220632 562874 220688
rect 562930 220632 576766 220688
rect 576822 220632 576827 220688
rect 562869 220630 576827 220632
rect 562869 220627 562935 220630
rect 576761 220627 576827 220630
rect 675886 220628 675892 220692
rect 675956 220690 675962 220692
rect 675956 220630 676292 220690
rect 675956 220628 675962 220630
rect 675017 220554 675083 220557
rect 663750 220552 675083 220554
rect 663750 220496 675022 220552
rect 675078 220496 675083 220552
rect 663750 220494 675083 220496
rect 140773 220418 140839 220421
rect 142245 220418 142311 220421
rect 140773 220416 142311 220418
rect 140773 220360 140778 220416
rect 140834 220360 142250 220416
rect 142306 220360 142311 220416
rect 140773 220358 142311 220360
rect 140773 220355 140839 220358
rect 142245 220355 142311 220358
rect 160829 220418 160895 220421
rect 166533 220418 166599 220421
rect 160829 220416 166599 220418
rect 160829 220360 160834 220416
rect 160890 220360 166538 220416
rect 166594 220360 166599 220416
rect 160829 220358 166599 220360
rect 160829 220355 160895 220358
rect 166533 220355 166599 220358
rect 565629 220418 565695 220421
rect 567377 220418 567443 220421
rect 565629 220416 567443 220418
rect 565629 220360 565634 220416
rect 565690 220360 567382 220416
rect 567438 220360 567443 220416
rect 565629 220358 567443 220360
rect 565629 220355 565695 220358
rect 567377 220355 567443 220358
rect 567653 220418 567719 220421
rect 568941 220418 569007 220421
rect 567653 220416 569007 220418
rect 567653 220360 567658 220416
rect 567714 220360 568946 220416
rect 569002 220360 569007 220416
rect 567653 220358 569007 220360
rect 567653 220355 567719 220358
rect 568941 220355 569007 220358
rect 644749 220418 644815 220421
rect 663750 220418 663810 220494
rect 675017 220491 675083 220494
rect 644749 220416 663810 220418
rect 644749 220360 644754 220416
rect 644810 220360 663810 220416
rect 644749 220358 663810 220360
rect 644749 220355 644815 220358
rect 166901 220282 166967 220285
rect 167085 220282 167151 220285
rect 166901 220280 167151 220282
rect 166901 220224 166906 220280
rect 166962 220224 167090 220280
rect 167146 220224 167151 220280
rect 166901 220222 167151 220224
rect 166901 220219 166967 220222
rect 167085 220219 167151 220222
rect 573357 220282 573423 220285
rect 582465 220282 582531 220285
rect 573357 220280 582531 220282
rect 573357 220224 573362 220280
rect 573418 220224 582470 220280
rect 582526 220224 582531 220280
rect 573357 220222 582531 220224
rect 573357 220219 573423 220222
rect 582465 220219 582531 220222
rect 673913 220282 673979 220285
rect 673913 220280 676292 220282
rect 673913 220224 673918 220280
rect 673974 220224 676292 220280
rect 673913 220222 676292 220224
rect 673913 220219 673979 220222
rect 180517 220146 180583 220149
rect 185761 220146 185827 220149
rect 180517 220144 185827 220146
rect 180517 220088 180522 220144
rect 180578 220088 185766 220144
rect 185822 220088 185827 220144
rect 180517 220086 185827 220088
rect 180517 220083 180583 220086
rect 185761 220083 185827 220086
rect 551185 220146 551251 220149
rect 552841 220146 552907 220149
rect 551185 220144 552907 220146
rect 551185 220088 551190 220144
rect 551246 220088 552846 220144
rect 552902 220088 552907 220144
rect 551185 220086 552907 220088
rect 551185 220083 551251 220086
rect 552841 220083 552907 220086
rect 566825 220146 566891 220149
rect 567837 220146 567903 220149
rect 566825 220144 567903 220146
rect 566825 220088 566830 220144
rect 566886 220088 567842 220144
rect 567898 220088 567903 220144
rect 566825 220086 567903 220088
rect 566825 220083 566891 220086
rect 567837 220083 567903 220086
rect 653029 220146 653095 220149
rect 668025 220146 668091 220149
rect 653029 220144 668091 220146
rect 653029 220088 653034 220144
rect 653090 220088 668030 220144
rect 668086 220088 668091 220144
rect 653029 220086 668091 220088
rect 653029 220083 653095 220086
rect 668025 220083 668091 220086
rect 576577 220010 576643 220013
rect 581821 220010 581887 220013
rect 576577 220008 581887 220010
rect 576577 219952 576582 220008
rect 576638 219952 581826 220008
rect 581882 219952 581887 220008
rect 576577 219950 581887 219952
rect 576577 219947 576643 219950
rect 581821 219947 581887 219950
rect 683389 219874 683455 219877
rect 683389 219872 683468 219874
rect 683389 219816 683394 219872
rect 683450 219816 683468 219872
rect 683389 219814 683468 219816
rect 683389 219811 683455 219814
rect 141969 219738 142035 219741
rect 144177 219738 144243 219741
rect 141969 219736 144243 219738
rect 141969 219680 141974 219736
rect 142030 219680 144182 219736
rect 144238 219680 144243 219736
rect 141969 219678 144243 219680
rect 141969 219675 142035 219678
rect 144177 219675 144243 219678
rect 202413 219738 202479 219741
rect 203149 219738 203215 219741
rect 611629 219738 611695 219741
rect 202413 219736 203215 219738
rect 202413 219680 202418 219736
rect 202474 219680 203154 219736
rect 203210 219680 203215 219736
rect 202413 219678 203215 219680
rect 202413 219675 202479 219678
rect 203149 219675 203215 219678
rect 489870 219736 611695 219738
rect 489870 219680 611634 219736
rect 611690 219680 611695 219736
rect 489870 219678 611695 219680
rect 195881 219602 195947 219605
rect 196341 219602 196407 219605
rect 195881 219600 196407 219602
rect 195881 219544 195886 219600
rect 195942 219544 196346 219600
rect 196402 219544 196407 219600
rect 195881 219542 196407 219544
rect 195881 219539 195947 219542
rect 196341 219539 196407 219542
rect 486969 219466 487035 219469
rect 489870 219466 489930 219678
rect 611629 219675 611695 219678
rect 486969 219464 489930 219466
rect 486969 219408 486974 219464
rect 487030 219408 489930 219464
rect 486969 219406 489930 219408
rect 515213 219466 515279 219469
rect 617241 219466 617307 219469
rect 515213 219464 617307 219466
rect 515213 219408 515218 219464
rect 515274 219408 617246 219464
rect 617302 219408 617307 219464
rect 515213 219406 617307 219408
rect 486969 219403 487035 219406
rect 515213 219403 515279 219406
rect 617241 219403 617307 219406
rect 667749 219466 667815 219469
rect 667749 219464 676292 219466
rect 667749 219408 667754 219464
rect 667810 219408 676292 219464
rect 667749 219406 676292 219408
rect 667749 219403 667815 219406
rect 552289 219194 552355 219197
rect 556521 219194 556587 219197
rect 552289 219192 556587 219194
rect 552289 219136 552294 219192
rect 552350 219136 556526 219192
rect 556582 219136 556587 219192
rect 552289 219134 556587 219136
rect 552289 219131 552355 219134
rect 556521 219131 556587 219134
rect 561622 219132 561628 219196
rect 561692 219194 561698 219196
rect 562317 219194 562383 219197
rect 561692 219192 562383 219194
rect 561692 219136 562322 219192
rect 562378 219136 562383 219192
rect 561692 219134 562383 219136
rect 561692 219132 561698 219134
rect 562317 219131 562383 219134
rect 569217 219194 569283 219197
rect 572621 219194 572687 219197
rect 569217 219192 572687 219194
rect 569217 219136 569222 219192
rect 569278 219136 572626 219192
rect 572682 219136 572687 219192
rect 569217 219134 572687 219136
rect 569217 219131 569283 219134
rect 572621 219131 572687 219134
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 494697 218922 494763 218925
rect 655421 218922 655487 218925
rect 670785 218922 670851 218925
rect 494697 218920 596190 218922
rect 494697 218864 494702 218920
rect 494758 218864 596190 218920
rect 494697 218862 596190 218864
rect 494697 218859 494763 218862
rect 490373 218650 490439 218653
rect 594793 218650 594859 218653
rect 490373 218648 594859 218650
rect 490373 218592 490378 218648
rect 490434 218592 594798 218648
rect 594854 218592 594859 218648
rect 490373 218590 594859 218592
rect 596130 218650 596190 218862
rect 655421 218920 670851 218922
rect 655421 218864 655426 218920
rect 655482 218864 670790 218920
rect 670846 218864 670851 218920
rect 655421 218862 670851 218864
rect 655421 218859 655487 218862
rect 670785 218859 670851 218862
rect 648521 218650 648587 218653
rect 675201 218650 675267 218653
rect 683297 218650 683363 218653
rect 596130 218590 605850 218650
rect 490373 218587 490439 218590
rect 594793 218587 594859 218590
rect 169569 218514 169635 218517
rect 172881 218514 172947 218517
rect 169569 218512 172947 218514
rect 169569 218456 169574 218512
rect 169630 218456 172886 218512
rect 172942 218456 172947 218512
rect 169569 218454 172947 218456
rect 169569 218451 169635 218454
rect 172881 218451 172947 218454
rect 492673 218378 492739 218381
rect 493777 218378 493843 218381
rect 492673 218376 493843 218378
rect 492673 218320 492678 218376
rect 492734 218320 493782 218376
rect 493838 218320 493843 218376
rect 492673 218318 493843 218320
rect 492673 218315 492739 218318
rect 493777 218315 493843 218318
rect 496905 218378 496971 218381
rect 603257 218378 603323 218381
rect 496905 218376 603323 218378
rect 496905 218320 496910 218376
rect 496966 218320 603262 218376
rect 603318 218320 603323 218376
rect 496905 218318 603323 218320
rect 605790 218378 605850 218590
rect 648521 218648 675267 218650
rect 648521 218592 648526 218648
rect 648582 218592 675206 218648
rect 675262 218592 675267 218648
rect 648521 218590 675267 218592
rect 683284 218648 683363 218650
rect 683284 218592 683302 218648
rect 683358 218592 683363 218648
rect 683284 218590 683363 218592
rect 648521 218587 648587 218590
rect 675201 218587 675267 218590
rect 683297 218587 683363 218590
rect 631133 218378 631199 218381
rect 605790 218376 631199 218378
rect 605790 218320 631138 218376
rect 631194 218320 631199 218376
rect 605790 218318 631199 218320
rect 496905 218315 496971 218318
rect 603257 218315 603323 218318
rect 631133 218315 631199 218318
rect 675886 218316 675892 218380
rect 675956 218378 675962 218380
rect 675956 218318 676230 218378
rect 675956 218316 675962 218318
rect 676170 218242 676230 218318
rect 676170 218182 676292 218242
rect 487797 218106 487863 218109
rect 627453 218106 627519 218109
rect 487797 218104 627519 218106
rect 487797 218048 487802 218104
rect 487858 218048 627458 218104
rect 627514 218048 627519 218104
rect 487797 218046 627519 218048
rect 487797 218043 487863 218046
rect 627453 218043 627519 218046
rect 35801 217970 35867 217973
rect 61285 217970 61351 217973
rect 35801 217968 61351 217970
rect 35801 217912 35806 217968
rect 35862 217912 61290 217968
rect 61346 217912 61351 217968
rect 35801 217910 61351 217912
rect 35801 217907 35867 217910
rect 61285 217907 61351 217910
rect 508497 217834 508563 217837
rect 510153 217836 510219 217837
rect 509182 217834 509188 217836
rect 508497 217832 509188 217834
rect 508497 217776 508502 217832
rect 508558 217776 509188 217832
rect 508497 217774 509188 217776
rect 508497 217771 508563 217774
rect 509182 217772 509188 217774
rect 509252 217772 509258 217836
rect 510102 217834 510108 217836
rect 510062 217774 510108 217834
rect 510172 217832 510219 217836
rect 522573 217836 522639 217837
rect 522573 217834 522620 217836
rect 510214 217776 510219 217832
rect 510102 217772 510108 217774
rect 510172 217772 510219 217776
rect 522528 217832 522620 217834
rect 522528 217776 522578 217832
rect 522528 217774 522620 217776
rect 510153 217771 510219 217772
rect 522573 217772 522620 217774
rect 522684 217772 522690 217836
rect 555693 217834 555759 217837
rect 562685 217834 562751 217837
rect 555693 217832 562751 217834
rect 555693 217776 555698 217832
rect 555754 217776 562690 217832
rect 562746 217776 562751 217832
rect 555693 217774 562751 217776
rect 522573 217771 522639 217772
rect 555693 217771 555759 217774
rect 562685 217771 562751 217774
rect 562961 217834 563027 217837
rect 574093 217834 574159 217837
rect 562961 217832 574159 217834
rect 562961 217776 562966 217832
rect 563022 217776 574098 217832
rect 574154 217776 574159 217832
rect 562961 217774 574159 217776
rect 562961 217771 563027 217774
rect 574093 217771 574159 217774
rect 574318 217772 574324 217836
rect 574388 217834 574394 217836
rect 574829 217834 574895 217837
rect 574388 217832 574895 217834
rect 574388 217776 574834 217832
rect 574890 217776 574895 217832
rect 574388 217774 574895 217776
rect 574388 217772 574394 217774
rect 574829 217771 574895 217774
rect 675017 217834 675083 217837
rect 675017 217832 676292 217834
rect 675017 217776 675022 217832
rect 675078 217776 676292 217832
rect 675017 217774 676292 217776
rect 675017 217771 675083 217774
rect 505645 217562 505711 217565
rect 595161 217562 595227 217565
rect 505645 217560 595227 217562
rect 505645 217504 505650 217560
rect 505706 217504 595166 217560
rect 595222 217504 595227 217560
rect 505645 217502 595227 217504
rect 505645 217499 505711 217502
rect 595161 217499 595227 217502
rect 662045 217562 662111 217565
rect 675569 217562 675635 217565
rect 662045 217560 675635 217562
rect 662045 217504 662050 217560
rect 662106 217504 675574 217560
rect 675630 217504 675635 217560
rect 662045 217502 675635 217504
rect 662045 217499 662111 217502
rect 675569 217499 675635 217502
rect 675702 217364 675708 217428
rect 675772 217426 675778 217428
rect 675772 217366 676292 217426
rect 675772 217364 675778 217366
rect 493777 217292 493843 217293
rect 493726 217228 493732 217292
rect 493796 217290 493843 217292
rect 495341 217290 495407 217293
rect 498469 217290 498535 217293
rect 596357 217290 596423 217293
rect 493796 217288 493888 217290
rect 493838 217232 493888 217288
rect 493796 217230 493888 217232
rect 495341 217288 495450 217290
rect 495341 217232 495346 217288
rect 495402 217232 495450 217288
rect 493796 217228 493843 217230
rect 493777 217227 493843 217228
rect 495341 217227 495450 217232
rect 498469 217288 596423 217290
rect 498469 217232 498474 217288
rect 498530 217232 596362 217288
rect 596418 217232 596423 217288
rect 498469 217230 596423 217232
rect 498469 217227 498535 217230
rect 596357 217227 596423 217230
rect 656801 217290 656867 217293
rect 670785 217290 670851 217293
rect 656801 217288 670851 217290
rect 656801 217232 656806 217288
rect 656862 217232 670790 217288
rect 670846 217232 670851 217288
rect 656801 217230 670851 217232
rect 656801 217227 656867 217230
rect 670785 217227 670851 217230
rect 488671 217154 488737 217157
rect 488671 217152 489930 217154
rect 488671 217096 488676 217152
rect 488732 217096 489930 217152
rect 488671 217094 489930 217096
rect 488671 217091 488737 217094
rect 489870 216746 489930 217094
rect 495390 217018 495450 217227
rect 595713 217018 595779 217021
rect 495390 217016 595779 217018
rect 495390 216960 595718 217016
rect 595774 216960 595779 217016
rect 495390 216958 595779 216960
rect 595713 216955 595779 216958
rect 674649 217018 674715 217021
rect 674649 217016 676292 217018
rect 674649 216960 674654 217016
rect 674710 216960 676292 217016
rect 674649 216958 676292 216960
rect 674649 216955 674715 216958
rect 574093 216746 574159 216749
rect 574369 216748 574435 216749
rect 489870 216744 574159 216746
rect 489870 216688 574098 216744
rect 574154 216688 574159 216744
rect 489870 216686 574159 216688
rect 574093 216683 574159 216686
rect 574318 216684 574324 216748
rect 574388 216746 574435 216748
rect 574388 216744 574480 216746
rect 574430 216688 574480 216744
rect 574388 216686 574480 216688
rect 574388 216684 574435 216686
rect 574369 216683 574435 216684
rect 670969 216610 671035 216613
rect 670969 216608 676292 216610
rect 670969 216552 670974 216608
rect 671030 216552 676292 216608
rect 670969 216550 676292 216552
rect 670969 216547 671035 216550
rect 561622 216140 561628 216204
rect 561692 216202 561698 216204
rect 627913 216202 627979 216205
rect 561692 216200 627979 216202
rect 561692 216144 627918 216200
rect 627974 216144 627979 216200
rect 561692 216142 627979 216144
rect 561692 216140 561698 216142
rect 627913 216139 627979 216142
rect 665541 216202 665607 216205
rect 674833 216202 674899 216205
rect 665541 216200 671354 216202
rect 665541 216144 665546 216200
rect 665602 216144 671354 216200
rect 665541 216142 671354 216144
rect 665541 216139 665607 216142
rect 509182 215868 509188 215932
rect 509252 215930 509258 215932
rect 598473 215930 598539 215933
rect 509252 215928 598539 215930
rect 509252 215872 598478 215928
rect 598534 215872 598539 215928
rect 509252 215870 598539 215872
rect 509252 215868 509258 215870
rect 598473 215867 598539 215870
rect 652845 215930 652911 215933
rect 670693 215930 670759 215933
rect 652845 215928 670759 215930
rect 652845 215872 652850 215928
rect 652906 215872 670698 215928
rect 670754 215872 670759 215928
rect 652845 215870 670759 215872
rect 652845 215867 652911 215870
rect 670693 215867 670759 215870
rect 671294 215522 671354 216142
rect 674833 216200 676292 216202
rect 674833 216144 674838 216200
rect 674894 216144 676292 216200
rect 674833 216142 676292 216144
rect 674833 216139 674899 216142
rect 673177 215794 673243 215797
rect 673177 215792 676292 215794
rect 673177 215736 673182 215792
rect 673238 215736 676292 215792
rect 673177 215734 676292 215736
rect 673177 215731 673243 215734
rect 675937 215522 676003 215525
rect 671294 215520 676003 215522
rect 671294 215464 675942 215520
rect 675998 215464 676003 215520
rect 671294 215462 676003 215464
rect 675937 215459 676003 215462
rect 522614 215324 522620 215388
rect 522684 215386 522690 215388
rect 618897 215386 618963 215389
rect 522684 215384 618963 215386
rect 522684 215328 618902 215384
rect 618958 215328 618963 215384
rect 522684 215326 618963 215328
rect 522684 215324 522690 215326
rect 618897 215323 618963 215326
rect 676262 215310 676322 215356
rect 675886 215188 675892 215252
rect 675956 215250 675962 215252
rect 676078 215250 676322 215310
rect 675956 215190 676138 215250
rect 675956 215188 675962 215190
rect 47761 214978 47827 214981
rect 41492 214976 47827 214978
rect 41492 214920 47766 214976
rect 47822 214920 47827 214976
rect 41492 214918 47827 214920
rect 47761 214915 47827 214918
rect 673545 214978 673611 214981
rect 673545 214976 676292 214978
rect 673545 214920 673550 214976
rect 673606 214920 676292 214976
rect 673545 214918 676292 214920
rect 673545 214915 673611 214918
rect 35801 214706 35867 214709
rect 675937 214706 676003 214709
rect 35758 214704 35867 214706
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214643 35867 214648
rect 663750 214704 676003 214706
rect 663750 214648 675942 214704
rect 675998 214648 676003 214704
rect 663750 214646 676003 214648
rect 35758 214540 35818 214643
rect 658733 214570 658799 214573
rect 663750 214570 663810 214646
rect 675937 214643 676003 214646
rect 658733 214568 663810 214570
rect 658733 214512 658738 214568
rect 658794 214512 663810 214568
rect 658733 214510 663810 214512
rect 676170 214510 676292 214570
rect 658733 214507 658799 214510
rect 35801 214298 35867 214301
rect 35758 214296 35867 214298
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214235 35867 214240
rect 35758 214132 35818 214235
rect 575982 214026 576042 214404
rect 675886 214372 675892 214436
rect 675956 214434 675962 214436
rect 676170 214434 676230 214510
rect 675956 214374 676230 214434
rect 675956 214372 675962 214374
rect 674465 214162 674531 214165
rect 674465 214160 676292 214162
rect 674465 214104 674470 214160
rect 674526 214104 676292 214160
rect 674465 214102 676292 214104
rect 674465 214099 674531 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 670182 213890 670188 213892
rect 669270 213830 670188 213890
rect 44633 213754 44699 213757
rect 669270 213754 669330 213830
rect 670182 213828 670188 213830
rect 670252 213828 670258 213892
rect 41492 213752 44699 213754
rect 41492 213696 44638 213752
rect 44694 213696 44699 213752
rect 41492 213694 44699 213696
rect 44633 213691 44699 213694
rect 663750 213694 669330 213754
rect 673361 213754 673427 213757
rect 673361 213752 676292 213754
rect 673361 213696 673366 213752
rect 673422 213696 676292 213752
rect 673361 213694 676292 213696
rect 661493 213482 661559 213485
rect 663750 213482 663810 213694
rect 673361 213691 673427 213694
rect 672993 213618 673059 213621
rect 669454 213616 673059 213618
rect 669454 213560 672998 213616
rect 673054 213560 673059 213616
rect 669454 213558 673059 213560
rect 669454 213482 669514 213558
rect 672993 213555 673059 213558
rect 661493 213480 663810 213482
rect 661493 213424 661498 213480
rect 661554 213424 663810 213480
rect 661493 213422 663810 213424
rect 668534 213422 669514 213482
rect 661493 213419 661559 213422
rect 47761 213346 47827 213349
rect 41492 213344 47827 213346
rect 41492 213288 47766 213344
rect 47822 213288 47827 213344
rect 41492 213286 47827 213288
rect 47761 213283 47827 213286
rect 45553 212938 45619 212941
rect 41492 212936 45619 212938
rect 41492 212880 45558 212936
rect 45614 212880 45619 212936
rect 41492 212878 45619 212880
rect 45553 212875 45619 212878
rect 656525 212938 656591 212941
rect 668534 212938 668594 213422
rect 672901 213346 672967 213349
rect 672901 213344 676292 213346
rect 672901 213288 672906 213344
rect 672962 213288 676292 213344
rect 672901 213286 676292 213288
rect 672901 213283 672967 213286
rect 670182 213012 670188 213076
rect 670252 213074 670258 213076
rect 674097 213074 674163 213077
rect 670252 213072 674163 213074
rect 670252 213016 674102 213072
rect 674158 213016 674163 213072
rect 670252 213014 674163 213016
rect 670252 213012 670258 213014
rect 674097 213011 674163 213014
rect 683113 212938 683179 212941
rect 656525 212936 668594 212938
rect 656525 212880 656530 212936
rect 656586 212880 668594 212936
rect 682916 212936 683179 212938
rect 682916 212908 683118 212936
rect 656525 212878 668594 212880
rect 682886 212880 683118 212908
rect 683174 212880 683179 212936
rect 682886 212878 683179 212880
rect 656525 212875 656591 212878
rect 682886 212500 682946 212878
rect 683113 212875 683179 212878
rect 35390 212261 35450 212500
rect 35390 212256 35499 212261
rect 35390 212200 35438 212256
rect 35494 212200 35499 212256
rect 35390 212198 35499 212200
rect 35433 212195 35499 212198
rect 44265 212122 44331 212125
rect 41492 212120 44331 212122
rect 41492 212064 44270 212120
rect 44326 212064 44331 212120
rect 41492 212062 44331 212064
rect 44265 212059 44331 212062
rect 35617 211850 35683 211853
rect 35574 211848 35683 211850
rect 35574 211792 35622 211848
rect 35678 211792 35683 211848
rect 35574 211787 35683 211792
rect 39573 211850 39639 211853
rect 42793 211850 42859 211853
rect 39573 211848 42859 211850
rect 39573 211792 39578 211848
rect 39634 211792 42798 211848
rect 42854 211792 42859 211848
rect 39573 211790 42859 211792
rect 39573 211787 39639 211790
rect 42793 211787 42859 211790
rect 35574 211684 35634 211787
rect 575982 211714 576042 212228
rect 675845 212122 675911 212125
rect 675845 212120 676292 212122
rect 675845 212064 675850 212120
rect 675906 212064 676292 212120
rect 675845 212062 676292 212064
rect 675845 212059 675911 212062
rect 578325 211714 578391 211717
rect 575982 211712 578391 211714
rect 575982 211656 578330 211712
rect 578386 211656 578391 211712
rect 575982 211654 578391 211656
rect 578325 211651 578391 211654
rect 679022 211445 679082 211684
rect 35801 211442 35867 211445
rect 35758 211440 35867 211442
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211379 35867 211384
rect 678973 211440 679082 211445
rect 678973 211384 678978 211440
rect 679034 211384 679082 211440
rect 678973 211382 679082 211384
rect 678973 211379 679039 211382
rect 35758 211276 35818 211379
rect 47945 210898 48011 210901
rect 41492 210896 48011 210898
rect 41492 210840 47950 210896
rect 48006 210840 48011 210896
rect 41492 210838 48011 210840
rect 47945 210835 48011 210838
rect 676254 210836 676260 210900
rect 676324 210898 676330 210900
rect 676622 210898 676628 210900
rect 676324 210838 676628 210898
rect 676324 210836 676330 210838
rect 676622 210836 676628 210838
rect 676692 210836 676698 210900
rect 675886 210564 675892 210628
rect 675956 210626 675962 210628
rect 680353 210626 680419 210629
rect 675956 210624 680419 210626
rect 675956 210568 680358 210624
rect 680414 210568 680419 210624
rect 675956 210566 680419 210568
rect 675956 210564 675962 210566
rect 680353 210563 680419 210566
rect 35758 210221 35818 210460
rect 670734 210428 670740 210492
rect 670804 210490 670810 210492
rect 671981 210490 672047 210493
rect 670804 210488 672047 210490
rect 670804 210432 671986 210488
rect 672042 210432 672047 210488
rect 670804 210430 672047 210432
rect 670804 210428 670810 210430
rect 671981 210427 672047 210430
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 575982 209810 576042 210052
rect 671981 209946 672047 209949
rect 678930 209946 678990 210294
rect 683297 210291 683363 210294
rect 671981 209944 678990 209946
rect 671981 209888 671986 209944
rect 672042 209888 678990 209944
rect 671981 209886 678990 209888
rect 671981 209883 672047 209886
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 46933 209674 46999 209677
rect 41492 209672 46999 209674
rect 41492 209616 46938 209672
rect 46994 209616 46999 209672
rect 41492 209614 46999 209616
rect 46933 209611 46999 209614
rect 674097 209674 674163 209677
rect 675845 209674 675911 209677
rect 674097 209672 675911 209674
rect 674097 209616 674102 209672
rect 674158 209616 675850 209672
rect 675906 209616 675911 209672
rect 674097 209614 675911 209616
rect 674097 209611 674163 209614
rect 675845 209611 675911 209614
rect 35574 208997 35634 209236
rect 35574 208992 35683 208997
rect 35574 208936 35622 208992
rect 35678 208936 35683 208992
rect 35574 208934 35683 208936
rect 35617 208931 35683 208934
rect 35758 208589 35818 208828
rect 35758 208584 35867 208589
rect 35758 208528 35806 208584
rect 35862 208528 35867 208584
rect 35758 208526 35867 208528
rect 35801 208523 35867 208526
rect 44357 208450 44423 208453
rect 41492 208448 44423 208450
rect 41492 208392 44362 208448
rect 44418 208392 44423 208448
rect 41492 208390 44423 208392
rect 44357 208387 44423 208390
rect 672625 208316 672691 208317
rect 672574 208252 672580 208316
rect 672644 208314 672691 208316
rect 672644 208312 672736 208314
rect 672686 208256 672736 208312
rect 672644 208254 672736 208256
rect 672644 208252 672691 208254
rect 672625 208251 672691 208252
rect 40033 208178 40099 208181
rect 41638 208178 41644 208180
rect 40033 208176 41644 208178
rect 40033 208120 40038 208176
rect 40094 208120 41644 208176
rect 40033 208118 41644 208120
rect 40033 208115 40099 208118
rect 41638 208116 41644 208118
rect 41708 208116 41714 208180
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 35758 207773 35818 208012
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 35758 207768 35867 207773
rect 35758 207712 35806 207768
rect 35862 207712 35867 207768
rect 35758 207710 35867 207712
rect 35801 207707 35867 207710
rect 41689 207770 41755 207773
rect 49509 207770 49575 207773
rect 41689 207768 49575 207770
rect 41689 207712 41694 207768
rect 41750 207712 49514 207768
rect 49570 207712 49575 207768
rect 41689 207710 49575 207712
rect 41689 207707 41755 207710
rect 49509 207707 49575 207710
rect 40542 207364 40602 207604
rect 575982 207498 576042 207876
rect 668025 207634 668091 207637
rect 678973 207634 679039 207637
rect 668025 207632 679039 207634
rect 668025 207576 668030 207632
rect 668086 207576 678978 207632
rect 679034 207576 679039 207632
rect 668025 207574 679039 207576
rect 668025 207571 668091 207574
rect 678973 207571 679039 207574
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40534 207300 40540 207364
rect 40604 207300 40610 207364
rect 44173 207226 44239 207229
rect 41492 207224 44239 207226
rect 41492 207168 44178 207224
rect 44234 207168 44239 207224
rect 41492 207166 44239 207168
rect 44173 207163 44239 207166
rect 40677 206954 40743 206957
rect 42885 206954 42951 206957
rect 40677 206952 42951 206954
rect 40677 206896 40682 206952
rect 40738 206896 42890 206952
rect 42946 206896 42951 206952
rect 40677 206894 42951 206896
rect 40677 206891 40743 206894
rect 42885 206891 42951 206894
rect 676070 206892 676076 206956
rect 676140 206954 676146 206956
rect 676857 206954 676923 206957
rect 676140 206952 676923 206954
rect 676140 206896 676862 206952
rect 676918 206896 676923 206952
rect 676140 206894 676923 206896
rect 676140 206892 676146 206894
rect 676857 206891 676923 206894
rect 40726 206548 40786 206788
rect 40718 206484 40724 206548
rect 40788 206484 40794 206548
rect 41321 206546 41387 206549
rect 48773 206546 48839 206549
rect 41321 206544 48839 206546
rect 41321 206488 41326 206544
rect 41382 206488 48778 206544
rect 48834 206488 48839 206544
rect 41321 206486 48839 206488
rect 41321 206483 41387 206486
rect 48773 206483 48839 206486
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 35801 206138 35867 206141
rect 40910 206140 40970 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 35758 206136 35867 206138
rect 35758 206080 35806 206136
rect 35862 206080 35867 206136
rect 35758 206075 35867 206080
rect 40902 206076 40908 206140
rect 40972 206076 40978 206140
rect 41137 206138 41203 206141
rect 43161 206138 43227 206141
rect 41137 206136 43227 206138
rect 41137 206080 41142 206136
rect 41198 206080 43166 206136
rect 43222 206080 43227 206136
rect 41137 206078 43227 206080
rect 41137 206075 41203 206078
rect 43161 206075 43227 206078
rect 35758 205972 35818 206075
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 40309 205730 40375 205733
rect 41454 205730 41460 205732
rect 40309 205728 41460 205730
rect 40309 205672 40314 205728
rect 40370 205672 41460 205728
rect 40309 205670 41460 205672
rect 40309 205667 40375 205670
rect 41454 205668 41460 205670
rect 41524 205668 41530 205732
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 675753 205594 675819 205597
rect 676438 205594 676444 205596
rect 675753 205592 676444 205594
rect 41462 205322 41522 205564
rect 675753 205536 675758 205592
rect 675814 205536 676444 205592
rect 675753 205534 676444 205536
rect 675753 205531 675819 205534
rect 676438 205532 676444 205534
rect 676508 205532 676514 205596
rect 44633 205322 44699 205325
rect 41462 205320 44699 205322
rect 41462 205264 44638 205320
rect 44694 205264 44699 205320
rect 41462 205262 44699 205264
rect 44633 205259 44699 205262
rect 35758 204917 35818 205156
rect 35758 204912 35867 204917
rect 35758 204856 35806 204912
rect 35862 204856 35867 204912
rect 35758 204854 35867 204856
rect 35801 204851 35867 204854
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 35801 204506 35867 204509
rect 35758 204504 35867 204506
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35758 204443 35867 204448
rect 41689 204506 41755 204509
rect 43989 204506 44055 204509
rect 41689 204504 44055 204506
rect 41689 204448 41694 204504
rect 41750 204448 43994 204504
rect 44050 204448 44055 204504
rect 41689 204446 44055 204448
rect 41689 204443 41755 204446
rect 43989 204443 44055 204446
rect 35758 204340 35818 204443
rect 675753 204234 675819 204237
rect 676070 204234 676076 204236
rect 675753 204232 676076 204234
rect 675753 204176 675758 204232
rect 675814 204176 676076 204232
rect 675753 204174 676076 204176
rect 675753 204171 675819 204174
rect 676070 204172 676076 204174
rect 676140 204172 676146 204236
rect 41689 204098 41755 204101
rect 43805 204098 43871 204101
rect 668025 204098 668091 204101
rect 41689 204096 43871 204098
rect 41689 204040 41694 204096
rect 41750 204040 43810 204096
rect 43866 204040 43871 204096
rect 41689 204038 43871 204040
rect 41689 204035 41755 204038
rect 43805 204035 43871 204038
rect 666694 204096 668091 204098
rect 666694 204040 668030 204096
rect 668086 204040 668091 204096
rect 666694 204038 668091 204040
rect 666694 204030 666754 204038
rect 668025 204035 668091 204038
rect 666356 203970 666754 204030
rect 28582 203693 28642 203932
rect 672809 203826 672875 203829
rect 28533 203688 28642 203693
rect 28533 203632 28538 203688
rect 28594 203632 28642 203688
rect 28533 203630 28642 203632
rect 672766 203824 672875 203826
rect 672766 203768 672814 203824
rect 672870 203768 672875 203824
rect 672766 203763 672875 203768
rect 28533 203627 28599 203630
rect 46197 203554 46263 203557
rect 41492 203552 46263 203554
rect 41492 203496 46202 203552
rect 46258 203496 46263 203552
rect 41492 203494 46263 203496
rect 46197 203491 46263 203494
rect 40677 203282 40743 203285
rect 43069 203282 43135 203285
rect 40677 203280 43135 203282
rect 40677 203224 40682 203280
rect 40738 203224 43074 203280
rect 43130 203224 43135 203280
rect 40677 203222 43135 203224
rect 575982 203282 576042 203524
rect 672766 203421 672826 203763
rect 672717 203416 672826 203421
rect 672717 203360 672722 203416
rect 672778 203360 672826 203416
rect 672717 203358 672826 203360
rect 672717 203355 672783 203358
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 40677 203219 40743 203222
rect 43069 203219 43135 203222
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 670785 202874 670851 202877
rect 675201 202874 675267 202877
rect 670785 202872 675267 202874
rect 670785 202816 670790 202872
rect 670846 202816 675206 202872
rect 675262 202816 675267 202872
rect 670785 202814 675267 202816
rect 670785 202811 670851 202814
rect 675201 202811 675267 202814
rect 672574 202540 672580 202604
rect 672644 202602 672650 202604
rect 672809 202602 672875 202605
rect 672644 202600 672875 202602
rect 672644 202544 672814 202600
rect 672870 202544 672875 202600
rect 672644 202542 672875 202544
rect 672644 202540 672650 202542
rect 672809 202539 672875 202542
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 674465 201378 674531 201381
rect 675293 201378 675359 201381
rect 674465 201376 675359 201378
rect 575982 200834 576042 201348
rect 674465 201320 674470 201376
rect 674526 201320 675298 201376
rect 675354 201320 675359 201376
rect 674465 201318 675359 201320
rect 674465 201315 674531 201318
rect 675293 201315 675359 201318
rect 673545 201106 673611 201109
rect 675109 201106 675175 201109
rect 673545 201104 675175 201106
rect 673545 201048 673550 201104
rect 673606 201048 675114 201104
rect 675170 201048 675175 201104
rect 673545 201046 675175 201048
rect 673545 201043 673611 201046
rect 675109 201043 675175 201046
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 673177 200834 673243 200837
rect 675477 200834 675543 200837
rect 673177 200832 675543 200834
rect 673177 200776 673182 200832
rect 673238 200776 675482 200832
rect 675538 200776 675543 200832
rect 673177 200774 675543 200776
rect 673177 200771 673243 200774
rect 675477 200771 675543 200774
rect 675753 200834 675819 200837
rect 676254 200834 676260 200836
rect 675753 200832 676260 200834
rect 675753 200776 675758 200832
rect 675814 200776 676260 200832
rect 675753 200774 676260 200776
rect 675753 200771 675819 200774
rect 676254 200772 676260 200774
rect 676324 200772 676330 200836
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 28533 199338 28599 199341
rect 42241 199338 42307 199341
rect 28533 199336 42307 199338
rect 28533 199280 28538 199336
rect 28594 199280 42246 199336
rect 42302 199280 42307 199336
rect 28533 199278 42307 199280
rect 28533 199275 28599 199278
rect 42241 199275 42307 199278
rect 667933 199202 667999 199205
rect 666694 199200 667999 199202
rect 575982 198930 576042 199172
rect 666694 199144 667938 199200
rect 667994 199144 667999 199200
rect 666694 199142 667999 199144
rect 666694 199134 666754 199142
rect 667933 199139 667999 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 675753 198388 675819 198389
rect 675702 198386 675708 198388
rect 675662 198326 675708 198386
rect 675772 198384 675819 198388
rect 675814 198328 675819 198384
rect 675702 198324 675708 198326
rect 675772 198324 675819 198328
rect 675753 198323 675819 198324
rect 590377 198250 590443 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 590377 198187 590443 198190
rect 42057 197026 42123 197029
rect 44357 197026 44423 197029
rect 42057 197024 44423 197026
rect 42057 196968 42062 197024
rect 42118 196968 44362 197024
rect 44418 196968 44423 197024
rect 42057 196966 44423 196968
rect 42057 196963 42123 196966
rect 44357 196963 44423 196966
rect 49509 196482 49575 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49509 196480 52164 196482
rect 49509 196424 49514 196480
rect 49570 196424 52164 196480
rect 49509 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49509 196419 49575 196422
rect 578509 196419 578575 196422
rect 676622 196210 676628 196212
rect 675342 196150 676628 196210
rect 673361 196074 673427 196077
rect 675109 196074 675175 196077
rect 673361 196072 675175 196074
rect 673361 196016 673366 196072
rect 673422 196016 675114 196072
rect 675170 196016 675175 196072
rect 673361 196014 675175 196016
rect 673361 196011 673427 196014
rect 675109 196011 675175 196014
rect 675342 195990 675402 196150
rect 676622 196148 676628 196150
rect 676692 196148 676698 196212
rect 675296 195941 675402 195990
rect 675293 195936 675402 195941
rect 675293 195880 675298 195936
rect 675354 195930 675402 195936
rect 675354 195880 675359 195930
rect 675293 195875 675359 195880
rect 41873 195260 41939 195261
rect 41822 195258 41828 195260
rect 41782 195198 41828 195258
rect 41892 195256 41939 195260
rect 41934 195200 41939 195256
rect 41822 195196 41828 195198
rect 41892 195196 41939 195200
rect 41873 195195 41939 195196
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 48313 194442 48379 194445
rect 48313 194440 52164 194442
rect 48313 194384 48318 194440
rect 48374 194384 52164 194440
rect 48313 194382 52164 194384
rect 48313 194379 48379 194382
rect 666356 194178 666754 194238
rect 666694 194170 666754 194178
rect 667933 194170 667999 194173
rect 666694 194168 667999 194170
rect 666694 194112 667938 194168
rect 667994 194112 667999 194168
rect 666694 194110 667999 194112
rect 667933 194107 667999 194110
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 40718 193156 40724 193220
rect 40788 193218 40794 193220
rect 41781 193218 41847 193221
rect 40788 193216 41847 193218
rect 40788 193160 41786 193216
rect 41842 193160 41847 193216
rect 40788 193158 41847 193160
rect 40788 193156 40794 193158
rect 41781 193155 41847 193158
rect 671981 193218 672047 193221
rect 675109 193218 675175 193221
rect 671981 193216 675175 193218
rect 671981 193160 671986 193216
rect 672042 193160 675114 193216
rect 675170 193160 675175 193216
rect 671981 193158 675175 193160
rect 671981 193155 672047 193158
rect 675109 193155 675175 193158
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 48773 192402 48839 192405
rect 48773 192400 52164 192402
rect 48773 192344 48778 192400
rect 48834 192344 52164 192400
rect 48773 192342 52164 192344
rect 48773 192339 48839 192342
rect 575982 192266 576042 192644
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 42057 191586 42123 191589
rect 43989 191586 44055 191589
rect 42057 191584 44055 191586
rect 42057 191528 42062 191584
rect 42118 191528 43994 191584
rect 44050 191528 44055 191584
rect 42057 191526 44055 191528
rect 42057 191523 42123 191526
rect 43989 191523 44055 191526
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 44633 190498 44699 190501
rect 42425 190496 44699 190498
rect 42425 190440 42430 190496
rect 42486 190440 44638 190496
rect 44694 190440 44699 190496
rect 42425 190438 44699 190440
rect 42425 190435 42491 190438
rect 44633 190435 44699 190438
rect 47761 190498 47827 190501
rect 47761 190496 52164 190498
rect 47761 190440 47766 190496
rect 47822 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47761 190438 52164 190440
rect 47761 190435 47827 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 667933 189682 667999 189685
rect 676857 189682 676923 189685
rect 666878 189680 676923 189682
rect 666878 189624 667938 189680
rect 667994 189624 676862 189680
rect 676918 189624 676923 189680
rect 666878 189622 676923 189624
rect 666878 189342 666938 189622
rect 667933 189619 667999 189622
rect 676857 189619 676923 189622
rect 666356 189282 666938 189342
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 186826 42491 186829
rect 44173 186826 44239 186829
rect 42425 186824 44239 186826
rect 42425 186768 42430 186824
rect 42486 186768 44178 186824
rect 44234 186768 44239 186824
rect 42425 186766 44239 186768
rect 42425 186763 42491 186766
rect 44173 186763 44239 186766
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 40534 186356 40540 186420
rect 40604 186418 40610 186420
rect 41781 186418 41847 186421
rect 40604 186416 41847 186418
rect 40604 186360 41786 186416
rect 41842 186360 41847 186416
rect 40604 186358 41847 186360
rect 40604 186356 40610 186358
rect 41781 186355 41847 186358
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41781 186012 41847 186013
rect 41781 186008 41828 186012
rect 41892 186010 41898 186012
rect 41781 185952 41786 186008
rect 41781 185948 41828 185952
rect 41892 185950 41938 186010
rect 41892 185948 41898 185950
rect 41781 185947 41847 185948
rect 673361 185602 673427 185605
rect 683113 185602 683179 185605
rect 673361 185600 683179 185602
rect 673361 185544 673366 185600
rect 673422 185544 683118 185600
rect 683174 185544 683179 185600
rect 673361 185542 683179 185544
rect 673361 185539 673427 185542
rect 683113 185539 683179 185542
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 666694 184378 666754 184386
rect 668025 184378 668091 184381
rect 666694 184376 668091 184378
rect 666694 184320 668030 184376
rect 668086 184320 668091 184376
rect 666694 184318 668091 184320
rect 41454 184044 41460 184108
rect 41524 184106 41530 184108
rect 41781 184106 41847 184109
rect 41524 184104 41847 184106
rect 41524 184048 41786 184104
rect 41842 184048 41847 184104
rect 41524 184046 41847 184048
rect 41524 184044 41530 184046
rect 41781 184043 41847 184046
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 668025 184315 668091 184318
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 42425 180706 42491 180709
rect 46933 180706 46999 180709
rect 42425 180704 46999 180706
rect 42425 180648 42430 180704
rect 42486 180648 46938 180704
rect 46994 180648 46999 180704
rect 42425 180646 46999 180648
rect 42425 180643 42491 180646
rect 46933 180643 46999 180646
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 666356 179490 666754 179550
rect 666694 179482 666754 179490
rect 668025 179482 668091 179485
rect 666694 179480 668091 179482
rect 666694 179424 668030 179480
rect 668086 179424 668091 179480
rect 666694 179422 668091 179424
rect 668025 179419 668091 179422
rect 42057 179346 42123 179349
rect 50705 179346 50771 179349
rect 42057 179344 50771 179346
rect 42057 179288 42062 179344
rect 42118 179288 50710 179344
rect 50766 179288 50771 179344
rect 42057 179286 50771 179288
rect 42057 179283 42123 179286
rect 50705 179283 50771 179286
rect 683113 178802 683179 178805
rect 683070 178800 683179 178802
rect 683070 178744 683118 178800
rect 683174 178744 683179 178800
rect 683070 178739 683179 178744
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 683070 178500 683130 178739
rect 674281 178122 674347 178125
rect 674281 178120 676292 178122
rect 674281 178064 674286 178120
rect 674342 178064 676292 178120
rect 674281 178062 676292 178064
rect 674281 178059 674347 178062
rect 671153 177986 671219 177989
rect 666694 177984 671219 177986
rect 666694 177928 671158 177984
rect 671214 177928 671219 177984
rect 666694 177926 671219 177928
rect 666694 177918 666754 177926
rect 671153 177923 671219 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 672441 177714 672507 177717
rect 672441 177712 676292 177714
rect 672441 177656 672446 177712
rect 672502 177656 676292 177712
rect 672441 177654 676292 177656
rect 672441 177651 672507 177654
rect 667565 177306 667631 177309
rect 667565 177304 676292 177306
rect 667565 177248 667570 177304
rect 667626 177248 676292 177304
rect 667565 177246 676292 177248
rect 667565 177243 667631 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 674281 176898 674347 176901
rect 674281 176896 676292 176898
rect 674281 176840 674286 176896
rect 674342 176840 676292 176896
rect 674281 176838 676292 176840
rect 674281 176835 674347 176838
rect 667013 176490 667079 176493
rect 667013 176488 676292 176490
rect 667013 176432 667018 176488
rect 667074 176432 676292 176488
rect 667013 176430 676292 176432
rect 667013 176427 667079 176430
rect 674465 176082 674531 176085
rect 674465 176080 676292 176082
rect 674465 176024 674470 176080
rect 674526 176024 676292 176080
rect 674465 176022 676292 176024
rect 674465 176019 674531 176022
rect 673913 175674 673979 175677
rect 673913 175672 676292 175674
rect 673913 175616 673918 175672
rect 673974 175616 676292 175672
rect 673913 175614 676292 175616
rect 673913 175611 673979 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674649 175266 674715 175269
rect 674649 175264 676292 175266
rect 575982 175130 576042 175236
rect 674649 175208 674654 175264
rect 674710 175208 676292 175264
rect 674649 175206 676292 175208
rect 674649 175203 674715 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 667749 174994 667815 174997
rect 667749 174992 672826 174994
rect 667749 174936 667754 174992
rect 667810 174936 672826 174992
rect 667749 174934 672826 174936
rect 667749 174931 667815 174934
rect 672766 174858 672826 174934
rect 672766 174798 676292 174858
rect 669405 174722 669471 174725
rect 666694 174720 669471 174722
rect 666694 174664 669410 174720
rect 669466 174664 669471 174720
rect 666694 174662 669471 174664
rect 666694 174654 666754 174662
rect 669405 174659 669471 174662
rect 666356 174594 666754 174654
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 674925 174042 674991 174045
rect 674925 174040 676292 174042
rect 674925 173984 674930 174040
rect 674986 173984 676292 174040
rect 674925 173982 676292 173984
rect 674925 173979 674991 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675518 173572 675524 173636
rect 675588 173634 675594 173636
rect 675588 173574 676292 173634
rect 675588 173572 675594 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 668209 173090 668275 173093
rect 666694 173088 668275 173090
rect 666694 173032 668214 173088
rect 668270 173032 668275 173088
rect 666694 173030 668275 173032
rect 666694 173022 666754 173030
rect 668209 173027 668275 173030
rect 666356 172962 666754 173022
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 675702 172348 675708 172412
rect 675772 172410 675778 172412
rect 675772 172350 676292 172410
rect 675772 172348 675778 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 669405 172002 669471 172005
rect 669405 172000 676292 172002
rect 669405 171944 669410 172000
rect 669466 171944 676292 172000
rect 669405 171942 676292 171944
rect 669405 171939 669471 171942
rect 678237 171594 678303 171597
rect 678237 171592 678316 171594
rect 678237 171536 678242 171592
rect 678298 171536 678316 171592
rect 678237 171534 678316 171536
rect 678237 171531 678303 171534
rect 675334 171124 675340 171188
rect 675404 171186 675410 171188
rect 675404 171126 676292 171186
rect 675404 171124 675410 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 673913 170778 673979 170781
rect 673913 170776 676292 170778
rect 673913 170720 673918 170776
rect 673974 170720 676292 170776
rect 673913 170718 676292 170720
rect 673913 170715 673979 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 671981 170370 672047 170373
rect 671981 170368 676292 170370
rect 671981 170312 671986 170368
rect 672042 170312 676292 170368
rect 671981 170310 676292 170312
rect 671981 170307 672047 170310
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 675940 169698 676230 169758
rect 668393 169690 668459 169693
rect 666694 169688 668459 169690
rect 666694 169632 668398 169688
rect 668454 169632 668459 169688
rect 666694 169630 668459 169632
rect 668393 169627 668459 169630
rect 669446 169628 669452 169692
rect 669516 169690 669522 169692
rect 670601 169690 670667 169693
rect 675940 169692 676000 169698
rect 669516 169688 670667 169690
rect 669516 169632 670606 169688
rect 670662 169632 670667 169688
rect 669516 169630 670667 169632
rect 669516 169628 669522 169630
rect 670601 169627 670667 169630
rect 675886 169628 675892 169692
rect 675956 169630 676000 169692
rect 675956 169628 675962 169630
rect 676170 169554 676230 169698
rect 676170 169494 676292 169554
rect 675109 169418 675175 169421
rect 675937 169418 676003 169421
rect 675109 169416 676003 169418
rect 675109 169360 675114 169416
rect 675170 169360 675942 169416
rect 675998 169360 676003 169416
rect 675109 169358 676003 169360
rect 675109 169355 675175 169358
rect 675937 169355 676003 169358
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 670509 169146 670575 169149
rect 670509 169144 676292 169146
rect 670509 169088 670514 169144
rect 670570 169088 676292 169144
rect 670509 169086 676292 169088
rect 670509 169083 670575 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673177 168738 673243 168741
rect 673177 168736 676292 168738
rect 673177 168680 673182 168736
rect 673238 168680 676292 168736
rect 673177 168678 676292 168680
rect 673177 168675 673243 168678
rect 673545 168330 673611 168333
rect 673545 168328 676292 168330
rect 673545 168272 673550 168328
rect 673606 168272 676292 168328
rect 673545 168270 676292 168272
rect 673545 168267 673611 168270
rect 672257 168194 672323 168197
rect 666694 168192 672323 168194
rect 666694 168136 672262 168192
rect 672318 168136 672323 168192
rect 666694 168134 672323 168136
rect 666694 168126 666754 168134
rect 672257 168131 672323 168134
rect 666356 168066 666754 168126
rect 672257 167922 672323 167925
rect 672257 167920 676292 167922
rect 672257 167864 672262 167920
rect 672318 167864 676292 167920
rect 672257 167862 676292 167864
rect 672257 167859 672323 167862
rect 675702 167452 675708 167516
rect 675772 167514 675778 167516
rect 675772 167454 676292 167514
rect 675772 167452 675778 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 676814 166429 676874 166668
rect 676581 166428 676647 166429
rect 676581 166426 676628 166428
rect 676536 166424 676628 166426
rect 676536 166368 676586 166424
rect 676536 166366 676628 166368
rect 676581 166364 676628 166366
rect 676692 166364 676698 166428
rect 676814 166424 676923 166429
rect 676814 166368 676862 166424
rect 676918 166368 676923 166424
rect 676814 166366 676923 166368
rect 676581 166363 676647 166364
rect 676857 166363 676923 166366
rect 672349 166290 672415 166293
rect 673545 166290 673611 166293
rect 672349 166288 673611 166290
rect 672349 166232 672354 166288
rect 672410 166232 673550 166288
rect 673606 166232 673611 166288
rect 672349 166230 673611 166232
rect 672349 166227 672415 166230
rect 673545 166227 673611 166230
rect 589457 165610 589523 165613
rect 672165 165610 672231 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 672165 165608 676095 165610
rect 672165 165552 672170 165608
rect 672226 165552 676034 165608
rect 676090 165552 676095 165608
rect 672165 165550 676095 165552
rect 589457 165547 589523 165550
rect 672165 165547 672231 165550
rect 676029 165547 676095 165550
rect 668209 164930 668275 164933
rect 666694 164928 668275 164930
rect 666694 164872 668214 164928
rect 668270 164872 668275 164928
rect 666694 164870 668275 164872
rect 666694 164862 666754 164870
rect 668209 164867 668275 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668209 163298 668275 163301
rect 666694 163296 668275 163298
rect 666694 163240 668214 163296
rect 668270 163240 668275 163296
rect 666694 163238 668275 163240
rect 666694 163230 666754 163238
rect 668209 163235 668275 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675518 162148 675524 162212
rect 675588 162210 675594 162212
rect 676070 162210 676076 162212
rect 675588 162150 676076 162210
rect 675588 162148 675594 162150
rect 676070 162148 676076 162150
rect 676140 162148 676146 162212
rect 672717 161394 672783 161397
rect 675477 161394 675543 161397
rect 672717 161392 675543 161394
rect 672717 161336 672722 161392
rect 672778 161336 675482 161392
rect 675538 161336 675543 161392
rect 672717 161334 675543 161336
rect 672717 161331 672783 161334
rect 675477 161331 675543 161334
rect 675661 161258 675727 161261
rect 675661 161256 675770 161258
rect 675661 161200 675666 161256
rect 675722 161200 675770 161256
rect 675661 161195 675770 161200
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 675710 160037 675770 161195
rect 668209 160034 668275 160037
rect 666694 160032 668275 160034
rect 575982 159898 576042 160004
rect 666694 159976 668214 160032
rect 668270 159976 668275 160032
rect 666694 159974 668275 159976
rect 675710 160032 675819 160037
rect 675710 159976 675758 160032
rect 675814 159976 675819 160032
rect 675710 159974 675819 159976
rect 666694 159966 666754 159974
rect 668209 159971 668275 159974
rect 675753 159971 675819 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 674925 159490 674991 159493
rect 675477 159490 675543 159493
rect 674925 159488 675543 159490
rect 674925 159432 674930 159488
rect 674986 159432 675482 159488
rect 675538 159432 675543 159488
rect 674925 159430 675543 159432
rect 674925 159427 674991 159430
rect 675477 159427 675543 159430
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 668577 158402 668643 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 668643 158402
rect 666694 158344 668582 158400
rect 668638 158344 668643 158400
rect 666694 158342 668643 158344
rect 666694 158334 666754 158342
rect 668577 158339 668643 158342
rect 666356 158274 666754 158334
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675385 157044 675451 157045
rect 675334 157042 675340 157044
rect 675294 156982 675340 157042
rect 675404 157040 675451 157044
rect 675446 156984 675451 157040
rect 675334 156980 675340 156982
rect 675404 156980 675451 156984
rect 675385 156979 675451 156980
rect 675753 157042 675819 157045
rect 676438 157042 676444 157044
rect 675753 157040 676444 157042
rect 675753 156984 675758 157040
rect 675814 156984 676444 157040
rect 675753 156982 676444 156984
rect 675753 156979 675819 156982
rect 676438 156980 676444 156982
rect 676508 156980 676514 157044
rect 673913 156498 673979 156501
rect 675109 156498 675175 156501
rect 673913 156496 675175 156498
rect 673913 156440 673918 156496
rect 673974 156440 675114 156496
rect 675170 156440 675175 156496
rect 673913 156438 675175 156440
rect 673913 156435 673979 156438
rect 675109 156435 675175 156438
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 675753 155818 675819 155821
rect 676254 155818 676260 155820
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 675753 155816 676260 155818
rect 675753 155760 675758 155816
rect 675814 155760 676260 155816
rect 675753 155758 676260 155760
rect 589457 155755 589523 155758
rect 675753 155755 675819 155758
rect 676254 155756 676260 155758
rect 676324 155756 676330 155820
rect 668301 155138 668367 155141
rect 666694 155136 668367 155138
rect 666694 155080 668306 155136
rect 668362 155080 668367 155136
rect 666694 155078 668367 155080
rect 666694 155070 666754 155078
rect 668301 155075 668367 155078
rect 666356 155010 666754 155070
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 666878 153310 673470 153370
rect 673410 153234 673470 153310
rect 673729 153234 673795 153237
rect 673410 153232 673795 153234
rect 673410 153176 673734 153232
rect 673790 153176 673795 153232
rect 673410 153174 673795 153176
rect 673729 153171 673795 153174
rect 675661 153098 675727 153101
rect 675886 153098 675892 153100
rect 675661 153096 675892 153098
rect 675661 153040 675666 153096
rect 675722 153040 675892 153096
rect 675661 153038 675892 153040
rect 675661 153035 675727 153038
rect 675886 153036 675892 153038
rect 675956 153036 675962 153100
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675753 151466 675819 151469
rect 676622 151466 676628 151468
rect 675753 151464 676628 151466
rect 675753 151408 675758 151464
rect 675814 151408 676628 151464
rect 675753 151406 676628 151408
rect 675753 151403 675819 151406
rect 676622 151404 676628 151406
rect 676692 151404 676698 151468
rect 673177 151330 673243 151333
rect 675109 151330 675175 151333
rect 673177 151328 675175 151330
rect 673177 151272 673182 151328
rect 673238 151272 675114 151328
rect 675170 151272 675175 151328
rect 673177 151270 675175 151272
rect 673177 151267 673243 151270
rect 675109 151267 675175 151270
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 671705 150378 671771 150381
rect 666878 150376 671771 150378
rect 666878 150320 671710 150376
rect 671766 150320 671771 150376
rect 666878 150318 671771 150320
rect 666878 150174 666938 150318
rect 671705 150315 671771 150318
rect 671981 150378 672047 150381
rect 675109 150378 675175 150381
rect 671981 150376 675175 150378
rect 671981 150320 671986 150376
rect 672042 150320 675114 150376
rect 675170 150320 675175 150376
rect 671981 150318 675175 150320
rect 671981 150315 672047 150318
rect 675109 150315 675175 150318
rect 666356 150114 666938 150174
rect 670509 150106 670575 150109
rect 674925 150106 674991 150109
rect 670509 150104 674991 150106
rect 670509 150048 670514 150104
rect 670570 150048 674930 150104
rect 674986 150048 674991 150104
rect 670509 150046 674991 150048
rect 670509 150043 670575 150046
rect 674925 150043 674991 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 669405 149018 669471 149021
rect 675293 149018 675359 149021
rect 669405 149016 675359 149018
rect 669405 148960 669410 149016
rect 669466 148960 675298 149016
rect 675354 148960 675359 149016
rect 669405 148958 675359 148960
rect 669405 148955 669471 148958
rect 675293 148955 675359 148958
rect 668209 148610 668275 148613
rect 666694 148608 668275 148610
rect 666694 148552 668214 148608
rect 668270 148552 668275 148608
rect 666694 148550 668275 148552
rect 666694 148542 666754 148550
rect 668209 148547 668275 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 675661 147660 675727 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 588537 147595 588603 147598
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 671521 145346 671587 145349
rect 666694 145344 671587 145346
rect 666694 145288 671526 145344
rect 671582 145288 671587 145344
rect 666694 145286 671587 145288
rect 666694 145278 666754 145286
rect 671521 145283 671587 145286
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669221 143714 669287 143717
rect 666694 143712 669287 143714
rect 666694 143656 669226 143712
rect 669282 143656 669287 143712
rect 666694 143654 669287 143656
rect 666694 143646 666754 143654
rect 669221 143651 669287 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 669262 140450 669268 140452
rect 666694 140390 669268 140450
rect 666694 140382 666754 140390
rect 669262 140388 669268 140390
rect 669332 140388 669338 140452
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668945 138818 669011 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 669011 138818
rect 666694 138760 668950 138816
rect 669006 138760 669011 138816
rect 666694 138758 669011 138760
rect 666694 138750 666754 138758
rect 668945 138755 669011 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 668209 135554 668275 135557
rect 666694 135552 668275 135554
rect 666694 135496 668214 135552
rect 668270 135496 668275 135552
rect 666694 135494 668275 135496
rect 666694 135486 666754 135494
rect 668209 135491 668275 135494
rect 666356 135426 666754 135486
rect 590377 134602 590443 134605
rect 667381 134602 667447 134605
rect 676029 134602 676095 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 667381 134600 676095 134602
rect 667381 134544 667386 134600
rect 667442 134544 676034 134600
rect 676090 134544 676095 134600
rect 667381 134542 676095 134544
rect 590377 134539 590443 134542
rect 667381 134539 667447 134542
rect 676029 134539 676095 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 669221 133786 669287 133789
rect 666694 133784 669287 133786
rect 666694 133728 669226 133784
rect 669282 133728 669287 133784
rect 666694 133726 669287 133728
rect 669221 133723 669287 133726
rect 672942 133316 672948 133380
rect 673012 133378 673018 133380
rect 673012 133318 676292 133378
rect 673012 133316 673018 133318
rect 667197 133242 667263 133245
rect 667197 133240 672826 133242
rect 667197 133184 667202 133240
rect 667258 133184 672826 133240
rect 667197 133182 672826 133184
rect 667197 133179 667263 133182
rect 672766 133106 672826 133182
rect 672766 133046 676322 133106
rect 589457 132970 589523 132973
rect 669221 132970 669287 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 669221 132968 669330 132970
rect 669221 132912 669226 132968
rect 669282 132912 669330 132968
rect 676262 132940 676322 133046
rect 589457 132907 589523 132910
rect 669221 132907 669330 132912
rect 669270 132834 669330 132907
rect 673494 132834 673500 132836
rect 669270 132774 673500 132834
rect 673494 132772 673500 132774
rect 673564 132772 673570 132836
rect 676029 132562 676095 132565
rect 676029 132560 676292 132562
rect 676029 132504 676034 132560
rect 676090 132504 676292 132560
rect 676029 132502 676292 132504
rect 676029 132499 676095 132502
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 674281 132154 674347 132157
rect 674281 132152 676292 132154
rect 674281 132096 674286 132152
rect 674342 132096 676292 132152
rect 674281 132094 676292 132096
rect 674281 132091 674347 132094
rect 672717 131746 672783 131749
rect 672717 131744 676292 131746
rect 672717 131688 672722 131744
rect 672778 131688 676292 131744
rect 672717 131686 676292 131688
rect 672717 131683 672783 131686
rect 589457 131338 589523 131341
rect 674465 131338 674531 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674465 131336 676292 131338
rect 674465 131280 674470 131336
rect 674526 131280 676292 131336
rect 674465 131278 676292 131280
rect 589457 131275 589523 131278
rect 674465 131275 674531 131278
rect 668945 131202 669011 131205
rect 672349 131202 672415 131205
rect 668945 131200 672415 131202
rect 668945 131144 668950 131200
rect 669006 131144 672354 131200
rect 672410 131144 672415 131200
rect 668945 131142 672415 131144
rect 668945 131139 669011 131142
rect 672349 131139 672415 131142
rect 669957 130930 670023 130933
rect 669957 130928 676292 130930
rect 669957 130872 669962 130928
rect 670018 130872 676292 130928
rect 669957 130870 676292 130872
rect 669957 130867 670023 130870
rect 668761 130658 668827 130661
rect 666694 130656 668827 130658
rect 666694 130600 668766 130656
rect 668822 130600 668827 130656
rect 666694 130598 668827 130600
rect 666694 130590 666754 130598
rect 668761 130595 668827 130598
rect 666356 130530 666754 130590
rect 674649 130522 674715 130525
rect 674649 130520 676292 130522
rect 674649 130464 674654 130520
rect 674710 130464 676292 130520
rect 674649 130462 676292 130464
rect 674649 130459 674715 130462
rect 675845 130114 675911 130117
rect 675845 130112 676292 130114
rect 675845 130056 675850 130112
rect 675906 130056 676292 130112
rect 675845 130054 676292 130056
rect 675845 130051 675911 130054
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588721 129706 588787 129709
rect 673361 129706 673427 129709
rect 588721 129704 592572 129706
rect 588721 129648 588726 129704
rect 588782 129648 592572 129704
rect 588721 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 588721 129643 588787 129646
rect 673361 129643 673427 129646
rect 676262 129029 676322 129268
rect 668577 129026 668643 129029
rect 666694 129024 668643 129026
rect 666694 128968 668582 129024
rect 668638 128968 668643 129024
rect 666694 128966 668643 128968
rect 666694 128958 666754 128966
rect 668577 128963 668643 128966
rect 676213 129024 676322 129029
rect 676213 128968 676218 129024
rect 676274 128968 676322 129024
rect 676213 128966 676322 128968
rect 676213 128963 676279 128966
rect 666356 128898 666754 128958
rect 676446 128620 676506 128860
rect 676438 128556 676444 128620
rect 676508 128556 676514 128620
rect 671337 128346 671403 128349
rect 676029 128346 676095 128349
rect 671337 128344 676095 128346
rect 671337 128288 671342 128344
rect 671398 128288 676034 128344
rect 676090 128288 676095 128344
rect 671337 128286 676095 128288
rect 671337 128283 671403 128286
rect 676029 128283 676095 128286
rect 676262 128212 676322 128452
rect 676254 128148 676260 128212
rect 676324 128148 676330 128212
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676262 127805 676322 128044
rect 676213 127800 676322 127805
rect 676213 127744 676218 127800
rect 676274 127744 676322 127800
rect 676213 127742 676322 127744
rect 676213 127739 676279 127742
rect 674833 127394 674899 127397
rect 676446 127394 676506 127636
rect 674833 127392 676506 127394
rect 674833 127336 674838 127392
rect 674894 127336 676506 127392
rect 674833 127334 676506 127336
rect 674833 127331 674899 127334
rect 668577 126986 668643 126989
rect 675845 126986 675911 126989
rect 668577 126984 675911 126986
rect 668577 126928 668582 126984
rect 668638 126928 675850 126984
rect 675906 126928 675911 126984
rect 668577 126926 675911 126928
rect 668577 126923 668643 126926
rect 675845 126923 675911 126926
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 673361 126578 673427 126581
rect 676262 126578 676322 126820
rect 673361 126576 676322 126578
rect 673361 126520 673366 126576
rect 673422 126520 676322 126576
rect 673361 126518 676322 126520
rect 673361 126515 673427 126518
rect 589917 126442 589983 126445
rect 589917 126440 592572 126442
rect 589917 126384 589922 126440
rect 589978 126384 592572 126440
rect 589917 126382 592572 126384
rect 589917 126379 589983 126382
rect 682334 126173 682394 126412
rect 682334 126168 682443 126173
rect 682334 126112 682382 126168
rect 682438 126112 682443 126168
rect 682334 126110 682443 126112
rect 682377 126107 682443 126110
rect 683070 125765 683130 126004
rect 670734 125762 670740 125764
rect 666694 125702 670740 125762
rect 666694 125694 666754 125702
rect 670734 125700 670740 125702
rect 670804 125700 670810 125764
rect 676213 125762 676279 125765
rect 676213 125760 676322 125762
rect 676213 125704 676218 125760
rect 676274 125704 676322 125760
rect 676213 125699 676322 125704
rect 683070 125760 683179 125765
rect 683070 125704 683118 125760
rect 683174 125704 683179 125760
rect 683070 125702 683179 125704
rect 683113 125699 683179 125702
rect 666356 125634 666754 125694
rect 676262 125596 676322 125699
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 668025 125354 668091 125357
rect 678973 125354 679039 125357
rect 668025 125352 679039 125354
rect 668025 125296 668030 125352
rect 668086 125296 678978 125352
rect 679034 125296 679039 125352
rect 668025 125294 679039 125296
rect 668025 125291 668091 125294
rect 678973 125291 679039 125294
rect 683254 124949 683314 125188
rect 683254 124944 683363 124949
rect 683254 124888 683302 124944
rect 683358 124888 683363 124944
rect 683254 124886 683363 124888
rect 683297 124883 683363 124886
rect 589365 124810 589431 124813
rect 672349 124810 672415 124813
rect 589365 124808 592572 124810
rect 589365 124752 589370 124808
rect 589426 124752 592572 124808
rect 589365 124750 592572 124752
rect 672349 124808 676292 124810
rect 672349 124752 672354 124808
rect 672410 124752 676292 124808
rect 672349 124750 676292 124752
rect 589365 124747 589431 124750
rect 672349 124747 672415 124750
rect 674465 124402 674531 124405
rect 674465 124400 676292 124402
rect 674465 124344 674470 124400
rect 674526 124344 676292 124400
rect 674465 124342 676292 124344
rect 674465 124339 674531 124342
rect 672901 124130 672967 124133
rect 666694 124128 672967 124130
rect 666694 124072 672906 124128
rect 672962 124072 672967 124128
rect 666694 124070 672967 124072
rect 666694 124062 666754 124070
rect 672901 124067 672967 124070
rect 666356 124002 666754 124062
rect 673177 123994 673243 123997
rect 673177 123992 676292 123994
rect 673177 123936 673182 123992
rect 673238 123936 676292 123992
rect 673177 123934 676292 123936
rect 673177 123931 673243 123934
rect 578693 123586 578759 123589
rect 575798 123584 578759 123586
rect 575798 123528 578698 123584
rect 578754 123528 578759 123584
rect 575798 123526 578759 123528
rect 575798 123012 575858 123526
rect 578693 123523 578759 123526
rect 674649 123586 674715 123589
rect 674649 123584 676292 123586
rect 674649 123528 674654 123584
rect 674710 123528 676292 123584
rect 674649 123526 676292 123528
rect 674649 123523 674715 123526
rect 589549 123178 589615 123181
rect 673453 123178 673519 123181
rect 589549 123176 592572 123178
rect 589549 123120 589554 123176
rect 589610 123120 592572 123176
rect 589549 123118 592572 123120
rect 673453 123176 676292 123178
rect 673453 123120 673458 123176
rect 673514 123120 676292 123176
rect 673453 123118 676292 123120
rect 589549 123115 589615 123118
rect 673453 123115 673519 123118
rect 675702 122844 675708 122908
rect 675772 122906 675778 122908
rect 675937 122906 676003 122909
rect 675772 122904 676003 122906
rect 675772 122848 675942 122904
rect 675998 122848 676003 122904
rect 675772 122846 676003 122848
rect 675772 122844 675778 122846
rect 675937 122843 676003 122846
rect 676170 122710 676292 122770
rect 668761 122634 668827 122637
rect 676170 122634 676230 122710
rect 668761 122632 676230 122634
rect 668761 122576 668766 122632
rect 668822 122576 676230 122632
rect 668761 122574 676230 122576
rect 668761 122571 668827 122574
rect 676170 122302 676292 122362
rect 673913 122226 673979 122229
rect 676170 122226 676230 122302
rect 673913 122224 676230 122226
rect 673913 122168 673918 122224
rect 673974 122168 676230 122224
rect 673913 122166 676230 122168
rect 673913 122163 673979 122166
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589549 121546 589615 121549
rect 589549 121544 592572 121546
rect 589549 121488 589554 121544
rect 589610 121488 592572 121544
rect 589549 121486 592572 121488
rect 589549 121483 589615 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 671521 121410 671587 121413
rect 675894 121410 675954 121622
rect 676806 121620 676812 121684
rect 676876 121682 676882 121684
rect 683113 121682 683179 121685
rect 676876 121680 683179 121682
rect 676876 121624 683118 121680
rect 683174 121624 683179 121680
rect 676876 121622 683179 121624
rect 676876 121620 676882 121622
rect 683113 121619 683179 121622
rect 671521 121408 675954 121410
rect 671521 121352 671526 121408
rect 671582 121352 675954 121408
rect 671521 121350 675954 121352
rect 671521 121347 671587 121350
rect 679022 121277 679082 121516
rect 678973 121272 679082 121277
rect 678973 121216 678978 121272
rect 679034 121216 679082 121272
rect 678973 121214 679082 121216
rect 678973 121211 679039 121214
rect 666356 120738 666938 120798
rect 666878 120458 666938 120738
rect 674097 120458 674163 120461
rect 666878 120456 674163 120458
rect 666878 120400 674102 120456
rect 674158 120400 674163 120456
rect 666878 120398 674163 120400
rect 674097 120395 674163 120398
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 669221 119642 669287 119645
rect 673453 119642 673519 119645
rect 669221 119640 673519 119642
rect 669221 119584 669226 119640
rect 669282 119584 673458 119640
rect 673514 119584 673519 119640
rect 669221 119582 673519 119584
rect 669221 119579 669287 119582
rect 673453 119579 673519 119582
rect 668945 119234 669011 119237
rect 666694 119232 669011 119234
rect 666694 119176 668950 119232
rect 669006 119176 669011 119232
rect 666694 119174 669011 119176
rect 666694 119166 666754 119174
rect 668945 119171 669011 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 672533 117602 672599 117605
rect 666694 117600 672599 117602
rect 666694 117544 672538 117600
rect 672594 117544 672599 117600
rect 666694 117542 672599 117544
rect 666694 117534 666754 117542
rect 672533 117539 672599 117542
rect 666356 117474 666754 117534
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 675109 116786 675175 116789
rect 675845 116786 675911 116789
rect 675109 116784 675911 116786
rect 675109 116728 675114 116784
rect 675170 116728 675850 116784
rect 675906 116728 675911 116784
rect 675109 116726 675911 116728
rect 675109 116723 675175 116726
rect 675845 116723 675911 116726
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 675886 116452 675892 116516
rect 675956 116514 675962 116516
rect 683297 116514 683363 116517
rect 675956 116512 683363 116514
rect 675956 116456 683302 116512
rect 683358 116456 683363 116512
rect 675956 116454 683363 116456
rect 675956 116452 675962 116454
rect 683297 116451 683363 116454
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 672165 115834 672231 115837
rect 666694 115832 672231 115834
rect 666694 115776 672170 115832
rect 672226 115776 672231 115832
rect 666694 115774 672231 115776
rect 672165 115771 672231 115774
rect 674046 115772 674052 115836
rect 674116 115834 674122 115836
rect 675477 115834 675543 115837
rect 674116 115832 675543 115834
rect 674116 115776 675482 115832
rect 675538 115776 675543 115832
rect 674116 115774 675543 115776
rect 674116 115772 674122 115774
rect 675477 115771 675543 115774
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669221 114338 669287 114341
rect 666694 114336 669287 114338
rect 666694 114280 669226 114336
rect 669282 114280 669287 114336
rect 666694 114278 669287 114280
rect 666694 114270 666754 114278
rect 669221 114275 669287 114278
rect 666356 114210 666754 114270
rect 675753 114202 675819 114205
rect 676438 114202 676444 114204
rect 675753 114200 676444 114202
rect 675753 114144 675758 114200
rect 675814 114144 676444 114200
rect 675753 114142 676444 114144
rect 675753 114139 675819 114142
rect 676438 114140 676444 114142
rect 676508 114140 676514 114204
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 668945 112706 669011 112709
rect 666694 112704 669011 112706
rect 666694 112648 668950 112704
rect 669006 112648 669011 112704
rect 666694 112646 669011 112648
rect 666694 112638 666754 112646
rect 668945 112643 669011 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 589457 111754 589523 111757
rect 675753 111754 675819 111757
rect 676806 111754 676812 111756
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 675753 111752 676812 111754
rect 675753 111696 675758 111752
rect 675814 111696 676812 111752
rect 675753 111694 676812 111696
rect 589457 111691 589523 111694
rect 675753 111691 675819 111694
rect 676806 111692 676812 111694
rect 676876 111692 676882 111756
rect 675661 111348 675727 111349
rect 675661 111344 675708 111348
rect 675772 111346 675778 111348
rect 675661 111288 675666 111344
rect 675661 111284 675708 111288
rect 675772 111286 675818 111346
rect 675772 111284 675778 111286
rect 675661 111283 675727 111284
rect 671521 111074 671587 111077
rect 666694 111072 671587 111074
rect 666694 111016 671526 111072
rect 671582 111016 671587 111072
rect 666694 111014 671587 111016
rect 666694 111006 666754 111014
rect 671521 111011 671587 111014
rect 666356 110946 666754 111006
rect 674465 110394 674531 110397
rect 675109 110394 675175 110397
rect 674465 110392 675175 110394
rect 674465 110336 674470 110392
rect 674526 110336 675114 110392
rect 675170 110336 675175 110392
rect 674465 110334 675175 110336
rect 674465 110331 674531 110334
rect 675109 110331 675175 110334
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589457 110122 589523 110125
rect 589457 110120 592572 110122
rect 589457 110064 589462 110120
rect 589518 110064 592572 110120
rect 589457 110062 592572 110064
rect 589457 110059 589523 110062
rect 666645 109374 666711 109377
rect 666356 109372 666711 109374
rect 666356 109316 666650 109372
rect 666706 109316 666711 109372
rect 666356 109314 666711 109316
rect 666645 109311 666711 109314
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 667933 107810 667999 107813
rect 666694 107808 667999 107810
rect 666694 107752 667938 107808
rect 667994 107752 667999 107808
rect 666694 107750 667999 107752
rect 666694 107742 666754 107750
rect 667933 107747 667999 107750
rect 666356 107682 666754 107742
rect 672349 106994 672415 106997
rect 675385 106994 675451 106997
rect 672349 106992 675451 106994
rect 672349 106936 672354 106992
rect 672410 106936 675390 106992
rect 675446 106936 675451 106992
rect 672349 106934 675451 106936
rect 672349 106931 672415 106934
rect 675385 106931 675451 106934
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 673177 106314 673243 106317
rect 675109 106314 675175 106317
rect 673177 106312 675175 106314
rect 673177 106256 673182 106312
rect 673238 106256 675114 106312
rect 675170 106256 675175 106312
rect 673177 106254 675175 106256
rect 673177 106251 673243 106254
rect 675109 106251 675175 106254
rect 668025 106178 668091 106181
rect 672717 106178 672783 106181
rect 666694 106176 672783 106178
rect 666694 106120 668030 106176
rect 668086 106120 672722 106176
rect 672778 106120 672783 106176
rect 666694 106118 672783 106120
rect 666694 106110 666754 106118
rect 668025 106115 668091 106118
rect 672717 106115 672783 106118
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589825 105226 589891 105229
rect 589825 105224 592572 105226
rect 589825 105168 589830 105224
rect 589886 105168 592572 105224
rect 589825 105166 592572 105168
rect 589825 105163 589891 105166
rect 675661 104818 675727 104821
rect 675886 104818 675892 104820
rect 675661 104816 675892 104818
rect 675661 104760 675666 104816
rect 675722 104760 675892 104816
rect 675661 104758 675892 104760
rect 675661 104755 675727 104758
rect 675886 104756 675892 104758
rect 675956 104756 675962 104820
rect 666356 104418 666754 104478
rect 666694 104410 666754 104418
rect 668209 104410 668275 104413
rect 666694 104408 668275 104410
rect 666694 104352 668214 104408
rect 668270 104352 668275 104408
rect 666694 104350 668275 104352
rect 668209 104347 668275 104350
rect 588537 103594 588603 103597
rect 588537 103592 592572 103594
rect 588537 103536 588542 103592
rect 588598 103536 592572 103592
rect 588537 103534 592572 103536
rect 588537 103531 588603 103534
rect 575982 103186 576042 103428
rect 578509 103186 578575 103189
rect 575982 103184 578575 103186
rect 575982 103128 578514 103184
rect 578570 103128 578575 103184
rect 575982 103126 578575 103128
rect 578509 103123 578575 103126
rect 675753 103186 675819 103189
rect 676254 103186 676260 103188
rect 675753 103184 676260 103186
rect 675753 103128 675758 103184
rect 675814 103128 676260 103184
rect 675753 103126 676260 103128
rect 675753 103123 675819 103126
rect 676254 103124 676260 103126
rect 676324 103124 676330 103188
rect 666356 102786 666754 102846
rect 666694 102778 666754 102786
rect 667933 102778 667999 102781
rect 668577 102778 668643 102781
rect 666694 102776 668643 102778
rect 666694 102720 667938 102776
rect 667994 102720 668582 102776
rect 668638 102720 668643 102776
rect 666694 102718 668643 102720
rect 667933 102715 667999 102718
rect 668577 102715 668643 102718
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579153 101690 579219 101693
rect 575798 101688 579219 101690
rect 575798 101632 579158 101688
rect 579214 101632 579219 101688
rect 575798 101630 579219 101632
rect 575798 101252 575858 101630
rect 579153 101627 579219 101630
rect 673361 101010 673427 101013
rect 675109 101010 675175 101013
rect 673361 101008 675175 101010
rect 673361 100952 673366 101008
rect 673422 100952 675114 101008
rect 675170 100952 675175 101008
rect 673361 100950 675175 100952
rect 673361 100947 673427 100950
rect 675109 100947 675175 100950
rect 579521 99242 579587 99245
rect 575798 99240 579587 99242
rect 575798 99184 579526 99240
rect 579582 99184 579587 99240
rect 575798 99182 579587 99184
rect 575798 99076 575858 99182
rect 579521 99179 579587 99182
rect 578601 97474 578667 97477
rect 575798 97472 578667 97474
rect 575798 97416 578606 97472
rect 578662 97416 578667 97472
rect 575798 97414 578667 97416
rect 575798 96900 575858 97414
rect 578601 97411 578667 97414
rect 635549 96930 635615 96933
rect 635774 96930 635780 96932
rect 635549 96928 635780 96930
rect 635549 96872 635554 96928
rect 635610 96872 635780 96928
rect 635549 96870 635780 96872
rect 635549 96867 635615 96870
rect 635774 96868 635780 96870
rect 635844 96868 635850 96932
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 648061 96522 648127 96525
rect 649257 96522 649323 96525
rect 648061 96520 649323 96522
rect 648061 96464 648066 96520
rect 648122 96464 649262 96520
rect 649318 96464 649323 96520
rect 648061 96462 649323 96464
rect 648061 96459 648127 96462
rect 649257 96459 649323 96462
rect 645577 96114 645643 96117
rect 648797 96114 648863 96117
rect 645577 96112 648863 96114
rect 645577 96056 645582 96112
rect 645638 96056 648802 96112
rect 648858 96056 648863 96112
rect 645577 96054 648863 96056
rect 645577 96051 645643 96054
rect 648797 96051 648863 96054
rect 633934 95916 633940 95980
rect 634004 95978 634010 95980
rect 635733 95978 635799 95981
rect 634004 95976 635799 95978
rect 634004 95920 635738 95976
rect 635794 95920 635799 95976
rect 634004 95918 635799 95920
rect 634004 95916 634010 95918
rect 635733 95915 635799 95918
rect 647877 95842 647943 95845
rect 656341 95842 656407 95845
rect 647877 95840 656407 95842
rect 647877 95784 647882 95840
rect 647938 95784 656346 95840
rect 656402 95784 656407 95840
rect 647877 95782 656407 95784
rect 647877 95779 647943 95782
rect 656341 95779 656407 95782
rect 578325 95026 578391 95029
rect 575798 95024 578391 95026
rect 575798 94968 578330 95024
rect 578386 94968 578391 95024
rect 575798 94966 578391 94968
rect 575798 94724 575858 94966
rect 578325 94963 578391 94966
rect 647325 95026 647391 95029
rect 647325 95024 647434 95026
rect 647325 94968 647330 95024
rect 647386 94968 647434 95024
rect 647325 94963 647434 94968
rect 625429 94482 625495 94485
rect 625429 94480 628268 94482
rect 625429 94424 625434 94480
rect 625490 94424 628268 94480
rect 647374 94452 647434 94963
rect 625429 94422 628268 94424
rect 625429 94419 625495 94422
rect 655053 94210 655119 94213
rect 655053 94208 656788 94210
rect 655053 94152 655058 94208
rect 655114 94152 656788 94208
rect 655053 94150 656788 94152
rect 655053 94147 655119 94150
rect 626349 93666 626415 93669
rect 626349 93664 628268 93666
rect 626349 93608 626354 93664
rect 626410 93608 628268 93664
rect 626349 93606 628268 93608
rect 626349 93603 626415 93606
rect 654685 93394 654751 93397
rect 665357 93394 665423 93397
rect 654685 93392 656788 93394
rect 654685 93336 654690 93392
rect 654746 93336 656788 93392
rect 654685 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 654685 93331 654751 93334
rect 665357 93331 665423 93334
rect 579245 93122 579311 93125
rect 575798 93120 579311 93122
rect 575798 93064 579250 93120
rect 579306 93064 579311 93120
rect 575798 93062 579311 93064
rect 575798 92548 575858 93062
rect 579245 93059 579311 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626165 92850 626231 92853
rect 626165 92848 628268 92850
rect 626165 92792 626170 92848
rect 626226 92792 628268 92848
rect 626165 92790 628268 92792
rect 626165 92787 626231 92790
rect 656758 92548 656818 93062
rect 663977 92578 664043 92581
rect 663596 92576 664043 92578
rect 663596 92520 663982 92576
rect 664038 92520 664043 92576
rect 663596 92518 664043 92520
rect 663977 92515 664043 92518
rect 625797 92034 625863 92037
rect 648613 92034 648679 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648679 92034
rect 648140 91976 648618 92032
rect 648674 91976 648679 92032
rect 648140 91974 648679 91976
rect 625797 91971 625863 91974
rect 648613 91971 648679 91974
rect 664161 91762 664227 91765
rect 663596 91760 664227 91762
rect 663596 91704 664166 91760
rect 664222 91704 664227 91760
rect 663596 91702 664227 91704
rect 664161 91699 664227 91702
rect 655421 91490 655487 91493
rect 655421 91488 656788 91490
rect 655421 91432 655426 91488
rect 655482 91432 656788 91488
rect 655421 91430 656788 91432
rect 655421 91427 655487 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 663793 91082 663859 91085
rect 663566 91080 663859 91082
rect 663566 91024 663798 91080
rect 663854 91024 663859 91080
rect 663566 91022 663859 91024
rect 578693 90946 578759 90949
rect 575798 90944 578759 90946
rect 575798 90888 578698 90944
rect 578754 90888 578759 90944
rect 575798 90886 578759 90888
rect 575798 90372 575858 90886
rect 578693 90883 578759 90886
rect 655421 90674 655487 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 663566 90644 663626 91022
rect 663793 91019 663859 91022
rect 655421 90614 656788 90616
rect 655421 90611 655487 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664529 89858 664595 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664595 89858
rect 663596 89800 664534 89856
rect 664590 89800 664595 89856
rect 663596 89798 664595 89800
rect 655789 89795 655855 89798
rect 664529 89795 664595 89798
rect 625245 89586 625311 89589
rect 648245 89586 648311 89589
rect 625245 89584 628268 89586
rect 625245 89528 625250 89584
rect 625306 89528 628268 89584
rect 625245 89526 628268 89528
rect 648140 89584 648311 89586
rect 648140 89528 648250 89584
rect 648306 89528 648311 89584
rect 648140 89526 648311 89528
rect 625245 89523 625311 89526
rect 648245 89523 648311 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 625429 88770 625495 88773
rect 625429 88768 628268 88770
rect 625429 88712 625434 88768
rect 625490 88712 628268 88768
rect 625429 88710 628268 88712
rect 625429 88707 625495 88710
rect 624969 88634 625035 88637
rect 625245 88634 625311 88637
rect 624969 88632 625311 88634
rect 624969 88576 624974 88632
rect 625030 88576 625250 88632
rect 625306 88576 625311 88632
rect 624969 88574 625311 88576
rect 624969 88571 625035 88574
rect 625245 88571 625311 88574
rect 575982 88090 576042 88196
rect 579245 88090 579311 88093
rect 575982 88088 579311 88090
rect 575982 88032 579250 88088
rect 579306 88032 579311 88088
rect 575982 88030 579311 88032
rect 579245 88027 579311 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 625613 87138 625679 87141
rect 650545 87138 650611 87141
rect 625613 87136 628268 87138
rect 625613 87080 625618 87136
rect 625674 87080 628268 87136
rect 625613 87078 628268 87080
rect 648140 87136 650611 87138
rect 648140 87080 650550 87136
rect 650606 87080 650611 87136
rect 648140 87078 650611 87080
rect 625613 87075 625679 87078
rect 650545 87075 650611 87078
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 625337 85506 625403 85509
rect 625337 85504 628268 85506
rect 625337 85448 625342 85504
rect 625398 85448 628268 85504
rect 625337 85446 628268 85448
rect 625337 85443 625403 85446
rect 626441 84690 626507 84693
rect 648613 84690 648679 84693
rect 626441 84688 628268 84690
rect 626441 84632 626446 84688
rect 626502 84632 628268 84688
rect 626441 84630 628268 84632
rect 648140 84688 648679 84690
rect 648140 84632 648618 84688
rect 648674 84632 648679 84688
rect 648140 84630 648679 84632
rect 626441 84627 626507 84630
rect 648613 84627 648679 84630
rect 579245 84010 579311 84013
rect 575798 84008 579311 84010
rect 575798 83952 579250 84008
rect 579306 83952 579311 84008
rect 575798 83950 579311 83952
rect 575798 83844 575858 83950
rect 579245 83947 579311 83950
rect 625797 83874 625863 83877
rect 625797 83872 628268 83874
rect 625797 83816 625802 83872
rect 625858 83816 628268 83872
rect 625797 83814 628268 83816
rect 625797 83811 625863 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 578693 82242 578759 82245
rect 650269 82242 650335 82245
rect 575798 82240 578759 82242
rect 575798 82184 578698 82240
rect 578754 82184 578759 82240
rect 648140 82240 650335 82242
rect 575798 82182 578759 82184
rect 575798 81668 575858 82182
rect 578693 82179 578759 82182
rect 628790 81698 628850 82212
rect 648140 82184 650274 82240
rect 650330 82184 650335 82240
rect 648140 82182 650335 82184
rect 650269 82179 650335 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 579429 80066 579495 80069
rect 575798 80064 579495 80066
rect 575798 80008 579434 80064
rect 579490 80008 579495 80064
rect 575798 80006 579495 80008
rect 575798 79492 575858 80006
rect 579429 80003 579495 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 635774 78100 635780 78164
rect 635844 78162 635850 78164
rect 647509 78162 647575 78165
rect 635844 78160 647575 78162
rect 635844 78104 647514 78160
rect 647570 78104 647575 78160
rect 635844 78102 647575 78104
rect 635844 78100 635850 78102
rect 647509 78099 647575 78102
rect 578509 77890 578575 77893
rect 575798 77888 578575 77890
rect 575798 77832 578514 77888
rect 578570 77832 578575 77888
rect 575798 77830 578575 77832
rect 575798 77316 575858 77830
rect 578509 77827 578575 77830
rect 580441 77890 580507 77893
rect 580441 77888 625170 77890
rect 580441 77832 580446 77888
rect 580502 77832 625170 77888
rect 580441 77830 625170 77832
rect 580441 77827 580507 77830
rect 625110 77618 625170 77830
rect 637062 77618 637068 77620
rect 625110 77558 637068 77618
rect 637062 77556 637068 77558
rect 637132 77618 637138 77620
rect 639597 77618 639663 77621
rect 637132 77616 639663 77618
rect 637132 77560 639602 77616
rect 639658 77560 639663 77616
rect 637132 77558 639663 77560
rect 637132 77556 637138 77558
rect 639597 77555 639663 77558
rect 623037 77346 623103 77349
rect 633893 77346 633959 77349
rect 623037 77344 633959 77346
rect 623037 77288 623042 77344
rect 623098 77288 633898 77344
rect 633954 77288 633959 77344
rect 623037 77286 633959 77288
rect 623037 77283 623103 77286
rect 633893 77283 633959 77286
rect 579061 75714 579127 75717
rect 575798 75712 579127 75714
rect 575798 75656 579066 75712
rect 579122 75656 579127 75712
rect 575798 75654 579127 75656
rect 575798 75140 575858 75654
rect 579061 75651 579127 75654
rect 646313 74218 646379 74221
rect 646270 74216 646379 74218
rect 646270 74160 646318 74216
rect 646374 74160 646379 74216
rect 646270 74155 646379 74160
rect 646270 73848 646330 74155
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 646497 71770 646563 71773
rect 646454 71768 646563 71770
rect 646454 71712 646502 71768
rect 646558 71712 646563 71768
rect 646454 71707 646563 71712
rect 646454 71400 646514 71707
rect 578509 71226 578575 71229
rect 575798 71224 578575 71226
rect 575798 71168 578514 71224
rect 578570 71168 578575 71224
rect 575798 71166 578575 71168
rect 575798 70788 575858 71166
rect 578509 71163 578575 71166
rect 646129 69186 646195 69189
rect 646086 69184 646195 69186
rect 646086 69128 646134 69184
rect 646190 69128 646195 69184
rect 646086 69123 646195 69128
rect 646086 68952 646146 69123
rect 575798 66874 575858 68612
rect 646129 67146 646195 67149
rect 646086 67144 646195 67146
rect 646086 67088 646134 67144
rect 646190 67088 646195 67144
rect 646086 67083 646195 67088
rect 579521 66874 579587 66877
rect 575798 66872 579587 66874
rect 575798 66816 579526 66872
rect 579582 66816 579587 66872
rect 575798 66814 579587 66816
rect 575798 66436 575858 66814
rect 579521 66811 579587 66814
rect 646086 66504 646146 67083
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 647325 64426 647391 64429
rect 646638 64424 647391 64426
rect 646638 64368 647330 64424
rect 647386 64368 647391 64424
rect 646638 64366 647391 64368
rect 646638 64056 646698 64366
rect 647325 64363 647391 64366
rect 648981 62114 649047 62117
rect 646638 62112 649047 62114
rect 575982 61842 576042 62084
rect 646638 62056 648986 62112
rect 649042 62056 649047 62112
rect 646638 62054 649047 62056
rect 579521 61842 579587 61845
rect 575982 61840 579587 61842
rect 575982 61784 579526 61840
rect 579582 61784 579587 61840
rect 575982 61782 579587 61784
rect 579521 61779 579587 61782
rect 646638 61608 646698 62054
rect 648981 62051 649047 62054
rect 578877 60482 578943 60485
rect 575798 60480 578943 60482
rect 575798 60424 578882 60480
rect 578938 60424 578943 60480
rect 575798 60422 578943 60424
rect 575798 59908 575858 60422
rect 578877 60419 578943 60422
rect 648613 59258 648679 59261
rect 646638 59256 648679 59258
rect 646638 59200 648618 59256
rect 648674 59200 648679 59256
rect 646638 59198 648679 59200
rect 646638 59160 646698 59198
rect 648613 59195 648679 59198
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 647509 57354 647575 57357
rect 646638 57352 647575 57354
rect 646638 57296 647514 57352
rect 647570 57296 647575 57352
rect 646638 57294 647575 57296
rect 646638 56712 646698 57294
rect 647509 57291 647575 57294
rect 578325 56130 578391 56133
rect 575798 56128 578391 56130
rect 575798 56072 578330 56128
rect 578386 56072 578391 56128
rect 575798 56070 578391 56072
rect 575798 55556 575858 56070
rect 578325 56067 578391 56070
rect 461710 54980 461716 55044
rect 461780 55042 461786 55044
rect 576117 55042 576183 55045
rect 461780 55040 576183 55042
rect 461780 54984 576122 55040
rect 576178 54984 576183 55040
rect 461780 54982 576183 54984
rect 461780 54980 461786 54982
rect 576117 54979 576183 54982
rect 462630 54708 462636 54772
rect 462700 54770 462706 54772
rect 577681 54770 577747 54773
rect 462700 54768 577747 54770
rect 462700 54712 577686 54768
rect 577742 54712 577747 54768
rect 462700 54710 577747 54712
rect 462700 54708 462706 54710
rect 577681 54707 577747 54710
rect 591297 54498 591363 54501
rect 460798 54496 591363 54498
rect 460798 54440 591302 54496
rect 591358 54440 591363 54496
rect 460798 54438 591363 54440
rect 460798 53685 460858 54438
rect 591297 54435 591363 54438
rect 461710 53892 461716 53956
rect 461780 53892 461786 53956
rect 462630 53892 462636 53956
rect 462700 53892 462706 53956
rect 461718 53685 461778 53892
rect 462638 53685 462698 53892
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462589 53680 462698 53685
rect 462589 53624 462594 53680
rect 462650 53624 462698 53680
rect 462589 53622 462698 53624
rect 463141 53682 463207 53685
rect 473905 53682 473971 53685
rect 463141 53680 473971 53682
rect 463141 53624 463146 53680
rect 463202 53624 473910 53680
rect 473966 53624 473971 53680
rect 463141 53622 473971 53624
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53619 462655 53622
rect 463141 53619 463207 53622
rect 473905 53619 473971 53622
rect 564525 53682 564591 53685
rect 574737 53682 574803 53685
rect 564525 53680 574803 53682
rect 564525 53624 564530 53680
rect 564586 53624 574742 53680
rect 574798 53624 574803 53680
rect 564525 53622 574803 53624
rect 564525 53619 564591 53622
rect 574737 53619 574803 53622
rect 461945 53138 462011 53141
rect 472801 53138 472867 53141
rect 461945 53136 472867 53138
rect 461945 53080 461950 53136
rect 462006 53080 472806 53136
rect 472862 53080 472867 53136
rect 461945 53078 472867 53080
rect 461945 53075 462011 53078
rect 472801 53075 472867 53078
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661769 47791 661835 47794
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47789 661835 47791
rect 661388 47733 661774 47789
rect 661830 47733 661835 47789
rect 661388 47731 661835 47733
rect 661769 47728 661835 47731
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 458214 44372 458220 44436
rect 458284 44434 458290 44436
rect 459185 44434 459251 44437
rect 458284 44432 459251 44434
rect 458284 44376 459190 44432
rect 459246 44376 459251 44432
rect 458284 44374 459251 44376
rect 458284 44372 458290 44374
rect 459185 44371 459251 44374
rect 461342 44372 461348 44436
rect 461412 44434 461418 44436
rect 461945 44434 462011 44437
rect 461412 44432 462011 44434
rect 461412 44376 461950 44432
rect 462006 44376 462011 44432
rect 461412 44374 462011 44376
rect 461412 44372 461418 44374
rect 461945 44371 462011 44374
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462497 44434 462563 44437
rect 462332 44432 462563 44434
rect 462332 44376 462502 44432
rect 462558 44376 462563 44432
rect 462332 44374 462563 44376
rect 462332 44372 462338 44374
rect 462497 44371 462563 44374
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 255865 44162 255931 44165
rect 460105 44162 460171 44165
rect 463877 44162 463943 44165
rect 255865 44160 460171 44162
rect 255865 44104 255870 44160
rect 255926 44104 460110 44160
rect 460166 44104 460171 44160
rect 255865 44102 460171 44104
rect 255865 44099 255931 44102
rect 460105 44099 460171 44102
rect 460890 44160 463943 44162
rect 460890 44104 463882 44160
rect 463938 44104 463943 44160
rect 460890 44102 463943 44104
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 307293 43890 307359 43893
rect 440233 43890 440299 43893
rect 307293 43888 440299 43890
rect 307293 43832 307298 43888
rect 307354 43832 440238 43888
rect 440294 43832 440299 43888
rect 307293 43830 440299 43832
rect 307293 43827 307359 43830
rect 440233 43827 440299 43830
rect 441061 43890 441127 43893
rect 460890 43890 460950 44102
rect 463877 44099 463943 44102
rect 441061 43888 460950 43890
rect 441061 43832 441066 43888
rect 441122 43832 460950 43888
rect 441061 43830 460950 43832
rect 441061 43827 441127 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 446213 42258 446279 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 405641 41852 405707 41853
rect 405590 41850 405596 41852
rect 405550 41790 405596 41850
rect 405660 41848 405707 41852
rect 405702 41792 405707 41848
rect 405590 41788 405596 41790
rect 405660 41788 405707 41792
rect 405641 41787 405707 41788
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446213 42256 461183 42258
rect 446213 42200 446218 42256
rect 446274 42200 461122 42256
rect 461178 42200 461183 42256
rect 446213 42198 461183 42200
rect 446213 42195 446279 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 446213 41578 446279 41581
rect 427770 41576 446279 41578
rect 427770 41520 446218 41576
rect 446274 41520 446279 41576
rect 427770 41518 446279 41520
rect 446213 41515 446279 41518
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 675708 892196 675772 892260
rect 675892 887708 675956 887772
rect 675524 887436 675588 887500
rect 676628 882600 676692 882604
rect 676628 882544 676678 882600
rect 676678 882544 676692 882600
rect 676628 882540 676692 882544
rect 675708 881860 675772 881924
rect 675524 876480 675588 876484
rect 675524 876424 675538 876480
rect 675538 876424 675588 876480
rect 675524 876420 675588 876424
rect 675524 873488 675588 873492
rect 675524 873432 675574 873488
rect 675574 873432 675588 873488
rect 675524 873428 675588 873432
rect 676260 869756 676324 869820
rect 676628 868668 676692 868732
rect 675708 867172 675772 867236
rect 675892 865676 675956 865740
rect 676076 865404 676140 865468
rect 41828 813180 41892 813244
rect 41828 811956 41892 812020
rect 41828 809296 41892 809300
rect 41828 809240 41842 809296
rect 41842 809240 41892 809296
rect 41828 809236 41892 809240
rect 40724 805564 40788 805628
rect 40908 805156 40972 805220
rect 40540 804884 40604 804948
rect 42012 801484 42076 801548
rect 41276 801212 41340 801276
rect 41092 800804 41156 800868
rect 40356 800532 40420 800596
rect 41092 796860 41156 796924
rect 41276 796180 41340 796244
rect 42012 794472 42076 794476
rect 42012 794416 42062 794472
rect 42062 794416 42076 794472
rect 42012 794412 42076 794416
rect 40356 793052 40420 793116
rect 40908 790604 40972 790668
rect 41644 790196 41708 790260
rect 40540 789380 40604 789444
rect 41828 789108 41892 789172
rect 40724 788700 40788 788764
rect 41460 788156 41524 788220
rect 675340 788080 675404 788084
rect 675340 788024 675390 788080
rect 675390 788024 675404 788080
rect 675340 788020 675404 788024
rect 675524 786720 675588 786724
rect 675524 786664 675538 786720
rect 675538 786664 675588 786720
rect 675524 786660 675588 786664
rect 674236 783804 674300 783868
rect 676996 779860 677060 779924
rect 41460 769796 41524 769860
rect 40724 766532 40788 766596
rect 40540 765308 40604 765372
rect 40908 764900 40972 764964
rect 41644 759052 41708 759116
rect 40356 757692 40420 757756
rect 41828 757692 41892 757756
rect 40356 755108 40420 755172
rect 40908 754836 40972 754900
rect 42012 754836 42076 754900
rect 40724 752116 40788 752180
rect 42380 752116 42444 752180
rect 42012 750408 42076 750412
rect 42012 750352 42026 750408
rect 42026 750352 42076 750408
rect 42012 750348 42076 750352
rect 42380 749592 42444 749596
rect 42380 749536 42430 749592
rect 42430 749536 42444 749592
rect 42380 749532 42444 749536
rect 40540 749396 40604 749460
rect 41644 745588 41708 745652
rect 41460 745316 41524 745380
rect 41828 744908 41892 744972
rect 674420 742460 674484 742524
rect 674788 742248 674852 742252
rect 674788 742192 674838 742248
rect 674838 742192 674852 742248
rect 674788 742188 674852 742192
rect 674604 738108 674668 738172
rect 674788 734980 674852 735044
rect 676812 732940 676876 733004
rect 675524 728316 675588 728380
rect 675340 728044 675404 728108
rect 674236 726412 674300 726476
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 675156 723148 675220 723212
rect 40724 721708 40788 721772
rect 674972 721712 675036 721716
rect 674972 721656 675022 721712
rect 675022 721656 675036 721712
rect 674972 721652 675036 721656
rect 40540 718524 40604 718588
rect 41644 718252 41708 718316
rect 41828 716076 41892 716140
rect 41276 714232 41340 714236
rect 41276 714176 41290 714232
rect 41290 714176 41340 714232
rect 41276 714172 41340 714176
rect 41276 712132 41340 712196
rect 677180 707950 677244 708014
rect 40724 707100 40788 707164
rect 40540 704244 40604 704308
rect 41828 702068 41892 702132
rect 41644 701796 41708 701860
rect 41460 700436 41524 700500
rect 674236 696628 674300 696692
rect 675340 686156 675404 686220
rect 41460 684626 41524 684690
rect 41828 683844 41892 683908
rect 41828 683572 41892 683636
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 676076 678948 676140 679012
rect 41828 678872 41892 678876
rect 41828 678816 41842 678872
rect 41842 678816 41892 678872
rect 41828 678812 41892 678816
rect 40908 677750 40972 677754
rect 40908 677694 40958 677750
rect 40958 677694 40972 677750
rect 40908 677690 40972 677694
rect 41828 672692 41892 672756
rect 41092 672420 41156 672484
rect 40356 671468 40420 671532
rect 41092 669020 41156 669084
rect 40356 666300 40420 666364
rect 40908 665212 40972 665276
rect 674420 664396 674484 664460
rect 40724 664124 40788 664188
rect 676812 663308 676876 663372
rect 40540 662764 40604 662828
rect 674604 662356 674668 662420
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 41460 657188 41524 657252
rect 675340 644812 675404 644876
rect 44220 642228 44284 642292
rect 41460 640596 41524 640660
rect 675340 640384 675404 640388
rect 675340 640328 675354 640384
rect 675354 640328 675404 640384
rect 675340 640324 675404 640328
rect 41644 639372 41708 639436
rect 40540 637332 40604 637396
rect 674236 636788 674300 636852
rect 40724 635292 40788 635356
rect 40908 634884 40972 634948
rect 675156 631348 675220 631412
rect 41828 629852 41892 629916
rect 676076 629716 676140 629780
rect 42380 624744 42444 624748
rect 42380 624688 42430 624744
rect 42430 624688 42444 624744
rect 42380 624684 42444 624688
rect 40908 623732 40972 623796
rect 40724 620740 40788 620804
rect 42380 620740 42444 620804
rect 40540 619788 40604 619852
rect 41460 616252 41524 616316
rect 673868 616116 673932 616180
rect 41828 615980 41892 616044
rect 41644 615436 41708 615500
rect 676812 604692 676876 604756
rect 674236 602924 674300 602988
rect 44220 599660 44284 599724
rect 43116 599252 43180 599316
rect 42012 597212 42076 597276
rect 43116 597000 43180 597004
rect 43116 596944 43130 597000
rect 43130 596944 43180 597000
rect 43116 596940 43180 596944
rect 41828 593948 41892 594012
rect 675156 592860 675220 592924
rect 40724 592486 40788 592550
rect 41828 592316 41892 592380
rect 42196 591228 42260 591292
rect 676076 590548 676140 590612
rect 675892 586196 675956 586260
rect 42012 586120 42076 586124
rect 42012 586064 42026 586120
rect 42026 586064 42076 586120
rect 42012 586060 42076 586064
rect 41828 585108 41892 585172
rect 41092 584836 41156 584900
rect 40356 584564 40420 584628
rect 676076 584564 676140 584628
rect 40356 581572 40420 581636
rect 41092 580212 41156 580276
rect 40908 577764 40972 577828
rect 40540 575724 40604 575788
rect 40724 574636 40788 574700
rect 41460 572732 41524 572796
rect 42012 572248 42076 572252
rect 42012 572192 42026 572248
rect 42026 572192 42076 572248
rect 42012 572188 42076 572192
rect 41644 571508 41708 571572
rect 676812 570692 676876 570756
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675340 563136 675404 563140
rect 675340 563080 675390 563136
rect 675390 563080 675404 563136
rect 675340 563076 675404 563080
rect 674420 558996 674484 559060
rect 41092 558724 41156 558788
rect 41092 557488 41156 557552
rect 41828 553964 41892 554028
rect 676812 553964 676876 554028
rect 41828 552740 41892 552804
rect 41828 550624 41892 550628
rect 41828 550568 41842 550624
rect 41842 550568 41892 550624
rect 41828 550564 41892 550568
rect 676996 550292 677060 550356
rect 675892 547572 675956 547636
rect 674236 547028 674300 547092
rect 676076 546756 676140 546820
rect 40724 545668 40788 545732
rect 675340 545532 675404 545596
rect 40540 545396 40604 545460
rect 40540 537372 40604 537436
rect 40724 536964 40788 537028
rect 41460 530708 41524 530772
rect 41828 529484 41892 529548
rect 41644 529212 41708 529276
rect 676996 503644 677060 503708
rect 675892 488820 675956 488884
rect 675892 487868 675956 487932
rect 674420 484740 674484 484804
rect 675892 483516 675956 483580
rect 673868 455228 673932 455292
rect 675340 447748 675404 447812
rect 41828 426396 41892 426460
rect 42012 424764 42076 424828
rect 42196 424220 42260 424284
rect 41828 422724 41892 422788
rect 41828 421908 41892 421972
rect 41460 418780 41524 418844
rect 41644 413340 41708 413404
rect 42196 413340 42260 413404
rect 675340 410484 675404 410548
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40908 405588 40972 405652
rect 41828 401840 41892 401844
rect 41828 401784 41842 401840
rect 41842 401784 41892 401840
rect 41828 401780 41892 401784
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 40540 400012 40604 400076
rect 41460 398788 41524 398852
rect 676076 398788 676140 398852
rect 676628 396748 676692 396812
rect 676444 396340 676508 396404
rect 676260 395116 676324 395180
rect 675892 392804 675956 392868
rect 675708 388452 675772 388516
rect 676628 385324 676692 385388
rect 676444 382196 676508 382260
rect 40540 380564 40604 380628
rect 41460 379808 41524 379812
rect 41460 379752 41510 379808
rect 41510 379752 41524 379808
rect 41460 379748 41524 379752
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40724 378116 40788 378180
rect 676260 377436 676324 377500
rect 41276 374580 41340 374644
rect 676076 373628 676140 373692
rect 41644 372676 41708 372740
rect 675892 372948 675956 373012
rect 41828 371860 41892 371924
rect 41276 368460 41340 368524
rect 40724 363700 40788 363764
rect 41828 360088 41892 360092
rect 41828 360032 41842 360088
rect 41842 360032 41892 360088
rect 41828 360028 41892 360032
rect 41644 359484 41708 359548
rect 41460 358668 41524 358732
rect 40540 356084 40604 356148
rect 675524 353364 675588 353428
rect 675708 352956 675772 353020
rect 675938 352140 676002 352204
rect 675892 351928 675956 351932
rect 675892 351872 675906 351928
rect 675906 351872 675956 351928
rect 675892 351868 675956 351872
rect 676444 346624 676508 346628
rect 676444 346568 676494 346624
rect 676494 346568 676508 346624
rect 676444 346564 676508 346568
rect 676812 346156 676876 346220
rect 44404 342892 44468 342956
rect 44220 341532 44284 341596
rect 675524 340776 675588 340780
rect 675524 340720 675574 340776
rect 675574 340720 675588 340776
rect 675524 340716 675588 340720
rect 42748 340444 42812 340508
rect 44588 340172 44652 340236
rect 676444 340172 676508 340236
rect 41644 338132 41708 338196
rect 675892 337724 675956 337788
rect 42932 337588 42996 337652
rect 43116 337180 43180 337244
rect 40724 336908 40788 336972
rect 42012 336500 42076 336564
rect 41828 335684 41892 335748
rect 40540 335276 40604 335340
rect 40908 333644 40972 333708
rect 676076 328340 676140 328404
rect 676260 325484 676324 325548
rect 40908 325348 40972 325412
rect 676812 325212 676876 325276
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 41828 319968 41892 319972
rect 41828 319912 41878 319968
rect 41878 319912 41892 319968
rect 41828 319908 41892 319912
rect 40724 318956 40788 319020
rect 40540 317324 40604 317388
rect 43116 315964 43180 316028
rect 42012 313712 42076 313716
rect 42012 313656 42062 313712
rect 42062 313656 42076 313712
rect 42012 313652 42076 313656
rect 42932 312700 42996 312764
rect 675708 309028 675772 309092
rect 675708 308756 675772 308820
rect 675892 307124 675956 307188
rect 676628 304506 676692 304570
rect 676444 300596 676508 300660
rect 44404 300052 44468 300116
rect 675708 299372 675772 299436
rect 44588 299236 44652 299300
rect 44220 298420 44284 298484
rect 42748 297604 42812 297668
rect 675524 297332 675588 297396
rect 42012 296788 42076 296852
rect 676260 294476 676324 294540
rect 40540 292528 40604 292592
rect 675524 292224 675588 292228
rect 675524 292168 675574 292224
rect 675574 292168 675588 292224
rect 675524 292164 675588 292168
rect 41828 291484 41892 291548
rect 676444 291484 676508 291548
rect 676628 290804 676692 290868
rect 40724 289172 40788 289236
rect 41644 284820 41708 284884
rect 42012 284276 42076 284340
rect 675892 283596 675956 283660
rect 675708 282840 675772 282844
rect 675708 282784 675722 282840
rect 675722 282784 675772 282840
rect 675708 282780 675772 282784
rect 676076 281148 676140 281212
rect 40908 278428 40972 278492
rect 40724 277068 40788 277132
rect 40540 274212 40604 274276
rect 42012 272368 42076 272372
rect 42012 272312 42026 272368
rect 42026 272312 42076 272368
rect 42012 272308 42076 272312
rect 41460 270404 41524 270468
rect 41828 270056 41892 270060
rect 41828 270000 41878 270056
rect 41878 270000 41892 270056
rect 41828 269996 41892 270000
rect 674972 264148 675036 264212
rect 676076 263604 676140 263668
rect 676812 261564 676876 261628
rect 676996 259932 677060 259996
rect 40540 250140 40604 250204
rect 676812 250140 676876 250204
rect 40724 249732 40788 249796
rect 674972 249732 675036 249796
rect 676076 249596 676140 249660
rect 676996 242252 677060 242316
rect 676812 241980 676876 242044
rect 674972 241708 675036 241772
rect 42012 237356 42076 237420
rect 40724 236540 40788 236604
rect 40540 230420 40604 230484
rect 674972 230148 675036 230212
rect 674052 229740 674116 229804
rect 42012 228984 42076 228988
rect 42012 228928 42026 228984
rect 42026 228928 42076 228984
rect 42012 228924 42076 228928
rect 672948 227020 673012 227084
rect 673500 223620 673564 223684
rect 561628 222184 561692 222188
rect 561628 222128 561678 222184
rect 561678 222128 561692 222184
rect 561628 222124 561692 222128
rect 675892 220628 675956 220692
rect 561628 219132 561692 219196
rect 675892 218316 675956 218380
rect 509188 217772 509252 217836
rect 510108 217832 510172 217836
rect 510108 217776 510158 217832
rect 510158 217776 510172 217832
rect 510108 217772 510172 217776
rect 522620 217832 522684 217836
rect 522620 217776 522634 217832
rect 522634 217776 522684 217832
rect 522620 217772 522684 217776
rect 574324 217772 574388 217836
rect 675708 217364 675772 217428
rect 493732 217288 493796 217292
rect 493732 217232 493782 217288
rect 493782 217232 493796 217288
rect 493732 217228 493796 217232
rect 574324 216744 574388 216748
rect 574324 216688 574374 216744
rect 574374 216688 574388 216744
rect 574324 216684 574388 216688
rect 561628 216140 561692 216204
rect 509188 215868 509252 215932
rect 522620 215324 522684 215388
rect 675892 215188 675956 215252
rect 675892 214372 675956 214436
rect 670188 213828 670252 213892
rect 670188 213012 670252 213076
rect 676260 210836 676324 210900
rect 676628 210836 676692 210900
rect 675892 210564 675956 210628
rect 670740 210428 670804 210492
rect 41828 210020 41892 210084
rect 672580 208312 672644 208316
rect 672580 208256 672630 208312
rect 672630 208256 672644 208312
rect 672580 208252 672644 208256
rect 41644 208116 41708 208180
rect 40540 207300 40604 207364
rect 676076 206892 676140 206956
rect 40724 206484 40788 206548
rect 40908 206076 40972 206140
rect 41460 205668 41524 205732
rect 676444 205532 676508 205596
rect 676076 204172 676140 204236
rect 672580 202540 672644 202604
rect 676260 200772 676324 200836
rect 675708 198384 675772 198388
rect 675708 198328 675758 198384
rect 675758 198328 675772 198384
rect 675708 198324 675772 198328
rect 676628 196148 676692 196212
rect 41828 195256 41892 195260
rect 41828 195200 41878 195256
rect 41878 195200 41892 195256
rect 41828 195196 41892 195200
rect 40908 194924 40972 194988
rect 40724 193156 40788 193220
rect 675892 192748 675956 192812
rect 40540 186356 40604 186420
rect 41828 186008 41892 186012
rect 41828 185952 41842 186008
rect 41842 185952 41892 186008
rect 41828 185948 41892 185952
rect 41460 184044 41524 184108
rect 675524 173572 675588 173636
rect 675892 172756 675956 172820
rect 675708 172348 675772 172412
rect 675340 171124 675404 171188
rect 669452 169628 669516 169692
rect 675892 169628 675956 169692
rect 675708 167452 675772 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 675524 162148 675588 162212
rect 676076 162148 676140 162212
rect 675340 157040 675404 157044
rect 675340 156984 675390 157040
rect 675390 156984 675404 157040
rect 675340 156980 675404 156984
rect 676444 156980 676508 157044
rect 676260 155756 676324 155820
rect 675892 153036 675956 153100
rect 676628 151404 676692 151468
rect 676076 148412 676140 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 669268 140388 669332 140452
rect 672948 133316 673012 133380
rect 673500 132772 673564 132836
rect 676444 128556 676508 128620
rect 676260 128148 676324 128212
rect 676076 126924 676140 126988
rect 670740 125700 670804 125764
rect 675708 122844 675772 122908
rect 676812 121620 676876 121684
rect 675892 116452 675956 116516
rect 674052 115772 674116 115836
rect 676444 114140 676508 114204
rect 676812 111692 676876 111756
rect 675708 111344 675772 111348
rect 675708 111288 675722 111344
rect 675722 111288 675772 111344
rect 675708 111284 675772 111288
rect 676076 108156 676140 108220
rect 675892 104756 675956 104820
rect 676260 103124 676324 103188
rect 635780 96868 635844 96932
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95916 634004 95980
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 635780 78100 635844 78164
rect 637068 77556 637132 77620
rect 461716 54980 461780 55044
rect 462636 54708 462700 54772
rect 461716 53892 461780 53956
rect 462636 53892 462700 53956
rect 194364 50220 194428 50284
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 458220 44372 458284 44436
rect 461348 44372 461412 44436
rect 462268 44372 462332 44436
rect 141740 43964 141804 44028
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 405596 41848 405660 41852
rect 405596 41792 405646 41848
rect 405646 41792 405660 41848
rect 405596 41788 405660 41792
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 675707 892260 675773 892261
rect 675707 892196 675708 892260
rect 675772 892196 675773 892260
rect 675707 892195 675773 892196
rect 675523 887500 675589 887501
rect 675523 887436 675524 887500
rect 675588 887436 675589 887500
rect 675523 887435 675589 887436
rect 675526 882330 675586 887435
rect 675710 886410 675770 892195
rect 675891 887772 675957 887773
rect 675891 887708 675892 887772
rect 675956 887708 675957 887772
rect 675891 887707 675957 887708
rect 675894 887090 675954 887707
rect 675894 887030 676322 887090
rect 675710 886350 676138 886410
rect 675526 882270 675954 882330
rect 675707 881924 675773 881925
rect 675707 881860 675708 881924
rect 675772 881860 675773 881924
rect 675707 881859 675773 881860
rect 675523 876484 675589 876485
rect 675523 876420 675524 876484
rect 675588 876420 675589 876484
rect 675523 876419 675589 876420
rect 675526 873493 675586 876419
rect 675523 873492 675589 873493
rect 675523 873428 675524 873492
rect 675588 873428 675589 873492
rect 675523 873427 675589 873428
rect 675710 867237 675770 881859
rect 675707 867236 675773 867237
rect 675707 867172 675708 867236
rect 675772 867172 675773 867236
rect 675707 867171 675773 867172
rect 675894 865741 675954 882270
rect 675891 865740 675957 865741
rect 675891 865676 675892 865740
rect 675956 865676 675957 865740
rect 675891 865675 675957 865676
rect 676078 865469 676138 886350
rect 676262 869821 676322 887030
rect 676627 882604 676693 882605
rect 676627 882540 676628 882604
rect 676692 882540 676693 882604
rect 676627 882539 676693 882540
rect 676259 869820 676325 869821
rect 676259 869756 676260 869820
rect 676324 869756 676325 869820
rect 676259 869755 676325 869756
rect 676630 868733 676690 882539
rect 676627 868732 676693 868733
rect 676627 868668 676628 868732
rect 676692 868668 676693 868732
rect 676627 868667 676693 868668
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40723 805628 40789 805629
rect 40723 805564 40724 805628
rect 40788 805564 40789 805628
rect 40723 805563 40789 805564
rect 40539 804948 40605 804949
rect 40539 804884 40540 804948
rect 40604 804884 40605 804948
rect 40539 804883 40605 804884
rect 40355 800596 40421 800597
rect 40355 800532 40356 800596
rect 40420 800532 40421 800596
rect 40355 800531 40421 800532
rect 40358 793117 40418 800531
rect 40355 793116 40421 793117
rect 40355 793052 40356 793116
rect 40420 793052 40421 793116
rect 40355 793051 40421 793052
rect 40542 789445 40602 804883
rect 40539 789444 40605 789445
rect 40539 789380 40540 789444
rect 40604 789380 40605 789444
rect 40539 789379 40605 789380
rect 40726 788765 40786 805563
rect 40907 805220 40973 805221
rect 40907 805156 40908 805220
rect 40972 805156 40973 805220
rect 40907 805155 40973 805156
rect 40910 790669 40970 805155
rect 41275 801276 41341 801277
rect 41275 801212 41276 801276
rect 41340 801212 41341 801276
rect 41275 801211 41341 801212
rect 41091 800868 41157 800869
rect 41091 800804 41092 800868
rect 41156 800804 41157 800868
rect 41091 800803 41157 800804
rect 41094 796925 41154 800803
rect 41091 796924 41157 796925
rect 41091 796860 41092 796924
rect 41156 796860 41157 796924
rect 41091 796859 41157 796860
rect 41278 796245 41338 801211
rect 41275 796244 41341 796245
rect 41275 796180 41276 796244
rect 41340 796180 41341 796244
rect 41275 796179 41341 796180
rect 40907 790668 40973 790669
rect 40907 790604 40908 790668
rect 40972 790604 40973 790668
rect 40907 790603 40973 790604
rect 40723 788764 40789 788765
rect 40723 788700 40724 788764
rect 40788 788700 40789 788764
rect 40723 788699 40789 788700
rect 41462 788221 41522 812910
rect 41827 812020 41893 812021
rect 41827 811956 41828 812020
rect 41892 811956 41893 812020
rect 41827 811955 41893 811956
rect 41830 811610 41890 811955
rect 41646 811550 41890 811610
rect 41646 790261 41706 811550
rect 41827 809300 41893 809301
rect 41827 809236 41828 809300
rect 41892 809236 41893 809300
rect 41827 809235 41893 809236
rect 41643 790260 41709 790261
rect 41643 790196 41644 790260
rect 41708 790196 41709 790260
rect 41643 790195 41709 790196
rect 41830 789173 41890 809235
rect 42011 801548 42077 801549
rect 42011 801484 42012 801548
rect 42076 801484 42077 801548
rect 42011 801483 42077 801484
rect 42014 794477 42074 801483
rect 42011 794476 42077 794477
rect 42011 794412 42012 794476
rect 42076 794412 42077 794476
rect 42011 794411 42077 794412
rect 41827 789172 41893 789173
rect 41827 789108 41828 789172
rect 41892 789108 41893 789172
rect 41827 789107 41893 789108
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 675339 788084 675405 788085
rect 675339 788020 675340 788084
rect 675404 788020 675405 788084
rect 675339 788019 675405 788020
rect 674235 783868 674301 783869
rect 674235 783804 674236 783868
rect 674300 783804 674301 783868
rect 674235 783803 674301 783804
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40723 766596 40789 766597
rect 40723 766532 40724 766596
rect 40788 766532 40789 766596
rect 40723 766531 40789 766532
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757756 40421 757757
rect 40355 757692 40356 757756
rect 40420 757692 40421 757756
rect 40355 757691 40421 757692
rect 40358 755173 40418 757691
rect 40355 755172 40421 755173
rect 40355 755108 40356 755172
rect 40420 755108 40421 755172
rect 40355 755107 40421 755108
rect 40542 749461 40602 765307
rect 40726 752181 40786 766531
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40910 754901 40970 764899
rect 40907 754900 40973 754901
rect 40907 754836 40908 754900
rect 40972 754836 40973 754900
rect 40907 754835 40973 754836
rect 40723 752180 40789 752181
rect 40723 752116 40724 752180
rect 40788 752116 40789 752180
rect 40723 752115 40789 752116
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 745381 41522 769795
rect 41643 759116 41709 759117
rect 41643 759052 41644 759116
rect 41708 759052 41709 759116
rect 41643 759051 41709 759052
rect 41646 745653 41706 759051
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41643 745652 41709 745653
rect 41643 745588 41644 745652
rect 41708 745588 41709 745652
rect 41643 745587 41709 745588
rect 41459 745380 41525 745381
rect 41459 745316 41460 745380
rect 41524 745316 41525 745380
rect 41459 745315 41525 745316
rect 41830 744973 41890 757691
rect 42011 754900 42077 754901
rect 42011 754836 42012 754900
rect 42076 754836 42077 754900
rect 42011 754835 42077 754836
rect 42014 750413 42074 754835
rect 42379 752180 42445 752181
rect 42379 752116 42380 752180
rect 42444 752116 42445 752180
rect 42379 752115 42445 752116
rect 42011 750412 42077 750413
rect 42011 750348 42012 750412
rect 42076 750348 42077 750412
rect 42011 750347 42077 750348
rect 42382 749597 42442 752115
rect 42379 749596 42445 749597
rect 42379 749532 42380 749596
rect 42444 749532 42445 749596
rect 42379 749531 42445 749532
rect 41827 744972 41893 744973
rect 41827 744908 41828 744972
rect 41892 744908 41893 744972
rect 41827 744907 41893 744908
rect 674238 726477 674298 783803
rect 674419 742524 674485 742525
rect 674419 742460 674420 742524
rect 674484 742460 674485 742524
rect 674419 742459 674485 742460
rect 674235 726476 674301 726477
rect 674235 726412 674236 726476
rect 674300 726412 674301 726476
rect 674235 726411 674301 726412
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 704309 40602 718523
rect 40726 707165 40786 721707
rect 41275 714236 41341 714237
rect 41275 714172 41276 714236
rect 41340 714172 41341 714236
rect 41275 714171 41341 714172
rect 41278 712197 41338 714171
rect 41275 712196 41341 712197
rect 41275 712132 41276 712196
rect 41340 712132 41341 712196
rect 41275 712131 41341 712132
rect 40723 707164 40789 707165
rect 40723 707100 40724 707164
rect 40788 707100 40789 707164
rect 40723 707099 40789 707100
rect 40539 704308 40605 704309
rect 40539 704244 40540 704308
rect 40604 704244 40605 704308
rect 40539 704243 40605 704244
rect 41462 700501 41522 725190
rect 41643 718316 41709 718317
rect 41643 718252 41644 718316
rect 41708 718252 41709 718316
rect 41643 718251 41709 718252
rect 41646 701861 41706 718251
rect 41827 716140 41893 716141
rect 41827 716076 41828 716140
rect 41892 716076 41893 716140
rect 41827 716075 41893 716076
rect 41830 702133 41890 716075
rect 41827 702132 41893 702133
rect 41827 702068 41828 702132
rect 41892 702068 41893 702132
rect 41827 702067 41893 702068
rect 41643 701860 41709 701861
rect 41643 701796 41644 701860
rect 41708 701796 41709 701860
rect 41643 701795 41709 701796
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 674235 696692 674301 696693
rect 674235 696628 674236 696692
rect 674300 696628 674301 696692
rect 674235 696627 674301 696628
rect 41459 684690 41525 684691
rect 41459 684626 41460 684690
rect 41524 684626 41525 684690
rect 41459 684625 41525 684626
rect 41462 684450 41522 684625
rect 41462 684390 41890 684450
rect 41830 683909 41890 684390
rect 41827 683908 41893 683909
rect 41827 683844 41828 683908
rect 41892 683844 41893 683908
rect 41827 683843 41893 683844
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683090 41890 683571
rect 41646 683030 41890 683090
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 41646 678990 41706 683030
rect 40723 678927 40789 678928
rect 41462 678930 41706 678990
rect 40355 671532 40421 671533
rect 40355 671468 40356 671532
rect 40420 671468 40421 671532
rect 40355 671467 40421 671468
rect 40358 666365 40418 671467
rect 40355 666364 40421 666365
rect 40355 666300 40356 666364
rect 40420 666300 40421 666364
rect 40355 666299 40421 666300
rect 40542 662829 40602 678927
rect 40726 664189 40786 678927
rect 40907 677754 40973 677755
rect 40907 677690 40908 677754
rect 40972 677690 40973 677754
rect 40907 677689 40973 677690
rect 40910 665277 40970 677689
rect 41091 672484 41157 672485
rect 41091 672420 41092 672484
rect 41156 672420 41157 672484
rect 41091 672419 41157 672420
rect 41094 669085 41154 672419
rect 41091 669084 41157 669085
rect 41091 669020 41092 669084
rect 41156 669020 41157 669084
rect 41091 669019 41157 669020
rect 40907 665276 40973 665277
rect 40907 665212 40908 665276
rect 40972 665212 40973 665276
rect 40907 665211 40973 665212
rect 40723 664188 40789 664189
rect 40723 664124 40724 664188
rect 40788 664124 40789 664188
rect 40723 664123 40789 664124
rect 40539 662828 40605 662829
rect 40539 662764 40540 662828
rect 40604 662764 40605 662828
rect 40539 662763 40605 662764
rect 41462 657253 41522 678930
rect 41827 678876 41893 678877
rect 41827 678812 41828 678876
rect 41892 678812 41893 678876
rect 41827 678811 41893 678812
rect 41830 678330 41890 678811
rect 41646 678270 41890 678330
rect 41646 658613 41706 678270
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 44219 642292 44285 642293
rect 44219 642228 44220 642292
rect 44284 642228 44285 642292
rect 44219 642227 44285 642228
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 637396 40605 637397
rect 40539 637332 40540 637396
rect 40604 637332 40605 637396
rect 40539 637331 40605 637332
rect 40542 619853 40602 637331
rect 40723 635356 40789 635357
rect 40723 635292 40724 635356
rect 40788 635292 40789 635356
rect 40723 635291 40789 635292
rect 40726 620805 40786 635291
rect 40907 634948 40973 634949
rect 40907 634884 40908 634948
rect 40972 634884 40973 634948
rect 40907 634883 40973 634884
rect 40910 623797 40970 634883
rect 40907 623796 40973 623797
rect 40907 623732 40908 623796
rect 40972 623732 40973 623796
rect 40907 623731 40973 623732
rect 40723 620804 40789 620805
rect 40723 620740 40724 620804
rect 40788 620740 40789 620804
rect 40723 620739 40789 620740
rect 40539 619852 40605 619853
rect 40539 619788 40540 619852
rect 40604 619788 40605 619852
rect 40539 619787 40605 619788
rect 41462 616317 41522 640595
rect 41643 639436 41709 639437
rect 41643 639372 41644 639436
rect 41708 639372 41709 639436
rect 41643 639371 41709 639372
rect 41459 616316 41525 616317
rect 41459 616252 41460 616316
rect 41524 616252 41525 616316
rect 41459 616251 41525 616252
rect 41646 615501 41706 639371
rect 41827 629916 41893 629917
rect 41827 629852 41828 629916
rect 41892 629852 41893 629916
rect 41827 629851 41893 629852
rect 41830 616045 41890 629851
rect 42379 624748 42445 624749
rect 42379 624684 42380 624748
rect 42444 624684 42445 624748
rect 42379 624683 42445 624684
rect 42382 620805 42442 624683
rect 42379 620804 42445 620805
rect 42379 620740 42380 620804
rect 42444 620740 42445 620804
rect 42379 620739 42445 620740
rect 41827 616044 41893 616045
rect 41827 615980 41828 616044
rect 41892 615980 41893 616044
rect 41827 615979 41893 615980
rect 41643 615500 41709 615501
rect 41643 615436 41644 615500
rect 41708 615436 41709 615500
rect 41643 615435 41709 615436
rect 44222 599725 44282 642227
rect 674238 636853 674298 696627
rect 674422 664461 674482 742459
rect 674787 742252 674853 742253
rect 674787 742188 674788 742252
rect 674852 742188 674853 742252
rect 674787 742187 674853 742188
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674419 664460 674485 664461
rect 674419 664396 674420 664460
rect 674484 664396 674485 664460
rect 674419 664395 674485 664396
rect 674606 662421 674666 738107
rect 674790 735045 674850 742187
rect 674787 735044 674853 735045
rect 674787 734980 674788 735044
rect 674852 734980 674853 735044
rect 674787 734979 674853 734980
rect 675342 728109 675402 788019
rect 675523 786724 675589 786725
rect 675523 786660 675524 786724
rect 675588 786660 675589 786724
rect 675523 786659 675589 786660
rect 675526 728381 675586 786659
rect 676995 779924 677061 779925
rect 676995 779860 676996 779924
rect 677060 779860 677061 779924
rect 676995 779859 677061 779860
rect 676811 733004 676877 733005
rect 676811 732940 676812 733004
rect 676876 732940 676877 733004
rect 676811 732939 676877 732940
rect 675523 728380 675589 728381
rect 675523 728316 675524 728380
rect 675588 728316 675589 728380
rect 675523 728315 675589 728316
rect 675339 728108 675405 728109
rect 675339 728044 675340 728108
rect 675404 728044 675405 728108
rect 675339 728043 675405 728044
rect 675155 723212 675221 723213
rect 675155 723148 675156 723212
rect 675220 723148 675221 723212
rect 675155 723147 675221 723148
rect 674971 721716 675037 721717
rect 674971 721652 674972 721716
rect 675036 721652 675037 721716
rect 674971 721651 675037 721652
rect 674974 717630 675034 721651
rect 675158 721170 675218 723147
rect 675158 721110 675586 721170
rect 675526 717630 675586 721110
rect 674974 717570 675402 717630
rect 675526 717570 676138 717630
rect 675342 686221 675402 717570
rect 675339 686220 675405 686221
rect 675339 686156 675340 686220
rect 675404 686156 675405 686220
rect 675339 686155 675405 686156
rect 676078 679013 676138 717570
rect 676075 679012 676141 679013
rect 676075 678948 676076 679012
rect 676140 678948 676141 679012
rect 676075 678947 676141 678948
rect 676814 663373 676874 732939
rect 676998 727290 677058 779859
rect 676998 727230 677242 727290
rect 677182 708015 677242 727230
rect 677179 708014 677245 708015
rect 677179 707950 677180 708014
rect 677244 707950 677245 708014
rect 677179 707949 677245 707950
rect 676811 663372 676877 663373
rect 676811 663308 676812 663372
rect 676876 663308 676877 663372
rect 676811 663307 676877 663308
rect 674603 662420 674669 662421
rect 674603 662356 674604 662420
rect 674668 662356 674669 662420
rect 674603 662355 674669 662356
rect 675339 644876 675405 644877
rect 675339 644812 675340 644876
rect 675404 644812 675405 644876
rect 675339 644811 675405 644812
rect 675342 640389 675402 644811
rect 675339 640388 675405 640389
rect 675339 640324 675340 640388
rect 675404 640324 675405 640388
rect 675339 640323 675405 640324
rect 674235 636852 674301 636853
rect 674235 636788 674236 636852
rect 674300 636788 674301 636852
rect 674235 636787 674301 636788
rect 675155 631412 675221 631413
rect 675155 631348 675156 631412
rect 675220 631348 675221 631412
rect 675155 631347 675221 631348
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 44219 599724 44285 599725
rect 44219 599660 44220 599724
rect 44284 599660 44285 599724
rect 44219 599659 44285 599660
rect 43115 599316 43181 599317
rect 43115 599252 43116 599316
rect 43180 599252 43181 599316
rect 43115 599251 43181 599252
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 594012 41893 594013
rect 41827 594010 41828 594012
rect 40542 593950 41828 594010
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 581637 40418 584563
rect 40355 581636 40421 581637
rect 40355 581572 40356 581636
rect 40420 581572 40421 581636
rect 40355 581571 40421 581572
rect 40542 575789 40602 593950
rect 41827 593948 41828 593950
rect 41892 593948 41893 594012
rect 41827 593947 41893 593948
rect 40723 592550 40789 592551
rect 40723 592486 40724 592550
rect 40788 592486 40789 592550
rect 40723 592485 40789 592486
rect 40539 575788 40605 575789
rect 40539 575724 40540 575788
rect 40604 575724 40605 575788
rect 40539 575723 40605 575724
rect 40726 574701 40786 592485
rect 41827 592380 41893 592381
rect 41827 592316 41828 592380
rect 41892 592316 41893 592380
rect 41827 592315 41893 592316
rect 41830 592050 41890 592315
rect 41462 591990 41890 592050
rect 41462 591970 41522 591990
rect 40910 591910 41522 591970
rect 40910 577829 40970 591910
rect 42014 587210 42074 597211
rect 43118 597005 43178 599251
rect 43115 597004 43181 597005
rect 43115 596940 43116 597004
rect 43180 596940 43181 597004
rect 43115 596939 43181 596940
rect 42195 591292 42261 591293
rect 42195 591228 42196 591292
rect 42260 591228 42261 591292
rect 42195 591227 42261 591228
rect 41462 587150 42074 587210
rect 41091 584900 41157 584901
rect 41091 584836 41092 584900
rect 41156 584836 41157 584900
rect 41091 584835 41157 584836
rect 41094 580277 41154 584835
rect 41091 580276 41157 580277
rect 41091 580212 41092 580276
rect 41156 580212 41157 580276
rect 41091 580211 41157 580212
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 41462 572797 41522 587150
rect 42198 586530 42258 591227
rect 41646 586470 42258 586530
rect 41459 572796 41525 572797
rect 41459 572732 41460 572796
rect 41524 572732 41525 572796
rect 41459 572731 41525 572732
rect 41646 571573 41706 586470
rect 42011 586124 42077 586125
rect 42011 586060 42012 586124
rect 42076 586060 42077 586124
rect 42011 586059 42077 586060
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41643 571572 41709 571573
rect 41643 571508 41644 571572
rect 41708 571508 41709 571572
rect 41643 571507 41709 571508
rect 41830 570213 41890 585107
rect 42014 572253 42074 586059
rect 42011 572252 42077 572253
rect 42011 572188 42012 572252
rect 42076 572188 42077 572252
rect 42011 572187 42077 572188
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41091 558788 41157 558789
rect 41091 558724 41092 558788
rect 41156 558724 41157 558788
rect 41091 558723 41157 558724
rect 41094 557553 41154 558723
rect 41091 557552 41157 557553
rect 41091 557488 41092 557552
rect 41156 557488 41157 557552
rect 41091 557487 41157 557488
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 537437 40602 545395
rect 40539 537436 40605 537437
rect 40539 537372 40540 537436
rect 40604 537372 40605 537436
rect 40539 537371 40605 537372
rect 40726 537029 40786 545667
rect 40723 537028 40789 537029
rect 40723 536964 40724 537028
rect 40788 536964 40789 537028
rect 40723 536963 40789 536964
rect 41462 530773 41522 553350
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41830 552530 41890 552739
rect 41646 552470 41890 552530
rect 41459 530772 41525 530773
rect 41459 530708 41460 530772
rect 41524 530708 41525 530772
rect 41459 530707 41525 530708
rect 41646 529277 41706 552470
rect 41827 550628 41893 550629
rect 41827 550564 41828 550628
rect 41892 550564 41893 550628
rect 41827 550563 41893 550564
rect 41830 529549 41890 550563
rect 41827 529548 41893 529549
rect 41827 529484 41828 529548
rect 41892 529484 41893 529548
rect 41827 529483 41893 529484
rect 41643 529276 41709 529277
rect 41643 529212 41644 529276
rect 41708 529212 41709 529276
rect 41643 529211 41709 529212
rect 673870 455293 673930 616115
rect 674235 602988 674301 602989
rect 674235 602924 674236 602988
rect 674300 602924 674301 602988
rect 674235 602923 674301 602924
rect 674238 547093 674298 602923
rect 675158 592925 675218 631347
rect 676075 629780 676141 629781
rect 676075 629716 676076 629780
rect 676140 629716 676141 629780
rect 676075 629715 676141 629716
rect 675155 592924 675221 592925
rect 675155 592860 675156 592924
rect 675220 592860 675221 592924
rect 675155 592859 675221 592860
rect 676078 590613 676138 629715
rect 676811 604756 676877 604757
rect 676811 604692 676812 604756
rect 676876 604692 676877 604756
rect 676811 604691 676877 604692
rect 676075 590612 676141 590613
rect 676075 590548 676076 590612
rect 676140 590548 676141 590612
rect 676075 590547 676141 590548
rect 675891 586260 675957 586261
rect 675891 586196 675892 586260
rect 675956 586196 675957 586260
rect 675891 586195 675957 586196
rect 675339 563140 675405 563141
rect 675339 563076 675340 563140
rect 675404 563076 675405 563140
rect 675339 563075 675405 563076
rect 674419 559060 674485 559061
rect 674419 558996 674420 559060
rect 674484 558996 674485 559060
rect 674419 558995 674485 558996
rect 674235 547092 674301 547093
rect 674235 547028 674236 547092
rect 674300 547028 674301 547092
rect 674235 547027 674301 547028
rect 674422 484805 674482 558995
rect 675342 545597 675402 563075
rect 675894 547637 675954 586195
rect 676075 584628 676141 584629
rect 676075 584564 676076 584628
rect 676140 584564 676141 584628
rect 676075 584563 676141 584564
rect 675891 547636 675957 547637
rect 675891 547572 675892 547636
rect 675956 547572 675957 547636
rect 675891 547571 675957 547572
rect 676078 546821 676138 584563
rect 676814 570757 676874 604691
rect 676811 570756 676877 570757
rect 676811 570692 676812 570756
rect 676876 570692 676877 570756
rect 676811 570691 676877 570692
rect 676811 554028 676877 554029
rect 676811 553964 676812 554028
rect 676876 553964 676877 554028
rect 676811 553963 676877 553964
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 675339 545596 675405 545597
rect 675339 545532 675340 545596
rect 675404 545532 675405 545596
rect 675339 545531 675405 545532
rect 676814 495450 676874 553963
rect 676995 550356 677061 550357
rect 676995 550292 676996 550356
rect 677060 550292 677061 550356
rect 676995 550291 677061 550292
rect 676998 503709 677058 550291
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676262 495390 676874 495450
rect 676262 489970 676322 495390
rect 675710 489910 676322 489970
rect 675710 485790 675770 489910
rect 675894 489230 676138 489290
rect 675894 488885 675954 489230
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 676078 488610 676138 489230
rect 676078 488550 676506 488610
rect 675891 487932 675957 487933
rect 675891 487868 675892 487932
rect 675956 487930 675957 487932
rect 676446 487930 676506 488550
rect 675956 487870 676322 487930
rect 676446 487870 677058 487930
rect 675956 487868 675957 487870
rect 675891 487867 675957 487868
rect 675710 485730 675954 485790
rect 674419 484804 674485 484805
rect 674419 484740 674420 484804
rect 674484 484740 674485 484804
rect 674419 484739 674485 484740
rect 675894 483581 675954 485730
rect 675891 483580 675957 483581
rect 675891 483516 675892 483580
rect 675956 483516 675957 483580
rect 675891 483515 675957 483516
rect 676262 483030 676322 487870
rect 676998 483030 677058 487870
rect 676262 482970 676874 483030
rect 676998 482970 677242 483030
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 675339 447812 675405 447813
rect 675339 447748 675340 447812
rect 675404 447748 675405 447812
rect 675339 447747 675405 447748
rect 41827 426460 41893 426461
rect 41827 426396 41828 426460
rect 41892 426396 41893 426460
rect 41827 426395 41893 426396
rect 41830 426050 41890 426395
rect 40542 425990 41890 426050
rect 40542 400077 40602 425990
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41827 422788 41893 422789
rect 41827 422724 41828 422788
rect 41892 422724 41893 422788
rect 41827 422723 41893 422724
rect 41830 422310 41890 422723
rect 40726 422250 41890 422310
rect 40726 409461 40786 422250
rect 41827 421972 41893 421973
rect 41827 421970 41828 421972
rect 40910 421910 41828 421970
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40910 405653 40970 421910
rect 41827 421908 41828 421910
rect 41892 421908 41893 421972
rect 41827 421907 41893 421908
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40907 405652 40973 405653
rect 40907 405588 40908 405652
rect 40972 405588 40973 405652
rect 40907 405587 40973 405588
rect 40539 400076 40605 400077
rect 40539 400012 40540 400076
rect 40604 400012 40605 400076
rect 40539 400011 40605 400012
rect 41462 398853 41522 418779
rect 41643 413404 41709 413405
rect 41643 413340 41644 413404
rect 41708 413340 41709 413404
rect 41643 413339 41709 413340
rect 41646 402990 41706 413339
rect 42014 408510 42074 424763
rect 42195 424284 42261 424285
rect 42195 424220 42196 424284
rect 42260 424220 42261 424284
rect 42195 424219 42261 424220
rect 42198 413405 42258 424219
rect 42195 413404 42261 413405
rect 42195 413340 42196 413404
rect 42260 413340 42261 413404
rect 42195 413339 42261 413340
rect 675342 410549 675402 447747
rect 675339 410548 675405 410549
rect 675339 410484 675340 410548
rect 675404 410484 675405 410548
rect 675339 410483 675405 410484
rect 41830 408450 42074 408510
rect 41830 406333 41890 408450
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401845 41890 402930
rect 41827 401844 41893 401845
rect 41827 401780 41828 401844
rect 41892 401780 41893 401844
rect 41827 401779 41893 401780
rect 676814 400485 676874 482970
rect 677182 401301 677242 482970
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 392868 675957 392869
rect 675891 392804 675892 392868
rect 675956 392804 675957 392868
rect 675891 392803 675957 392804
rect 675707 388516 675773 388517
rect 675707 388452 675708 388516
rect 675772 388452 675773 388516
rect 675707 388451 675773 388452
rect 40539 380628 40605 380629
rect 40539 380564 40540 380628
rect 40604 380564 40605 380628
rect 40539 380563 40605 380564
rect 40542 356149 40602 380563
rect 41459 379812 41525 379813
rect 41459 379748 41460 379812
rect 41524 379748 41525 379812
rect 41459 379747 41525 379748
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363765 40786 378115
rect 41275 374644 41341 374645
rect 41275 374580 41276 374644
rect 41340 374580 41341 374644
rect 41275 374579 41341 374580
rect 41278 368525 41338 374579
rect 41275 368524 41341 368525
rect 41275 368460 41276 368524
rect 41340 368460 41341 368524
rect 41275 368459 41341 368460
rect 40723 363764 40789 363765
rect 40723 363700 40724 363764
rect 40788 363700 40789 363764
rect 40723 363699 40789 363700
rect 41462 358733 41522 379747
rect 675710 378725 675770 388451
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 675894 373013 675954 392803
rect 676078 373693 676138 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676443 396404 676509 396405
rect 676443 396340 676444 396404
rect 676508 396340 676509 396404
rect 676443 396339 676509 396340
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676262 377501 676322 395115
rect 676446 382261 676506 396339
rect 676630 385389 676690 396747
rect 676627 385388 676693 385389
rect 676627 385324 676628 385388
rect 676692 385324 676693 385388
rect 676627 385323 676693 385324
rect 676443 382260 676509 382261
rect 676443 382196 676444 382260
rect 676508 382196 676509 382260
rect 676443 382195 676509 382196
rect 676259 377500 676325 377501
rect 676259 377436 676260 377500
rect 676324 377436 676325 377500
rect 676259 377435 676325 377436
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675891 373012 675957 373013
rect 675891 372948 675892 373012
rect 675956 372948 675957 373012
rect 675891 372947 675957 372948
rect 41643 372740 41709 372741
rect 41643 372676 41644 372740
rect 41708 372676 41709 372740
rect 41643 372675 41709 372676
rect 41646 359549 41706 372675
rect 41827 371924 41893 371925
rect 41827 371860 41828 371924
rect 41892 371860 41893 371924
rect 41827 371859 41893 371860
rect 41830 360093 41890 371859
rect 41827 360092 41893 360093
rect 41827 360028 41828 360092
rect 41892 360028 41893 360092
rect 41827 360027 41893 360028
rect 41643 359548 41709 359549
rect 41643 359484 41644 359548
rect 41708 359484 41709 359548
rect 41643 359483 41709 359484
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 40539 356148 40605 356149
rect 40539 356084 40540 356148
rect 40604 356084 40605 356148
rect 40539 356083 40605 356084
rect 675523 353428 675589 353429
rect 675523 353364 675524 353428
rect 675588 353364 675589 353428
rect 675523 353363 675589 353364
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 341596 44285 341597
rect 44219 341532 44220 341596
rect 44284 341532 44285 341596
rect 44219 341531 44285 341532
rect 42747 340508 42813 340509
rect 42747 340444 42748 340508
rect 42812 340444 42813 340508
rect 42747 340443 42813 340444
rect 41643 338196 41709 338197
rect 41643 338132 41644 338196
rect 41708 338132 41709 338196
rect 41643 338131 41709 338132
rect 40723 336972 40789 336973
rect 40723 336908 40724 336972
rect 40788 336908 40789 336972
rect 40723 336907 40789 336908
rect 40539 335340 40605 335341
rect 40539 335276 40540 335340
rect 40604 335276 40605 335340
rect 40539 335275 40605 335276
rect 40542 317389 40602 335275
rect 40726 319021 40786 336907
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40910 325413 40970 333643
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 41646 319970 41706 338131
rect 42011 336564 42077 336565
rect 42011 336500 42012 336564
rect 42076 336500 42077 336564
rect 42011 336499 42077 336500
rect 41827 335748 41893 335749
rect 41827 335684 41828 335748
rect 41892 335684 41893 335748
rect 41827 335683 41893 335684
rect 41830 324869 41890 335683
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41827 319972 41893 319973
rect 41827 319970 41828 319972
rect 41646 319910 41828 319970
rect 41827 319908 41828 319910
rect 41892 319908 41893 319972
rect 41827 319907 41893 319908
rect 40723 319020 40789 319021
rect 40723 318956 40724 319020
rect 40788 318956 40789 319020
rect 40723 318955 40789 318956
rect 40539 317388 40605 317389
rect 40539 317324 40540 317388
rect 40604 317324 40605 317388
rect 40539 317323 40605 317324
rect 42014 313717 42074 336499
rect 42011 313716 42077 313717
rect 42011 313652 42012 313716
rect 42076 313652 42077 313716
rect 42011 313651 42077 313652
rect 42750 297669 42810 340443
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 42934 312765 42994 337587
rect 43115 337244 43181 337245
rect 43115 337180 43116 337244
rect 43180 337180 43181 337244
rect 43115 337179 43181 337180
rect 43118 316029 43178 337179
rect 43115 316028 43181 316029
rect 43115 315964 43116 316028
rect 43180 315964 43181 316028
rect 43115 315963 43181 315964
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 44222 298485 44282 341531
rect 44406 300117 44466 342891
rect 675526 340781 675586 353363
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 349210 675770 352955
rect 675937 352204 676003 352205
rect 675937 352140 675938 352204
rect 676002 352202 676003 352204
rect 676002 352142 676322 352202
rect 676002 352140 676003 352142
rect 675937 352139 676003 352140
rect 675891 351932 675957 351933
rect 675891 351868 675892 351932
rect 675956 351930 675957 351932
rect 675956 351870 676138 351930
rect 675956 351868 675957 351870
rect 675891 351867 675957 351868
rect 675710 349150 675954 349210
rect 675523 340780 675589 340781
rect 675523 340716 675524 340780
rect 675588 340716 675589 340780
rect 675523 340715 675589 340716
rect 44587 340236 44653 340237
rect 44587 340172 44588 340236
rect 44652 340172 44653 340236
rect 44587 340171 44653 340172
rect 44403 300116 44469 300117
rect 44403 300052 44404 300116
rect 44468 300052 44469 300116
rect 44403 300051 44469 300052
rect 44590 299301 44650 340171
rect 675894 337789 675954 349150
rect 675891 337788 675957 337789
rect 675891 337724 675892 337788
rect 675956 337724 675957 337788
rect 675891 337723 675957 337724
rect 676078 328405 676138 351870
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 676262 325549 676322 352142
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676446 340237 676506 346563
rect 676811 346220 676877 346221
rect 676811 346156 676812 346220
rect 676876 346156 676877 346220
rect 676811 346155 676877 346156
rect 676443 340236 676509 340237
rect 676443 340172 676444 340236
rect 676508 340172 676509 340236
rect 676443 340171 676509 340172
rect 676259 325548 676325 325549
rect 676259 325484 676260 325548
rect 676324 325484 676325 325548
rect 676259 325483 676325 325484
rect 676814 325277 676874 346155
rect 676811 325276 676877 325277
rect 676811 325212 676812 325276
rect 676876 325212 676877 325276
rect 676811 325211 676877 325212
rect 675707 309092 675773 309093
rect 675707 309028 675708 309092
rect 675772 309090 675773 309092
rect 675772 309030 675954 309090
rect 675772 309028 675773 309030
rect 675707 309027 675773 309028
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 302250 675770 308755
rect 675894 307770 675954 309030
rect 675894 307710 676506 307770
rect 675891 307188 675957 307189
rect 675891 307124 675892 307188
rect 675956 307124 675957 307188
rect 675891 307123 675957 307124
rect 675894 303650 675954 307123
rect 675894 303590 676138 303650
rect 675710 302190 675954 302250
rect 675707 299436 675773 299437
rect 675707 299372 675708 299436
rect 675772 299372 675773 299436
rect 675707 299371 675773 299372
rect 44587 299300 44653 299301
rect 44587 299236 44588 299300
rect 44652 299236 44653 299300
rect 44587 299235 44653 299236
rect 44219 298484 44285 298485
rect 44219 298420 44220 298484
rect 44284 298420 44285 298484
rect 44219 298419 44285 298420
rect 42747 297668 42813 297669
rect 42747 297604 42748 297668
rect 42812 297604 42813 297668
rect 42747 297603 42813 297604
rect 675523 297396 675589 297397
rect 675523 297332 675524 297396
rect 675588 297332 675589 297396
rect 675523 297331 675589 297332
rect 42011 296852 42077 296853
rect 42011 296788 42012 296852
rect 42076 296788 42077 296852
rect 42011 296787 42077 296788
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 41827 291548 41893 291549
rect 41827 291484 41828 291548
rect 41892 291484 41893 291548
rect 41827 291483 41893 291484
rect 41830 289830 41890 291483
rect 40910 289770 41890 289830
rect 40723 289236 40789 289237
rect 40723 289172 40724 289236
rect 40788 289172 40789 289236
rect 40723 289171 40789 289172
rect 40726 277133 40786 289171
rect 40910 278493 40970 289770
rect 42014 288010 42074 296787
rect 675526 292229 675586 297331
rect 675523 292228 675589 292229
rect 675523 292164 675524 292228
rect 675588 292164 675589 292228
rect 675523 292163 675589 292164
rect 41462 287950 42074 288010
rect 40907 278492 40973 278493
rect 40907 278428 40908 278492
rect 40972 278428 40973 278492
rect 40907 278427 40973 278428
rect 40723 277132 40789 277133
rect 40723 277068 40724 277132
rect 40788 277068 40789 277132
rect 40723 277067 40789 277068
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 287950
rect 41643 284884 41709 284885
rect 41643 284820 41644 284884
rect 41708 284820 41709 284884
rect 41643 284819 41709 284820
rect 41646 273730 41706 284819
rect 42011 284340 42077 284341
rect 42011 284276 42012 284340
rect 42076 284276 42077 284340
rect 42011 284275 42077 284276
rect 41646 273670 41890 273730
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 270061 41890 273670
rect 42014 272373 42074 284275
rect 675710 282845 675770 299371
rect 675894 283661 675954 302190
rect 675891 283660 675957 283661
rect 675891 283596 675892 283660
rect 675956 283596 675957 283660
rect 675891 283595 675957 283596
rect 675707 282844 675773 282845
rect 675707 282780 675708 282844
rect 675772 282780 675773 282844
rect 675707 282779 675773 282780
rect 676078 281213 676138 303590
rect 676446 302970 676506 307710
rect 676627 304570 676693 304571
rect 676627 304506 676628 304570
rect 676692 304506 676693 304570
rect 676627 304505 676693 304506
rect 676262 302910 676506 302970
rect 676262 294541 676322 302910
rect 676443 300660 676509 300661
rect 676443 300596 676444 300660
rect 676508 300596 676509 300660
rect 676443 300595 676509 300596
rect 676259 294540 676325 294541
rect 676259 294476 676260 294540
rect 676324 294476 676325 294540
rect 676259 294475 676325 294476
rect 676446 291549 676506 300595
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676630 290869 676690 304505
rect 676627 290868 676693 290869
rect 676627 290804 676628 290868
rect 676692 290804 676693 290868
rect 676627 290803 676693 290804
rect 676075 281212 676141 281213
rect 676075 281148 676076 281212
rect 676140 281148 676141 281212
rect 676075 281147 676141 281148
rect 42011 272372 42077 272373
rect 42011 272308 42012 272372
rect 42076 272308 42077 272372
rect 42011 272307 42077 272308
rect 41827 270060 41893 270061
rect 41827 269996 41828 270060
rect 41892 269996 41893 270060
rect 41827 269995 41893 269996
rect 674971 264212 675037 264213
rect 674971 264148 674972 264212
rect 675036 264148 675037 264212
rect 674971 264147 675037 264148
rect 40539 250204 40605 250205
rect 40539 250140 40540 250204
rect 40604 250140 40605 250204
rect 40539 250139 40605 250140
rect 40542 230485 40602 250139
rect 674974 249797 675034 264147
rect 676075 263668 676141 263669
rect 676075 263604 676076 263668
rect 676140 263604 676141 263668
rect 676075 263603 676141 263604
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 674971 249796 675037 249797
rect 674971 249732 674972 249796
rect 675036 249732 675037 249796
rect 674971 249731 675037 249732
rect 40726 236605 40786 249731
rect 676078 249661 676138 263603
rect 676811 261628 676877 261629
rect 676811 261564 676812 261628
rect 676876 261564 676877 261628
rect 676811 261563 676877 261564
rect 676814 250205 676874 261563
rect 676995 259996 677061 259997
rect 676995 259932 676996 259996
rect 677060 259932 677061 259996
rect 676995 259931 677061 259932
rect 676811 250204 676877 250205
rect 676811 250140 676812 250204
rect 676876 250140 676877 250204
rect 676811 250139 676877 250140
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 676998 242317 677058 259931
rect 676995 242316 677061 242317
rect 676995 242252 676996 242316
rect 677060 242252 677061 242316
rect 676995 242251 677061 242252
rect 676811 242044 676877 242045
rect 676811 241980 676812 242044
rect 676876 241980 676877 242044
rect 676811 241979 676877 241980
rect 674971 241772 675037 241773
rect 674971 241708 674972 241772
rect 675036 241708 675037 241772
rect 674971 241707 675037 241708
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 40723 236604 40789 236605
rect 40723 236540 40724 236604
rect 40788 236540 40789 236604
rect 40723 236539 40789 236540
rect 40539 230484 40605 230485
rect 40539 230420 40540 230484
rect 40604 230420 40605 230484
rect 40539 230419 40605 230420
rect 42014 228989 42074 237355
rect 674974 230213 675034 241707
rect 674971 230212 675037 230213
rect 674971 230148 674972 230212
rect 675036 230148 675037 230212
rect 674971 230147 675037 230148
rect 674051 229804 674117 229805
rect 674051 229740 674052 229804
rect 674116 229740 674117 229804
rect 674051 229739 674117 229740
rect 42011 228988 42077 228989
rect 42011 228924 42012 228988
rect 42076 228924 42077 228988
rect 42011 228923 42077 228924
rect 672947 227084 673013 227085
rect 672947 227020 672948 227084
rect 673012 227020 673013 227084
rect 672947 227019 673013 227020
rect 561627 222188 561693 222189
rect 561627 222124 561628 222188
rect 561692 222124 561693 222188
rect 561627 222123 561693 222124
rect 561630 219197 561690 222123
rect 561627 219196 561693 219197
rect 561627 219132 561628 219196
rect 561692 219132 561693 219196
rect 561627 219131 561693 219132
rect 509187 217836 509253 217837
rect 509187 217772 509188 217836
rect 509252 217772 509253 217836
rect 522619 217836 522685 217837
rect 509187 217771 509253 217772
rect 510107 217772 510108 217822
rect 510172 217772 510173 217822
rect 510107 217771 510173 217772
rect 522619 217772 522620 217836
rect 522684 217772 522685 217836
rect 522619 217771 522685 217772
rect 509190 215933 509250 217771
rect 509187 215932 509253 215933
rect 509187 215868 509188 215932
rect 509252 215868 509253 215932
rect 509187 215867 509253 215868
rect 522622 215389 522682 217771
rect 561630 216205 561690 219131
rect 574323 217772 574324 217822
rect 574388 217772 574389 217822
rect 574323 217771 574389 217772
rect 574326 216749 574386 217142
rect 574323 216748 574389 216749
rect 574323 216684 574324 216748
rect 574388 216684 574389 216748
rect 574323 216683 574389 216684
rect 561627 216204 561693 216205
rect 561627 216140 561628 216204
rect 561692 216140 561693 216204
rect 561627 216139 561693 216140
rect 522619 215388 522685 215389
rect 522619 215324 522620 215388
rect 522684 215324 522685 215388
rect 522619 215323 522685 215324
rect 670187 213892 670253 213893
rect 670187 213828 670188 213892
rect 670252 213828 670253 213892
rect 670187 213827 670253 213828
rect 670190 213077 670250 213827
rect 670187 213076 670253 213077
rect 670187 213012 670188 213076
rect 670252 213012 670253 213076
rect 670187 213011 670253 213012
rect 670739 210492 670805 210493
rect 670739 210428 670740 210492
rect 670804 210428 670805 210492
rect 670739 210427 670805 210428
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 41643 208180 41709 208181
rect 41643 208116 41644 208180
rect 41708 208116 41709 208180
rect 41643 208115 41709 208116
rect 40539 207364 40605 207365
rect 40539 207300 40540 207364
rect 40604 207300 40605 207364
rect 40539 207299 40605 207300
rect 40542 186421 40602 207299
rect 40723 206548 40789 206549
rect 40723 206484 40724 206548
rect 40788 206484 40789 206548
rect 40723 206483 40789 206484
rect 40726 193221 40786 206483
rect 40907 206140 40973 206141
rect 40907 206076 40908 206140
rect 40972 206076 40973 206140
rect 40907 206075 40973 206076
rect 40910 194989 40970 206075
rect 41459 205732 41525 205733
rect 41459 205668 41460 205732
rect 41524 205668 41525 205732
rect 41459 205667 41525 205668
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 193220 40789 193221
rect 40723 193156 40724 193220
rect 40788 193156 40789 193220
rect 40723 193155 40789 193156
rect 40539 186420 40605 186421
rect 40539 186356 40540 186420
rect 40604 186356 40605 186420
rect 40539 186355 40605 186356
rect 41462 184109 41522 205667
rect 41646 190470 41706 208115
rect 41830 195261 41890 210019
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 41646 190410 41890 190470
rect 41830 186013 41890 190410
rect 41827 186012 41893 186013
rect 41827 185948 41828 186012
rect 41892 185948 41893 186012
rect 41827 185947 41893 185948
rect 41459 184108 41525 184109
rect 41459 184044 41460 184108
rect 41524 184044 41525 184108
rect 41459 184043 41525 184044
rect 669451 169692 669517 169693
rect 669451 169628 669452 169692
rect 669516 169628 669517 169692
rect 669451 169627 669517 169628
rect 669454 157350 669514 169627
rect 669270 157290 669514 157350
rect 669270 140453 669330 157290
rect 669267 140452 669333 140453
rect 669267 140388 669268 140452
rect 669332 140388 669333 140452
rect 669267 140387 669333 140388
rect 670742 125765 670802 210427
rect 672579 208316 672645 208317
rect 672579 208252 672580 208316
rect 672644 208252 672645 208316
rect 672579 208251 672645 208252
rect 672582 202605 672642 208251
rect 672579 202604 672645 202605
rect 672579 202540 672580 202604
rect 672644 202540 672645 202604
rect 672579 202539 672645 202540
rect 672950 133381 673010 227019
rect 673499 223684 673565 223685
rect 673499 223620 673500 223684
rect 673564 223620 673565 223684
rect 673499 223619 673565 223620
rect 672947 133380 673013 133381
rect 672947 133316 672948 133380
rect 673012 133316 673013 133380
rect 672947 133315 673013 133316
rect 673502 132837 673562 223619
rect 673499 132836 673565 132837
rect 673499 132772 673500 132836
rect 673564 132772 673565 132836
rect 673499 132771 673565 132772
rect 670739 125764 670805 125765
rect 670739 125700 670740 125764
rect 670804 125700 670805 125764
rect 670739 125699 670805 125700
rect 674054 115837 674114 229739
rect 675891 220692 675957 220693
rect 675891 220628 675892 220692
rect 675956 220690 675957 220692
rect 676814 220690 676874 241979
rect 675956 220630 676874 220690
rect 675956 220628 675957 220630
rect 675891 220627 675957 220628
rect 675894 218590 676506 218650
rect 675894 218381 675954 218590
rect 675891 218380 675957 218381
rect 675891 218316 675892 218380
rect 675956 218316 675957 218380
rect 675891 218315 675957 218316
rect 675707 217428 675773 217429
rect 675707 217364 675708 217428
rect 675772 217364 675773 217428
rect 675707 217363 675773 217364
rect 675710 198389 675770 217363
rect 675891 215252 675957 215253
rect 675891 215188 675892 215252
rect 675956 215250 675957 215252
rect 675956 215190 676322 215250
rect 675956 215188 675957 215190
rect 675891 215187 675957 215188
rect 675891 214436 675957 214437
rect 675891 214372 675892 214436
rect 675956 214372 675957 214436
rect 675891 214371 675957 214372
rect 675894 211170 675954 214371
rect 675894 211110 676138 211170
rect 675891 210628 675957 210629
rect 675891 210564 675892 210628
rect 675956 210564 675957 210628
rect 675891 210563 675957 210564
rect 675707 198388 675773 198389
rect 675707 198324 675708 198388
rect 675772 198324 675773 198388
rect 675707 198323 675773 198324
rect 675894 192813 675954 210563
rect 676078 210490 676138 211110
rect 676262 210901 676322 215190
rect 676259 210900 676325 210901
rect 676259 210836 676260 210900
rect 676324 210836 676325 210900
rect 676259 210835 676325 210836
rect 676078 210430 676322 210490
rect 676075 206956 676141 206957
rect 676075 206892 676076 206956
rect 676140 206892 676141 206956
rect 676075 206891 676141 206892
rect 676078 204237 676138 206891
rect 676075 204236 676141 204237
rect 676075 204172 676076 204236
rect 676140 204172 676141 204236
rect 676075 204171 676141 204172
rect 676262 200837 676322 210430
rect 676446 205597 676506 218590
rect 676627 210900 676693 210901
rect 676627 210836 676628 210900
rect 676692 210836 676693 210900
rect 676627 210835 676693 210836
rect 676443 205596 676509 205597
rect 676443 205532 676444 205596
rect 676508 205532 676509 205596
rect 676443 205531 676509 205532
rect 676259 200836 676325 200837
rect 676259 200772 676260 200836
rect 676324 200772 676325 200836
rect 676259 200771 676325 200772
rect 676630 196213 676690 210835
rect 676627 196212 676693 196213
rect 676627 196148 676628 196212
rect 676692 196148 676693 196212
rect 676627 196147 676693 196148
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 675523 173636 675589 173637
rect 675523 173572 675524 173636
rect 675588 173572 675589 173636
rect 675523 173571 675589 173572
rect 675339 171188 675405 171189
rect 675339 171124 675340 171188
rect 675404 171124 675405 171188
rect 675339 171123 675405 171124
rect 675342 157045 675402 171123
rect 675526 162213 675586 173571
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 675707 172412 675773 172413
rect 675707 172348 675708 172412
rect 675772 172348 675773 172412
rect 675894 172410 675954 172755
rect 675894 172350 676506 172410
rect 675707 172347 675773 172348
rect 675710 169010 675770 172347
rect 675891 169692 675957 169693
rect 675891 169628 675892 169692
rect 675956 169690 675957 169692
rect 675956 169630 676322 169690
rect 675956 169628 675957 169630
rect 675891 169627 675957 169628
rect 675710 168950 675954 169010
rect 675707 167516 675773 167517
rect 675707 167452 675708 167516
rect 675772 167452 675773 167516
rect 675707 167451 675773 167452
rect 675523 162212 675589 162213
rect 675523 162148 675524 162212
rect 675588 162148 675589 162212
rect 675523 162147 675589 162148
rect 675339 157044 675405 157045
rect 675339 156980 675340 157044
rect 675404 156980 675405 157044
rect 675339 156979 675405 156980
rect 675710 147661 675770 167451
rect 675894 153101 675954 168950
rect 676075 162212 676141 162213
rect 676075 162148 676076 162212
rect 676140 162148 676141 162212
rect 676075 162147 676141 162148
rect 675891 153100 675957 153101
rect 675891 153036 675892 153100
rect 675956 153036 675957 153100
rect 675891 153035 675957 153036
rect 676078 148477 676138 162147
rect 676262 155821 676322 169630
rect 676446 157045 676506 172350
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 157044 676509 157045
rect 676443 156980 676444 157044
rect 676508 156980 676509 157044
rect 676443 156979 676509 156980
rect 676259 155820 676325 155821
rect 676259 155756 676260 155820
rect 676324 155756 676325 155820
rect 676259 155755 676325 155756
rect 676630 151469 676690 166363
rect 676627 151468 676693 151469
rect 676627 151404 676628 151468
rect 676692 151404 676693 151468
rect 676627 151403 676693 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 676443 128620 676509 128621
rect 676443 128556 676444 128620
rect 676508 128556 676509 128620
rect 676443 128555 676509 128556
rect 676259 128212 676325 128213
rect 676259 128148 676260 128212
rect 676324 128148 676325 128212
rect 676259 128147 676325 128148
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675707 122908 675773 122909
rect 675707 122844 675708 122908
rect 675772 122844 675773 122908
rect 675707 122843 675773 122844
rect 674051 115836 674117 115837
rect 674051 115772 674052 115836
rect 674116 115772 674117 115836
rect 674051 115771 674117 115772
rect 675710 111349 675770 122843
rect 675891 116516 675957 116517
rect 675891 116452 675892 116516
rect 675956 116452 675957 116516
rect 675891 116451 675957 116452
rect 675707 111348 675773 111349
rect 675707 111284 675708 111348
rect 675772 111284 675773 111348
rect 675707 111283 675773 111284
rect 675894 104821 675954 116451
rect 676078 108221 676138 126923
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675891 104820 675957 104821
rect 675891 104756 675892 104820
rect 675956 104756 675957 104820
rect 675891 104755 675957 104756
rect 676262 103189 676322 128147
rect 676446 114205 676506 128555
rect 676811 121684 676877 121685
rect 676811 121620 676812 121684
rect 676876 121620 676877 121684
rect 676811 121619 676877 121620
rect 676443 114204 676509 114205
rect 676443 114140 676444 114204
rect 676508 114140 676509 114204
rect 676443 114139 676509 114140
rect 676814 111757 676874 121619
rect 676811 111756 676877 111757
rect 676811 111692 676812 111756
rect 676876 111692 676877 111756
rect 676811 111691 676877 111692
rect 676259 103188 676325 103189
rect 676259 103124 676260 103188
rect 676324 103124 676325 103188
rect 676259 103123 676325 103124
rect 635779 96932 635845 96933
rect 635779 96868 635780 96932
rect 635844 96868 635845 96932
rect 635779 96867 635845 96868
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95980 634005 95981
rect 633939 95916 633940 95980
rect 634004 95916 634005 95980
rect 633939 95915 634005 95916
rect 633942 78573 634002 95915
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 635782 78165 635842 96867
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 635779 78164 635845 78165
rect 635779 78100 635780 78164
rect 635844 78100 635845 78164
rect 635779 78099 635845 78100
rect 637070 77621 637130 84150
rect 637067 77620 637133 77621
rect 637067 77556 637068 77620
rect 637132 77556 637133 77620
rect 637067 77555 637133 77556
rect 461715 55044 461781 55045
rect 461715 54980 461716 55044
rect 461780 54980 461781 55044
rect 461715 54979 461781 54980
rect 461718 53957 461778 54979
rect 462635 54772 462701 54773
rect 462635 54708 462636 54772
rect 462700 54708 462701 54772
rect 462635 54707 462701 54708
rect 462638 53957 462698 54707
rect 461715 53956 461781 53957
rect 461715 53892 461716 53956
rect 461780 53892 461781 53956
rect 461715 53891 461781 53892
rect 462635 53956 462701 53957
rect 462635 53892 462636 53956
rect 462700 53892 462701 53956
rect 462635 53891 462701 53892
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 194366 42125 194426 50219
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 458219 44436 458285 44437
rect 458219 44372 458220 44436
rect 458284 44372 458285 44436
rect 458219 44371 458285 44372
rect 461347 44436 461413 44437
rect 461347 44372 461348 44436
rect 461412 44372 461413 44436
rect 461347 44371 461413 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 405595 41852 405661 41853
rect 405595 41788 405596 41852
rect 405660 41788 405661 41852
rect 405595 41787 405661 41788
rect 421974 41850 422034 42059
rect 421974 41790 422162 41850
rect 405598 40578 405658 41787
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 458222 40578 458282 44371
rect 461350 41938 461410 44371
rect 462270 41938 462330 44371
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 510022 217836 510258 218058
rect 510022 217822 510108 217836
rect 510108 217822 510172 217836
rect 510172 217822 510258 217836
rect 493646 217292 493882 217378
rect 493646 217228 493732 217292
rect 493732 217228 493796 217292
rect 493796 217228 493882 217292
rect 493646 217142 493882 217228
rect 574238 217836 574474 218058
rect 574238 217822 574324 217836
rect 574324 217822 574388 217836
rect 574388 217822 574474 217836
rect 574238 217142 574474 217378
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
rect 405510 40342 405746 40578
rect 458134 40342 458370 40578
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 509980 218058 574516 218100
rect 509980 217822 510022 218058
rect 510258 217822 574238 218058
rect 574474 217822 574516 218058
rect 509980 217780 574516 217822
rect 493604 217378 574516 217420
rect 493604 217142 493646 217378
rect 493882 217142 574238 217378
rect 574474 217142 574516 217378
rect 493604 217100 574516 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 405468 40578 458412 40620
rect 405468 40342 405510 40578
rect 405746 40342 458134 40578
rect 458370 40342 458412 40578
rect 405468 40300 458412 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 0
transform 1 0 255300 0 1 6032
box 0 0 1 1
use caravan_motto  caravan_motto
timestamp 0
transform 1 0 -54560 0 1 -52
box 0 0 1 1
use copyright_block_a  copyright_block_a
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206074 0 1 2336
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1666432150
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1666432150
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1666432150
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666432150
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1666432150
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666432150
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1666432150
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1666432150
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1666432150
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1666432150
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666432150
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666432150
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666432150
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666432150
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666432150
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666432150
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1666432150
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666432150
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666432150
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666432150
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1666432150
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1666432150
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666432150
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666432150
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666432150
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666432150
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666432150
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666432150
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666432150
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666432150
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666432150
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666432150
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666432150
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666432150
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666432150
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666432150
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666432150
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666432150
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666432150
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666432150
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666432150
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666432150
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666432150
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666432150
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666432150
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666432150
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666432150
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666432150
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666432150
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666432150
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666432150
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666432150
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666432150
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666432150
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666432150
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666432150
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666432150
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666432150
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666432150
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666432150
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666432150
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666432150
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666432150
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666432150
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666432150
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666432150
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666432150
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use caravan_power_routing  caravan_power_routing
timestamp 1666432150
transform 1 0 0 0 1 0
box 6022 30806 711814 997678
use caravan_signal_routing  caravan_signal_routing
timestamp 1666432150
transform 1 0 0 0 1 0
box 39764 415548 677806 997846
use user_analog_project_wrapper  mprj
timestamp 1666432150
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use chip_io_alt  padframe
timestamp 1666432150
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering_alt  sigbuf
timestamp 1666432150
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 953022 710789 965190 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030789 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030789 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030789 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386210 1018624 398378 1030789 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284410 1018624 296578 1030789 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030789 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030789 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030789 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030789 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18976 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
