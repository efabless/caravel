// This is the unpowered netlist.
module housekeeping_alt (debug_in,
    debug_mode,
    debug_oeb,
    debug_out,
    pad_flash_clk,
    pad_flash_clk_oeb,
    pad_flash_csb,
    pad_flash_csb_oeb,
    pad_flash_io0_di,
    pad_flash_io0_do,
    pad_flash_io0_ieb,
    pad_flash_io0_oeb,
    pad_flash_io1_di,
    pad_flash_io1_do,
    pad_flash_io1_ieb,
    pad_flash_io1_oeb,
    pll_bypass,
    pll_dco_ena,
    pll_ena,
    porb,
    qspi_enabled,
    reset,
    ser_rx,
    ser_tx,
    serial_clock,
    serial_data_1,
    serial_data_2,
    serial_load,
    serial_resetn,
    spi_csb,
    spi_enabled,
    spi_sck,
    spi_sdi,
    spi_sdo,
    spi_sdoenb,
    spimemio_flash_clk,
    spimemio_flash_csb,
    spimemio_flash_io0_di,
    spimemio_flash_io0_do,
    spimemio_flash_io0_oeb,
    spimemio_flash_io1_di,
    spimemio_flash_io1_do,
    spimemio_flash_io1_oeb,
    spimemio_flash_io2_di,
    spimemio_flash_io2_do,
    spimemio_flash_io2_oeb,
    spimemio_flash_io3_di,
    spimemio_flash_io3_do,
    spimemio_flash_io3_oeb,
    trap,
    uart_enabled,
    user_clock,
    usr1_vcc_pwrgood,
    usr1_vdd_pwrgood,
    usr2_vcc_pwrgood,
    usr2_vdd_pwrgood,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rstn_i,
    wb_stb_i,
    wb_we_i,
    irq,
    mask_rev_in,
    mgmt_gpio_in,
    mgmt_gpio_oeb,
    mgmt_gpio_out,
    pll90_sel,
    pll_div,
    pll_sel,
    pll_trim,
    pwr_ctrl_out,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o,
    wb_sel_i);
 output debug_in;
 input debug_mode;
 input debug_oeb;
 input debug_out;
 output pad_flash_clk;
 output pad_flash_clk_oeb;
 output pad_flash_csb;
 output pad_flash_csb_oeb;
 input pad_flash_io0_di;
 output pad_flash_io0_do;
 output pad_flash_io0_ieb;
 output pad_flash_io0_oeb;
 input pad_flash_io1_di;
 output pad_flash_io1_do;
 output pad_flash_io1_ieb;
 output pad_flash_io1_oeb;
 output pll_bypass;
 output pll_dco_ena;
 output pll_ena;
 input porb;
 input qspi_enabled;
 output reset;
 output ser_rx;
 input ser_tx;
 output serial_clock;
 output serial_data_1;
 output serial_data_2;
 output serial_load;
 output serial_resetn;
 input spi_csb;
 input spi_enabled;
 input spi_sck;
 output spi_sdi;
 input spi_sdo;
 input spi_sdoenb;
 input spimemio_flash_clk;
 input spimemio_flash_csb;
 output spimemio_flash_io0_di;
 input spimemio_flash_io0_do;
 input spimemio_flash_io0_oeb;
 output spimemio_flash_io1_di;
 input spimemio_flash_io1_do;
 input spimemio_flash_io1_oeb;
 output spimemio_flash_io2_di;
 input spimemio_flash_io2_do;
 input spimemio_flash_io2_oeb;
 output spimemio_flash_io3_di;
 input spimemio_flash_io3_do;
 input spimemio_flash_io3_oeb;
 input trap;
 input uart_enabled;
 input user_clock;
 input usr1_vcc_pwrgood;
 input usr1_vdd_pwrgood;
 input usr2_vcc_pwrgood;
 input usr2_vdd_pwrgood;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rstn_i;
 input wb_stb_i;
 input wb_we_i;
 output [2:0] irq;
 input [31:0] mask_rev_in;
 input [37:0] mgmt_gpio_in;
 output [37:0] mgmt_gpio_oeb;
 output [37:0] mgmt_gpio_out;
 output [2:0] pll90_sel;
 output [4:0] pll_div;
 output [2:0] pll_sel;
 output [25:0] pll_trim;
 output [3:0] pwr_ctrl_out;
 input [31:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 input [3:0] wb_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire \clk1_output_dest[0] ;
 wire \clk1_output_dest[1] ;
 wire \clk2_output_dest[0] ;
 wire \clk2_output_dest[1] ;
 wire clknet_0__1111_;
 wire clknet_0_csclk;
 wire clknet_0_user_clock;
 wire clknet_0_wb_clk_i;
 wire clknet_0_wbbd_sck;
 wire clknet_1_0__leaf__1111_;
 wire clknet_1_0__leaf_user_clock;
 wire clknet_1_0__leaf_wbbd_sck;
 wire clknet_1_1__leaf__1111_;
 wire clknet_1_1__leaf_user_clock;
 wire clknet_1_1__leaf_wbbd_sck;
 wire clknet_3_0_0_csclk;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_csclk;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_csclk;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_csclk;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_csclk;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_csclk;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_csclk;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_csclk;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_csclk;
 wire clknet_leaf_10_csclk;
 wire clknet_leaf_11_csclk;
 wire clknet_leaf_12_csclk;
 wire clknet_leaf_13_csclk;
 wire clknet_leaf_14_csclk;
 wire clknet_leaf_15_csclk;
 wire clknet_leaf_16_csclk;
 wire clknet_leaf_17_csclk;
 wire clknet_leaf_18_csclk;
 wire clknet_leaf_19_csclk;
 wire clknet_leaf_1_csclk;
 wire clknet_leaf_20_csclk;
 wire clknet_leaf_21_csclk;
 wire clknet_leaf_22_csclk;
 wire clknet_leaf_23_csclk;
 wire clknet_leaf_24_csclk;
 wire clknet_leaf_25_csclk;
 wire clknet_leaf_26_csclk;
 wire clknet_leaf_27_csclk;
 wire clknet_leaf_28_csclk;
 wire clknet_leaf_29_csclk;
 wire clknet_leaf_2_csclk;
 wire clknet_leaf_30_csclk;
 wire clknet_leaf_31_csclk;
 wire clknet_leaf_32_csclk;
 wire clknet_leaf_33_csclk;
 wire clknet_leaf_35_csclk;
 wire clknet_leaf_36_csclk;
 wire clknet_leaf_37_csclk;
 wire clknet_leaf_38_csclk;
 wire clknet_leaf_39_csclk;
 wire clknet_leaf_3_csclk;
 wire clknet_leaf_40_csclk;
 wire clknet_leaf_41_csclk;
 wire clknet_leaf_42_csclk;
 wire clknet_leaf_43_csclk;
 wire clknet_leaf_44_csclk;
 wire clknet_leaf_45_csclk;
 wire clknet_leaf_46_csclk;
 wire clknet_leaf_47_csclk;
 wire clknet_leaf_48_csclk;
 wire clknet_leaf_49_csclk;
 wire clknet_leaf_4_csclk;
 wire clknet_leaf_50_csclk;
 wire clknet_leaf_51_csclk;
 wire clknet_leaf_52_csclk;
 wire clknet_leaf_53_csclk;
 wire clknet_leaf_54_csclk;
 wire clknet_leaf_55_csclk;
 wire clknet_leaf_56_csclk;
 wire clknet_leaf_57_csclk;
 wire clknet_leaf_58_csclk;
 wire clknet_leaf_59_csclk;
 wire clknet_leaf_5_csclk;
 wire clknet_leaf_60_csclk;
 wire clknet_leaf_61_csclk;
 wire clknet_leaf_62_csclk;
 wire clknet_leaf_63_csclk;
 wire clknet_leaf_64_csclk;
 wire clknet_leaf_66_csclk;
 wire clknet_leaf_67_csclk;
 wire clknet_leaf_68_csclk;
 wire clknet_leaf_69_csclk;
 wire clknet_leaf_6_csclk;
 wire clknet_leaf_70_csclk;
 wire clknet_leaf_71_csclk;
 wire clknet_leaf_72_csclk;
 wire clknet_leaf_73_csclk;
 wire clknet_leaf_74_csclk;
 wire clknet_leaf_75_csclk;
 wire clknet_leaf_76_csclk;
 wire clknet_leaf_77_csclk;
 wire clknet_leaf_7_csclk;
 wire clknet_leaf_8_csclk;
 wire clknet_leaf_9_csclk;
 wire csclk;
 wire \gpio_configure[0][0] ;
 wire \gpio_configure[0][10] ;
 wire \gpio_configure[0][11] ;
 wire \gpio_configure[0][12] ;
 wire \gpio_configure[0][1] ;
 wire \gpio_configure[0][2] ;
 wire \gpio_configure[0][3] ;
 wire \gpio_configure[0][4] ;
 wire \gpio_configure[0][5] ;
 wire \gpio_configure[0][6] ;
 wire \gpio_configure[0][7] ;
 wire \gpio_configure[0][8] ;
 wire \gpio_configure[0][9] ;
 wire \gpio_configure[10][0] ;
 wire \gpio_configure[10][10] ;
 wire \gpio_configure[10][11] ;
 wire \gpio_configure[10][12] ;
 wire \gpio_configure[10][1] ;
 wire \gpio_configure[10][2] ;
 wire \gpio_configure[10][3] ;
 wire \gpio_configure[10][4] ;
 wire \gpio_configure[10][5] ;
 wire \gpio_configure[10][6] ;
 wire \gpio_configure[10][7] ;
 wire \gpio_configure[10][8] ;
 wire \gpio_configure[10][9] ;
 wire \gpio_configure[11][0] ;
 wire \gpio_configure[11][10] ;
 wire \gpio_configure[11][11] ;
 wire \gpio_configure[11][12] ;
 wire \gpio_configure[11][1] ;
 wire \gpio_configure[11][2] ;
 wire \gpio_configure[11][3] ;
 wire \gpio_configure[11][4] ;
 wire \gpio_configure[11][5] ;
 wire \gpio_configure[11][6] ;
 wire \gpio_configure[11][7] ;
 wire \gpio_configure[11][8] ;
 wire \gpio_configure[11][9] ;
 wire \gpio_configure[12][0] ;
 wire \gpio_configure[12][10] ;
 wire \gpio_configure[12][11] ;
 wire \gpio_configure[12][12] ;
 wire \gpio_configure[12][1] ;
 wire \gpio_configure[12][2] ;
 wire \gpio_configure[12][3] ;
 wire \gpio_configure[12][4] ;
 wire \gpio_configure[12][5] ;
 wire \gpio_configure[12][6] ;
 wire \gpio_configure[12][7] ;
 wire \gpio_configure[12][8] ;
 wire \gpio_configure[12][9] ;
 wire \gpio_configure[13][0] ;
 wire \gpio_configure[13][10] ;
 wire \gpio_configure[13][11] ;
 wire \gpio_configure[13][12] ;
 wire \gpio_configure[13][1] ;
 wire \gpio_configure[13][2] ;
 wire \gpio_configure[13][3] ;
 wire \gpio_configure[13][4] ;
 wire \gpio_configure[13][5] ;
 wire \gpio_configure[13][6] ;
 wire \gpio_configure[13][7] ;
 wire \gpio_configure[13][8] ;
 wire \gpio_configure[13][9] ;
 wire \gpio_configure[14][0] ;
 wire \gpio_configure[14][10] ;
 wire \gpio_configure[14][11] ;
 wire \gpio_configure[14][12] ;
 wire \gpio_configure[14][1] ;
 wire \gpio_configure[14][2] ;
 wire \gpio_configure[14][3] ;
 wire \gpio_configure[14][4] ;
 wire \gpio_configure[14][5] ;
 wire \gpio_configure[14][6] ;
 wire \gpio_configure[14][7] ;
 wire \gpio_configure[14][8] ;
 wire \gpio_configure[14][9] ;
 wire \gpio_configure[15][0] ;
 wire \gpio_configure[15][10] ;
 wire \gpio_configure[15][11] ;
 wire \gpio_configure[15][12] ;
 wire \gpio_configure[15][1] ;
 wire \gpio_configure[15][2] ;
 wire \gpio_configure[15][3] ;
 wire \gpio_configure[15][4] ;
 wire \gpio_configure[15][5] ;
 wire \gpio_configure[15][6] ;
 wire \gpio_configure[15][7] ;
 wire \gpio_configure[15][8] ;
 wire \gpio_configure[15][9] ;
 wire \gpio_configure[16][0] ;
 wire \gpio_configure[16][10] ;
 wire \gpio_configure[16][11] ;
 wire \gpio_configure[16][12] ;
 wire \gpio_configure[16][1] ;
 wire \gpio_configure[16][2] ;
 wire \gpio_configure[16][3] ;
 wire \gpio_configure[16][4] ;
 wire \gpio_configure[16][5] ;
 wire \gpio_configure[16][6] ;
 wire \gpio_configure[16][7] ;
 wire \gpio_configure[16][8] ;
 wire \gpio_configure[16][9] ;
 wire \gpio_configure[17][0] ;
 wire \gpio_configure[17][10] ;
 wire \gpio_configure[17][11] ;
 wire \gpio_configure[17][12] ;
 wire \gpio_configure[17][1] ;
 wire \gpio_configure[17][2] ;
 wire \gpio_configure[17][3] ;
 wire \gpio_configure[17][4] ;
 wire \gpio_configure[17][5] ;
 wire \gpio_configure[17][6] ;
 wire \gpio_configure[17][7] ;
 wire \gpio_configure[17][8] ;
 wire \gpio_configure[17][9] ;
 wire \gpio_configure[18][0] ;
 wire \gpio_configure[18][10] ;
 wire \gpio_configure[18][11] ;
 wire \gpio_configure[18][12] ;
 wire \gpio_configure[18][1] ;
 wire \gpio_configure[18][2] ;
 wire \gpio_configure[18][3] ;
 wire \gpio_configure[18][4] ;
 wire \gpio_configure[18][5] ;
 wire \gpio_configure[18][6] ;
 wire \gpio_configure[18][7] ;
 wire \gpio_configure[18][8] ;
 wire \gpio_configure[18][9] ;
 wire \gpio_configure[19][0] ;
 wire \gpio_configure[19][10] ;
 wire \gpio_configure[19][11] ;
 wire \gpio_configure[19][12] ;
 wire \gpio_configure[19][1] ;
 wire \gpio_configure[19][2] ;
 wire \gpio_configure[19][3] ;
 wire \gpio_configure[19][4] ;
 wire \gpio_configure[19][5] ;
 wire \gpio_configure[19][6] ;
 wire \gpio_configure[19][7] ;
 wire \gpio_configure[19][8] ;
 wire \gpio_configure[19][9] ;
 wire \gpio_configure[1][0] ;
 wire \gpio_configure[1][10] ;
 wire \gpio_configure[1][11] ;
 wire \gpio_configure[1][12] ;
 wire \gpio_configure[1][1] ;
 wire \gpio_configure[1][2] ;
 wire \gpio_configure[1][3] ;
 wire \gpio_configure[1][4] ;
 wire \gpio_configure[1][5] ;
 wire \gpio_configure[1][6] ;
 wire \gpio_configure[1][7] ;
 wire \gpio_configure[1][8] ;
 wire \gpio_configure[1][9] ;
 wire \gpio_configure[20][0] ;
 wire \gpio_configure[20][10] ;
 wire \gpio_configure[20][11] ;
 wire \gpio_configure[20][12] ;
 wire \gpio_configure[20][1] ;
 wire \gpio_configure[20][2] ;
 wire \gpio_configure[20][3] ;
 wire \gpio_configure[20][4] ;
 wire \gpio_configure[20][5] ;
 wire \gpio_configure[20][6] ;
 wire \gpio_configure[20][7] ;
 wire \gpio_configure[20][8] ;
 wire \gpio_configure[20][9] ;
 wire \gpio_configure[21][0] ;
 wire \gpio_configure[21][10] ;
 wire \gpio_configure[21][11] ;
 wire \gpio_configure[21][12] ;
 wire \gpio_configure[21][1] ;
 wire \gpio_configure[21][2] ;
 wire \gpio_configure[21][3] ;
 wire \gpio_configure[21][4] ;
 wire \gpio_configure[21][5] ;
 wire \gpio_configure[21][6] ;
 wire \gpio_configure[21][7] ;
 wire \gpio_configure[21][8] ;
 wire \gpio_configure[21][9] ;
 wire \gpio_configure[22][0] ;
 wire \gpio_configure[22][10] ;
 wire \gpio_configure[22][11] ;
 wire \gpio_configure[22][12] ;
 wire \gpio_configure[22][1] ;
 wire \gpio_configure[22][2] ;
 wire \gpio_configure[22][3] ;
 wire \gpio_configure[22][4] ;
 wire \gpio_configure[22][5] ;
 wire \gpio_configure[22][6] ;
 wire \gpio_configure[22][7] ;
 wire \gpio_configure[22][8] ;
 wire \gpio_configure[22][9] ;
 wire \gpio_configure[23][0] ;
 wire \gpio_configure[23][10] ;
 wire \gpio_configure[23][11] ;
 wire \gpio_configure[23][12] ;
 wire \gpio_configure[23][1] ;
 wire \gpio_configure[23][2] ;
 wire \gpio_configure[23][3] ;
 wire \gpio_configure[23][4] ;
 wire \gpio_configure[23][5] ;
 wire \gpio_configure[23][6] ;
 wire \gpio_configure[23][7] ;
 wire \gpio_configure[23][8] ;
 wire \gpio_configure[23][9] ;
 wire \gpio_configure[24][0] ;
 wire \gpio_configure[24][10] ;
 wire \gpio_configure[24][11] ;
 wire \gpio_configure[24][12] ;
 wire \gpio_configure[24][1] ;
 wire \gpio_configure[24][2] ;
 wire \gpio_configure[24][3] ;
 wire \gpio_configure[24][4] ;
 wire \gpio_configure[24][5] ;
 wire \gpio_configure[24][6] ;
 wire \gpio_configure[24][7] ;
 wire \gpio_configure[24][8] ;
 wire \gpio_configure[24][9] ;
 wire \gpio_configure[25][0] ;
 wire \gpio_configure[25][10] ;
 wire \gpio_configure[25][11] ;
 wire \gpio_configure[25][12] ;
 wire \gpio_configure[25][1] ;
 wire \gpio_configure[25][2] ;
 wire \gpio_configure[25][3] ;
 wire \gpio_configure[25][4] ;
 wire \gpio_configure[25][5] ;
 wire \gpio_configure[25][6] ;
 wire \gpio_configure[25][7] ;
 wire \gpio_configure[25][8] ;
 wire \gpio_configure[25][9] ;
 wire \gpio_configure[26][0] ;
 wire \gpio_configure[26][10] ;
 wire \gpio_configure[26][11] ;
 wire \gpio_configure[26][12] ;
 wire \gpio_configure[26][1] ;
 wire \gpio_configure[26][2] ;
 wire \gpio_configure[26][3] ;
 wire \gpio_configure[26][4] ;
 wire \gpio_configure[26][5] ;
 wire \gpio_configure[26][6] ;
 wire \gpio_configure[26][7] ;
 wire \gpio_configure[26][8] ;
 wire \gpio_configure[26][9] ;
 wire \gpio_configure[27][0] ;
 wire \gpio_configure[27][10] ;
 wire \gpio_configure[27][11] ;
 wire \gpio_configure[27][12] ;
 wire \gpio_configure[27][1] ;
 wire \gpio_configure[27][2] ;
 wire \gpio_configure[27][3] ;
 wire \gpio_configure[27][4] ;
 wire \gpio_configure[27][5] ;
 wire \gpio_configure[27][6] ;
 wire \gpio_configure[27][7] ;
 wire \gpio_configure[27][8] ;
 wire \gpio_configure[27][9] ;
 wire \gpio_configure[28][0] ;
 wire \gpio_configure[28][10] ;
 wire \gpio_configure[28][11] ;
 wire \gpio_configure[28][12] ;
 wire \gpio_configure[28][1] ;
 wire \gpio_configure[28][2] ;
 wire \gpio_configure[28][3] ;
 wire \gpio_configure[28][4] ;
 wire \gpio_configure[28][5] ;
 wire \gpio_configure[28][6] ;
 wire \gpio_configure[28][7] ;
 wire \gpio_configure[28][8] ;
 wire \gpio_configure[28][9] ;
 wire \gpio_configure[29][0] ;
 wire \gpio_configure[29][10] ;
 wire \gpio_configure[29][11] ;
 wire \gpio_configure[29][12] ;
 wire \gpio_configure[29][1] ;
 wire \gpio_configure[29][2] ;
 wire \gpio_configure[29][3] ;
 wire \gpio_configure[29][4] ;
 wire \gpio_configure[29][5] ;
 wire \gpio_configure[29][6] ;
 wire \gpio_configure[29][7] ;
 wire \gpio_configure[29][8] ;
 wire \gpio_configure[29][9] ;
 wire \gpio_configure[2][0] ;
 wire \gpio_configure[2][10] ;
 wire \gpio_configure[2][11] ;
 wire \gpio_configure[2][12] ;
 wire \gpio_configure[2][1] ;
 wire \gpio_configure[2][2] ;
 wire \gpio_configure[2][3] ;
 wire \gpio_configure[2][4] ;
 wire \gpio_configure[2][5] ;
 wire \gpio_configure[2][6] ;
 wire \gpio_configure[2][7] ;
 wire \gpio_configure[2][8] ;
 wire \gpio_configure[2][9] ;
 wire \gpio_configure[30][0] ;
 wire \gpio_configure[30][10] ;
 wire \gpio_configure[30][11] ;
 wire \gpio_configure[30][12] ;
 wire \gpio_configure[30][1] ;
 wire \gpio_configure[30][2] ;
 wire \gpio_configure[30][3] ;
 wire \gpio_configure[30][4] ;
 wire \gpio_configure[30][5] ;
 wire \gpio_configure[30][6] ;
 wire \gpio_configure[30][7] ;
 wire \gpio_configure[30][8] ;
 wire \gpio_configure[30][9] ;
 wire \gpio_configure[31][0] ;
 wire \gpio_configure[31][10] ;
 wire \gpio_configure[31][11] ;
 wire \gpio_configure[31][12] ;
 wire \gpio_configure[31][1] ;
 wire \gpio_configure[31][2] ;
 wire \gpio_configure[31][3] ;
 wire \gpio_configure[31][4] ;
 wire \gpio_configure[31][5] ;
 wire \gpio_configure[31][6] ;
 wire \gpio_configure[31][7] ;
 wire \gpio_configure[31][8] ;
 wire \gpio_configure[31][9] ;
 wire \gpio_configure[32][0] ;
 wire \gpio_configure[32][10] ;
 wire \gpio_configure[32][11] ;
 wire \gpio_configure[32][12] ;
 wire \gpio_configure[32][1] ;
 wire \gpio_configure[32][2] ;
 wire \gpio_configure[32][3] ;
 wire \gpio_configure[32][4] ;
 wire \gpio_configure[32][5] ;
 wire \gpio_configure[32][6] ;
 wire \gpio_configure[32][7] ;
 wire \gpio_configure[32][8] ;
 wire \gpio_configure[32][9] ;
 wire \gpio_configure[33][0] ;
 wire \gpio_configure[33][10] ;
 wire \gpio_configure[33][11] ;
 wire \gpio_configure[33][12] ;
 wire \gpio_configure[33][1] ;
 wire \gpio_configure[33][2] ;
 wire \gpio_configure[33][3] ;
 wire \gpio_configure[33][4] ;
 wire \gpio_configure[33][5] ;
 wire \gpio_configure[33][6] ;
 wire \gpio_configure[33][7] ;
 wire \gpio_configure[33][8] ;
 wire \gpio_configure[33][9] ;
 wire \gpio_configure[34][0] ;
 wire \gpio_configure[34][10] ;
 wire \gpio_configure[34][11] ;
 wire \gpio_configure[34][12] ;
 wire \gpio_configure[34][1] ;
 wire \gpio_configure[34][2] ;
 wire \gpio_configure[34][3] ;
 wire \gpio_configure[34][4] ;
 wire \gpio_configure[34][5] ;
 wire \gpio_configure[34][6] ;
 wire \gpio_configure[34][7] ;
 wire \gpio_configure[34][8] ;
 wire \gpio_configure[34][9] ;
 wire \gpio_configure[35][0] ;
 wire \gpio_configure[35][10] ;
 wire \gpio_configure[35][11] ;
 wire \gpio_configure[35][12] ;
 wire \gpio_configure[35][1] ;
 wire \gpio_configure[35][2] ;
 wire \gpio_configure[35][3] ;
 wire \gpio_configure[35][4] ;
 wire \gpio_configure[35][5] ;
 wire \gpio_configure[35][6] ;
 wire \gpio_configure[35][7] ;
 wire \gpio_configure[35][8] ;
 wire \gpio_configure[35][9] ;
 wire \gpio_configure[36][0] ;
 wire \gpio_configure[36][10] ;
 wire \gpio_configure[36][11] ;
 wire \gpio_configure[36][12] ;
 wire \gpio_configure[36][1] ;
 wire \gpio_configure[36][2] ;
 wire \gpio_configure[36][3] ;
 wire \gpio_configure[36][4] ;
 wire \gpio_configure[36][5] ;
 wire \gpio_configure[36][6] ;
 wire \gpio_configure[36][7] ;
 wire \gpio_configure[36][8] ;
 wire \gpio_configure[36][9] ;
 wire \gpio_configure[37][0] ;
 wire \gpio_configure[37][10] ;
 wire \gpio_configure[37][11] ;
 wire \gpio_configure[37][12] ;
 wire \gpio_configure[37][1] ;
 wire \gpio_configure[37][2] ;
 wire \gpio_configure[37][3] ;
 wire \gpio_configure[37][4] ;
 wire \gpio_configure[37][5] ;
 wire \gpio_configure[37][6] ;
 wire \gpio_configure[37][7] ;
 wire \gpio_configure[37][8] ;
 wire \gpio_configure[37][9] ;
 wire \gpio_configure[3][0] ;
 wire \gpio_configure[3][10] ;
 wire \gpio_configure[3][11] ;
 wire \gpio_configure[3][12] ;
 wire \gpio_configure[3][1] ;
 wire \gpio_configure[3][2] ;
 wire \gpio_configure[3][3] ;
 wire \gpio_configure[3][4] ;
 wire \gpio_configure[3][5] ;
 wire \gpio_configure[3][6] ;
 wire \gpio_configure[3][7] ;
 wire \gpio_configure[3][8] ;
 wire \gpio_configure[3][9] ;
 wire \gpio_configure[4][0] ;
 wire \gpio_configure[4][10] ;
 wire \gpio_configure[4][11] ;
 wire \gpio_configure[4][12] ;
 wire \gpio_configure[4][1] ;
 wire \gpio_configure[4][2] ;
 wire \gpio_configure[4][3] ;
 wire \gpio_configure[4][4] ;
 wire \gpio_configure[4][5] ;
 wire \gpio_configure[4][6] ;
 wire \gpio_configure[4][7] ;
 wire \gpio_configure[4][8] ;
 wire \gpio_configure[4][9] ;
 wire \gpio_configure[5][0] ;
 wire \gpio_configure[5][10] ;
 wire \gpio_configure[5][11] ;
 wire \gpio_configure[5][12] ;
 wire \gpio_configure[5][1] ;
 wire \gpio_configure[5][2] ;
 wire \gpio_configure[5][3] ;
 wire \gpio_configure[5][4] ;
 wire \gpio_configure[5][5] ;
 wire \gpio_configure[5][6] ;
 wire \gpio_configure[5][7] ;
 wire \gpio_configure[5][8] ;
 wire \gpio_configure[5][9] ;
 wire \gpio_configure[6][0] ;
 wire \gpio_configure[6][10] ;
 wire \gpio_configure[6][11] ;
 wire \gpio_configure[6][12] ;
 wire \gpio_configure[6][1] ;
 wire \gpio_configure[6][2] ;
 wire \gpio_configure[6][3] ;
 wire \gpio_configure[6][4] ;
 wire \gpio_configure[6][5] ;
 wire \gpio_configure[6][6] ;
 wire \gpio_configure[6][7] ;
 wire \gpio_configure[6][8] ;
 wire \gpio_configure[6][9] ;
 wire \gpio_configure[7][0] ;
 wire \gpio_configure[7][10] ;
 wire \gpio_configure[7][11] ;
 wire \gpio_configure[7][12] ;
 wire \gpio_configure[7][1] ;
 wire \gpio_configure[7][2] ;
 wire \gpio_configure[7][3] ;
 wire \gpio_configure[7][4] ;
 wire \gpio_configure[7][5] ;
 wire \gpio_configure[7][6] ;
 wire \gpio_configure[7][7] ;
 wire \gpio_configure[7][8] ;
 wire \gpio_configure[7][9] ;
 wire \gpio_configure[8][0] ;
 wire \gpio_configure[8][10] ;
 wire \gpio_configure[8][11] ;
 wire \gpio_configure[8][12] ;
 wire \gpio_configure[8][1] ;
 wire \gpio_configure[8][2] ;
 wire \gpio_configure[8][3] ;
 wire \gpio_configure[8][4] ;
 wire \gpio_configure[8][5] ;
 wire \gpio_configure[8][6] ;
 wire \gpio_configure[8][7] ;
 wire \gpio_configure[8][8] ;
 wire \gpio_configure[8][9] ;
 wire \gpio_configure[9][0] ;
 wire \gpio_configure[9][10] ;
 wire \gpio_configure[9][11] ;
 wire \gpio_configure[9][12] ;
 wire \gpio_configure[9][1] ;
 wire \gpio_configure[9][2] ;
 wire \gpio_configure[9][3] ;
 wire \gpio_configure[9][4] ;
 wire \gpio_configure[9][5] ;
 wire \gpio_configure[9][6] ;
 wire \gpio_configure[9][7] ;
 wire \gpio_configure[9][8] ;
 wire \gpio_configure[9][9] ;
 wire \hkspi.SDO ;
 wire \hkspi.addr[0] ;
 wire \hkspi.addr[1] ;
 wire \hkspi.addr[2] ;
 wire \hkspi.addr[3] ;
 wire \hkspi.addr[4] ;
 wire \hkspi.addr[5] ;
 wire \hkspi.addr[6] ;
 wire \hkspi.addr[7] ;
 wire \hkspi.count[0] ;
 wire \hkspi.count[1] ;
 wire \hkspi.count[2] ;
 wire \hkspi.fixed[0] ;
 wire \hkspi.fixed[1] ;
 wire \hkspi.fixed[2] ;
 wire \hkspi.ldata[0] ;
 wire \hkspi.ldata[1] ;
 wire \hkspi.ldata[2] ;
 wire \hkspi.ldata[3] ;
 wire \hkspi.ldata[4] ;
 wire \hkspi.ldata[5] ;
 wire \hkspi.ldata[6] ;
 wire \hkspi.odata[1] ;
 wire \hkspi.odata[2] ;
 wire \hkspi.odata[3] ;
 wire \hkspi.odata[4] ;
 wire \hkspi.odata[5] ;
 wire \hkspi.odata[6] ;
 wire \hkspi.odata[7] ;
 wire \hkspi.pass_thru_mgmt ;
 wire \hkspi.pass_thru_mgmt_delay ;
 wire \hkspi.pass_thru_user ;
 wire \hkspi.pass_thru_user_delay ;
 wire \hkspi.pre_pass_thru_mgmt ;
 wire \hkspi.pre_pass_thru_user ;
 wire \hkspi.rdstb ;
 wire \hkspi.readmode ;
 wire \hkspi.sdoenb ;
 wire \hkspi.state[0] ;
 wire \hkspi.state[1] ;
 wire \hkspi.state[2] ;
 wire \hkspi.state[3] ;
 wire \hkspi.state[4] ;
 wire \hkspi.writemode ;
 wire \hkspi.wrstb ;
 wire hkspi_disable;
 wire irq_1_inputsrc;
 wire irq_2_inputsrc;
 wire irq_spi;
 wire \mgmt_gpio_data[0] ;
 wire \mgmt_gpio_data[10] ;
 wire \mgmt_gpio_data[11] ;
 wire \mgmt_gpio_data[12] ;
 wire \mgmt_gpio_data[13] ;
 wire \mgmt_gpio_data[14] ;
 wire \mgmt_gpio_data[15] ;
 wire \mgmt_gpio_data[16] ;
 wire \mgmt_gpio_data[17] ;
 wire \mgmt_gpio_data[18] ;
 wire \mgmt_gpio_data[19] ;
 wire \mgmt_gpio_data[1] ;
 wire \mgmt_gpio_data[20] ;
 wire \mgmt_gpio_data[21] ;
 wire \mgmt_gpio_data[22] ;
 wire \mgmt_gpio_data[23] ;
 wire \mgmt_gpio_data[24] ;
 wire \mgmt_gpio_data[25] ;
 wire \mgmt_gpio_data[26] ;
 wire \mgmt_gpio_data[27] ;
 wire \mgmt_gpio_data[28] ;
 wire \mgmt_gpio_data[29] ;
 wire \mgmt_gpio_data[2] ;
 wire \mgmt_gpio_data[30] ;
 wire \mgmt_gpio_data[31] ;
 wire \mgmt_gpio_data[32] ;
 wire \mgmt_gpio_data[33] ;
 wire \mgmt_gpio_data[34] ;
 wire \mgmt_gpio_data[35] ;
 wire \mgmt_gpio_data[36] ;
 wire \mgmt_gpio_data[37] ;
 wire \mgmt_gpio_data[3] ;
 wire \mgmt_gpio_data[4] ;
 wire \mgmt_gpio_data[5] ;
 wire \mgmt_gpio_data[6] ;
 wire \mgmt_gpio_data[7] ;
 wire \mgmt_gpio_data[8] ;
 wire \mgmt_gpio_data[9] ;
 wire \mgmt_gpio_data_buf[0] ;
 wire \mgmt_gpio_data_buf[10] ;
 wire \mgmt_gpio_data_buf[11] ;
 wire \mgmt_gpio_data_buf[12] ;
 wire \mgmt_gpio_data_buf[13] ;
 wire \mgmt_gpio_data_buf[14] ;
 wire \mgmt_gpio_data_buf[15] ;
 wire \mgmt_gpio_data_buf[16] ;
 wire \mgmt_gpio_data_buf[17] ;
 wire \mgmt_gpio_data_buf[18] ;
 wire \mgmt_gpio_data_buf[19] ;
 wire \mgmt_gpio_data_buf[1] ;
 wire \mgmt_gpio_data_buf[20] ;
 wire \mgmt_gpio_data_buf[21] ;
 wire \mgmt_gpio_data_buf[22] ;
 wire \mgmt_gpio_data_buf[23] ;
 wire \mgmt_gpio_data_buf[2] ;
 wire \mgmt_gpio_data_buf[3] ;
 wire \mgmt_gpio_data_buf[4] ;
 wire \mgmt_gpio_data_buf[5] ;
 wire \mgmt_gpio_data_buf[6] ;
 wire \mgmt_gpio_data_buf[7] ;
 wire \mgmt_gpio_data_buf[8] ;
 wire \mgmt_gpio_data_buf[9] ;
 wire mgmt_gpio_out_14_prebuff;
 wire mgmt_gpio_out_15_prebuff;
 wire mgmt_gpio_out_30_prebuff;
 wire mgmt_gpio_out_31_prebuff;
 wire mgmt_gpio_out_9_prebuff;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net375;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net376;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net377;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net378;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net379;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net380;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net381;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net382;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net383;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net384;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net385;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net386;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net387;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net388;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net389;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net39;
 wire net390;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \pad_count_1[0] ;
 wire \pad_count_1[1] ;
 wire \pad_count_1[2] ;
 wire \pad_count_1[3] ;
 wire \pad_count_1[4] ;
 wire \pad_count_2[0] ;
 wire \pad_count_2[1] ;
 wire \pad_count_2[2] ;
 wire \pad_count_2[3] ;
 wire \pad_count_2[4] ;
 wire \pad_count_2[5] ;
 wire pad_flash_clk_prebuff;
 wire reset_reg;
 wire serial_bb_clock;
 wire serial_bb_data_1;
 wire serial_bb_data_2;
 wire serial_bb_enable;
 wire serial_bb_load;
 wire serial_bb_resetn;
 wire serial_busy;
 wire serial_clock_pre;
 wire \serial_data_staging_1[0] ;
 wire \serial_data_staging_1[10] ;
 wire \serial_data_staging_1[11] ;
 wire \serial_data_staging_1[12] ;
 wire \serial_data_staging_1[1] ;
 wire \serial_data_staging_1[2] ;
 wire \serial_data_staging_1[3] ;
 wire \serial_data_staging_1[4] ;
 wire \serial_data_staging_1[5] ;
 wire \serial_data_staging_1[6] ;
 wire \serial_data_staging_1[7] ;
 wire \serial_data_staging_1[8] ;
 wire \serial_data_staging_1[9] ;
 wire \serial_data_staging_2[0] ;
 wire \serial_data_staging_2[10] ;
 wire \serial_data_staging_2[11] ;
 wire \serial_data_staging_2[12] ;
 wire \serial_data_staging_2[1] ;
 wire \serial_data_staging_2[2] ;
 wire \serial_data_staging_2[3] ;
 wire \serial_data_staging_2[4] ;
 wire \serial_data_staging_2[5] ;
 wire \serial_data_staging_2[6] ;
 wire \serial_data_staging_2[7] ;
 wire \serial_data_staging_2[8] ;
 wire \serial_data_staging_2[9] ;
 wire serial_load_pre;
 wire serial_resetn_pre;
 wire serial_xfer;
 wire trap_output_dest;
 wire \wbbd_addr[0] ;
 wire \wbbd_addr[1] ;
 wire \wbbd_addr[2] ;
 wire \wbbd_addr[3] ;
 wire \wbbd_addr[4] ;
 wire \wbbd_addr[5] ;
 wire \wbbd_addr[6] ;
 wire wbbd_busy;
 wire \wbbd_data[0] ;
 wire \wbbd_data[1] ;
 wire \wbbd_data[2] ;
 wire \wbbd_data[3] ;
 wire \wbbd_data[4] ;
 wire \wbbd_data[5] ;
 wire \wbbd_data[6] ;
 wire \wbbd_data[7] ;
 wire wbbd_sck;
 wire \wbbd_state[0] ;
 wire \wbbd_state[10] ;
 wire \wbbd_state[1] ;
 wire \wbbd_state[2] ;
 wire \wbbd_state[3] ;
 wire \wbbd_state[4] ;
 wire \wbbd_state[5] ;
 wire \wbbd_state[6] ;
 wire \wbbd_state[7] ;
 wire \wbbd_state[8] ;
 wire \wbbd_state[9] ;
 wire wbbd_write;
 wire \xfer_count[0] ;
 wire \xfer_count[1] ;
 wire \xfer_count[2] ;
 wire \xfer_count[3] ;
 wire \xfer_state[0] ;
 wire \xfer_state[1] ;
 wire \xfer_state[2] ;
 wire \xfer_state[3] ;
 wire [4:0] \xfer_sta ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_3114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_3189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_3224_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_3302_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_3338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1084_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_1861_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A (.DIODE(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A (.DIODE(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A (.DIODE(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A (.DIODE(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A (.DIODE(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A (.DIODE(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A (.DIODE(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A (.DIODE(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A (.DIODE(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A (.DIODE(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A (.DIODE(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A (.DIODE(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A (.DIODE(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A (.DIODE(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A (.DIODE(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A (.DIODE(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A (.DIODE(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A (.DIODE(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A_N (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A_N (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B1_N (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__C (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__C (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__C (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__C (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__C (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A1 (.DIODE(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__C1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__C (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__C (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__C (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__C (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__C (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__C (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A2 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__B1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A2 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B1 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B1 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B2 (.DIODE(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A2 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__C (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__C (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__C (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A1 (.DIODE(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__C (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__C (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__B (.DIODE(net2070));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__B (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A1 (.DIODE(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B2 (.DIODE(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A2 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B2 (.DIODE(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B2 (.DIODE(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__C (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__C (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A1 (.DIODE(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__B1 (.DIODE(_0941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A2 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A (.DIODE(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__B (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__C (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__C (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A1 (.DIODE(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B2 (.DIODE(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A1 (.DIODE(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A (.DIODE(net2070));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A_N (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B2 (.DIODE(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__C1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A3 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B1 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A2 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B2 (.DIODE(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__B1 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A2 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__C (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A3 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B2 (.DIODE(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A2 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B2 (.DIODE(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B1 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B1 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B2 (.DIODE(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A1 (.DIODE(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B2 (.DIODE(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B2 (.DIODE(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A1 (.DIODE(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A2 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__B1 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__B2 (.DIODE(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A2 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B2 (.DIODE(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__S (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A3 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__B1 (.DIODE(_0941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B2 (.DIODE(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B2 (.DIODE(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__B1 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B1 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B2 (.DIODE(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__B2 (.DIODE(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B2 (.DIODE(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B2 (.DIODE(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A2 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__C (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__C (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__D (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__B (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__C (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__C (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__C (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A1 (.DIODE(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A3 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A4 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A1 (.DIODE(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A2 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A1 (.DIODE(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B2 (.DIODE(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A1 (.DIODE(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__B1 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A1 (.DIODE(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A1 (.DIODE(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B1 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B2 (.DIODE(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A2 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__B2 (.DIODE(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A1 (.DIODE(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B2 (.DIODE(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A3 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A2 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B1 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B2 (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A1 (.DIODE(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A1 (.DIODE(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__B2 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B1 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B2 (.DIODE(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B2 (.DIODE(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A3 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A4 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A3 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A1 (.DIODE(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__B2 (.DIODE(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A2 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B2 (.DIODE(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A1 (.DIODE(\clk1_output_dest[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A1 (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B2 (.DIODE(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__C1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A3 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A4 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A3 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A2 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B1 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A1 (.DIODE(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A1 (.DIODE(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A1 (.DIODE(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A4 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A1 (.DIODE(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A1 (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A1 (.DIODE(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B2 (.DIODE(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A1 (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A3 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__B2 (.DIODE(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A1 (.DIODE(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A2 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B2 (.DIODE(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A2 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B2 (.DIODE(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A1 (.DIODE(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B2 (.DIODE(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B2 (.DIODE(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B2 (.DIODE(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B1 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B2 (.DIODE(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A1 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B2 (.DIODE(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A1 (.DIODE(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B2 (.DIODE(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B2 (.DIODE(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__C1 (.DIODE(_1139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B1 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A1 (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A3 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A1 (.DIODE(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__B2 (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A1 (.DIODE(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A2 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B2 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A1 (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B2 (.DIODE(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A2 (.DIODE(_0941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B2 (.DIODE(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A3 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B2 (.DIODE(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A3 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__C1 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__B1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A_N (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A1 (.DIODE(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A3 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__B2 (.DIODE(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A1 (.DIODE(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A3 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B1 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A1 (.DIODE(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B2 (.DIODE(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__C1 (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A2 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B1 (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A1 (.DIODE(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B2 (.DIODE(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A3 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B2 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B2 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A2 (.DIODE(_0941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B2 (.DIODE(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B2 (.DIODE(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A2 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A2 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A3 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A2 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B1 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A1 (.DIODE(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A3 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B2 (.DIODE(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A1 (.DIODE(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B2 (.DIODE(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A1 (.DIODE(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__B2 (.DIODE(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A1 (.DIODE(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A3 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B2 (.DIODE(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A1 (.DIODE(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B2 (.DIODE(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A3 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A3 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(_1222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A2 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__D1 (.DIODE(_1228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B (.DIODE(_1231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A (.DIODE(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__D (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__C (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__D (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__C (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__D (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__C (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__B (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__C (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__D (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__B2 (.DIODE(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A2 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A1 (.DIODE(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B2 (.DIODE(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B2 (.DIODE(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A1 (.DIODE(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A2 (.DIODE(_0881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A1 (.DIODE(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A3 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A4 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A1 (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A3 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__B2 (.DIODE(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A1 (.DIODE(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__B2 (.DIODE(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1 (.DIODE(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A3 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B2 (.DIODE(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A1 (.DIODE(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__B1 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A1 (.DIODE(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B2 (.DIODE(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__B1 (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A1 (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A1 (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A1 (.DIODE(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B2 (.DIODE(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A2 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A2 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B2 (.DIODE(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B2 (.DIODE(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B1 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__B2 (.DIODE(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A2 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B1 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A3 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__C1 (.DIODE(_1292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A2 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__B2 (.DIODE(\clk2_output_dest[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A1 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__C (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__D (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__C (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__D (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__D (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__B (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__D (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A2 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A3 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B1 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B2 (.DIODE(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__A3 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A1 (.DIODE(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A3 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A3 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A4 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A1 (.DIODE(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A3 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B1 (.DIODE(_0884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A2 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A2 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A1 (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__C1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A2 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A3 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A3 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A3 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A2 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__B2 (.DIODE(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A1 (.DIODE(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A3 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__B1 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A1 (.DIODE(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B2 (.DIODE(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B1 (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B2 (.DIODE(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B2 (.DIODE(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A1 (.DIODE(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A3 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A3 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A1 (.DIODE(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A2 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B1 (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B2 (.DIODE(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A1 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B2 (.DIODE(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A2 (.DIODE(_0908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A2 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A3 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A2 (.DIODE(_0941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__B1 (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A3 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A3 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A3 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__B1 (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A1 (.DIODE(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B2 (.DIODE(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A3 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A2 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A1 (.DIODE(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A2 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B1 (.DIODE(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A3 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B2 (.DIODE(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A2 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A2 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B2 (.DIODE(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A1 (.DIODE(irq_spi));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A3 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B2 (.DIODE(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A1 (.DIODE(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A2 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A3 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A4 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B1 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B2 (.DIODE(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A3 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__B2 (.DIODE(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A1 (.DIODE(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A3 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B1 (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__B2 (.DIODE(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__C1 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A0 (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B (.DIODE(net2388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__C (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__S (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A1 (.DIODE(\hkspi.rdstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A2 (.DIODE(\hkspi.wrstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A1 (.DIODE(\hkspi.rdstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A2 (.DIODE(\hkspi.wrstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A_N (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A_N (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A2 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A3 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A1 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__C1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__S (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1 (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__S (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A_N (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__S (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A_N (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A_N (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A1 (.DIODE(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A1 (.DIODE(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B1 (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__S (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1 (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__S (.DIODE(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A0 (.DIODE(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A1 (.DIODE(\hkspi.SDO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__S (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__S (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__S (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A1 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A2 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__B1 (.DIODE(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A1 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A2 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A4 (.DIODE(\hkspi.sdoenb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B1 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__S (.DIODE(\clk2_output_dest[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A1 (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A1 (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__S (.DIODE(\clk1_output_dest[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__S (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__S (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__C (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__D (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__B (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A0 (.DIODE(\hkspi.wrstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A2 (.DIODE(net2388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(net2017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__S (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__B1 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__C1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__S (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__C1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(net2017));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__B (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A2 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A0 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A2 (.DIODE(_1231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A0 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A0 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A0 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A2 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A0 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__A (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A2 (.DIODE(_1231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A0 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__S (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A0 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A0 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A2 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A0 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A2 (.DIODE(_1231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A0 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__S (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A0 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__S (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A0 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__S (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A0 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__D (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__C (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__C (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A (.DIODE(_1040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__C (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__C (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__B (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__C (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__D (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A_N (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__B (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__C (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__C (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__D (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A0 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__C (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__D (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__C (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__D (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__D (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A0 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A0 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__B (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__C (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__C (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__D (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__C (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__D (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__D (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__D (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__B (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__D (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__D (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__D (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__C (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A_N (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A_N (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A_N (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A_N (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__D (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__B (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__C1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__C1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__C1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__D1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__B (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__B (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__B (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__B1_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B1_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__B (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__C (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__C (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__C (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B1_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A3 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A4 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__D (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__D (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A4 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__D (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__B (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A4 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A3 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B1_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__D (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A2 (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__C (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B1_N (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__C (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__C (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__C (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__C (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__C (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__C (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__D (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__B (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__C (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__C (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__D_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B_N (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__D (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A_N (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__D (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A_N (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A_N (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__D (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__C (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A2 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__C (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__C (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__C (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__D (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A_N (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__C (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__D (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__D (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__C (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__C (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__C (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__C (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A_N (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__C (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__C (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__D (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__C (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__B (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__C (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__D (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A_N (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__D (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__C (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__C (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A3 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__D (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B1 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A3 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A3 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__C (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A_N (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B_N (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__D (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__B2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__C (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A_N (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__C (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__D (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__C (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__C (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A_N (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__D (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__B (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__C1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__C (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__D (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A_N (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__C (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__D (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__C (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__D (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__D (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__C (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__B (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__C (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__B (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__D (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__C (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__C (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__B (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__D (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__D (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__D (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A2 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A3 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B2 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A2 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A3 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A3 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__C (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A4 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A4 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__C (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B1 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__C (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__C1 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__B (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__D (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__C (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__C (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__C (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__D (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__C (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__C (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__C1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__D1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__C1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__D1 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A3 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B1 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__C (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B1 (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__C1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__D1 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__C1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__D1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__C1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__D1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__C (.DIODE(_2001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__D1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__C (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__D1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__B (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__C (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__B2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A_N (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__B2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__C (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__C (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__C (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__C (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A3 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__C (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__B2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B1 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__D (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A2 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__C (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__B (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__C (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__C (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__C (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A3 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B1 (.DIODE(_2001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B2 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__D (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A_N (.DIODE(_2017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A3 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A3 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A3 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A3 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A3 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__B2 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A3 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A3 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__C (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A3 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__C (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A2 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A2 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A3 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__D1 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A_N (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B2 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A3 (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__D (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A2 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A3 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__C (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A2 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B2 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__C1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A3 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__D (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A3 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B1 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__C1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A3 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A2 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A3 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__D1 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__C1 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__B1 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A2 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__C1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A2 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__C1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A2 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B2 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A3 (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B1 (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A2 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A2 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A3 (.DIODE(_1949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A2 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A3 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__C1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A3 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__C1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A3 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A4 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A_N (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__C (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A4 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A2 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A3 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A4 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A3 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A4 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A2 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__C (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B2 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__D (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A3 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B2 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A2 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A3 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A2 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A3 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B1 (.DIODE(_1868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A3 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A3 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__C (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A3 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A1 (.DIODE(_1604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A1 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A3 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B1 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A1 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A3 (.DIODE(_1975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A1 (.DIODE(_1707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A2 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__C1 (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A1 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A2 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A3 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__C1 (.DIODE(_1609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__C1 (.DIODE(_1881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A3 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A3 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A1 (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A3 (.DIODE(_1950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B2 (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A2 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A3 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(_1629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(_1628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A3 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A1 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B1 (.DIODE(_1661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_1883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_1726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A0 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A0 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A0 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__C (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__B (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__C (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__C1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__C (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__B (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A0 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__D (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A0 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A0 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__S (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A3 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__B1 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__C1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A0 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__D (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__S (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__S (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__S (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__B (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__S (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A (.DIODE(_0938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__S (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__B (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__S (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(_0865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A0 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A0 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__S (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__C (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__S (.DIODE(_2611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__C (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__S (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__C (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__S (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A0 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S (.DIODE(_2615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__B (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A0 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__S (.DIODE(_2616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__C (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__S (.DIODE(_2618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__S (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A0 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A0 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A0 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__S (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A0 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A0 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A0 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A0 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__C (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__C (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__S (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A0 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A0 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A0 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A0 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A0 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A0 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__C (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__S (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__S (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__B1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__C (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__B1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__B (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A2 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__B (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__D (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A2 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__C (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__B1 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__C1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__C1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A_N (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__C (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__C (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__C (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__C (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A1 (.DIODE(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A1 (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A_N (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__B_N (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__C (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__C (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B_N (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__C (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B1 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B2 (.DIODE(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__B (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__C (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B2 (.DIODE(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__C (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__C (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__D (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__C (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__D (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__C (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__D (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A1 (.DIODE(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B2 (.DIODE(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A2 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__B1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__B2 (.DIODE(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__B2 (.DIODE(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A_N (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__C (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__D (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__C (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__D (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__B1 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B1 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B2 (.DIODE(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A1 (.DIODE(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B2 (.DIODE(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__B (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__C (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B2 (.DIODE(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__B1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__C (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__D (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__C (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B_N (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__C (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__D (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A1 (.DIODE(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A1 (.DIODE(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B2 (.DIODE(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__C (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B2 (.DIODE(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__C (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__D (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A2 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__B1 (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A1 (.DIODE(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B2 (.DIODE(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B2 (.DIODE(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B2 (.DIODE(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A1 (.DIODE(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B2 (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__B2 (.DIODE(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A1 (.DIODE(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__B2 (.DIODE(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B2 (.DIODE(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A1 (.DIODE(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A3 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B2 (.DIODE(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A1 (.DIODE(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B2 (.DIODE(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__C (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A2 (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B2 (.DIODE(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A1 (.DIODE(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A3 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__B2 (.DIODE(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A3 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A4 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A4 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B2 (.DIODE(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A3 (.DIODE(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B2 (.DIODE(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B1 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A1 (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B2 (.DIODE(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A2 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B2 (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A1 (.DIODE(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__B1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A3 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A1 (.DIODE(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B1 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B2 (.DIODE(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A1 (.DIODE(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B2 (.DIODE(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A1 (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B2 (.DIODE(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A1 (.DIODE(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B2 (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A1 (.DIODE(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A3 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A1 (.DIODE(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B2 (.DIODE(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A1 (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B2 (.DIODE(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A1 (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B2 (.DIODE(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A1 (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A3 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B1 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B2 (.DIODE(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A1 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B2 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B1 (.DIODE(_2788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B2 (.DIODE(_2799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A3 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__B2 (.DIODE(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A1 (.DIODE(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__B2 (.DIODE(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A1 (.DIODE(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B2 (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A1 (.DIODE(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A1 (.DIODE(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B2 (.DIODE(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A1 (.DIODE(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A1 (.DIODE(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A2 (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A2 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__B1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1 (.DIODE(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B2 (.DIODE(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A1 (.DIODE(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A2 (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A3 (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__B1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A3 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__B1 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__B1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A2_N (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A1 (.DIODE(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__B2 (.DIODE(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__B1 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A1 (.DIODE(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A3 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A3 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B2 (.DIODE(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A1 (.DIODE(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__B2 (.DIODE(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A1 (.DIODE(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__B1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__B1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A1 (.DIODE(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A4 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B2 (.DIODE(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A3 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A2 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B1 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__B2 (.DIODE(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__A2 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A4 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A3 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__B1 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A2 (.DIODE(_2729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B2 (.DIODE(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A3 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__B2 (.DIODE(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B2 (.DIODE(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__B2 (.DIODE(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A3 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B1 (.DIODE(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A1 (.DIODE(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__C1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B2 (.DIODE(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A1 (.DIODE(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__B1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__B2 (.DIODE(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B2 (.DIODE(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A3 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__C1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A3 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B2 (.DIODE(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A2 (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A3 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A1 (.DIODE(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B1 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B2 (.DIODE(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A3 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B2 (.DIODE(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A1 (.DIODE(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A1 (.DIODE(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B1 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__B1 (.DIODE(_2887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A1 (.DIODE(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B2 (.DIODE(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B2 (.DIODE(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A1 (.DIODE(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B2 (.DIODE(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A1 (.DIODE(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1 (.DIODE(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A3 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A4 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__B1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A1 (.DIODE(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__B1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A3 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__B1 (.DIODE(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__B2 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__B2 (.DIODE(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A2 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B2 (.DIODE(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__B2 (.DIODE(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__B2 (.DIODE(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A1 (.DIODE(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B2 (.DIODE(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B1 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__C1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B2 (.DIODE(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__B (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__C (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__B1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__B2 (.DIODE(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A1 (.DIODE(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A1 (.DIODE(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A1 (.DIODE(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A1 (.DIODE(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__B1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A2 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A3 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__B1 (.DIODE(_2707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B2 (.DIODE(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__B1 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__C (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__B1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__C1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B2 (.DIODE(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B2 (.DIODE(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A2 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A3 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B2 (.DIODE(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A2 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B2 (.DIODE(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B1 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B2 (.DIODE(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A1 (.DIODE(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A2 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A3 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B1 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B2 (.DIODE(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A1 (.DIODE(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B2 (.DIODE(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A2 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A1 (.DIODE(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A1 (.DIODE(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A3 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A1 (.DIODE(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A2 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A3 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B2 (.DIODE(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B2 (.DIODE(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A2 (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A1 (.DIODE(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__B2 (.DIODE(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B1 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B2 (.DIODE(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B2 (.DIODE(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A2 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A3 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B2 (.DIODE(_2713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A3 (.DIODE(_2704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__B1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__C1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A1_N (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A2 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__B1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A2 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A3 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A3 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A2 (.DIODE(_2687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A3 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A4 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A2 (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__B1 (.DIODE(_2694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A1 (.DIODE(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B2 (.DIODE(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A1 (.DIODE(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__C1 (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A3 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B1 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A2 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A2 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A3 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B1 (.DIODE(_2688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B1 (.DIODE(_2723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A3 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__B1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__B1 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A2 (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A3 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A2 (.DIODE(_2683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B2 (.DIODE(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A1 (.DIODE(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A2 (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__C (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__B (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__C (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__D (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__C (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__D1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__C (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B_N (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__C (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__C (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__D (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__C (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__B (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__C (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__C (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__C (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__D (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__C (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A1 (.DIODE(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A1 (.DIODE(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A2 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B2 (.DIODE(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B1 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__B2 (.DIODE(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A1 (.DIODE(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A1 (.DIODE(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A2 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B2 (.DIODE(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__C (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A1 (.DIODE(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A2 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B1 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B1 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__C (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__C (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A1 (.DIODE(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__B2 (.DIODE(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A1 (.DIODE(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A1 (.DIODE(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B2 (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__B (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A1 (.DIODE(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A2 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__B1 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__C (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A3 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__C (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__C (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A2 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__B (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__C (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__D (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A1 (.DIODE(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B2 (.DIODE(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__B1 (.DIODE(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__B2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A2 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__B1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__B2 (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A2 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A3 (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__B2 (.DIODE(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B2 (.DIODE(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A1 (.DIODE(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B2 (.DIODE(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A1 (.DIODE(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A3 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A3 (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B2 (.DIODE(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A1 (.DIODE(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A1 (.DIODE(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B2 (.DIODE(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B2 (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A1 (.DIODE(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A2 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__B2 (.DIODE(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B1 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B2 (.DIODE(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__B1 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__B2 (.DIODE(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A1 (.DIODE(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A2 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__B1 (.DIODE(_3094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A1 (.DIODE(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__B2 (.DIODE(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B1 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B2 (.DIODE(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__B2 (.DIODE(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B1 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__B2 (.DIODE(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A2 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A3 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A4 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A2 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A1 (.DIODE(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B2 (.DIODE(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A1 (.DIODE(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__B2 (.DIODE(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A1 (.DIODE(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B2 (.DIODE(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A1 (.DIODE(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A2 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A2 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__B1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B1 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A1 (.DIODE(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__B2 (.DIODE(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A1 (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__B2 (.DIODE(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A1 (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__B2 (.DIODE(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1 (.DIODE(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B1 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B2 (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A1 (.DIODE(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A1 (.DIODE(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A2 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A1 (.DIODE(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__B2 (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A1 (.DIODE(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A2 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B2 (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B2 (.DIODE(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A1 (.DIODE(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A1 (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A1 (.DIODE(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A3 (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B2 (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A1 (.DIODE(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A2 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__B2 (.DIODE(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A1 (.DIODE(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A2 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__B1 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__B2 (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A1 (.DIODE(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B2 (.DIODE(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A1 (.DIODE(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A1 (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B2 (.DIODE(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A1 (.DIODE(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B2 (.DIODE(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A1 (.DIODE(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B2 (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__B1 (.DIODE(_3142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__B1 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A1 (.DIODE(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A2 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A1 (.DIODE(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B2 (.DIODE(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A3 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B1 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B2 (.DIODE(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A1 (.DIODE(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A1 (.DIODE(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A2 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B2 (.DIODE(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A1 (.DIODE(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B2 (.DIODE(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B2 (.DIODE(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A1 (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B2 (.DIODE(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B1 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B2 (.DIODE(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A1 (.DIODE(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B1 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B2 (.DIODE(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__B2 (.DIODE(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B1 (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__B1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A (.DIODE(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__C (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B1 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B2 (.DIODE(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__B2 (.DIODE(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A1 (.DIODE(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A2 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B2 (.DIODE(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__B1 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A1 (.DIODE(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A3 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B1 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B2 (.DIODE(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A1 (.DIODE(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__C1 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A1 (.DIODE(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A2 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B2 (.DIODE(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1 (.DIODE(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A3 (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B2 (.DIODE(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A2 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__B1 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__C (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A1 (.DIODE(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A2 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B2 (.DIODE(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A1 (.DIODE(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B2 (.DIODE(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A2 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B1 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A2 (.DIODE(_1439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A3 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A4 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A1 (.DIODE(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A1 (.DIODE(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B2 (.DIODE(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__B1 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A2 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A2 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B2 (.DIODE(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A1 (.DIODE(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__B2 (.DIODE(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A2 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B1 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A2 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B2 (.DIODE(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A1 (.DIODE(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A2 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B2 (.DIODE(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A1 (.DIODE(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A2 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A2 (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__B1 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__B2 (.DIODE(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A2 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B2 (.DIODE(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__B2 (.DIODE(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A3 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__B1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__C (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A2 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__B2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__C (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A1 (.DIODE(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__B2 (.DIODE(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A1 (.DIODE(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__B1 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__B2 (.DIODE(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__B2 (.DIODE(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B2 (.DIODE(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A1 (.DIODE(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A1 (.DIODE(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A1 (.DIODE(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B1 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A1 (.DIODE(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A1 (.DIODE(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A1 (.DIODE(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B2 (.DIODE(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A2 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__C1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A1 (.DIODE(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A1 (.DIODE(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B2 (.DIODE(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A2 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B2 (.DIODE(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A1 (.DIODE(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A2 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__B1 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A2 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B2 (.DIODE(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B2 (.DIODE(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B2 (.DIODE(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A2 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B1 (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A1 (.DIODE(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A1 (.DIODE(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A1 (.DIODE(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B1 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__B2 (.DIODE(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__B2 (.DIODE(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__B1 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B1 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B2 (.DIODE(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A3 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A4 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B2 (.DIODE(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A1 (.DIODE(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A1 (.DIODE(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A1 (.DIODE(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B2 (.DIODE(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A2 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B1 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A1 (.DIODE(\pad_count_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A2 (.DIODE(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A3 (.DIODE(_3006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B1 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A2 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B2 (.DIODE(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B1 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A2 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__B1 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B1 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B2 (.DIODE(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__B1 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A1 (.DIODE(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A1 (.DIODE(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B2 (.DIODE(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A2 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B1 (.DIODE(_3057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A1 (.DIODE(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A2 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A2 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__B2 (.DIODE(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A1 (.DIODE(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A2 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__B2 (.DIODE(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__B2 (.DIODE(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__C (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A1 (.DIODE(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A2 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__S (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(_3024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__B1 (.DIODE(_3027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A2 (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A3 (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__B1 (.DIODE(_3043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A2 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A3 (.DIODE(_3041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__B1 (.DIODE(_3018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A2 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A2 (.DIODE(_3009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__D1 (.DIODE(_3030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(_1441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A3 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__B1 (.DIODE(_3067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B1 (.DIODE(_3015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A2 (.DIODE(_3046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B2 (.DIODE(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B1 (.DIODE(_3068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B2 (.DIODE(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(_3003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(_3035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A1 (.DIODE(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(_3051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(_3013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B1 (.DIODE(_3060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B2 (.DIODE(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A2 (.DIODE(_3007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__B1 (.DIODE(_3054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A3 (.DIODE(_3028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__B1 (.DIODE(_3062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(_3005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B1 (.DIODE(_3025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A2 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A3 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(_3014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B1 (.DIODE(_3055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B2 (.DIODE(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A3 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B1 (.DIODE(_3017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B2 (.DIODE(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A2 (.DIODE(_3012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__B1 (.DIODE(_3022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A1 (.DIODE(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A2 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__B1 (.DIODE(_3362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__S (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A1 (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A2 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A0 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__S (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A1 (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A2 (.DIODE(_1231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A1 (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__A2 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A0 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__S (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A0 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__S (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A0 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__S (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__B1_N (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__B1_N (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__B2 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B2 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A1 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B2 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A1 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A1 (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__B2 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A4 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A (.DIODE(\wbbd_state[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1 (.DIODE(\wbbd_state[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A1 (.DIODE(\wbbd_state[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A2 (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__CLK (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__CLK (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__CLK (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__CLK (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__RESET_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__CLK (.DIODE(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__CLK (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__SET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__RESET_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__SET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__RESET_B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__CLK_N (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__CLK_N (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__CLK_N (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__CLK_N (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__CLK_N (.DIODE(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__RESET_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__RESET_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__CLK (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__RESET_B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7424__SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__SET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__RESET_B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__SET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__SET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__RESET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__CLK (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__SET_B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7509__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7512__SET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7517__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__SET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__7547__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__SET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7573__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__RESET_B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__RESET_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__RESET_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__RESET_B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__CLK (.DIODE(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7646__RESET_B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__A (.DIODE(irq_spi));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__7673__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__1111__A (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_csclk_A (.DIODE(csclk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_mgmt_gpio_in[4]_A  (.DIODE(mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock_A (.DIODE(user_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_2_0__f_mgmt_gpio_in[4]_A  (.DIODE(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_2_1__f_mgmt_gpio_in[4]_A  (.DIODE(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_2_2__f_mgmt_gpio_in[4]_A  (.DIODE(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_2_3__f_mgmt_gpio_in[4]_A  (.DIODE(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_csclk_A (.DIODE(clknet_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_csclk_A (.DIODE(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_csclk_A (.DIODE(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_csclk_A (.DIODE(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_csclk_A (.DIODE(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_csclk_A (.DIODE(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_csclk_A (.DIODE(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_csclk_A (.DIODE(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net2849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net2849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net2849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net2070));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(_3033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(_2663_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(_2647_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net2017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout473_A (.DIODE(net2017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net2696));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(net2696));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout481_A (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout482_A (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout485_A (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout486_A (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout487_A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout488_A (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout491_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout493_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout501_A (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout503_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout510_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout513_A (.DIODE(_0824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout516_A (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(\pad_count_1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout535_A (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout565_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout566_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout568_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout569_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout571_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout575_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout578_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout582_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout586_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout591_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout592_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout593_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout598_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold132_A (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1382_A (.DIODE(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1389_A (.DIODE(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1446_A (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1459_A (.DIODE(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1468_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1469_A (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1480_A (.DIODE(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1490_A (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1499_A (.DIODE(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1515_A (.DIODE(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1529_A (.DIODE(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1541_A (.DIODE(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1552_A (.DIODE(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1563_A (.DIODE(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1566_A (.DIODE(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1570_A (.DIODE(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1580_A (.DIODE(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1586_A (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1589_A (.DIODE(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1602_A (.DIODE(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1613_A (.DIODE(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1619_A (.DIODE(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1621_A (.DIODE(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1627_A (.DIODE(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1643_A (.DIODE(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1647_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1666_A (.DIODE(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1669_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1680_A (.DIODE(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1686_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1699_A (.DIODE(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1702_A (.DIODE(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1705_A (.DIODE(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1715_A (.DIODE(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1718_A (.DIODE(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1733_A (.DIODE(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1739_A (.DIODE(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1747_A (.DIODE(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1750_A (.DIODE(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1755_A (.DIODE(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold175_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1761_A (.DIODE(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1764_A (.DIODE(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1765_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1771_A (.DIODE(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1773_A (.DIODE(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1777_A (.DIODE(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1791_A (.DIODE(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1794_A (.DIODE(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1797_A (.DIODE(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1799_A (.DIODE(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1820_A (.DIODE(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1823_A (.DIODE(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1830_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1840_A (.DIODE(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1842_A (.DIODE(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1845_A (.DIODE(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1856_A (.DIODE(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1864_A (.DIODE(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1871_A (.DIODE(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold187_A (.DIODE(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1883_A (.DIODE(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1894_A (.DIODE(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1908_A (.DIODE(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1911_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1920_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1926_A (.DIODE(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1929_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1935_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1938_A (.DIODE(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1943_A (.DIODE(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1949_A (.DIODE(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1953_A (.DIODE(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold197_A (.DIODE(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1983_A (.DIODE(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1993_A (.DIODE(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2018_A (.DIODE(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2030_A (.DIODE(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2033_A (.DIODE(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2048_A (.DIODE(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2053_A (.DIODE(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2059_A (.DIODE(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2065_A (.DIODE(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2078_A (.DIODE(\clk1_output_dest[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2087_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2090_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2096_A (.DIODE(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2099_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2102_A (.DIODE(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold213_A (.DIODE(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2149_A (.DIODE(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2167_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2170_A (.DIODE(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2176_A (.DIODE(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2180_A (.DIODE(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2185_A (.DIODE(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2193_A (.DIODE(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2195_A (.DIODE(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2198_A (.DIODE(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2202_A (.DIODE(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2205_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2208_A (.DIODE(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2211_A (.DIODE(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2216_A (.DIODE(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2225_A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2236_A (.DIODE(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2256_A (.DIODE(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2258_A (.DIODE(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2268_A (.DIODE(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2281_A (.DIODE(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2286_A (.DIODE(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2288_A (.DIODE(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2298_A (.DIODE(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2301_A (.DIODE(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2312_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2316_A (.DIODE(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2323_A (.DIODE(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2331_A (.DIODE(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2333_A (.DIODE(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2350_A (.DIODE(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2353_A (.DIODE(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2357_A (.DIODE(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2359_A (.DIODE(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2364_A (.DIODE(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2367_A (.DIODE(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2371_A (.DIODE(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2374_A (.DIODE(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2403_A (.DIODE(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2406_A (.DIODE(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2412_A (.DIODE(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2416_A (.DIODE(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2418_A (.DIODE(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2420_A (.DIODE(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2428_A (.DIODE(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2431_A (.DIODE(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2436_A (.DIODE(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2441_A (.DIODE(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2446_A (.DIODE(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2450_A (.DIODE(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2452_A (.DIODE(serial_bb_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2457_A (.DIODE(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2462_A (.DIODE(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2467_A (.DIODE(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2469_A (.DIODE(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2473_A (.DIODE(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2475_A (.DIODE(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2487_A (.DIODE(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2489_A (.DIODE(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2504_A (.DIODE(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2517_A (.DIODE(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2519_A (.DIODE(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2521_A (.DIODE(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2523_A (.DIODE(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2533_A (.DIODE(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2537_A (.DIODE(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2539_A (.DIODE(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2553_A (.DIODE(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2591_A (.DIODE(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2598_A (.DIODE(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2603_A (.DIODE(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2608_A (.DIODE(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2654_A (.DIODE(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2658_A (.DIODE(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2674_A (.DIODE(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2695_A (.DIODE(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2697_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2720_A (.DIODE(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2734_A (.DIODE(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2737_A (.DIODE(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2741_A (.DIODE(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2751_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2758_A (.DIODE(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2770_A (.DIODE(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2772_A (.DIODE(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2777_A (.DIODE(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2792_A (.DIODE(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2798_A (.DIODE(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2803_A (.DIODE(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2811_A (.DIODE(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold281_A (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2821_A (.DIODE(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2829_A (.DIODE(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold282_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2832_A (.DIODE(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2841_A (.DIODE(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold284_A (.DIODE(net2388));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2854_A (.DIODE(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2866_A (.DIODE(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2884_A (.DIODE(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2887_A (.DIODE(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2889_A (.DIODE(\clk2_output_dest[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2892_A (.DIODE(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2902_A (.DIODE(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2907_A (.DIODE(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2909_A (.DIODE(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2931_A (.DIODE(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2933_A (.DIODE(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2939_A (.DIODE(irq_spi));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2949_A (.DIODE(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2955_A (.DIODE(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2957_A (.DIODE(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2960_A (.DIODE(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2964_A (.DIODE(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2978_A (.DIODE(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2987_A (.DIODE(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2991_A (.DIODE(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2996_A (.DIODE(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2998_A (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3003_A (.DIODE(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3006_A (.DIODE(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3023_A (.DIODE(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3025_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3040_A (.DIODE(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3050_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3053_A (.DIODE(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3055_A (.DIODE(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3082_A (.DIODE(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3093_A (.DIODE(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3148_A (.DIODE(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3150_A (.DIODE(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3155_A (.DIODE(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3157_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3160_A (.DIODE(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3164_A (.DIODE(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3172_A (.DIODE(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3187_A (.DIODE(_3366_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3210_A (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3247_A (.DIODE(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3249_A (.DIODE(\hkspi.SDO ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3250_A (.DIODE(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3252_A (.DIODE(\wbbd_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3259_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3264_A (.DIODE(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3279_A (.DIODE(\hkspi.wrstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3281_A (.DIODE(\hkspi.rdstb ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3282_A (.DIODE(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3285_A (.DIODE(hkspi_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold37_A (.DIODE(_2631_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold48_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold56_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold586_A (.DIODE(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold72_A (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold76_A (.DIODE(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(wb_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(wb_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(wb_adr_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(wb_adr_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(wb_adr_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(wb_adr_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(wb_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(wb_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(wb_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(wb_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(mask_rev_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(wb_adr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(wb_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(wb_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(wb_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(wb_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(wb_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(wb_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(wb_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(wb_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(wb_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(mask_rev_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(wb_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(wb_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(wb_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(wb_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(wb_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(wb_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(wb_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(wb_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(wb_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(wb_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(mask_rev_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(wb_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(wb_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(wb_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(wb_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(wb_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(wb_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(wb_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(wb_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(wb_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(wb_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(mask_rev_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(wb_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(wb_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(wb_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(wb_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(wb_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(wb_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(wb_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(wb_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(wb_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(wb_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(mask_rev_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(wb_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(wb_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(wb_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(wb_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(wb_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(wb_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(wb_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(wb_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(wb_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(wb_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(mask_rev_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(wb_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(wb_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(wb_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(wb_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(wb_rstn_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(wb_sel_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(wb_sel_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(wb_sel_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(wb_sel_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(wb_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(mask_rev_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(wb_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(mask_rev_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(mask_rev_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(mask_rev_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(debug_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(mask_rev_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(mask_rev_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(mask_rev_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(mask_rev_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(mask_rev_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(mask_rev_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(mask_rev_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(mask_rev_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(mask_rev_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(mask_rev_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(debug_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(mask_rev_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(mask_rev_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(mask_rev_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(mask_rev_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(mask_rev_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(mask_rev_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(mgmt_gpio_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(mgmt_gpio_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(mgmt_gpio_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(mgmt_gpio_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(debug_out));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(mgmt_gpio_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(mgmt_gpio_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(mgmt_gpio_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(mgmt_gpio_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(mgmt_gpio_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(mgmt_gpio_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(mgmt_gpio_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(mgmt_gpio_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(mgmt_gpio_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(mgmt_gpio_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(mask_rev_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(mgmt_gpio_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(mgmt_gpio_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(mgmt_gpio_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(mgmt_gpio_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(mgmt_gpio_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(mgmt_gpio_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(mgmt_gpio_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(mgmt_gpio_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(mgmt_gpio_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(mgmt_gpio_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(mask_rev_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(mgmt_gpio_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(mgmt_gpio_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(mgmt_gpio_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(mgmt_gpio_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(mgmt_gpio_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(mgmt_gpio_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(mgmt_gpio_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(mgmt_gpio_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(mgmt_gpio_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(mgmt_gpio_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(mask_rev_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(mgmt_gpio_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(mgmt_gpio_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(mgmt_gpio_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(pad_flash_io0_di));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(pad_flash_io1_di));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(porb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(qspi_enabled));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(ser_tx));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(spi_csb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(spi_enabled));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(mask_rev_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(spi_sck));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(spi_sdo));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(spi_sdoenb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(spimemio_flash_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(spimemio_flash_csb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(spimemio_flash_io0_do));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(spimemio_flash_io0_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(spimemio_flash_io1_do));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(spimemio_flash_io1_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(spimemio_flash_io2_do));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(mask_rev_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(spimemio_flash_io2_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(spimemio_flash_io3_do));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(spimemio_flash_io3_oeb));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(trap));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(uart_enabled));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(usr1_vcc_pwrgood));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(usr1_vdd_pwrgood));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(usr2_vcc_pwrgood));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(usr2_vdd_pwrgood));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(wb_adr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(mask_rev_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap400_A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap557_A (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_output234_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_output237_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_output243_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output273_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output311_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire365_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire507_A (.DIODE(net508));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3399_ (.A(\hkspi.addr[0] ),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _3400_ (.A(net3872),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _3401_ (.A(\hkspi.fixed[0] ),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_4 _3402_ (.A(\hkspi.state[0] ),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _3403_ (.A(net3860),
    .Y(_0820_));
 sky130_fd_sc_hd__inv_8 _3404_ (.A(net111),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(\gpio_configure[3][3] ),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _3406_ (.A(\xfer_count[1] ),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _3407_ (.A(\xfer_state[3] ),
    .Y(_0823_));
 sky130_fd_sc_hd__clkinv_4 _3408_ (.A(net527),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_2 _3409_ (.A(serial_xfer),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_2 _3410__1 (.A(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .Y(net623));
 sky130_fd_sc_hd__inv_2 _3411_ (.A(\gpio_configure[34][3] ),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _3412_ (.A(\gpio_configure[33][3] ),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _3413_ (.A(\gpio_configure[32][3] ),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _3414_ (.A(\gpio_configure[31][3] ),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _3415_ (.A(\gpio_configure[30][3] ),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _3416_ (.A(\gpio_configure[29][3] ),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(\gpio_configure[28][3] ),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _3418_ (.A(\gpio_configure[27][3] ),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _3419_ (.A(\gpio_configure[26][3] ),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(\gpio_configure[25][3] ),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _3421_ (.A(\gpio_configure[24][3] ),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(\gpio_configure[23][3] ),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _3423_ (.A(\gpio_configure[22][3] ),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _3424_ (.A(\gpio_configure[21][3] ),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _3425_ (.A(\gpio_configure[20][3] ),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _3426_ (.A(\gpio_configure[19][3] ),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(\gpio_configure[18][3] ),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _3428_ (.A(\gpio_configure[17][3] ),
    .Y(net183));
 sky130_fd_sc_hd__clkinv_2 _3429_ (.A(\gpio_configure[16][3] ),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _3430_ (.A(\gpio_configure[15][3] ),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _3431_ (.A(\gpio_configure[14][3] ),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _3432_ (.A(\gpio_configure[13][3] ),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _3433_ (.A(\gpio_configure[12][3] ),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _3434_ (.A(\gpio_configure[11][3] ),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(\gpio_configure[10][3] ),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _3436_ (.A(\gpio_configure[9][3] ),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _3437_ (.A(\gpio_configure[8][3] ),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _3438_ (.A(\gpio_configure[7][3] ),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _3439_ (.A(\gpio_configure[6][3] ),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _3440_ (.A(\gpio_configure[5][3] ),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _3441_ (.A(\gpio_configure[4][3] ),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _3442_ (.A(\gpio_configure[2][3] ),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _3443__2 (.A(clknet_1_0__leaf_wbbd_sck),
    .Y(net624));
 sky130_fd_sc_hd__inv_2 _3444_ (.A(net516),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_16 _3445_ (.A(net614),
    .Y(_0828_));
 sky130_fd_sc_hd__nor3_4 _3446_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _3447_ (.A(\hkspi.addr[4] ),
    .B(net525),
    .Y(_0830_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(net2449),
    .A1(\hkspi.addr[4] ),
    .S(net525),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(net2450),
    .A1(net903),
    .S(net524),
    .X(_0832_));
 sky130_fd_sc_hd__and2b_1 _3450_ (.A_N(net525),
    .B(net2846),
    .X(_0833_));
 sky130_fd_sc_hd__a21oi_1 _3451_ (.A1(net675),
    .A2(net525),
    .B1(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a21o_1 _3452_ (.A1(net2449),
    .A2(net525),
    .B1(net675),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(_0835_),
    .A1(net1152),
    .S(net524),
    .X(_0836_));
 sky130_fd_sc_hd__o21ba_1 _3454_ (.A1(net524),
    .A2(net676),
    .B1_N(net1153),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(\hkspi.addr[4] ),
    .A1(net1020),
    .S(net525),
    .X(_0838_));
 sky130_fd_sc_hd__and2b_1 _3456_ (.A_N(net524),
    .B(net1021),
    .X(_0839_));
 sky130_fd_sc_hd__a21o_1 _3457_ (.A1(net524),
    .A2(net2112),
    .B1(net1022),
    .X(_0840_));
 sky130_fd_sc_hd__a21oi_4 _3458_ (.A1(net524),
    .A2(net2112),
    .B1(_0839_),
    .Y(_0841_));
 sky130_fd_sc_hd__and3_4 _3459_ (.A(net2452),
    .B(net1154),
    .C(net1023),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_2 _3460_ (.A0(net1020),
    .A1(\hkspi.addr[2] ),
    .S(net525),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(_0843_),
    .A1(net2088),
    .S(net524),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\hkspi.addr[2] ),
    .A1(\hkspi.addr[1] ),
    .S(net525),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(_0845_),
    .A1(net2296),
    .S(net524),
    .X(_0846_));
 sky130_fd_sc_hd__and2b_1 _3464_ (.A_N(net658),
    .B(net2090),
    .X(_0847_));
 sky130_fd_sc_hd__nand2b_2 _3465_ (.A_N(net58),
    .B(net525),
    .Y(_0848_));
 sky130_fd_sc_hd__o21ba_1 _3466_ (.A1(net777),
    .A2(net525),
    .B1_N(net524),
    .X(_0849_));
 sky130_fd_sc_hd__a22oi_1 _3467_ (.A1(net524),
    .A2(net2067),
    .B1(net778),
    .B2(_0848_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _3468_ (.A1(net2936),
    .A2(net2067),
    .B1(net778),
    .B2(_0848_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\hkspi.addr[1] ),
    .A1(\hkspi.addr[0] ),
    .S(net525),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_4 _3470_ (.A0(_0852_),
    .A1(net2207),
    .S(net524),
    .X(_0853_));
 sky130_fd_sc_hd__and2_4 _3471_ (.A(net2069),
    .B(net644),
    .X(_0854_));
 sky130_fd_sc_hd__and3_2 _3472_ (.A(net420),
    .B(net2069),
    .C(net2209),
    .X(_0855_));
 sky130_fd_sc_hd__and3_1 _3473_ (.A(net391),
    .B(net420),
    .C(net419),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_1 _3474_ (.A(net2937),
    .B(net2209),
    .Y(_0857_));
 sky130_fd_sc_hd__o21a_1 _3475_ (.A1(net524),
    .A2(net676),
    .B1(_0836_),
    .X(_0858_));
 sky130_fd_sc_hd__nand2b_1 _3476_ (.A_N(net904),
    .B(net677),
    .Y(_0859_));
 sky130_fd_sc_hd__nor2_1 _3477_ (.A(net1023),
    .B(net678),
    .Y(_0860_));
 sky130_fd_sc_hd__and3_4 _3478_ (.A(net420),
    .B(net418),
    .C(net358),
    .X(_0861_));
 sky130_fd_sc_hd__a32o_4 _3479_ (.A1(\gpio_configure[14][7] ),
    .A2(net392),
    .A3(net389),
    .B1(_0861_),
    .B2(\gpio_configure[21][7] ),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _3480_ (.A(net2090),
    .B(net2298),
    .X(_0863_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(net417),
    .B(net416),
    .Y(_0864_));
 sky130_fd_sc_hd__and3_4 _3482_ (.A(net390),
    .B(net417),
    .C(net415),
    .X(_0865_));
 sky130_fd_sc_hd__and2b_1 _3483_ (.A_N(net2090),
    .B(net2298),
    .X(_0866_));
 sky130_fd_sc_hd__and3_4 _3484_ (.A(net2069),
    .B(net2209),
    .C(net414),
    .X(_0867_));
 sky130_fd_sc_hd__and3b_4 _3485_ (.A_N(net904),
    .B(net2848),
    .C(net755),
    .X(_0868_));
 sky130_fd_sc_hd__and3_4 _3486_ (.A(net419),
    .B(net413),
    .C(net385),
    .X(_0869_));
 sky130_fd_sc_hd__a221o_2 _3487_ (.A1(\gpio_configure[15][7] ),
    .A2(_0865_),
    .B1(_0869_),
    .B2(net10),
    .C1(_0862_),
    .X(_0870_));
 sky130_fd_sc_hd__and3_4 _3488_ (.A(net417),
    .B(net413),
    .C(net385),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_2 _3489_ (.A(net2069),
    .B(net2209),
    .Y(_0872_));
 sky130_fd_sc_hd__and3_4 _3490_ (.A(net413),
    .B(net385),
    .C(net410),
    .X(_0873_));
 sky130_fd_sc_hd__a221o_4 _3491_ (.A1(net28),
    .A2(_0871_),
    .B1(_0873_),
    .B2(net19),
    .C1(_0870_),
    .X(_0874_));
 sky130_fd_sc_hd__and3_4 _3492_ (.A(net2090),
    .B(net2298),
    .C(net419),
    .X(_0875_));
 sky130_fd_sc_hd__and3_2 _3493_ (.A(net390),
    .B(net419),
    .C(net415),
    .X(_0876_));
 sky130_fd_sc_hd__and3_4 _3494_ (.A(net419),
    .B(net359),
    .C(net416),
    .X(_0877_));
 sky130_fd_sc_hd__a32o_1 _3495_ (.A1(\gpio_configure[16][7] ),
    .A2(net391),
    .A3(net384),
    .B1(_0877_),
    .B2(\gpio_configure[24][7] ),
    .X(_0878_));
 sky130_fd_sc_hd__nor2_8 _3496_ (.A(net2113),
    .B(net678),
    .Y(_0879_));
 sky130_fd_sc_hd__and3_4 _3497_ (.A(net417),
    .B(net413),
    .C(net355),
    .X(_0880_));
 sky130_fd_sc_hd__and3_4 _3498_ (.A(net391),
    .B(net419),
    .C(net414),
    .X(_0881_));
 sky130_fd_sc_hd__a221o_1 _3499_ (.A1(\gpio_configure[27][7] ),
    .A2(_0880_),
    .B1(_0881_),
    .B2(\gpio_configure[12][7] ),
    .C1(_0878_),
    .X(_0882_));
 sky130_fd_sc_hd__and3_4 _3500_ (.A(net755),
    .B(net677),
    .C(net2451),
    .X(_0883_));
 sky130_fd_sc_hd__and3_4 _3501_ (.A(net420),
    .B(net417),
    .C(net380),
    .X(_0884_));
 sky130_fd_sc_hd__and2_4 _3502_ (.A(net2209),
    .B(net779),
    .X(_0885_));
 sky130_fd_sc_hd__and3_4 _3503_ (.A(net413),
    .B(net385),
    .C(net409),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_4 _3504_ (.A(net2090),
    .B(net658),
    .Y(_0887_));
 sky130_fd_sc_hd__nor4_1 _3505_ (.A(net779),
    .B(net2209),
    .C(net2090),
    .D(net2298),
    .Y(_0888_));
 sky130_fd_sc_hd__and3_4 _3506_ (.A(net391),
    .B(net418),
    .C(net407),
    .X(_0889_));
 sky130_fd_sc_hd__and3_4 _3507_ (.A(net2069),
    .B(net2208),
    .C(net408),
    .X(_0890_));
 sky130_fd_sc_hd__and3_4 _3508_ (.A(net419),
    .B(net380),
    .C(net407),
    .X(_0891_));
 sky130_fd_sc_hd__a32o_1 _3509_ (.A1(\gpio_configure[9][7] ),
    .A2(_0842_),
    .A3(net403),
    .B1(_0891_),
    .B2(\gpio_configure[34][7] ),
    .X(_0892_));
 sky130_fd_sc_hd__a221o_1 _3510_ (.A1(\gpio_configure[37][7] ),
    .A2(_0884_),
    .B1(_0886_),
    .B2(net33),
    .C1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__and3_2 _3511_ (.A(net755),
    .B(net1154),
    .C(net2452),
    .X(_0894_));
 sky130_fd_sc_hd__and3_4 _3512_ (.A(net417),
    .B(net413),
    .C(net377),
    .X(_0895_));
 sky130_fd_sc_hd__a32o_1 _3513_ (.A1(\gpio_configure[36][7] ),
    .A2(net387),
    .A3(net382),
    .B1(_0895_),
    .B2(\gpio_configure[3][7] ),
    .X(_0896_));
 sky130_fd_sc_hd__and3_2 _3514_ (.A(net416),
    .B(net779),
    .C(net2209),
    .X(_0897_));
 sky130_fd_sc_hd__and3_4 _3515_ (.A(net415),
    .B(net385),
    .C(net409),
    .X(_0898_));
 sky130_fd_sc_hd__and3_4 _3516_ (.A(net418),
    .B(net414),
    .C(net380),
    .X(_0899_));
 sky130_fd_sc_hd__a221o_1 _3517_ (.A1(net284),
    .A2(_0898_),
    .B1(_0899_),
    .B2(\gpio_configure[35][7] ),
    .C1(_0896_),
    .X(_0900_));
 sky130_fd_sc_hd__and3_4 _3518_ (.A(net392),
    .B(net418),
    .C(net414),
    .X(_0901_));
 sky130_fd_sc_hd__and3_2 _3519_ (.A(net418),
    .B(_0883_),
    .C(net408),
    .X(_0902_));
 sky130_fd_sc_hd__and3_4 _3520_ (.A(net419),
    .B(net357),
    .C(net413),
    .X(_0903_));
 sky130_fd_sc_hd__and3_4 _3521_ (.A(net419),
    .B(net413),
    .C(net377),
    .X(_0904_));
 sky130_fd_sc_hd__a32o_1 _3522_ (.A1(\gpio_configure[20][7] ),
    .A2(net359),
    .A3(net387),
    .B1(_0904_),
    .B2(\gpio_configure[4][7] ),
    .X(_0905_));
 sky130_fd_sc_hd__a221o_1 _3523_ (.A1(\gpio_configure[11][7] ),
    .A2(_0901_),
    .B1(_0902_),
    .B2(\gpio_configure[33][7] ),
    .C1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nor4_2 _3524_ (.A(_0882_),
    .B(_0893_),
    .C(_0900_),
    .D(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__and3_4 _3525_ (.A(net418),
    .B(net359),
    .C(net414),
    .X(_0908_));
 sky130_fd_sc_hd__and3_4 _3526_ (.A(_0854_),
    .B(net414),
    .C(net356),
    .X(_0909_));
 sky130_fd_sc_hd__and3_2 _3527_ (.A(net419),
    .B(net415),
    .C(net385),
    .X(_0910_));
 sky130_fd_sc_hd__a32o_4 _3528_ (.A1(\gpio_configure[28][7] ),
    .A2(net387),
    .A3(net355),
    .B1(_0910_),
    .B2(net275),
    .X(_0911_));
 sky130_fd_sc_hd__and3_4 _3529_ (.A(net418),
    .B(net416),
    .C(net356),
    .X(_0912_));
 sky130_fd_sc_hd__and3_4 _3530_ (.A(net660),
    .B(net419),
    .C(net357),
    .X(_0913_));
 sky130_fd_sc_hd__and3_4 _3531_ (.A(net417),
    .B(net415),
    .C(net377),
    .X(_0914_));
 sky130_fd_sc_hd__and3_1 _3532_ (.A(net420),
    .B(_0854_),
    .C(net382),
    .X(_0915_));
 sky130_fd_sc_hd__a32o_1 _3533_ (.A1(net60),
    .A2(net388),
    .A3(net382),
    .B1(_0914_),
    .B2(\gpio_configure[7][7] ),
    .X(_0916_));
 sky130_fd_sc_hd__a221o_1 _3534_ (.A1(\gpio_configure[31][7] ),
    .A2(_0912_),
    .B1(_0913_),
    .B2(\gpio_configure[22][7] ),
    .C1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__and3_4 _3535_ (.A(net418),
    .B(net356),
    .C(net407),
    .X(_0918_));
 sky130_fd_sc_hd__a32o_1 _3536_ (.A1(\gpio_configure[26][7] ),
    .A2(_0879_),
    .A3(_0890_),
    .B1(_0918_),
    .B2(\gpio_configure[25][7] ),
    .X(_0919_));
 sky130_fd_sc_hd__and3_4 _3537_ (.A(_0854_),
    .B(net357),
    .C(net408),
    .X(_0920_));
 sky130_fd_sc_hd__and3_4 _3538_ (.A(net420),
    .B(net2070),
    .C(net356),
    .X(_0921_));
 sky130_fd_sc_hd__a221o_1 _3539_ (.A1(\gpio_configure[18][7] ),
    .A2(_0920_),
    .B1(_0921_),
    .B2(\gpio_configure[30][7] ),
    .C1(_0919_),
    .X(_0922_));
 sky130_fd_sc_hd__a2111o_1 _3540_ (.A1(\gpio_configure[19][7] ),
    .A2(_0908_),
    .B1(_0911_),
    .C1(_0917_),
    .D1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _3541_ (.A(net416),
    .B(net412),
    .Y(_0924_));
 sky130_fd_sc_hd__and3_4 _3542_ (.A(net415),
    .B(net385),
    .C(net410),
    .X(_0925_));
 sky130_fd_sc_hd__and3_4 _3543_ (.A(net417),
    .B(net2092),
    .C(net377),
    .X(_0926_));
 sky130_fd_sc_hd__and3_4 _3544_ (.A(net417),
    .B(net357),
    .C(net407),
    .X(_0927_));
 sky130_fd_sc_hd__and3_4 _3545_ (.A(net419),
    .B(net415),
    .C(net377),
    .X(_0928_));
 sky130_fd_sc_hd__a32o_1 _3546_ (.A1(\gpio_configure[17][7] ),
    .A2(net357),
    .A3(net403),
    .B1(_0928_),
    .B2(\gpio_configure[8][7] ),
    .X(_0929_));
 sky130_fd_sc_hd__a221o_4 _3547_ (.A1(net292),
    .A2(_0925_),
    .B1(_0926_),
    .B2(\gpio_configure[1][7] ),
    .C1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__and3_2 _3548_ (.A(net420),
    .B(net779),
    .C(net2209),
    .X(_0931_));
 sky130_fd_sc_hd__and3_4 _3549_ (.A(net420),
    .B(net380),
    .C(net409),
    .X(_0932_));
 sky130_fd_sc_hd__and3_4 _3550_ (.A(net420),
    .B(net418),
    .C(net356),
    .X(_0933_));
 sky130_fd_sc_hd__a32o_4 _3551_ (.A1(net51),
    .A2(net381),
    .A3(net374),
    .B1(_0933_),
    .B2(\gpio_configure[29][7] ),
    .X(_0934_));
 sky130_fd_sc_hd__and3_4 _3552_ (.A(net415),
    .B(net410),
    .C(net756),
    .X(_0935_));
 sky130_fd_sc_hd__and3_4 _3553_ (.A(net418),
    .B(net416),
    .C(net380),
    .X(_0936_));
 sky130_fd_sc_hd__a221o_1 _3554_ (.A1(net70),
    .A2(_0935_),
    .B1(_0936_),
    .B2(net42),
    .C1(_0934_),
    .X(_0937_));
 sky130_fd_sc_hd__and3_4 _3555_ (.A(net392),
    .B(net420),
    .C(net418),
    .X(_0938_));
 sky130_fd_sc_hd__and3_4 _3556_ (.A(net660),
    .B(net417),
    .C(net377),
    .X(_0939_));
 sky130_fd_sc_hd__and3b_2 _3557_ (.A_N(net2452),
    .B(net1154),
    .C(net1023),
    .X(_0940_));
 sky130_fd_sc_hd__and3_4 _3558_ (.A(net419),
    .B(net415),
    .C(net372),
    .X(_0941_));
 sky130_fd_sc_hd__a32o_2 _3559_ (.A1(\gpio_configure[32][7] ),
    .A2(net383),
    .A3(net355),
    .B1(_0941_),
    .B2(\gpio_configure[0][7] ),
    .X(_0942_));
 sky130_fd_sc_hd__a221o_1 _3560_ (.A1(\gpio_configure[13][7] ),
    .A2(_0938_),
    .B1(_0939_),
    .B2(\gpio_configure[5][7] ),
    .C1(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__and3_4 _3561_ (.A(net660),
    .B(net419),
    .C(net377),
    .X(_0944_));
 sky130_fd_sc_hd__and3_2 _3562_ (.A(net419),
    .B(net407),
    .C(net377),
    .X(_0945_));
 sky130_fd_sc_hd__and3_1 _3563_ (.A(\gpio_configure[2][7] ),
    .B(_0890_),
    .C(net379),
    .X(_0946_));
 sky130_fd_sc_hd__and3_4 _3564_ (.A(_0842_),
    .B(net419),
    .C(net407),
    .X(_0947_));
 sky130_fd_sc_hd__and3_4 _3565_ (.A(net418),
    .B(net359),
    .C(net415),
    .X(_0948_));
 sky130_fd_sc_hd__a32o_1 _3566_ (.A1(\gpio_configure[10][7] ),
    .A2(net390),
    .A3(_0890_),
    .B1(_0948_),
    .B2(\gpio_configure[23][7] ),
    .X(_0949_));
 sky130_fd_sc_hd__a2111o_1 _3567_ (.A1(\gpio_configure[6][7] ),
    .A2(_0944_),
    .B1(_0946_),
    .C1(_0949_),
    .D1(_0943_),
    .X(_0950_));
 sky130_fd_sc_hd__nor4_2 _3568_ (.A(_0923_),
    .B(_0930_),
    .C(_0937_),
    .D(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__and3_4 _3569_ (.A(net2070),
    .B(net355),
    .C(net408),
    .X(_0952_));
 sky130_fd_sc_hd__nand3b_4 _3570_ (.A_N(_0874_),
    .B(_0907_),
    .C(_0951_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_8 _3571_ (.A(\hkspi.readmode ),
    .B(\hkspi.state[2] ),
    .Y(_0954_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(net3798),
    .A1(_0953_),
    .S(net509),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _3573_ (.A0(_0955_),
    .A1(net3873),
    .S(_0954_),
    .X(_0391_));
 sky130_fd_sc_hd__a32o_4 _3574_ (.A1(\gpio_configure[36][6] ),
    .A2(_0867_),
    .A3(net382),
    .B1(_0899_),
    .B2(\gpio_configure[35][6] ),
    .X(_0956_));
 sky130_fd_sc_hd__a221o_4 _3575_ (.A1(net27),
    .A2(_0871_),
    .B1(_0873_),
    .B2(net18),
    .C1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__and3_4 _3576_ (.A(net408),
    .B(net779),
    .C(net2209),
    .X(_0958_));
 sky130_fd_sc_hd__and3_1 _3577_ (.A(net409),
    .B(net2092),
    .C(net372),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_8 _3578_ (.A0(\serial_data_staging_2[12] ),
    .A1(serial_bb_data_2),
    .S(serial_bb_enable),
    .X(net303));
 sky130_fd_sc_hd__a32o_1 _3579_ (.A1(net372),
    .A2(net370),
    .A3(net303),
    .B1(_0935_),
    .B2(net69),
    .X(_0960_));
 sky130_fd_sc_hd__a221o_1 _3580_ (.A1(\gpio_configure[27][6] ),
    .A2(_0880_),
    .B1(_0925_),
    .B2(net291),
    .C1(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a32o_1 _3581_ (.A1(\gpio_configure[26][6] ),
    .A2(net355),
    .A3(_0890_),
    .B1(_0932_),
    .B2(net50),
    .X(_0962_));
 sky130_fd_sc_hd__a221o_1 _3582_ (.A1(\gpio_configure[12][6] ),
    .A2(_0881_),
    .B1(_0947_),
    .B2(\gpio_configure[10][6] ),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a32o_4 _3583_ (.A1(\gpio_configure[30][6] ),
    .A2(net388),
    .A3(net356),
    .B1(_0936_),
    .B2(net41),
    .X(_0964_));
 sky130_fd_sc_hd__a221o_1 _3584_ (.A1(\gpio_configure[15][6] ),
    .A2(_0865_),
    .B1(_0948_),
    .B2(\gpio_configure[23][6] ),
    .C1(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__a32o_1 _3585_ (.A1(\gpio_configure[0][6] ),
    .A2(net384),
    .A3(net373),
    .B1(_0913_),
    .B2(\gpio_configure[22][6] ),
    .X(_0966_));
 sky130_fd_sc_hd__a221o_1 _3586_ (.A1(\gpio_configure[9][6] ),
    .A2(_0889_),
    .B1(_0901_),
    .B2(\gpio_configure[11][6] ),
    .C1(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__nor4_2 _3587_ (.A(_0961_),
    .B(_0963_),
    .C(_0965_),
    .D(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__a32o_1 _3588_ (.A1(\gpio_configure[32][6] ),
    .A2(net384),
    .A3(net355),
    .B1(_0927_),
    .B2(\gpio_configure[17][6] ),
    .X(_0969_));
 sky130_fd_sc_hd__a221o_1 _3589_ (.A1(\gpio_configure[37][6] ),
    .A2(_0884_),
    .B1(_0938_),
    .B2(\gpio_configure[13][6] ),
    .C1(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__and3_1 _3590_ (.A(\gpio_configure[24][6] ),
    .B(net359),
    .C(net384),
    .X(_0971_));
 sky130_fd_sc_hd__a32o_1 _3591_ (.A1(net59),
    .A2(net389),
    .A3(_0883_),
    .B1(_0939_),
    .B2(\gpio_configure[5][6] ),
    .X(_0972_));
 sky130_fd_sc_hd__a2111o_1 _3592_ (.A1(\gpio_configure[19][6] ),
    .A2(_0908_),
    .B1(_0971_),
    .C1(_0972_),
    .D1(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__a32o_1 _3593_ (.A1(\gpio_configure[16][6] ),
    .A2(net390),
    .A3(net384),
    .B1(_0944_),
    .B2(\gpio_configure[6][6] ),
    .X(_0974_));
 sky130_fd_sc_hd__a32o_1 _3594_ (.A1(\gpio_configure[14][6] ),
    .A2(net390),
    .A3(net389),
    .B1(_0902_),
    .B2(\gpio_configure[33][6] ),
    .X(_0975_));
 sky130_fd_sc_hd__a221o_1 _3595_ (.A1(\gpio_configure[21][6] ),
    .A2(_0861_),
    .B1(_0912_),
    .B2(\gpio_configure[31][6] ),
    .C1(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__a2111o_1 _3596_ (.A1(\gpio_configure[1][6] ),
    .A2(_0926_),
    .B1(_0973_),
    .C1(_0974_),
    .D1(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a32o_4 _3597_ (.A1(\gpio_configure[28][6] ),
    .A2(net387),
    .A3(net356),
    .B1(_0918_),
    .B2(\gpio_configure[25][6] ),
    .X(_0978_));
 sky130_fd_sc_hd__and3_1 _3598_ (.A(net419),
    .B(net385),
    .C(net407),
    .X(_0979_));
 sky130_fd_sc_hd__a32o_1 _3599_ (.A1(\gpio_configure[4][6] ),
    .A2(net387),
    .A3(net377),
    .B1(_0886_),
    .B2(net32),
    .X(_0980_));
 sky130_fd_sc_hd__a221o_1 _3600_ (.A1(\gpio_configure[7][6] ),
    .A2(_0914_),
    .B1(_0928_),
    .B2(\gpio_configure[8][6] ),
    .C1(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__a2111o_1 _3601_ (.A1(net274),
    .A2(_0910_),
    .B1(_0978_),
    .C1(_0979_),
    .D1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__a32o_4 _3602_ (.A1(net283),
    .A2(net385),
    .A3(net376),
    .B1(_0895_),
    .B2(\gpio_configure[3][6] ),
    .X(_0983_));
 sky130_fd_sc_hd__a221o_1 _3603_ (.A1(\gpio_configure[20][6] ),
    .A2(_0903_),
    .B1(_0933_),
    .B2(\gpio_configure[29][6] ),
    .C1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a32o_1 _3604_ (.A1(\gpio_configure[18][6] ),
    .A2(net357),
    .A3(_0890_),
    .B1(_0945_),
    .B2(\gpio_configure[2][6] ),
    .X(_0985_));
 sky130_fd_sc_hd__a221o_1 _3605_ (.A1(net9),
    .A2(_0869_),
    .B1(_0891_),
    .B2(\gpio_configure[34][6] ),
    .C1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__nor4_2 _3606_ (.A(_0977_),
    .B(_0982_),
    .C(_0984_),
    .D(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand3b_4 _3607_ (.A_N(_0957_),
    .B(_0968_),
    .C(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\hkspi.ldata[5] ),
    .A1(_0988_),
    .S(net509),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _3609_ (.A0(_0989_),
    .A1(net3798),
    .S(_0954_),
    .X(_0390_));
 sky130_fd_sc_hd__a32o_2 _3610_ (.A1(\gpio_configure[9][5] ),
    .A2(net390),
    .A3(net403),
    .B1(_0877_),
    .B2(\gpio_configure[24][5] ),
    .X(_0990_));
 sky130_fd_sc_hd__a221o_4 _3611_ (.A1(net25),
    .A2(_0871_),
    .B1(_0873_),
    .B2(net17),
    .C1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__a32o_1 _3612_ (.A1(net282),
    .A2(_0868_),
    .A3(net376),
    .B1(_0908_),
    .B2(\gpio_configure[19][5] ),
    .X(_0992_));
 sky130_fd_sc_hd__a221o_1 _3613_ (.A1(\gpio_configure[34][5] ),
    .A2(_0891_),
    .B1(_0933_),
    .B2(\gpio_configure[29][5] ),
    .C1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a32o_4 _3614_ (.A1(\gpio_configure[33][5] ),
    .A2(net382),
    .A3(net403),
    .B1(_0899_),
    .B2(\gpio_configure[35][5] ),
    .X(_0994_));
 sky130_fd_sc_hd__a221o_1 _3615_ (.A1(\gpio_configure[1][5] ),
    .A2(_0926_),
    .B1(_0932_),
    .B2(net49),
    .C1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__and3_1 _3616_ (.A(\gpio_configure[8][5] ),
    .B(net383),
    .C(net377),
    .X(_0996_));
 sky130_fd_sc_hd__and3_4 _3617_ (.A(net412),
    .B(net407),
    .C(net373),
    .X(_0997_));
 sky130_fd_sc_hd__a32o_1 _3618_ (.A1(\gpio_configure[6][5] ),
    .A2(net389),
    .A3(net377),
    .B1(_0904_),
    .B2(\gpio_configure[4][5] ),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_8 _3619_ (.A0(\serial_data_staging_1[12] ),
    .A1(serial_bb_data_1),
    .S(serial_bb_enable),
    .X(net302));
 sky130_fd_sc_hd__a32o_1 _3620_ (.A1(net372),
    .A2(net370),
    .A3(net302),
    .B1(_0941_),
    .B2(\gpio_configure[0][5] ),
    .X(_0999_));
 sky130_fd_sc_hd__a221o_1 _3621_ (.A1(\gpio_configure[15][5] ),
    .A2(_0865_),
    .B1(_0925_),
    .B2(net290),
    .C1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__a2111o_4 _3622_ (.A1(net257),
    .A2(_0997_),
    .B1(_0998_),
    .C1(_0996_),
    .D1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__nor4_2 _3623_ (.A(_0991_),
    .B(_0993_),
    .C(_0995_),
    .D(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__a32o_1 _3624_ (.A1(\gpio_configure[2][5] ),
    .A2(_0890_),
    .A3(net378),
    .B1(_0938_),
    .B2(\gpio_configure[13][5] ),
    .X(_1003_));
 sky130_fd_sc_hd__a221o_1 _3625_ (.A1(\gpio_configure[22][5] ),
    .A2(_0913_),
    .B1(_0921_),
    .B2(\gpio_configure[30][5] ),
    .C1(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__a32o_1 _3626_ (.A1(\gpio_configure[18][5] ),
    .A2(net359),
    .A3(_0890_),
    .B1(_0939_),
    .B2(\gpio_configure[5][5] ),
    .X(_1005_));
 sky130_fd_sc_hd__a221o_1 _3627_ (.A1(\gpio_configure[7][5] ),
    .A2(_0914_),
    .B1(_0915_),
    .B2(net57),
    .C1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__a32o_1 _3628_ (.A1(\gpio_configure[32][5] ),
    .A2(net384),
    .A3(net355),
    .B1(_0927_),
    .B2(\gpio_configure[17][5] ),
    .X(_1007_));
 sky130_fd_sc_hd__a221o_1 _3629_ (.A1(\gpio_configure[16][5] ),
    .A2(_0876_),
    .B1(_0895_),
    .B2(\gpio_configure[3][5] ),
    .C1(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__a32o_1 _3630_ (.A1(\gpio_configure[12][5] ),
    .A2(net390),
    .A3(net387),
    .B1(_0886_),
    .B2(net31),
    .X(_1009_));
 sky130_fd_sc_hd__a221o_1 _3631_ (.A1(net68),
    .A2(_0935_),
    .B1(_0936_),
    .B2(net40),
    .C1(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__nor4_2 _3632_ (.A(_1004_),
    .B(_1006_),
    .C(_1008_),
    .D(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__a32o_1 _3633_ (.A1(\gpio_configure[25][5] ),
    .A2(net354),
    .A3(net403),
    .B1(_0903_),
    .B2(\gpio_configure[20][5] ),
    .X(_1012_));
 sky130_fd_sc_hd__a221o_1 _3634_ (.A1(\gpio_configure[27][5] ),
    .A2(_0880_),
    .B1(_0909_),
    .B2(\gpio_configure[28][5] ),
    .C1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__a32o_1 _3635_ (.A1(\gpio_configure[26][5] ),
    .A2(net355),
    .A3(_0890_),
    .B1(_0948_),
    .B2(\gpio_configure[23][5] ),
    .X(_1014_));
 sky130_fd_sc_hd__a221o_1 _3636_ (.A1(net8),
    .A2(_0869_),
    .B1(_0912_),
    .B2(\gpio_configure[31][5] ),
    .C1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and3_4 _3637_ (.A(net420),
    .B(net412),
    .C(net380),
    .X(_1016_));
 sky130_fd_sc_hd__a32o_1 _3638_ (.A1(\gpio_configure[36][5] ),
    .A2(net387),
    .A3(net380),
    .B1(\gpio_configure[21][5] ),
    .B2(_0861_),
    .X(_1017_));
 sky130_fd_sc_hd__a221o_4 _3639_ (.A1(\gpio_configure[37][5] ),
    .A2(_0884_),
    .B1(_1016_),
    .B2(net66),
    .C1(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__a32o_1 _3640_ (.A1(\gpio_configure[14][5] ),
    .A2(net390),
    .A3(net389),
    .B1(_0947_),
    .B2(\gpio_configure[10][5] ),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_1 _3641_ (.A1(\gpio_configure[11][5] ),
    .A2(_0901_),
    .B1(_0910_),
    .B2(net273),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__nor4_2 _3642_ (.A(_1013_),
    .B(_1015_),
    .C(_1018_),
    .D(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__nand3_4 _3643_ (.A(_1002_),
    .B(_1011_),
    .C(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(\hkspi.ldata[4] ),
    .A1(_1022_),
    .S(net509),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(_1023_),
    .A1(net3806),
    .S(_0954_),
    .X(_0389_));
 sky130_fd_sc_hd__and3_4 _3646_ (.A(net413),
    .B(net410),
    .C(net378),
    .X(_1024_));
 sky130_fd_sc_hd__and3_2 _3647_ (.A(net416),
    .B(net411),
    .C(net354),
    .X(_1025_));
 sky130_fd_sc_hd__and3_2 _3648_ (.A(net390),
    .B(net409),
    .C(net407),
    .X(_1026_));
 sky130_fd_sc_hd__and3_2 _3649_ (.A(net411),
    .B(net354),
    .C(net408),
    .X(_1027_));
 sky130_fd_sc_hd__and3_4 _3650_ (.A(net358),
    .B(net413),
    .C(net411),
    .X(_1028_));
 sky130_fd_sc_hd__and3_2 _3651_ (.A(net413),
    .B(net356),
    .C(net409),
    .X(_1029_));
 sky130_fd_sc_hd__and3_2 _3652_ (.A(net412),
    .B(net381),
    .C(net408),
    .X(_1030_));
 sky130_fd_sc_hd__and3_4 _3653_ (.A(net660),
    .B(net409),
    .C(net378),
    .X(_1031_));
 sky130_fd_sc_hd__and3_2 _3654_ (.A(net414),
    .B(net381),
    .C(net409),
    .X(_1032_));
 sky130_fd_sc_hd__and4_1 _3655_ (.A(net65),
    .B(net421),
    .C(net412),
    .D(net381),
    .X(_1033_));
 sky130_fd_sc_hd__and3_4 _3656_ (.A(net391),
    .B(net414),
    .C(net411),
    .X(_1034_));
 sky130_fd_sc_hd__and3_4 _3657_ (.A(net415),
    .B(net410),
    .C(net373),
    .X(_1035_));
 sky130_fd_sc_hd__and3_2 _3658_ (.A(net391),
    .B(net414),
    .C(net409),
    .X(_1036_));
 sky130_fd_sc_hd__and3_2 _3659_ (.A(net413),
    .B(net409),
    .C(net378),
    .X(_1037_));
 sky130_fd_sc_hd__and3_4 _3660_ (.A(net414),
    .B(net412),
    .C(net381),
    .X(_1038_));
 sky130_fd_sc_hd__and3_2 _3661_ (.A(net391),
    .B(net411),
    .C(net408),
    .X(_1039_));
 sky130_fd_sc_hd__and3_4 _3662_ (.A(net357),
    .B(net415),
    .C(net410),
    .X(_1040_));
 sky130_fd_sc_hd__and3_2 _3663_ (.A(net357),
    .B(net411),
    .C(net407),
    .X(_1041_));
 sky130_fd_sc_hd__and3_4 _3664_ (.A(net390),
    .B(net415),
    .C(net410),
    .X(_1042_));
 sky130_fd_sc_hd__and3_2 _3665_ (.A(net391),
    .B(net420),
    .C(net411),
    .X(_1043_));
 sky130_fd_sc_hd__and3_4 _3666_ (.A(net421),
    .B(net410),
    .C(net378),
    .X(_1044_));
 sky130_fd_sc_hd__and3_4 _3667_ (.A(net415),
    .B(net410),
    .C(net378),
    .X(_1045_));
 sky130_fd_sc_hd__and3_4 _3668_ (.A(net357),
    .B(net413),
    .C(net409),
    .X(_1046_));
 sky130_fd_sc_hd__and3_4 _3669_ (.A(net412),
    .B(net408),
    .C(net379),
    .X(_1047_));
 sky130_fd_sc_hd__and3_2 _3670_ (.A(net391),
    .B(net421),
    .C(net409),
    .X(_1048_));
 sky130_fd_sc_hd__and3_4 _3671_ (.A(net660),
    .B(net409),
    .C(net373),
    .X(_1049_));
 sky130_fd_sc_hd__and3_4 _3672_ (.A(net391),
    .B(net416),
    .C(net409),
    .X(_1050_));
 sky130_fd_sc_hd__and3_2 _3673_ (.A(net420),
    .B(net358),
    .C(net411),
    .X(_1051_));
 sky130_fd_sc_hd__and3_4 _3674_ (.A(net413),
    .B(net410),
    .C(net354),
    .X(_1052_));
 sky130_fd_sc_hd__and3_4 _3675_ (.A(net421),
    .B(net410),
    .C(net354),
    .X(_1053_));
 sky130_fd_sc_hd__a32o_1 _3676_ (.A1(\gpio_configure[27][12] ),
    .A2(net354),
    .A3(net371),
    .B1(_1024_),
    .B2(\gpio_configure[4][12] ),
    .X(_1054_));
 sky130_fd_sc_hd__a32o_1 _3677_ (.A1(\gpio_configure[32][4] ),
    .A2(net384),
    .A3(net355),
    .B1(_0952_),
    .B2(\gpio_configure[26][4] ),
    .X(_1055_));
 sky130_fd_sc_hd__a32o_1 _3678_ (.A1(\gpio_configure[31][12] ),
    .A2(net356),
    .A3(net374),
    .B1(_1025_),
    .B2(\gpio_configure[32][12] ),
    .X(_1056_));
 sky130_fd_sc_hd__a41o_1 _3679_ (.A1(\gpio_configure[30][12] ),
    .A2(net420),
    .A3(net411),
    .A4(net354),
    .B1(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__a221o_1 _3680_ (.A1(\gpio_configure[10][4] ),
    .A2(_0947_),
    .B1(_1026_),
    .B2(\gpio_configure[11][12] ),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__a2111o_1 _3681_ (.A1(\gpio_configure[24][12] ),
    .A2(_1040_),
    .B1(_1054_),
    .C1(_1055_),
    .D1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__and3_2 _3682_ (.A(net419),
    .B(net407),
    .C(net372),
    .X(_1060_));
 sky130_fd_sc_hd__a32o_2 _3683_ (.A1(net264),
    .A2(_0890_),
    .A3(net372),
    .B1(_0959_),
    .B2(serial_bb_clock),
    .X(_1061_));
 sky130_fd_sc_hd__a32o_1 _3684_ (.A1(\gpio_configure[0][4] ),
    .A2(net384),
    .A3(net373),
    .B1(_0861_),
    .B2(\gpio_configure[21][4] ),
    .X(_1062_));
 sky130_fd_sc_hd__a31o_1 _3685_ (.A1(\gpio_configure[33][12] ),
    .A2(net354),
    .A3(net375),
    .B1(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__a2111o_2 _3686_ (.A1(net256),
    .A2(_0997_),
    .B1(_1059_),
    .C1(_1061_),
    .D1(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__a32o_1 _3687_ (.A1(\gpio_configure[19][12] ),
    .A2(net359),
    .A3(net370),
    .B1(_0920_),
    .B2(\gpio_configure[18][4] ),
    .X(_1065_));
 sky130_fd_sc_hd__a31o_1 _3688_ (.A1(\gpio_configure[17][4] ),
    .A2(net359),
    .A3(net403),
    .B1(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a221o_1 _3689_ (.A1(\gpio_configure[19][4] ),
    .A2(_0908_),
    .B1(_1029_),
    .B2(\gpio_configure[29][12] ),
    .C1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__a32o_1 _3690_ (.A1(\gpio_configure[6][4] ),
    .A2(net389),
    .A3(net379),
    .B1(_1044_),
    .B2(\gpio_configure[6][12] ),
    .X(_1068_));
 sky130_fd_sc_hd__a32o_1 _3691_ (.A1(\gpio_configure[2][4] ),
    .A2(_0890_),
    .A3(net379),
    .B1(_0865_),
    .B2(\gpio_configure[15][4] ),
    .X(_1069_));
 sky130_fd_sc_hd__a32o_1 _3692_ (.A1(\gpio_configure[23][12] ),
    .A2(net358),
    .A3(net374),
    .B1(_1027_),
    .B2(\gpio_configure[26][12] ),
    .X(_1070_));
 sky130_fd_sc_hd__a32o_1 _3693_ (.A1(\gpio_configure[8][4] ),
    .A2(net384),
    .A3(net379),
    .B1(_1037_),
    .B2(\gpio_configure[5][12] ),
    .X(_1071_));
 sky130_fd_sc_hd__a31o_1 _3694_ (.A1(\gpio_configure[7][12] ),
    .A2(net379),
    .A3(net374),
    .B1(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__a211o_1 _3695_ (.A1(\gpio_configure[23][4] ),
    .A2(_0948_),
    .B1(_1070_),
    .C1(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a2111oi_1 _3696_ (.A1(\gpio_configure[21][12] ),
    .A2(_1046_),
    .B1(_1068_),
    .C1(_1069_),
    .D1(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__a32o_1 _3697_ (.A1(\gpio_configure[15][12] ),
    .A2(net391),
    .A3(net374),
    .B1(_1039_),
    .B2(\gpio_configure[10][12] ),
    .X(_1075_));
 sky130_fd_sc_hd__a221o_1 _3698_ (.A1(\gpio_configure[14][4] ),
    .A2(_0856_),
    .B1(_1028_),
    .B2(\gpio_configure[20][12] ),
    .C1(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__a32o_1 _3699_ (.A1(\gpio_configure[9][4] ),
    .A2(net392),
    .A3(net403),
    .B1(_0881_),
    .B2(\gpio_configure[12][4] ),
    .X(_1077_));
 sky130_fd_sc_hd__a32o_1 _3700_ (.A1(\gpio_configure[30][4] ),
    .A2(net388),
    .A3(net356),
    .B1(_1051_),
    .B2(\gpio_configure[22][12] ),
    .X(_1078_));
 sky130_fd_sc_hd__a221o_1 _3701_ (.A1(\gpio_configure[24][4] ),
    .A2(_0877_),
    .B1(_0912_),
    .B2(\gpio_configure[31][4] ),
    .C1(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__a2111o_2 _3702_ (.A1(\gpio_configure[11][4] ),
    .A2(_0901_),
    .B1(_1076_),
    .C1(_1077_),
    .D1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__a22o_1 _3703_ (.A1(\gpio_configure[13][4] ),
    .A2(_0938_),
    .B1(_1036_),
    .B2(\gpio_configure[13][12] ),
    .X(_1081_));
 sky130_fd_sc_hd__a31o_1 _3704_ (.A1(\gpio_configure[25][12] ),
    .A2(net359),
    .A3(net375),
    .B1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a22o_1 _3705_ (.A1(\gpio_configure[12][12] ),
    .A2(_1034_),
    .B1(_1043_),
    .B2(\gpio_configure[14][12] ),
    .X(_1083_));
 sky130_fd_sc_hd__a221o_4 _3706_ (.A1(\gpio_configure[28][4] ),
    .A2(_0909_),
    .B1(_0918_),
    .B2(\gpio_configure[25][4] ),
    .C1(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__a32o_1 _3707_ (.A1(\gpio_configure[33][4] ),
    .A2(net382),
    .A3(net403),
    .B1(_0891_),
    .B2(\gpio_configure[34][4] ),
    .X(_1085_));
 sky130_fd_sc_hd__a32o_1 _3708_ (.A1(net7),
    .A2(net387),
    .A3(_0868_),
    .B1(_0915_),
    .B2(net56),
    .X(_1086_));
 sky130_fd_sc_hd__a221o_1 _3709_ (.A1(\gpio_configure[34][12] ),
    .A2(_1030_),
    .B1(_1032_),
    .B2(\gpio_configure[37][12] ),
    .C1(_1033_),
    .X(_1087_));
 sky130_fd_sc_hd__a221o_2 _3710_ (.A1(\gpio_configure[37][4] ),
    .A2(_0884_),
    .B1(_0935_),
    .B2(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__a2111o_2 _3711_ (.A1(net24),
    .A2(_0871_),
    .B1(_1085_),
    .C1(_1086_),
    .D1(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__a2111o_2 _3712_ (.A1(\gpio_configure[29][4] ),
    .A2(_0933_),
    .B1(_1082_),
    .C1(_1084_),
    .D1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a32o_4 _3713_ (.A1(\gpio_configure[1][4] ),
    .A2(net403),
    .A3(net377),
    .B1(net30),
    .B2(_0886_),
    .X(_1091_));
 sky130_fd_sc_hd__a32o_2 _3714_ (.A1(\gpio_configure[1][12] ),
    .A2(net375),
    .A3(net373),
    .B1(_1041_),
    .B2(\gpio_configure[18][12] ),
    .X(_1092_));
 sky130_fd_sc_hd__a32o_2 _3715_ (.A1(net272),
    .A2(net385),
    .A3(net383),
    .B1(_0898_),
    .B2(net281),
    .X(_1093_));
 sky130_fd_sc_hd__a221o_2 _3716_ (.A1(\gpio_configure[16][4] ),
    .A2(_0876_),
    .B1(_0880_),
    .B2(\gpio_configure[27][4] ),
    .C1(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__a2111o_1 _3717_ (.A1(\gpio_configure[22][4] ),
    .A2(_0913_),
    .B1(_1091_),
    .C1(_1092_),
    .D1(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__a32o_1 _3718_ (.A1(\gpio_configure[9][12] ),
    .A2(net379),
    .A3(net375),
    .B1(_0903_),
    .B2(\gpio_configure[20][4] ),
    .X(_1096_));
 sky130_fd_sc_hd__a41o_1 _3719_ (.A1(\gpio_configure[16][12] ),
    .A2(net390),
    .A3(net416),
    .A4(net411),
    .B1(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__a32o_1 _3720_ (.A1(_0853_),
    .A2(_0868_),
    .A3(net408),
    .B1(_1047_),
    .B2(\gpio_configure[2][12] ),
    .X(_1098_));
 sky130_fd_sc_hd__a221o_1 _3721_ (.A1(net16),
    .A2(_0873_),
    .B1(_1052_),
    .B2(\gpio_configure[28][12] ),
    .C1(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__a2111o_1 _3722_ (.A1(\gpio_configure[0][12] ),
    .A2(_1035_),
    .B1(_1095_),
    .C1(_1097_),
    .D1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__a32o_1 _3723_ (.A1(\gpio_configure[3][12] ),
    .A2(net377),
    .A3(net370),
    .B1(_0914_),
    .B2(\gpio_configure[7][4] ),
    .X(_1101_));
 sky130_fd_sc_hd__a22o_1 _3724_ (.A1(net289),
    .A2(_0925_),
    .B1(_0939_),
    .B2(\gpio_configure[5][4] ),
    .X(_1102_));
 sky130_fd_sc_hd__a32o_4 _3725_ (.A1(\clk1_output_dest[1] ),
    .A2(net374),
    .A3(net373),
    .B1(_1050_),
    .B2(\gpio_configure[17][12] ),
    .X(_1103_));
 sky130_fd_sc_hd__a221o_1 _3726_ (.A1(\gpio_configure[3][4] ),
    .A2(_0895_),
    .B1(_1045_),
    .B2(\gpio_configure[8][12] ),
    .C1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a2111o_4 _3727_ (.A1(\gpio_configure[4][4] ),
    .A2(_0904_),
    .B1(_1101_),
    .C1(_1102_),
    .D1(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__a32o_1 _3728_ (.A1(\gpio_configure[35][12] ),
    .A2(net381),
    .A3(net371),
    .B1(_0899_),
    .B2(\gpio_configure[35][4] ),
    .X(_1106_));
 sky130_fd_sc_hd__a41o_1 _3729_ (.A1(\gpio_configure[36][12] ),
    .A2(net414),
    .A3(net412),
    .A4(net381),
    .B1(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__a32o_1 _3730_ (.A1(\gpio_configure[36][4] ),
    .A2(net387),
    .A3(net381),
    .B1(_0932_),
    .B2(net48),
    .X(_1108_));
 sky130_fd_sc_hd__a2111o_1 _3731_ (.A1(net39),
    .A2(_0936_),
    .B1(_1105_),
    .C1(_1107_),
    .D1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__nor4_2 _3732_ (.A(_1080_),
    .B(_1090_),
    .C(_1100_),
    .D(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__and4bb_2 _3733_ (.A_N(_1064_),
    .B_N(_1067_),
    .C(_1074_),
    .D(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_2 _3734_ (.A(net509),
    .B(clknet_1_1__leaf__1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__o211a_1 _3735_ (.A1(net3803),
    .A2(_0829_),
    .B1(\hkspi.state[2] ),
    .C1(\hkspi.readmode ),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_2 _3736_ (.A1(\hkspi.ldata[4] ),
    .A2(_0954_),
    .B1(_1112_),
    .B2(_1113_),
    .X(_0388_));
 sky130_fd_sc_hd__and3_1 _3737_ (.A(\gpio_configure[30][3] ),
    .B(net388),
    .C(net356),
    .X(_1114_));
 sky130_fd_sc_hd__and3_1 _3738_ (.A(\clk2_output_dest[1] ),
    .B(net374),
    .C(net373),
    .X(_1115_));
 sky130_fd_sc_hd__a32o_1 _3739_ (.A1(\gpio_configure[1][3] ),
    .A2(net403),
    .A3(net379),
    .B1(_1024_),
    .B2(\gpio_configure[4][11] ),
    .X(_1116_));
 sky130_fd_sc_hd__a32o_1 _3740_ (.A1(\gpio_configure[36][3] ),
    .A2(net387),
    .A3(net380),
    .B1(_1016_),
    .B2(net64),
    .X(_1117_));
 sky130_fd_sc_hd__a41o_1 _3741_ (.A1(\gpio_configure[37][11] ),
    .A2(net414),
    .A3(net380),
    .A4(_0885_),
    .B1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__a32o_1 _3742_ (.A1(\gpio_configure[35][11] ),
    .A2(net382),
    .A3(net371),
    .B1(_0914_),
    .B2(\gpio_configure[7][3] ),
    .X(_1119_));
 sky130_fd_sc_hd__a221o_1 _3743_ (.A1(\gpio_configure[35][3] ),
    .A2(_0899_),
    .B1(_0936_),
    .B2(net38),
    .C1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a311o_1 _3744_ (.A1(\gpio_configure[33][3] ),
    .A2(net380),
    .A3(net403),
    .B1(_1118_),
    .C1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__a22o_1 _3745_ (.A1(\gpio_configure[11][3] ),
    .A2(_0901_),
    .B1(_1034_),
    .B2(\gpio_configure[12][11] ),
    .X(_1122_));
 sky130_fd_sc_hd__a32o_1 _3746_ (.A1(\gpio_configure[14][3] ),
    .A2(net391),
    .A3(net388),
    .B1(_1043_),
    .B2(\gpio_configure[14][11] ),
    .X(_1123_));
 sky130_fd_sc_hd__a221o_1 _3747_ (.A1(\gpio_configure[20][11] ),
    .A2(_1028_),
    .B1(_1048_),
    .B2(\gpio_configure[15][11] ),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a221o_2 _3748_ (.A1(\gpio_configure[9][3] ),
    .A2(_0889_),
    .B1(_0938_),
    .B2(\gpio_configure[13][3] ),
    .C1(_1115_),
    .X(_1125_));
 sky130_fd_sc_hd__a221o_1 _3749_ (.A1(\gpio_configure[13][11] ),
    .A2(_1036_),
    .B1(_1039_),
    .B2(\gpio_configure[10][11] ),
    .C1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__a2111o_1 _3750_ (.A1(\gpio_configure[12][3] ),
    .A2(_0881_),
    .B1(_1122_),
    .C1(_1124_),
    .D1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__a32o_1 _3751_ (.A1(\gpio_configure[25][11] ),
    .A2(net358),
    .A3(net375),
    .B1(_1050_),
    .B2(\gpio_configure[17][11] ),
    .X(_1128_));
 sky130_fd_sc_hd__a221o_1 _3752_ (.A1(\gpio_configure[31][3] ),
    .A2(_0912_),
    .B1(_0918_),
    .B2(\gpio_configure[25][3] ),
    .C1(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__a32o_1 _3753_ (.A1(net95),
    .A2(net388),
    .A3(net373),
    .B1(_0909_),
    .B2(\gpio_configure[28][3] ),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _3754_ (.A1(\gpio_configure[29][3] ),
    .A2(_0933_),
    .B1(_1051_),
    .B2(\gpio_configure[22][11] ),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__a22o_1 _3755_ (.A1(net67),
    .A2(_0935_),
    .B1(_1030_),
    .B2(\gpio_configure[34][11] ),
    .X(_1132_));
 sky130_fd_sc_hd__a221o_1 _3756_ (.A1(\gpio_configure[34][3] ),
    .A2(_0891_),
    .B1(_0932_),
    .B2(net46),
    .C1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__a32o_1 _3757_ (.A1(net55),
    .A2(net388),
    .A3(net380),
    .B1(_0884_),
    .B2(\gpio_configure[37][3] ),
    .X(_1134_));
 sky130_fd_sc_hd__a221o_1 _3758_ (.A1(\gpio_configure[3][3] ),
    .A2(_0895_),
    .B1(_1038_),
    .B2(\gpio_configure[36][11] ),
    .C1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__nor4_2 _3759_ (.A(_1129_),
    .B(_1131_),
    .C(_1133_),
    .D(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__a32o_1 _3760_ (.A1(\gpio_configure[3][11] ),
    .A2(net378),
    .A3(net370),
    .B1(_1045_),
    .B2(\gpio_configure[8][11] ),
    .X(_1137_));
 sky130_fd_sc_hd__a32o_1 _3761_ (.A1(net6),
    .A2(net387),
    .A3(net385),
    .B1(_0925_),
    .B2(net288),
    .X(_1138_));
 sky130_fd_sc_hd__a221o_4 _3762_ (.A1(\gpio_configure[24][3] ),
    .A2(_0877_),
    .B1(_0939_),
    .B2(\gpio_configure[5][3] ),
    .C1(_1114_),
    .X(_1139_));
 sky130_fd_sc_hd__a221o_1 _3763_ (.A1(net23),
    .A2(_0871_),
    .B1(_0904_),
    .B2(\gpio_configure[4][3] ),
    .C1(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__a2111o_4 _3764_ (.A1(net14),
    .A2(_0873_),
    .B1(_1137_),
    .C1(_1138_),
    .D1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__a32o_1 _3765_ (.A1(\gpio_configure[33][11] ),
    .A2(net354),
    .A3(net375),
    .B1(_1040_),
    .B2(\gpio_configure[24][11] ),
    .X(_1142_));
 sky130_fd_sc_hd__a32o_1 _3766_ (.A1(\gpio_configure[22][3] ),
    .A2(net388),
    .A3(net358),
    .B1(_0920_),
    .B2(\gpio_configure[18][3] ),
    .X(_1143_));
 sky130_fd_sc_hd__a221o_1 _3767_ (.A1(\gpio_configure[6][3] ),
    .A2(_0944_),
    .B1(_0945_),
    .B2(\gpio_configure[2][3] ),
    .C1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__a32o_1 _3768_ (.A1(\gpio_configure[17][3] ),
    .A2(net358),
    .A3(net403),
    .B1(_1047_),
    .B2(\gpio_configure[2][11] ),
    .X(_1145_));
 sky130_fd_sc_hd__a221o_1 _3769_ (.A1(net29),
    .A2(_0886_),
    .B1(_0903_),
    .B2(\gpio_configure[20][3] ),
    .C1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__a32o_1 _3770_ (.A1(\gpio_configure[9][11] ),
    .A2(net379),
    .A3(net375),
    .B1(_1027_),
    .B2(\gpio_configure[26][11] ),
    .X(_1147_));
 sky130_fd_sc_hd__a221o_1 _3771_ (.A1(\gpio_configure[27][3] ),
    .A2(_0880_),
    .B1(_1052_),
    .B2(\gpio_configure[28][11] ),
    .C1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__a2111o_1 _3772_ (.A1(\gpio_configure[29][11] ),
    .A2(_1029_),
    .B1(_1144_),
    .C1(_1146_),
    .D1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__a211o_1 _3773_ (.A1(\gpio_configure[26][3] ),
    .A2(_0952_),
    .B1(_1142_),
    .C1(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__a32o_2 _3774_ (.A1(serial_bb_load),
    .A2(net372),
    .A3(net370),
    .B1(_1026_),
    .B2(\gpio_configure[11][11] ),
    .X(_1151_));
 sky130_fd_sc_hd__a221o_1 _3775_ (.A1(\gpio_configure[15][3] ),
    .A2(_0865_),
    .B1(_0947_),
    .B2(\gpio_configure[10][3] ),
    .C1(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a32o_1 _3776_ (.A1(\gpio_configure[1][11] ),
    .A2(net376),
    .A3(net372),
    .B1(_1035_),
    .B2(\gpio_configure[0][11] ),
    .X(_1153_));
 sky130_fd_sc_hd__a221o_4 _3777_ (.A1(\gpio_configure[0][3] ),
    .A2(_0941_),
    .B1(_1060_),
    .B2(net263),
    .C1(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__a31o_1 _3778_ (.A1(\gpio_configure[27][11] ),
    .A2(net354),
    .A3(net371),
    .B1(_1116_),
    .X(_1155_));
 sky130_fd_sc_hd__a22o_1 _3779_ (.A1(\gpio_configure[5][11] ),
    .A2(_1037_),
    .B1(_1042_),
    .B2(\gpio_configure[16][11] ),
    .X(_1156_));
 sky130_fd_sc_hd__a221o_1 _3780_ (.A1(\gpio_configure[21][3] ),
    .A2(_0861_),
    .B1(_1046_),
    .B2(\gpio_configure[21][11] ),
    .C1(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__a31o_1 _3781_ (.A1(\gpio_configure[16][3] ),
    .A2(net390),
    .A3(net384),
    .B1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__nor4_1 _3782_ (.A(_1152_),
    .B(_1154_),
    .C(_1155_),
    .D(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__a32o_4 _3783_ (.A1(net271),
    .A2(net386),
    .A3(net383),
    .B1(_0997_),
    .B2(net255),
    .X(_1160_));
 sky130_fd_sc_hd__a32o_2 _3784_ (.A1(\gpio_configure[32][3] ),
    .A2(net384),
    .A3(net356),
    .B1(_0948_),
    .B2(\gpio_configure[23][3] ),
    .X(_1161_));
 sky130_fd_sc_hd__a32o_1 _3785_ (.A1(\gpio_configure[31][11] ),
    .A2(net356),
    .A3(net374),
    .B1(_1053_),
    .B2(\gpio_configure[30][11] ),
    .X(_1162_));
 sky130_fd_sc_hd__a221o_1 _3786_ (.A1(\gpio_configure[18][11] ),
    .A2(_1041_),
    .B1(_1044_),
    .B2(\gpio_configure[6][11] ),
    .C1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__a32o_4 _3787_ (.A1(net298),
    .A2(net383),
    .A3(_0883_),
    .B1(_0898_),
    .B2(net279),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _3788_ (.A1(\gpio_configure[32][11] ),
    .A2(_1025_),
    .B1(_1031_),
    .B2(\gpio_configure[7][11] ),
    .C1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__a32o_2 _3789_ (.A1(\gpio_configure[8][3] ),
    .A2(net384),
    .A3(net379),
    .B1(_0908_),
    .B2(\gpio_configure[19][3] ),
    .X(_1166_));
 sky130_fd_sc_hd__a31o_1 _3790_ (.A1(\gpio_configure[19][11] ),
    .A2(net358),
    .A3(net371),
    .B1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__a311o_1 _3791_ (.A1(\gpio_configure[23][11] ),
    .A2(net357),
    .A3(net374),
    .B1(_1165_),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__nor4_1 _3792_ (.A(_1160_),
    .B(_1161_),
    .C(_1163_),
    .D(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__and4bb_4 _3793_ (.A_N(_1141_),
    .B_N(_1150_),
    .C(_1159_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__and4bb_4 _3794_ (.A_N(_1121_),
    .B_N(_1127_),
    .C(_1136_),
    .D(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(net509),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__o211a_1 _3796_ (.A1(\hkspi.ldata[2] ),
    .A2(_0829_),
    .B1(\hkspi.state[2] ),
    .C1(\hkspi.readmode ),
    .X(_1173_));
 sky130_fd_sc_hd__a22o_1 _3797_ (.A1(net3803),
    .A2(_0954_),
    .B1(_1172_),
    .B2(_1173_),
    .X(_0387_));
 sky130_fd_sc_hd__a32o_1 _3798_ (.A1(\gpio_configure[36][2] ),
    .A2(net387),
    .A3(net382),
    .B1(_1032_),
    .B2(\gpio_configure[37][10] ),
    .X(_1174_));
 sky130_fd_sc_hd__a32o_1 _3799_ (.A1(\gpio_configure[20][2] ),
    .A2(net357),
    .A3(net387),
    .B1(_1046_),
    .B2(\gpio_configure[21][10] ),
    .X(_1175_));
 sky130_fd_sc_hd__a31o_4 _3800_ (.A1(\gpio_configure[35][10] ),
    .A2(net382),
    .A3(net371),
    .B1(_1174_),
    .X(_1176_));
 sky130_fd_sc_hd__a32o_4 _3801_ (.A1(_0868_),
    .A2(net412),
    .A3(net407),
    .B1(_0884_),
    .B2(\gpio_configure[37][2] ),
    .X(_1177_));
 sky130_fd_sc_hd__a221o_2 _3802_ (.A1(net5),
    .A2(_0869_),
    .B1(_0873_),
    .B2(net13),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__a32o_1 _3803_ (.A1(\gpio_configure[9][2] ),
    .A2(net390),
    .A3(net403),
    .B1(_0901_),
    .B2(\gpio_configure[11][2] ),
    .X(_1179_));
 sky130_fd_sc_hd__a221o_1 _3804_ (.A1(\gpio_configure[30][2] ),
    .A2(_0921_),
    .B1(_0938_),
    .B2(\gpio_configure[13][2] ),
    .C1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__a32o_1 _3805_ (.A1(net97),
    .A2(net388),
    .A3(net373),
    .B1(_1049_),
    .B2(\clk1_output_dest[0] ),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_4 _3806_ (.A1(\gpio_configure[31][2] ),
    .A2(_0912_),
    .B1(_1048_),
    .B2(\gpio_configure[15][10] ),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a32o_1 _3807_ (.A1(\gpio_configure[3][10] ),
    .A2(net377),
    .A3(net370),
    .B1(_0914_),
    .B2(\gpio_configure[7][2] ),
    .X(_1183_));
 sky130_fd_sc_hd__a221o_1 _3808_ (.A1(\gpio_configure[3][2] ),
    .A2(_0895_),
    .B1(_0939_),
    .B2(\gpio_configure[5][2] ),
    .C1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__a2111o_1 _3809_ (.A1(\gpio_configure[4][2] ),
    .A2(_0904_),
    .B1(_1180_),
    .C1(_1182_),
    .D1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__a2111oi_2 _3810_ (.A1(\gpio_configure[34][2] ),
    .A2(_0891_),
    .B1(_1176_),
    .C1(_1178_),
    .D1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a32o_1 _3811_ (.A1(\gpio_configure[1][2] ),
    .A2(net403),
    .A3(net378),
    .B1(_1044_),
    .B2(\gpio_configure[6][10] ),
    .X(_1187_));
 sky130_fd_sc_hd__a221o_1 _3812_ (.A1(\gpio_configure[26][2] ),
    .A2(_0952_),
    .B1(_1047_),
    .B2(\gpio_configure[2][10] ),
    .C1(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__a32o_1 _3813_ (.A1(\gpio_configure[24][2] ),
    .A2(net357),
    .A3(net383),
    .B1(_0997_),
    .B2(net268),
    .X(_1189_));
 sky130_fd_sc_hd__a32o_1 _3814_ (.A1(\gpio_configure[2][2] ),
    .A2(_0890_),
    .A3(net377),
    .B1(net26),
    .B2(_0886_),
    .X(_1190_));
 sky130_fd_sc_hd__a221o_1 _3815_ (.A1(net270),
    .A2(_0910_),
    .B1(_1031_),
    .B2(\gpio_configure[7][10] ),
    .C1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__a32o_1 _3816_ (.A1(\gpio_configure[31][10] ),
    .A2(net355),
    .A3(net374),
    .B1(\gpio_configure[15][2] ),
    .B2(_0865_),
    .X(_1192_));
 sky130_fd_sc_hd__a221o_1 _3817_ (.A1(\gpio_configure[0][2] ),
    .A2(_0941_),
    .B1(_1037_),
    .B2(\gpio_configure[5][10] ),
    .C1(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__a2111o_1 _3818_ (.A1(\gpio_configure[4][10] ),
    .A2(_1024_),
    .B1(_1175_),
    .C1(_1191_),
    .D1(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__a2111oi_2 _3819_ (.A1(\gpio_configure[27][2] ),
    .A2(_0880_),
    .B1(_1188_),
    .C1(_1189_),
    .D1(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__a32o_1 _3820_ (.A1(\gpio_configure[25][10] ),
    .A2(net357),
    .A3(net376),
    .B1(_0947_),
    .B2(\gpio_configure[10][2] ),
    .X(_1196_));
 sky130_fd_sc_hd__a32o_1 _3821_ (.A1(\gpio_configure[9][10] ),
    .A2(net379),
    .A3(net376),
    .B1(_0861_),
    .B2(\gpio_configure[21][2] ),
    .X(_1197_));
 sky130_fd_sc_hd__a32o_1 _3822_ (.A1(\gpio_configure[33][10] ),
    .A2(net354),
    .A3(net375),
    .B1(_1025_),
    .B2(\gpio_configure[32][10] ),
    .X(_1198_));
 sky130_fd_sc_hd__a221o_1 _3823_ (.A1(\gpio_configure[23][2] ),
    .A2(_0948_),
    .B1(_1029_),
    .B2(\gpio_configure[29][10] ),
    .C1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__a32o_1 _3824_ (.A1(serial_bb_resetn),
    .A2(net372),
    .A3(net370),
    .B1(_1041_),
    .B2(\gpio_configure[18][10] ),
    .X(_1200_));
 sky130_fd_sc_hd__a32o_1 _3825_ (.A1(\gpio_configure[19][10] ),
    .A2(net357),
    .A3(net370),
    .B1(_1052_),
    .B2(\gpio_configure[28][10] ),
    .X(_1201_));
 sky130_fd_sc_hd__a221o_1 _3826_ (.A1(\gpio_configure[8][2] ),
    .A2(_0928_),
    .B1(_1027_),
    .B2(\gpio_configure[26][10] ),
    .C1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__a311o_1 _3827_ (.A1(\gpio_configure[11][10] ),
    .A2(net390),
    .A3(net370),
    .B1(_1200_),
    .C1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__nor4_1 _3828_ (.A(_1196_),
    .B(_1197_),
    .C(_1199_),
    .D(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(\gpio_configure[19][2] ),
    .A2(_0908_),
    .B1(_1042_),
    .B2(\gpio_configure[16][10] ),
    .X(_1205_));
 sky130_fd_sc_hd__a31o_1 _3830_ (.A1(\gpio_configure[1][10] ),
    .A2(net376),
    .A3(net372),
    .B1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a221o_1 _3831_ (.A1(\gpio_configure[16][2] ),
    .A2(_0876_),
    .B1(_1035_),
    .B2(\gpio_configure[0][10] ),
    .C1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__a32o_1 _3832_ (.A1(\gpio_configure[22][2] ),
    .A2(net389),
    .A3(net359),
    .B1(_0920_),
    .B2(\gpio_configure[18][2] ),
    .X(_1208_));
 sky130_fd_sc_hd__a32o_1 _3833_ (.A1(\gpio_configure[32][2] ),
    .A2(net384),
    .A3(net355),
    .B1(_1053_),
    .B2(\gpio_configure[30][10] ),
    .X(_1209_));
 sky130_fd_sc_hd__a32o_1 _3834_ (.A1(\gpio_configure[23][10] ),
    .A2(net357),
    .A3(net374),
    .B1(_0927_),
    .B2(\gpio_configure[17][2] ),
    .X(_1210_));
 sky130_fd_sc_hd__a31o_1 _3835_ (.A1(\gpio_configure[27][10] ),
    .A2(net354),
    .A3(net370),
    .B1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _3836_ (.A1(net278),
    .A2(_0898_),
    .B1(_1040_),
    .B2(\gpio_configure[24][10] ),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__nor4_1 _3837_ (.A(_1207_),
    .B(_1208_),
    .C(_1209_),
    .D(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__a32o_1 _3838_ (.A1(\gpio_configure[12][2] ),
    .A2(net391),
    .A3(net387),
    .B1(_1036_),
    .B2(\gpio_configure[13][10] ),
    .X(_1214_));
 sky130_fd_sc_hd__a22o_1 _3839_ (.A1(\gpio_configure[12][10] ),
    .A2(_1034_),
    .B1(_1051_),
    .B2(\gpio_configure[22][10] ),
    .X(_1215_));
 sky130_fd_sc_hd__a221o_1 _3840_ (.A1(\gpio_configure[20][10] ),
    .A2(_1028_),
    .B1(_1050_),
    .B2(\gpio_configure[17][10] ),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__a32o_1 _3841_ (.A1(\gpio_configure[14][2] ),
    .A2(net392),
    .A3(net389),
    .B1(_1043_),
    .B2(\gpio_configure[14][10] ),
    .X(_1217_));
 sky130_fd_sc_hd__a31o_1 _3842_ (.A1(\gpio_configure[28][2] ),
    .A2(net387),
    .A3(net356),
    .B1(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__a221o_1 _3843_ (.A1(\gpio_configure[25][2] ),
    .A2(_0918_),
    .B1(_1039_),
    .B2(\gpio_configure[10][10] ),
    .C1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__a2111oi_2 _3844_ (.A1(\gpio_configure[29][2] ),
    .A2(_0933_),
    .B1(_1214_),
    .C1(_1216_),
    .D1(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a32o_1 _3845_ (.A1(net54),
    .A2(net388),
    .A3(net381),
    .B1(_0899_),
    .B2(\gpio_configure[35][2] ),
    .X(_1221_));
 sky130_fd_sc_hd__a221o_4 _3846_ (.A1(net58),
    .A2(_0935_),
    .B1(_1030_),
    .B2(\gpio_configure[34][10] ),
    .C1(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__a31o_1 _3847_ (.A1(net297),
    .A2(net383),
    .A3(_0883_),
    .B1(_0979_),
    .X(_1223_));
 sky130_fd_sc_hd__a32o_1 _3848_ (.A1(net262),
    .A2(_0890_),
    .A3(net373),
    .B1(_0944_),
    .B2(\gpio_configure[6][2] ),
    .X(_1224_));
 sky130_fd_sc_hd__a2111o_1 _3849_ (.A1(net45),
    .A2(_0932_),
    .B1(_1222_),
    .C1(_1223_),
    .D1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__a22o_2 _3850_ (.A1(net22),
    .A2(_0871_),
    .B1(_0925_),
    .B2(net287),
    .X(_1226_));
 sky130_fd_sc_hd__a32o_1 _3851_ (.A1(\gpio_configure[33][2] ),
    .A2(net381),
    .A3(net403),
    .B1(_1016_),
    .B2(net63),
    .X(_1227_));
 sky130_fd_sc_hd__a221o_4 _3852_ (.A1(net37),
    .A2(_0936_),
    .B1(_1038_),
    .B2(\gpio_configure[36][10] ),
    .C1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__a2111oi_2 _3853_ (.A1(\gpio_configure[8][10] ),
    .A2(_1045_),
    .B1(_1225_),
    .C1(_1226_),
    .D1(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__and4_1 _3854_ (.A(_1204_),
    .B(_1213_),
    .C(net345),
    .D(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__and3_4 _3855_ (.A(_1186_),
    .B(_1195_),
    .C(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__nand2_1 _3856_ (.A(_0829_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__o211a_1 _3857_ (.A1(net3800),
    .A2(_0829_),
    .B1(\hkspi.state[2] ),
    .C1(\hkspi.readmode ),
    .X(_1233_));
 sky130_fd_sc_hd__a22o_1 _3858_ (.A1(net3812),
    .A2(_0954_),
    .B1(_1232_),
    .B2(_1233_),
    .X(_0386_));
 sky130_fd_sc_hd__and4_2 _3859_ (.A(net62),
    .B(net421),
    .C(net411),
    .D(net380),
    .X(_1234_));
 sky130_fd_sc_hd__and4_1 _3860_ (.A(\gpio_configure[20][9] ),
    .B(net359),
    .C(net413),
    .D(net411),
    .X(_1235_));
 sky130_fd_sc_hd__and4_1 _3861_ (.A(irq_2_inputsrc),
    .B(net417),
    .C(net415),
    .D(net372),
    .X(_1236_));
 sky130_fd_sc_hd__and3_2 _3862_ (.A(net277),
    .B(net385),
    .C(net376),
    .X(_1237_));
 sky130_fd_sc_hd__and4_2 _3863_ (.A(net21),
    .B(net417),
    .C(net413),
    .D(net385),
    .X(_1238_));
 sky130_fd_sc_hd__and3_1 _3864_ (.A(net421),
    .B(net417),
    .C(net386),
    .X(_1239_));
 sky130_fd_sc_hd__and4_2 _3865_ (.A(net259),
    .B(net421),
    .C(net417),
    .D(net386),
    .X(_1240_));
 sky130_fd_sc_hd__a32o_4 _3866_ (.A1(net53),
    .A2(net388),
    .A3(net380),
    .B1(_0932_),
    .B2(net44),
    .X(_1241_));
 sky130_fd_sc_hd__a221o_4 _3867_ (.A1(\gpio_configure[7][1] ),
    .A2(_0914_),
    .B1(_1045_),
    .B2(\gpio_configure[8][9] ),
    .C1(_1238_),
    .X(_1242_));
 sky130_fd_sc_hd__a221o_1 _3868_ (.A1(\gpio_configure[4][1] ),
    .A2(_0904_),
    .B1(_0936_),
    .B2(net72),
    .C1(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__a221o_1 _3869_ (.A1(\gpio_configure[34][9] ),
    .A2(_1030_),
    .B1(_1032_),
    .B2(\gpio_configure[37][9] ),
    .C1(_1234_),
    .X(_1244_));
 sky130_fd_sc_hd__a32o_1 _3870_ (.A1(\gpio_configure[35][9] ),
    .A2(net381),
    .A3(net371),
    .B1(_0899_),
    .B2(\gpio_configure[35][1] ),
    .X(_1245_));
 sky130_fd_sc_hd__a221o_1 _3871_ (.A1(net47),
    .A2(_0935_),
    .B1(_1038_),
    .B2(\gpio_configure[36][9] ),
    .C1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__a311o_2 _3872_ (.A1(\gpio_configure[36][1] ),
    .A2(net387),
    .A3(net380),
    .B1(_1244_),
    .C1(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__a2111o_4 _3873_ (.A1(\gpio_configure[33][1] ),
    .A2(_0902_),
    .B1(_1241_),
    .C1(_1243_),
    .D1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__a31o_2 _3874_ (.A1(\gpio_configure[0][1] ),
    .A2(net383),
    .A3(net373),
    .B1(_0979_),
    .X(_1249_));
 sky130_fd_sc_hd__a31o_1 _3875_ (.A1(net286),
    .A2(net403),
    .A3(net373),
    .B1(_1236_),
    .X(_1250_));
 sky130_fd_sc_hd__a31o_4 _3876_ (.A1(\gpio_configure[3][9] ),
    .A2(net378),
    .A3(net370),
    .B1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__a32o_1 _3877_ (.A1(\gpio_configure[9][9] ),
    .A2(net378),
    .A3(net376),
    .B1(_0926_),
    .B2(\gpio_configure[1][1] ),
    .X(_1252_));
 sky130_fd_sc_hd__a221o_1 _3878_ (.A1(\gpio_configure[11][9] ),
    .A2(_1026_),
    .B1(_1037_),
    .B2(\gpio_configure[5][9] ),
    .C1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__nor4_4 _3879_ (.A(_1248_),
    .B(_1249_),
    .C(_1251_),
    .D(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__a22o_1 _3880_ (.A1(\gpio_configure[12][1] ),
    .A2(_0881_),
    .B1(_1036_),
    .B2(\gpio_configure[13][9] ),
    .X(_1255_));
 sky130_fd_sc_hd__a31o_1 _3881_ (.A1(\gpio_configure[25][9] ),
    .A2(net358),
    .A3(net375),
    .B1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a32o_1 _3882_ (.A1(\gpio_configure[9][1] ),
    .A2(net391),
    .A3(net403),
    .B1(_1034_),
    .B2(\gpio_configure[12][9] ),
    .X(_1257_));
 sky130_fd_sc_hd__a41o_1 _3883_ (.A1(\gpio_configure[14][9] ),
    .A2(net391),
    .A3(net420),
    .A4(net411),
    .B1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__a221o_1 _3884_ (.A1(\gpio_configure[31][1] ),
    .A2(_0912_),
    .B1(_1039_),
    .B2(\gpio_configure[10][9] ),
    .C1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a32o_1 _3885_ (.A1(\gpio_configure[14][1] ),
    .A2(net392),
    .A3(net388),
    .B1(_0909_),
    .B2(\gpio_configure[28][1] ),
    .X(_1260_));
 sky130_fd_sc_hd__a221o_1 _3886_ (.A1(\gpio_configure[25][1] ),
    .A2(_0918_),
    .B1(_1051_),
    .B2(\gpio_configure[22][9] ),
    .C1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__a221o_2 _3887_ (.A1(\gpio_configure[15][9] ),
    .A2(_1048_),
    .B1(_1050_),
    .B2(\gpio_configure[17][9] ),
    .C1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__a2111oi_4 _3888_ (.A1(\gpio_configure[29][1] ),
    .A2(_0933_),
    .B1(_1256_),
    .C1(_1259_),
    .D1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__a32o_4 _3889_ (.A1(net296),
    .A2(net383),
    .A3(_0883_),
    .B1(_0944_),
    .B2(\gpio_configure[6][1] ),
    .X(_1264_));
 sky130_fd_sc_hd__a32o_1 _3890_ (.A1(\gpio_configure[31][9] ),
    .A2(net356),
    .A3(net374),
    .B1(_0908_),
    .B2(\gpio_configure[19][1] ),
    .X(_1265_));
 sky130_fd_sc_hd__a221o_1 _3891_ (.A1(\gpio_configure[21][9] ),
    .A2(_1046_),
    .B1(_1047_),
    .B2(\gpio_configure[2][9] ),
    .C1(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__a31o_1 _3892_ (.A1(\gpio_configure[10][1] ),
    .A2(net390),
    .A3(_0890_),
    .B1(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__a32o_1 _3893_ (.A1(\gpio_configure[32][1] ),
    .A2(net384),
    .A3(net355),
    .B1(_0948_),
    .B2(\gpio_configure[23][1] ),
    .X(_1268_));
 sky130_fd_sc_hd__a32o_2 _3894_ (.A1(\gpio_configure[27][9] ),
    .A2(net356),
    .A3(net371),
    .B1(_1041_),
    .B2(\gpio_configure[18][9] ),
    .X(_1269_));
 sky130_fd_sc_hd__a221o_1 _3895_ (.A1(\gpio_configure[24][1] ),
    .A2(_0877_),
    .B1(_0913_),
    .B2(\gpio_configure[22][1] ),
    .C1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__a2111o_1 _3896_ (.A1(\gpio_configure[18][1] ),
    .A2(_0920_),
    .B1(_1237_),
    .C1(_1268_),
    .D1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a2111o_1 _3897_ (.A1(\gpio_configure[4][9] ),
    .A2(_1024_),
    .B1(_1264_),
    .C1(_1267_),
    .D1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__a32o_1 _3898_ (.A1(\gpio_configure[19][9] ),
    .A2(net358),
    .A3(net371),
    .B1(_1025_),
    .B2(\gpio_configure[32][9] ),
    .X(_1273_));
 sky130_fd_sc_hd__a221o_1 _3899_ (.A1(\gpio_configure[26][1] ),
    .A2(_0952_),
    .B1(_1052_),
    .B2(\gpio_configure[28][9] ),
    .C1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a22o_1 _3900_ (.A1(\gpio_configure[26][9] ),
    .A2(_1027_),
    .B1(_1053_),
    .B2(\gpio_configure[30][9] ),
    .X(_1275_));
 sky130_fd_sc_hd__a31o_1 _3901_ (.A1(\gpio_configure[23][9] ),
    .A2(net357),
    .A3(_0931_),
    .B1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a32o_1 _3902_ (.A1(serial_bb_enable),
    .A2(_0940_),
    .A3(net371),
    .B1(_1031_),
    .B2(\gpio_configure[7][9] ),
    .X(_1277_));
 sky130_fd_sc_hd__a221o_1 _3903_ (.A1(\gpio_configure[21][1] ),
    .A2(_0861_),
    .B1(_0903_),
    .B2(\gpio_configure[20][1] ),
    .C1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__a2111o_1 _3904_ (.A1(\gpio_configure[24][9] ),
    .A2(_1040_),
    .B1(_1274_),
    .C1(_1276_),
    .D1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__a32o_1 _3905_ (.A1(\gpio_configure[33][9] ),
    .A2(net355),
    .A3(net375),
    .B1(_0927_),
    .B2(\gpio_configure[17][1] ),
    .X(_1280_));
 sky130_fd_sc_hd__a221o_1 _3906_ (.A1(net15),
    .A2(_0886_),
    .B1(_1044_),
    .B2(\gpio_configure[6][9] ),
    .C1(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__a32o_1 _3907_ (.A1(\gpio_configure[16][1] ),
    .A2(net390),
    .A3(net383),
    .B1(_1042_),
    .B2(\gpio_configure[16][9] ),
    .X(_1282_));
 sky130_fd_sc_hd__a221o_4 _3908_ (.A1(net267),
    .A2(_0997_),
    .B1(_1060_),
    .B2(net261),
    .C1(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__a32o_1 _3909_ (.A1(\gpio_configure[1][9] ),
    .A2(net375),
    .A3(net373),
    .B1(_0865_),
    .B2(\gpio_configure[15][1] ),
    .X(_1284_));
 sky130_fd_sc_hd__a221o_1 _3910_ (.A1(\gpio_configure[27][1] ),
    .A2(_0880_),
    .B1(_1029_),
    .B2(\gpio_configure[29][9] ),
    .C1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__a32o_2 _3911_ (.A1(net294),
    .A2(net385),
    .A3(net383),
    .B1(_1035_),
    .B2(\gpio_configure[0][9] ),
    .X(_1286_));
 sky130_fd_sc_hd__a221o_1 _3912_ (.A1(\gpio_configure[8][1] ),
    .A2(_0928_),
    .B1(_0945_),
    .B2(\gpio_configure[2][1] ),
    .C1(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__nor4_1 _3913_ (.A(_1281_),
    .B(_1283_),
    .C(_1285_),
    .D(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__a32o_1 _3914_ (.A1(\gpio_configure[34][1] ),
    .A2(net382),
    .A3(_0890_),
    .B1(_0884_),
    .B2(\gpio_configure[37][1] ),
    .X(_1289_));
 sky130_fd_sc_hd__a32o_4 _3915_ (.A1(net35),
    .A2(net387),
    .A3(net386),
    .B1(_0939_),
    .B2(\gpio_configure[5][1] ),
    .X(_1290_));
 sky130_fd_sc_hd__a221o_1 _3916_ (.A1(\gpio_configure[11][1] ),
    .A2(_0901_),
    .B1(_0938_),
    .B2(\gpio_configure[13][1] ),
    .C1(_1235_),
    .X(_1291_));
 sky130_fd_sc_hd__a221o_4 _3917_ (.A1(net12),
    .A2(_0873_),
    .B1(_0925_),
    .B2(net280),
    .C1(_1240_),
    .X(_1292_));
 sky130_fd_sc_hd__a311o_1 _3918_ (.A1(net96),
    .A2(net389),
    .A3(net373),
    .B1(_1291_),
    .C1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a2111o_4 _3919_ (.A1(\gpio_configure[3][1] ),
    .A2(_0895_),
    .B1(_1289_),
    .C1(_1290_),
    .D1(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__a221oi_4 _3920_ (.A1(\gpio_configure[30][1] ),
    .A2(_0921_),
    .B1(_1049_),
    .B2(\clk2_output_dest[0] ),
    .C1(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__and4bb_1 _3921_ (.A_N(_1272_),
    .B_N(_1279_),
    .C(_1288_),
    .D(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__nand3_4 _3922_ (.A(_1254_),
    .B(net344),
    .C(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__mux2_1 _3923_ (.A0(\hkspi.ldata[0] ),
    .A1(_1297_),
    .S(net509),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(_1298_),
    .A1(net3800),
    .S(_0954_),
    .X(_0385_));
 sky130_fd_sc_hd__and4_1 _3925_ (.A(\gpio_configure[29][8] ),
    .B(net414),
    .C(net355),
    .D(net409),
    .X(_1299_));
 sky130_fd_sc_hd__a32o_1 _3926_ (.A1(\gpio_configure[25][8] ),
    .A2(net359),
    .A3(net375),
    .B1(_0877_),
    .B2(\gpio_configure[24][0] ),
    .X(_1300_));
 sky130_fd_sc_hd__and4_2 _3927_ (.A(irq_1_inputsrc),
    .B(net417),
    .C(net415),
    .D(net372),
    .X(_1301_));
 sky130_fd_sc_hd__nor3_2 _3928_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .C(reset_reg),
    .Y(_1302_));
 sky130_fd_sc_hd__inv_2 _3929_ (.A(_1302_),
    .Y(net299));
 sky130_fd_sc_hd__and4_1 _3930_ (.A(net20),
    .B(net417),
    .C(net413),
    .D(net385),
    .X(_1303_));
 sky130_fd_sc_hd__and4_1 _3931_ (.A(\gpio_configure[18][8] ),
    .B(net357),
    .C(net410),
    .D(net407),
    .X(_1304_));
 sky130_fd_sc_hd__a32o_1 _3932_ (.A1(\gpio_configure[33][8] ),
    .A2(net354),
    .A3(net376),
    .B1(_0997_),
    .B2(net266),
    .X(_1305_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(net389),
    .B(net906),
    .Y(_1306_));
 sky130_fd_sc_hd__a22o_1 _3934_ (.A1(net36),
    .A2(_0935_),
    .B1(_1030_),
    .B2(\gpio_configure[34][8] ),
    .X(_1307_));
 sky130_fd_sc_hd__a32o_1 _3935_ (.A1(net52),
    .A2(net388),
    .A3(net381),
    .B1(_0899_),
    .B2(\gpio_configure[35][0] ),
    .X(_1308_));
 sky130_fd_sc_hd__a32o_1 _3936_ (.A1(\gpio_configure[33][0] ),
    .A2(net381),
    .A3(net403),
    .B1(_1032_),
    .B2(\gpio_configure[37][8] ),
    .X(_1309_));
 sky130_fd_sc_hd__a31o_1 _3937_ (.A1(\gpio_configure[4][0] ),
    .A2(net387),
    .A3(net379),
    .B1(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__a41o_1 _3938_ (.A1(net258),
    .A2(net420),
    .A3(_0868_),
    .A4(net411),
    .B1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__a32o_1 _3939_ (.A1(\gpio_configure[35][8] ),
    .A2(net381),
    .A3(net371),
    .B1(_1038_),
    .B2(\gpio_configure[36][8] ),
    .X(_1312_));
 sky130_fd_sc_hd__a32o_1 _3940_ (.A1(\gpio_configure[36][0] ),
    .A2(_0867_),
    .A3(net380),
    .B1(_0884_),
    .B2(\gpio_configure[37][0] ),
    .X(_1313_));
 sky130_fd_sc_hd__a221o_1 _3941_ (.A1(\gpio_configure[34][0] ),
    .A2(_0891_),
    .B1(_0932_),
    .B2(net43),
    .C1(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__a2111o_1 _3942_ (.A1(net61),
    .A2(_1016_),
    .B1(_1311_),
    .C1(_1312_),
    .D1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__a2111o_4 _3943_ (.A1(net71),
    .A2(_0936_),
    .B1(_1307_),
    .C1(_1308_),
    .D1(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__o311a_2 _3944_ (.A1(\hkspi.pass_thru_mgmt_delay ),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .A3(reset_reg),
    .B1(net386),
    .C1(net374),
    .X(_1317_));
 sky130_fd_sc_hd__a221o_1 _3945_ (.A1(\gpio_configure[7][0] ),
    .A2(_0914_),
    .B1(_1045_),
    .B2(\gpio_configure[8][8] ),
    .C1(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__a32o_1 _3946_ (.A1(\gpio_configure[2][0] ),
    .A2(_0890_),
    .A3(net378),
    .B1(_1044_),
    .B2(\gpio_configure[6][8] ),
    .X(_1319_));
 sky130_fd_sc_hd__a32o_1 _3947_ (.A1(net276),
    .A2(net386),
    .A3(net376),
    .B1(_0925_),
    .B2(net269),
    .X(_1320_));
 sky130_fd_sc_hd__a221o_2 _3948_ (.A1(net386),
    .A2(net370),
    .B1(_1239_),
    .B2(net265),
    .C1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__a31o_1 _3949_ (.A1(\gpio_configure[7][8] ),
    .A2(net378),
    .A3(net374),
    .B1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a311o_1 _3950_ (.A1(\gpio_configure[10][0] ),
    .A2(net390),
    .A3(_0890_),
    .B1(_1319_),
    .C1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a32o_1 _3951_ (.A1(\gpio_configure[17][8] ),
    .A2(net391),
    .A3(net375),
    .B1(_1039_),
    .B2(\gpio_configure[10][8] ),
    .X(_1324_));
 sky130_fd_sc_hd__a31o_1 _3952_ (.A1(\gpio_configure[14][0] ),
    .A2(net392),
    .A3(net388),
    .B1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__a32o_1 _3953_ (.A1(\gpio_configure[15][8] ),
    .A2(net392),
    .A3(net374),
    .B1(_0889_),
    .B2(\gpio_configure[9][0] ),
    .X(_1326_));
 sky130_fd_sc_hd__a221o_1 _3954_ (.A1(\gpio_configure[29][0] ),
    .A2(_0933_),
    .B1(_1028_),
    .B2(\gpio_configure[20][8] ),
    .C1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__a22o_1 _3955_ (.A1(\gpio_configure[31][0] ),
    .A2(_0912_),
    .B1(_0938_),
    .B2(\gpio_configure[13][0] ),
    .X(_1328_));
 sky130_fd_sc_hd__a32o_1 _3956_ (.A1(net98),
    .A2(net388),
    .A3(net373),
    .B1(_1034_),
    .B2(\gpio_configure[12][8] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _3957_ (.A1(\gpio_configure[25][0] ),
    .A2(_0918_),
    .B1(_1051_),
    .B2(\gpio_configure[22][8] ),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a31o_1 _3958_ (.A1(\gpio_configure[30][0] ),
    .A2(net388),
    .A3(_0879_),
    .B1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__a311o_1 _3959_ (.A1(\gpio_configure[28][0] ),
    .A2(_0867_),
    .A3(_0879_),
    .B1(_1328_),
    .C1(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__a2111o_4 _3960_ (.A1(\gpio_configure[14][8] ),
    .A2(_1043_),
    .B1(_1325_),
    .C1(_1327_),
    .D1(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nor4_1 _3961_ (.A(_1316_),
    .B(_1318_),
    .C(_1323_),
    .D(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__a32o_1 _3962_ (.A1(\gpio_configure[1][8] ),
    .A2(net375),
    .A3(net372),
    .B1(_0865_),
    .B2(\gpio_configure[15][0] ),
    .X(_1335_));
 sky130_fd_sc_hd__a32o_1 _3963_ (.A1(hkspi_disable),
    .A2(net382),
    .A3(net375),
    .B1(_1047_),
    .B2(\gpio_configure[2][8] ),
    .X(_1336_));
 sky130_fd_sc_hd__a221o_1 _3964_ (.A1(\gpio_configure[19][0] ),
    .A2(_0908_),
    .B1(_0920_),
    .B2(\gpio_configure[18][0] ),
    .C1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a31o_2 _3965_ (.A1(\gpio_configure[22][0] ),
    .A2(net388),
    .A3(net358),
    .B1(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__a32o_1 _3966_ (.A1(net293),
    .A2(net385),
    .A3(net383),
    .B1(_0944_),
    .B2(\gpio_configure[6][0] ),
    .X(_1339_));
 sky130_fd_sc_hd__a31o_1 _3967_ (.A1(\gpio_configure[23][8] ),
    .A2(net357),
    .A3(net374),
    .B1(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__a221o_1 _3968_ (.A1(\gpio_configure[0][0] ),
    .A2(_0941_),
    .B1(_1040_),
    .B2(\gpio_configure[24][8] ),
    .C1(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__a32o_1 _3969_ (.A1(\gpio_configure[9][8] ),
    .A2(net379),
    .A3(net375),
    .B1(_1037_),
    .B2(\gpio_configure[5][8] ),
    .X(_1342_));
 sky130_fd_sc_hd__a2111o_1 _3970_ (.A1(\gpio_configure[27][0] ),
    .A2(_0880_),
    .B1(_1342_),
    .C1(_1304_),
    .D1(_1341_),
    .X(_1343_));
 sky130_fd_sc_hd__a2111o_1 _3971_ (.A1(\gpio_configure[28][8] ),
    .A2(_1052_),
    .B1(_1335_),
    .C1(_1338_),
    .D1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__a32o_4 _3972_ (.A1(\gpio_configure[31][8] ),
    .A2(net354),
    .A3(net374),
    .B1(_1025_),
    .B2(\gpio_configure[32][8] ),
    .X(_1345_));
 sky130_fd_sc_hd__a31o_1 _3973_ (.A1(\gpio_configure[32][0] ),
    .A2(net383),
    .A3(net355),
    .B1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a22o_1 _3974_ (.A1(\gpio_configure[0][8] ),
    .A2(_1035_),
    .B1(_1042_),
    .B2(\gpio_configure[16][8] ),
    .X(_1347_));
 sky130_fd_sc_hd__a221o_1 _3975_ (.A1(\gpio_configure[16][0] ),
    .A2(_0876_),
    .B1(_1024_),
    .B2(\gpio_configure[4][8] ),
    .C1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a311o_1 _3976_ (.A1(serial_busy),
    .A2(net372),
    .A3(net370),
    .B1(_1346_),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a32o_2 _3977_ (.A1(net285),
    .A2(net403),
    .A3(net373),
    .B1(_1060_),
    .B2(net260),
    .X(_1350_));
 sky130_fd_sc_hd__a32o_1 _3978_ (.A1(\gpio_configure[19][8] ),
    .A2(net357),
    .A3(net370),
    .B1(_1027_),
    .B2(\gpio_configure[26][8] ),
    .X(_1351_));
 sky130_fd_sc_hd__a2111o_1 _3979_ (.A1(\gpio_configure[20][0] ),
    .A2(_0903_),
    .B1(_1305_),
    .C1(_1350_),
    .D1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__a221o_1 _3980_ (.A1(\gpio_configure[11][8] ),
    .A2(_1026_),
    .B1(_1046_),
    .B2(\gpio_configure[21][8] ),
    .C1(_1301_),
    .X(_1353_));
 sky130_fd_sc_hd__a32o_1 _3981_ (.A1(\gpio_configure[27][8] ),
    .A2(net355),
    .A3(net370),
    .B1(\gpio_configure[21][0] ),
    .B2(_0861_),
    .X(_1354_));
 sky130_fd_sc_hd__a32o_1 _3982_ (.A1(net295),
    .A2(net384),
    .A3(_0883_),
    .B1(_0952_),
    .B2(\gpio_configure[26][0] ),
    .X(_1355_));
 sky130_fd_sc_hd__a2111o_1 _3983_ (.A1(\gpio_configure[8][0] ),
    .A2(_0928_),
    .B1(_1353_),
    .C1(_1354_),
    .D1(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__a22o_1 _3984_ (.A1(net4),
    .A2(_0886_),
    .B1(_1053_),
    .B2(\gpio_configure[30][8] ),
    .X(_1357_));
 sky130_fd_sc_hd__a31o_1 _3985_ (.A1(irq_spi),
    .A2(net389),
    .A3(net385),
    .B1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__a221o_1 _3986_ (.A1(\gpio_configure[17][0] ),
    .A2(_0927_),
    .B1(_0948_),
    .B2(\gpio_configure[23][0] ),
    .C1(_1299_),
    .X(_1359_));
 sky130_fd_sc_hd__a2111o_1 _3987_ (.A1(\gpio_configure[1][0] ),
    .A2(_0926_),
    .B1(_1356_),
    .C1(_1358_),
    .D1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__nor4_1 _3988_ (.A(_1344_),
    .B(_1349_),
    .C(_1352_),
    .D(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__a41o_1 _3989_ (.A1(net93),
    .A2(net417),
    .A3(net416),
    .A4(net385),
    .B1(_1303_),
    .X(_1362_));
 sky130_fd_sc_hd__a221o_2 _3990_ (.A1(net11),
    .A2(_0873_),
    .B1(_0895_),
    .B2(\gpio_configure[3][0] ),
    .C1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__a32o_1 _3991_ (.A1(\gpio_configure[12][0] ),
    .A2(net392),
    .A3(_0867_),
    .B1(_1036_),
    .B2(\gpio_configure[13][8] ),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_4 _3992_ (.A1(\gpio_configure[11][0] ),
    .A2(_0901_),
    .B1(_1049_),
    .B2(trap_output_dest),
    .C1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__a32o_1 _3993_ (.A1(\gpio_configure[3][8] ),
    .A2(net377),
    .A3(net370),
    .B1(_0939_),
    .B2(\gpio_configure[5][0] ),
    .X(_1366_));
 sky130_fd_sc_hd__a2111oi_4 _3994_ (.A1(net34),
    .A2(_0869_),
    .B1(_1363_),
    .C1(_1365_),
    .D1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__and4b_4 _3995_ (.A_N(_1300_),
    .B(_1334_),
    .C(_1361_),
    .D(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__nor2_1 _3996_ (.A(_0954_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a22o_1 _3997_ (.A1(net3802),
    .A2(_0954_),
    .B1(_1369_),
    .B2(net509),
    .X(_0384_));
 sky130_fd_sc_hd__nor2_1 _3998_ (.A(\hkspi.state[3] ),
    .B(\hkspi.state[2] ),
    .Y(_1370_));
 sky130_fd_sc_hd__o31a_2 _3999_ (.A1(\hkspi.state[0] ),
    .A2(\hkspi.state[3] ),
    .A3(\hkspi.state[2] ),
    .B1(\hkspi.count[0] ),
    .X(_1371_));
 sky130_fd_sc_hd__a21oi_1 _4000_ (.A1(net3908),
    .A2(_1371_),
    .B1(\hkspi.count[2] ),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_2 _4001_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .Y(_1373_));
 sky130_fd_sc_hd__and3_1 _4002_ (.A(\hkspi.count[2] ),
    .B(net3908),
    .C(_1371_),
    .X(_1374_));
 sky130_fd_sc_hd__nor2_1 _4003_ (.A(_1372_),
    .B(_1374_),
    .Y(_0100_));
 sky130_fd_sc_hd__xor2_1 _4004_ (.A(net3890),
    .B(_1371_),
    .X(_0099_));
 sky130_fd_sc_hd__nor4_1 _4005_ (.A(net3898),
    .B(\hkspi.state[0] ),
    .C(net3899),
    .D(\hkspi.state[2] ),
    .Y(_1375_));
 sky130_fd_sc_hd__nor2_1 _4006_ (.A(_1371_),
    .B(_1375_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_4 _4007_ (.A(_0819_),
    .B(net525),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _4008_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[0] ),
    .Y(_1377_));
 sky130_fd_sc_hd__and3_2 _4009_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .X(_1378_));
 sky130_fd_sc_hd__nand3_1 _4010_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .Y(_1379_));
 sky130_fd_sc_hd__and4_2 _4011_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .D(\hkspi.state[2] ),
    .X(_1380_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(\hkspi.fixed[2] ),
    .B(\hkspi.fixed[1] ),
    .Y(_1381_));
 sky130_fd_sc_hd__o311ai_4 _4013_ (.A1(\hkspi.fixed[2] ),
    .A2(\hkspi.fixed[1] ),
    .A3(_0818_),
    .B1(_0819_),
    .C1(_1380_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_4 _4014_ (.A(_1376_),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__and4_2 _4015_ (.A(\hkspi.addr[3] ),
    .B(\hkspi.addr[2] ),
    .C(\hkspi.addr[1] ),
    .D(\hkspi.addr[0] ),
    .X(_1384_));
 sky130_fd_sc_hd__and3_1 _4016_ (.A(\hkspi.addr[5] ),
    .B(\hkspi.addr[4] ),
    .C(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(\hkspi.addr[6] ),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__a41o_1 _4018_ (.A1(\hkspi.addr[6] ),
    .A2(\hkspi.addr[5] ),
    .A3(\hkspi.addr[4] ),
    .A4(_1384_),
    .B1(_0834_),
    .X(_1387_));
 sky130_fd_sc_hd__o2bb2a_1 _4019_ (.A1_N(_1376_),
    .A2_N(_1382_),
    .B1(_0833_),
    .B2(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__o2bb2a_1 _4020_ (.A1_N(_1388_),
    .A2_N(_1387_),
    .B1(_1383_),
    .B2(net2846),
    .X(_0097_));
 sky130_fd_sc_hd__a31o_1 _4021_ (.A1(\hkspi.addr[5] ),
    .A2(\hkspi.addr[4] ),
    .A3(_1384_),
    .B1(\hkspi.addr[6] ),
    .X(_1389_));
 sky130_fd_sc_hd__o211a_1 _4022_ (.A1(_1382_),
    .A2(_1386_),
    .B1(_1389_),
    .C1(_1376_),
    .X(_1390_));
 sky130_fd_sc_hd__a21o_1 _4023_ (.A1(net2449),
    .A2(net525),
    .B1(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__o21a_1 _4024_ (.A1(net3848),
    .A2(_1383_),
    .B1(_1391_),
    .X(_0096_));
 sky130_fd_sc_hd__nor2_1 _4025_ (.A(net525),
    .B(_1384_),
    .Y(_1392_));
 sky130_fd_sc_hd__a21oi_1 _4026_ (.A1(\hkspi.addr[4] ),
    .A2(_1384_),
    .B1(\hkspi.addr[5] ),
    .Y(_1393_));
 sky130_fd_sc_hd__o31ai_1 _4027_ (.A1(net525),
    .A2(_1385_),
    .A3(_1393_),
    .B1(_0830_),
    .Y(_1394_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(net2449),
    .A1(_1394_),
    .S(_1383_),
    .X(_0095_));
 sky130_fd_sc_hd__a31o_1 _4029_ (.A1(\hkspi.addr[2] ),
    .A2(\hkspi.addr[1] ),
    .A3(\hkspi.addr[0] ),
    .B1(net525),
    .X(_1395_));
 sky130_fd_sc_hd__a21oi_1 _4030_ (.A1(\hkspi.addr[4] ),
    .A2(_1384_),
    .B1(net525),
    .Y(_1396_));
 sky130_fd_sc_hd__a41o_1 _4031_ (.A1(\hkspi.addr[3] ),
    .A2(\hkspi.addr[2] ),
    .A3(\hkspi.addr[1] ),
    .A4(\hkspi.addr[0] ),
    .B1(\hkspi.addr[4] ),
    .X(_1397_));
 sky130_fd_sc_hd__a22o_1 _4032_ (.A1(\hkspi.addr[3] ),
    .A2(\hkspi.state[3] ),
    .B1(_1396_),
    .B2(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(net3882),
    .A1(_1398_),
    .S(_1383_),
    .X(_0094_));
 sky130_fd_sc_hd__a31o_1 _4034_ (.A1(\hkspi.addr[2] ),
    .A2(\hkspi.addr[1] ),
    .A3(\hkspi.addr[0] ),
    .B1(\hkspi.addr[3] ),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _4035_ (.A1(\hkspi.addr[2] ),
    .A2(net525),
    .B1(_1392_),
    .B2(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(net3881),
    .A1(_1400_),
    .S(_1383_),
    .X(_0093_));
 sky130_fd_sc_hd__a21oi_1 _4037_ (.A1(\hkspi.addr[1] ),
    .A2(\hkspi.addr[0] ),
    .B1(\hkspi.addr[2] ),
    .Y(_1401_));
 sky130_fd_sc_hd__a2bb2o_1 _4038_ (.A1_N(_1401_),
    .A2_N(_1395_),
    .B1(net525),
    .B2(\hkspi.addr[1] ),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(net3885),
    .A1(_1402_),
    .S(_1383_),
    .X(_0092_));
 sky130_fd_sc_hd__and4_1 _4040_ (.A(_1383_),
    .B(\hkspi.addr[0] ),
    .C(\hkspi.addr[1] ),
    .D(_1376_),
    .X(_1403_));
 sky130_fd_sc_hd__a22oi_1 _4041_ (.A1(net3904),
    .A2(_1376_),
    .B1(_1383_),
    .B2(net3892),
    .Y(_1404_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(_1403_),
    .B(_1404_),
    .Y(_0091_));
 sky130_fd_sc_hd__o211a_1 _4043_ (.A1(_0816_),
    .A2(net525),
    .B1(_0848_),
    .C1(_1383_),
    .X(_1405_));
 sky130_fd_sc_hd__a31o_1 _4044_ (.A1(net3892),
    .A2(_1376_),
    .A3(_1382_),
    .B1(_1405_),
    .X(_0090_));
 sky130_fd_sc_hd__and3_1 _4045_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[0] ),
    .C(\hkspi.state[0] ),
    .X(_1406_));
 sky130_fd_sc_hd__and4_1 _4046_ (.A(\hkspi.count[2] ),
    .B(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .D(\hkspi.state[0] ),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(\hkspi.pass_thru_user_delay ),
    .A1(net3846),
    .S(_1407_),
    .X(_0089_));
 sky130_fd_sc_hd__a41o_1 _4048_ (.A1(_0819_),
    .A2(_1370_),
    .A3(_0820_),
    .A4(net3849),
    .B1(net3871),
    .X(_0088_));
 sky130_fd_sc_hd__and4b_1 _4049_ (.A_N(\hkspi.count[0] ),
    .B(\hkspi.state[0] ),
    .C(\hkspi.count[2] ),
    .D(\hkspi.count[1] ),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(net3888),
    .A1(net3872),
    .S(_1408_),
    .X(_0087_));
 sky130_fd_sc_hd__a31o_1 _4051_ (.A1(_1370_),
    .A2(_0819_),
    .A3(net3860),
    .B1(net3874),
    .X(_0086_));
 sky130_fd_sc_hd__o31a_1 _4052_ (.A1(\hkspi.state[0] ),
    .A2(\hkspi.state[3] ),
    .A3(\hkspi.state[2] ),
    .B1(\hkspi.readmode ),
    .X(_1409_));
 sky130_fd_sc_hd__o221a_1 _4053_ (.A1(_1370_),
    .A2(_1378_),
    .B1(_1409_),
    .B2(net3905),
    .C1(_0819_),
    .X(_0085_));
 sky130_fd_sc_hd__o41a_1 _4054_ (.A1(\hkspi.count[2] ),
    .A2(\hkspi.count[1] ),
    .A3(\hkspi.count[0] ),
    .A4(_0819_),
    .B1(net3886),
    .X(_1410_));
 sky130_fd_sc_hd__a31o_1 _4055_ (.A1(net58),
    .A2(\hkspi.state[0] ),
    .A3(_0829_),
    .B1(_1410_),
    .X(_0084_));
 sky130_fd_sc_hd__and4bb_1 _4056_ (.A_N(\hkspi.count[2] ),
    .B_N(\hkspi.count[1] ),
    .C(\hkspi.count[0] ),
    .D(\hkspi.state[0] ),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(net3891),
    .A1(net58),
    .S(_1411_),
    .X(_0083_));
 sky130_fd_sc_hd__nor3b_4 _4058_ (.A(\hkspi.state[0] ),
    .B(\hkspi.state[3] ),
    .C_N(\hkspi.state[2] ),
    .Y(_1412_));
 sky130_fd_sc_hd__o211a_1 _4059_ (.A1(\hkspi.fixed[2] ),
    .A2(\hkspi.fixed[1] ),
    .B1(_1378_),
    .C1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__a31oi_4 _4060_ (.A1(\hkspi.state[0] ),
    .A2(_1373_),
    .A3(_1377_),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__a211o_2 _4061_ (.A1(\hkspi.state[0] ),
    .A2(_0829_),
    .B1(_1411_),
    .C1(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__nor2_1 _4062_ (.A(_0819_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__a21oi_1 _4063_ (.A1(_0818_),
    .A2(\hkspi.fixed[2] ),
    .B1(\hkspi.state[0] ),
    .Y(_1417_));
 sky130_fd_sc_hd__o32a_1 _4064_ (.A1(net3887),
    .A2(_1417_),
    .A3(_1415_),
    .B1(net3880),
    .B2(_1416_),
    .X(_0082_));
 sky130_fd_sc_hd__o22ai_1 _4065_ (.A1(_1415_),
    .A2(net3878),
    .B1(\hkspi.fixed[1] ),
    .B2(_1416_),
    .Y(_1418_));
 sky130_fd_sc_hd__o41ai_1 _4066_ (.A1(\hkspi.fixed[1] ),
    .A2(net3878),
    .A3(\hkspi.state[0] ),
    .A4(_1414_),
    .B1(_1418_),
    .Y(_0081_));
 sky130_fd_sc_hd__nor3_1 _4067_ (.A(\hkspi.fixed[0] ),
    .B(\hkspi.state[0] ),
    .C(_1414_),
    .Y(_1419_));
 sky130_fd_sc_hd__a221o_1 _4068_ (.A1(net3878),
    .A2(_1415_),
    .B1(_1416_),
    .B2(net58),
    .C1(_1419_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(net2097),
    .A1(net2283),
    .S(net507),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4070_ (.A0(net2283),
    .A1(net2014),
    .S(net507),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(net2014),
    .A1(net2692),
    .S(net507),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(net2692),
    .A1(net2024),
    .S(net507),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(net2024),
    .A1(net2030),
    .S(net507),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(net2030),
    .A1(net2345),
    .S(net507),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(net2345),
    .A1(net58),
    .S(net507),
    .X(_0073_));
 sky130_fd_sc_hd__and4b_1 _4076_ (.A_N(\hkspi.count[1] ),
    .B(net58),
    .C(_1406_),
    .D(\hkspi.count[2] ),
    .X(_1420_));
 sky130_fd_sc_hd__o21bai_1 _4077_ (.A1(_0817_),
    .A2(_1406_),
    .B1_N(_1420_),
    .Y(_0072_));
 sky130_fd_sc_hd__nor3_2 _4078_ (.A(net3622),
    .B(net2388),
    .C(net67),
    .Y(_1421_));
 sky130_fd_sc_hd__and2_1 _4079_ (.A(net563),
    .B(net366),
    .X(_0021_));
 sky130_fd_sc_hd__a211o_1 _4080_ (.A1(\hkspi.count[0] ),
    .A2(\hkspi.pre_pass_thru_mgmt ),
    .B1(_0819_),
    .C1(_1373_),
    .X(_1422_));
 sky130_fd_sc_hd__a22o_1 _4081_ (.A1(net58),
    .A2(_1408_),
    .B1(_1422_),
    .B2(net3846),
    .X(_0071_));
 sky130_fd_sc_hd__o211a_1 _4082_ (.A1(\hkspi.writemode ),
    .A2(net3903),
    .B1(\hkspi.state[2] ),
    .C1(_1378_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_8 _4083_ (.A0(serial_clock_pre),
    .A1(serial_bb_clock),
    .S(serial_bb_enable),
    .X(net301));
 sky130_fd_sc_hd__o21a_2 _4084_ (.A1(\hkspi.rdstb ),
    .A2(\hkspi.wrstb ),
    .B1(net369),
    .X(_1423_));
 sky130_fd_sc_hd__o21ai_2 _4085_ (.A1(\hkspi.rdstb ),
    .A2(\hkspi.wrstb ),
    .B1(net369),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(net112),
    .B(net111),
    .Y(_1425_));
 sky130_fd_sc_hd__nor2_8 _4087_ (.A(net114),
    .B(net113),
    .Y(_1426_));
 sky130_fd_sc_hd__a211oi_4 _4088_ (.A1(net112),
    .A2(net111),
    .B1(net114),
    .C1(net113),
    .Y(_1427_));
 sky130_fd_sc_hd__and4bb_1 _4089_ (.A_N(net118),
    .B_N(net119),
    .C(net120),
    .D(net117),
    .X(_1428_));
 sky130_fd_sc_hd__nor4_1 _4090_ (.A(net101),
    .B(net100),
    .C(net103),
    .D(net102),
    .Y(_1429_));
 sky130_fd_sc_hd__nor4b_1 _4091_ (.A(net109),
    .B(net108),
    .C(net115),
    .D_N(net116),
    .Y(_1430_));
 sky130_fd_sc_hd__nor4_1 _4092_ (.A(net105),
    .B(net104),
    .C(net107),
    .D(net106),
    .Y(_1431_));
 sky130_fd_sc_hd__and4_1 _4093_ (.A(net131),
    .B(net169),
    .C(_1428_),
    .D(_1430_),
    .X(_1432_));
 sky130_fd_sc_hd__a211oi_1 _4094_ (.A1(net112),
    .A2(net111),
    .B1(net130),
    .C1(net129),
    .Y(_1433_));
 sky130_fd_sc_hd__and4_1 _4095_ (.A(_1426_),
    .B(_1429_),
    .C(_1431_),
    .D(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__and4bb_2 _4096_ (.A_N(net123),
    .B_N(net122),
    .C(_1432_),
    .D(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__a22o_1 _4097_ (.A1(net3834),
    .A2(_1423_),
    .B1(_1435_),
    .B2(net3875),
    .X(_0011_));
 sky130_fd_sc_hd__a32o_1 _4098_ (.A1(net3878),
    .A2(_1380_),
    .A3(_1381_),
    .B1(\hkspi.state[0] ),
    .B2(_1379_),
    .X(_0004_));
 sky130_fd_sc_hd__nor4_1 _4099_ (.A(net3894),
    .B(\xfer_count[2] ),
    .C(\xfer_count[3] ),
    .D(_0822_),
    .Y(_1436_));
 sky130_fd_sc_hd__o41a_1 _4100_ (.A1(\xfer_count[0] ),
    .A2(\xfer_count[2] ),
    .A3(\xfer_count[3] ),
    .A4(_0822_),
    .B1(\xfer_state[3] ),
    .X(_1437_));
 sky130_fd_sc_hd__and2b_4 _4101_ (.A_N(\pad_count_2[0] ),
    .B(\pad_count_2[1] ),
    .X(_1438_));
 sky130_fd_sc_hd__and2b_4 _4102_ (.A_N(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .X(_1439_));
 sky130_fd_sc_hd__and2b_4 _4103_ (.A_N(net514),
    .B(net515),
    .X(_1440_));
 sky130_fd_sc_hd__and4bb_4 _4104_ (.A_N(\pad_count_2[0] ),
    .B_N(net514),
    .C(net515),
    .D(\pad_count_2[1] ),
    .X(_1441_));
 sky130_fd_sc_hd__nand2_1 _4105_ (.A(_1439_),
    .B(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__nand4bb_4 _4106_ (.A_N(\xfer_count[1] ),
    .B_N(\xfer_count[0] ),
    .C(\xfer_count[2] ),
    .D(\xfer_count[3] ),
    .Y(_1443_));
 sky130_fd_sc_hd__nor2_1 _4107_ (.A(_1443_),
    .B(net301),
    .Y(_1444_));
 sky130_fd_sc_hd__a41o_1 _4108_ (.A1(net527),
    .A2(_1439_),
    .A3(_1441_),
    .A4(_1444_),
    .B1(_1437_),
    .X(_0017_));
 sky130_fd_sc_hd__a21o_1 _4109_ (.A1(\wbbd_state[8] ),
    .A2(_1423_),
    .B1(net3808),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_1 _4110_ (.A1(\wbbd_state[9] ),
    .A2(_1423_),
    .B1(net3809),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _4111_ (.A1(\wbbd_state[10] ),
    .A2(_1423_),
    .B1(net3805),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _4112_ (.A1(\xfer_state[0] ),
    .A2(_0825_),
    .B1(net3895),
    .B2(\xfer_state[3] ),
    .X(_0014_));
 sky130_fd_sc_hd__a31o_1 _4113_ (.A1(net3846),
    .A2(_1407_),
    .A3(_0817_),
    .B1(net3849),
    .X(_0005_));
 sky130_fd_sc_hd__nand2b_1 _4114_ (.A_N(_1435_),
    .B(net3875),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2b_1 _4115_ (.A_N(net3854),
    .B(_1445_),
    .Y(_0009_));
 sky130_fd_sc_hd__and2_4 _4116_ (.A(net527),
    .B(net301),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_2 _4117_ (.A(net527),
    .B(net301),
    .Y(_1447_));
 sky130_fd_sc_hd__a211o_1 _4118_ (.A1(_1443_),
    .A2(net527),
    .B1(net526),
    .C1(_1446_),
    .X(_0015_));
 sky130_fd_sc_hd__a32o_1 _4119_ (.A1(net527),
    .A2(_1444_),
    .A3(_1442_),
    .B1(serial_xfer),
    .B2(\xfer_state[0] ),
    .X(_0016_));
 sky130_fd_sc_hd__a31o_1 _4120_ (.A1(\hkspi.pre_pass_thru_mgmt ),
    .A2(\hkspi.state[0] ),
    .A3(_1378_),
    .B1(net3860),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(net3846),
    .B(\hkspi.pre_pass_thru_mgmt ),
    .Y(_1448_));
 sky130_fd_sc_hd__a32o_1 _4122_ (.A1(net3890),
    .A2(_1406_),
    .A3(_1448_),
    .B1(net3899),
    .B2(_1379_),
    .X(_0007_));
 sky130_fd_sc_hd__nand3_1 _4123_ (.A(\hkspi.fixed[0] ),
    .B(_1378_),
    .C(_1381_),
    .Y(_1449_));
 sky130_fd_sc_hd__a22o_1 _4124_ (.A1(net3899),
    .A2(_1378_),
    .B1(_1449_),
    .B2(net3902),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_2 _4125_ (.A0(net84),
    .A1(net67),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net247));
 sky130_fd_sc_hd__nor2_1 _4126_ (.A(\hkspi.pass_thru_mgmt_delay ),
    .B(net564),
    .Y(net248));
 sky130_fd_sc_hd__mux2_1 _4127_ (.A0(net83),
    .A1(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_mgmt ),
    .X(pad_flash_clk_prebuff));
 sky130_fd_sc_hd__nor2_1 _4128_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net564),
    .Y(net246));
 sky130_fd_sc_hd__nand2b_2 _4129_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net86),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(net250),
    .Y(net251));
 sky130_fd_sc_hd__nor2_2 _4131_ (.A(\hkspi.pass_thru_mgmt ),
    .B(net88),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _4132_ (.A(net253),
    .Y(net254));
 sky130_fd_sc_hd__mux2_2 _4133_ (.A0(net85),
    .A1(net58),
    .S(\hkspi.pass_thru_mgmt_delay ),
    .X(net249));
 sky130_fd_sc_hd__and2b_4 _4134_ (.A_N(\hkspi.pass_thru_mgmt_delay ),
    .B(net73),
    .X(net307));
 sky130_fd_sc_hd__and2b_4 _4135_ (.A_N(\hkspi.pass_thru_mgmt ),
    .B(net74),
    .X(net308));
 sky130_fd_sc_hd__nor2_1 _4136_ (.A(\hkspi.state[4] ),
    .B(\hkspi.state[1] ),
    .Y(_1450_));
 sky130_fd_sc_hd__o21a_1 _4137_ (.A1(\hkspi.state[2] ),
    .A2(_1450_),
    .B1(_0954_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_2 _4138_ (.A0(\mgmt_gpio_data[37] ),
    .A1(net91),
    .S(net76),
    .X(net239));
 sky130_fd_sc_hd__mux2_2 _4139_ (.A0(\mgmt_gpio_data[36] ),
    .A1(net89),
    .S(net76),
    .X(net238));
 sky130_fd_sc_hd__nand2_4 _4140_ (.A(net76),
    .B(net92),
    .Y(_1451_));
 sky130_fd_sc_hd__o21ai_4 _4141_ (.A1(\gpio_configure[37][3] ),
    .A2(net76),
    .B1(_1451_),
    .Y(net205));
 sky130_fd_sc_hd__nand2_4 _4142_ (.A(net76),
    .B(net90),
    .Y(_1452_));
 sky130_fd_sc_hd__o21ai_4 _4143_ (.A1(\gpio_configure[36][3] ),
    .A2(net76),
    .B1(_1452_),
    .Y(net204));
 sky130_fd_sc_hd__nand2_2 _4144_ (.A(net82),
    .B(net79),
    .Y(_1453_));
 sky130_fd_sc_hd__o21ai_4 _4145_ (.A1(\gpio_configure[35][3] ),
    .A2(net79),
    .B1(_1453_),
    .Y(net203));
 sky130_fd_sc_hd__mux2_8 _4146_ (.A0(\mgmt_gpio_data[32] ),
    .A1(net80),
    .S(net79),
    .X(net234));
 sky130_fd_sc_hd__mux2_8 _4147_ (.A0(\mgmt_gpio_data[33] ),
    .A1(net78),
    .S(net79),
    .X(net235));
 sky130_fd_sc_hd__mux2_8 _4148_ (.A0(\mgmt_gpio_data[35] ),
    .A1(net81),
    .S(net79),
    .X(net237));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(\mgmt_gpio_data[10] ),
    .A1(net58),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net214));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(\mgmt_gpio_data[9] ),
    .A1(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .S(\hkspi.pass_thru_user ),
    .X(mgmt_gpio_out_9_prebuff));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(\mgmt_gpio_data[8] ),
    .A1(net67),
    .S(\hkspi.pass_thru_user_delay ),
    .X(net245));
 sky130_fd_sc_hd__mux2_8 _4152_ (.A0(\mgmt_gpio_data[6] ),
    .A1(net77),
    .S(net94),
    .X(net243));
 sky130_fd_sc_hd__mux2_1 _4153_ (.A0(\mgmt_gpio_data[1] ),
    .A1(\hkspi.SDO ),
    .S(net369),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(_1454_),
    .A1(net38),
    .S(\hkspi.pass_thru_user ),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_2 _4155_ (.A0(_1455_),
    .A1(net74),
    .S(\hkspi.pass_thru_mgmt ),
    .X(net222));
 sky130_fd_sc_hd__mux2_4 _4156_ (.A0(\mgmt_gpio_data[0] ),
    .A1(net3),
    .S(net1),
    .X(net213));
 sky130_fd_sc_hd__o31ai_1 _4157_ (.A1(hkspi_disable),
    .A2(\gpio_configure[3][3] ),
    .A3(net67),
    .B1(\gpio_configure[1][3] ),
    .Y(_1456_));
 sky130_fd_sc_hd__o41a_2 _4158_ (.A1(hkspi_disable),
    .A2(\gpio_configure[3][3] ),
    .A3(net67),
    .A4(\hkspi.sdoenb ),
    .B1(_1456_),
    .X(net186));
 sky130_fd_sc_hd__nand2_4 _4159_ (.A(net1),
    .B(net2),
    .Y(_1457_));
 sky130_fd_sc_hd__o21ai_4 _4160_ (.A1(\gpio_configure[0][3] ),
    .A2(net1),
    .B1(_1457_),
    .Y(net175));
 sky130_fd_sc_hd__mux2_1 _4161_ (.A0(\mgmt_gpio_data[15] ),
    .A1(clknet_1_1__leaf_user_clock),
    .S(\clk2_output_dest[0] ),
    .X(mgmt_gpio_out_15_prebuff));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(\mgmt_gpio_data[14] ),
    .A1(clknet_4_13__leaf_wb_clk_i),
    .S(\clk1_output_dest[0] ),
    .X(mgmt_gpio_out_14_prebuff));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(\mgmt_gpio_data[31] ),
    .A1(clknet_1_0__leaf_user_clock),
    .S(\clk2_output_dest[1] ),
    .X(mgmt_gpio_out_31_prebuff));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(\mgmt_gpio_data[30] ),
    .A1(clknet_4_13__leaf_wb_clk_i),
    .S(\clk1_output_dest[1] ),
    .X(mgmt_gpio_out_30_prebuff));
 sky130_fd_sc_hd__mux2_2 _4165_ (.A0(\mgmt_gpio_data[13] ),
    .A1(net93),
    .S(trap_output_dest),
    .X(net217));
 sky130_fd_sc_hd__mux2_4 _4166_ (.A0(serial_resetn_pre),
    .A1(serial_bb_resetn),
    .S(serial_bb_enable),
    .X(net305));
 sky130_fd_sc_hd__mux2_8 _4167_ (.A0(serial_load_pre),
    .A1(serial_bb_load),
    .S(serial_bb_enable),
    .X(net304));
 sky130_fd_sc_hd__nor4_2 _4168_ (.A(wbbd_busy),
    .B(hkspi_disable),
    .C(\gpio_configure[3][3] ),
    .D(net67),
    .Y(_1458_));
 sky130_fd_sc_hd__a22o_2 _4169_ (.A1(wbbd_busy),
    .A2(clknet_1_1__leaf_wbbd_sck),
    .B1(_1458_),
    .B2(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .X(csclk));
 sky130_fd_sc_hd__and2_1 _4170_ (.A(_1424_),
    .B(\wbbd_state[8] ),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _4171_ (.A(_1424_),
    .B(net3834),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _4172_ (.A(_1424_),
    .B(\wbbd_state[9] ),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _4173_ (.A(net68),
    .B(net94),
    .X(net300));
 sky130_fd_sc_hd__and2_1 _4174_ (.A(net63),
    .B(net79),
    .X(net306));
 sky130_fd_sc_hd__and2_1 _4175_ (.A(net36),
    .B(net1),
    .X(net171));
 sky130_fd_sc_hd__and2_2 _4176_ (.A(irq_1_inputsrc),
    .B(net70),
    .X(net173));
 sky130_fd_sc_hd__and2_2 _4177_ (.A(irq_2_inputsrc),
    .B(net39),
    .X(net174));
 sky130_fd_sc_hd__and2_1 _4178_ (.A(_1424_),
    .B(\wbbd_state[10] ),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(\hkspi.wrstb ),
    .A1(net2040),
    .S(net524),
    .X(_1459_));
 sky130_fd_sc_hd__and4_4 _4180_ (.A(net358),
    .B(net416),
    .C(net409),
    .D(net503),
    .X(_1460_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(net58),
    .A1(net2661),
    .S(net524),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(net3466),
    .A1(net499),
    .S(_1460_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(net2346),
    .A1(\wbbd_data[1] ),
    .S(net524),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(net3609),
    .A1(net491),
    .S(_1460_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_4 _4185_ (.A0(net2031),
    .A1(\wbbd_data[2] ),
    .S(net524),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(net3114),
    .A1(net487),
    .S(_1460_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_8 _4187_ (.A0(net2025),
    .A1(\wbbd_data[3] ),
    .S(net524),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(net2571),
    .A1(net483),
    .S(_1460_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(net2693),
    .A1(net790),
    .S(wbbd_busy),
    .X(_1465_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(net2721),
    .A1(net478),
    .S(_1460_),
    .X(_0069_));
 sky130_fd_sc_hd__and3_4 _4191_ (.A(net906),
    .B(net383),
    .C(net501),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(net3791),
    .A1(net495),
    .S(_1466_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(net3168),
    .A1(net489),
    .S(_1466_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(net2548),
    .A1(net484),
    .S(_1466_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net3127),
    .A1(net479),
    .S(_1466_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4196_ (.A0(net3633),
    .A1(net474),
    .S(_1466_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_4 _4197_ (.A0(net2015),
    .A1(\wbbd_data[5] ),
    .S(net524),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(net2554),
    .A1(net472),
    .S(_1466_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net2284),
    .A1(\wbbd_data[6] ),
    .S(wbbd_busy),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(net2830),
    .A1(net468),
    .S(_1466_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net2098),
    .A1(\wbbd_data[7] ),
    .S(wbbd_busy),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _4202_ (.A0(net2724),
    .A1(net465),
    .S(_1466_),
    .X(_0108_));
 sky130_fd_sc_hd__and4_4 _4203_ (.A(net415),
    .B(net906),
    .C(net410),
    .D(net501),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _4204_ (.A0(net3795),
    .A1(net495),
    .S(_1470_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net3096),
    .A1(net489),
    .S(_1470_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(net2637),
    .A1(net484),
    .S(_1470_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(net3209),
    .A1(net479),
    .S(_1470_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(net3376),
    .A1(net474),
    .S(_1470_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net2293),
    .A1(net472),
    .S(_1470_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(net2792),
    .A1(net468),
    .S(_1470_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net2715),
    .A1(net465),
    .S(_1470_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _4212_ (.A(net403),
    .B(net372),
    .C(net501),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(net3758),
    .A1(net495),
    .S(_1471_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(net3084),
    .A1(net489),
    .S(_1471_),
    .X(_0118_));
 sky130_fd_sc_hd__o311a_2 _4215_ (.A1(net3622),
    .A2(net2388),
    .A3(net67),
    .B1(net388),
    .C1(net380),
    .X(_1472_));
 sky130_fd_sc_hd__o221a_4 _4216_ (.A1(net369),
    .A2(_0864_),
    .B1(_0936_),
    .B2(_1472_),
    .C1(net504),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(net2758),
    .A1(net1088),
    .S(_0936_),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(net3247),
    .A1(_1474_),
    .S(_1473_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(net3522),
    .A1(net492),
    .S(_0936_),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(net3692),
    .A1(_1475_),
    .S(_1473_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(net2249),
    .A1(net488),
    .S(_0936_),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _4222_ (.A0(net2740),
    .A1(_1476_),
    .S(_1473_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(net2513),
    .A1(net481),
    .S(_0936_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(net2789),
    .A1(_1477_),
    .S(_1473_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(net3252),
    .A1(net477),
    .S(_0936_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(net3592),
    .A1(_1478_),
    .S(_1473_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net1991),
    .A1(net2017),
    .S(_0936_),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _4228_ (.A0(net2021),
    .A1(_1479_),
    .S(_1473_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(net2542),
    .A1(net685),
    .S(_0936_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net2786),
    .A1(_1480_),
    .S(_1473_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(net2943),
    .A1(net466),
    .S(_0936_),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _4232_ (.A0(net3308),
    .A1(_1481_),
    .S(_1473_),
    .X(_0126_));
 sky130_fd_sc_hd__o221a_4 _4233_ (.A1(net369),
    .A2(_0924_),
    .B1(_0935_),
    .B2(_1472_),
    .C1(net672),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(net3373),
    .A1(net497),
    .S(_0935_),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(net3684),
    .A1(_1483_),
    .S(_1482_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(net2918),
    .A1(net490),
    .S(_0935_),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _4237_ (.A0(net3302),
    .A1(_1484_),
    .S(_1482_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(net2055),
    .A1(net486),
    .S(_0935_),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_1 _4239_ (.A0(net2687),
    .A1(_1485_),
    .S(_1482_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(net2460),
    .A1(net480),
    .S(_0935_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(net2777),
    .A1(_1486_),
    .S(_1482_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(net3173),
    .A1(net708),
    .S(_0935_),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(net3469),
    .A1(_1487_),
    .S(_1482_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net2355),
    .A1(net471),
    .S(_0935_),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(net3378),
    .A1(_1488_),
    .S(_1482_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(net3170),
    .A1(net468),
    .S(_0935_),
    .X(_1489_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(net3479),
    .A1(_1489_),
    .S(_1482_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(net2807),
    .A1(net465),
    .S(_0935_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(net3311),
    .A1(_1490_),
    .S(_1482_),
    .X(_0134_));
 sky130_fd_sc_hd__o311a_4 _4250_ (.A1(net3909),
    .A2(net908),
    .A3(net67),
    .B1(_0936_),
    .C1(net672),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(net2758),
    .A1(net1088),
    .S(_1491_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(net3522),
    .A1(net492),
    .S(_1491_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net2249),
    .A1(net488),
    .S(_1491_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(net2513),
    .A1(net481),
    .S(_1491_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(net3252),
    .A1(net477),
    .S(_1491_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(net1991),
    .A1(net2017),
    .S(_1491_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(net2542),
    .A1(net685),
    .S(_1491_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(net2943),
    .A1(net466),
    .S(_1491_),
    .X(_0142_));
 sky130_fd_sc_hd__and4_2 _4259_ (.A(net415),
    .B(net410),
    .C(net372),
    .D(net501),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(net3747),
    .A1(net495),
    .S(_1492_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net3104),
    .A1(net489),
    .S(_1492_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(net2601),
    .A1(net484),
    .S(_1492_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net3124),
    .A1(net479),
    .S(_1492_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(net3665),
    .A1(net474),
    .S(_1492_),
    .X(_0147_));
 sky130_fd_sc_hd__and3_4 _4265_ (.A(net375),
    .B(net373),
    .C(net503),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(net3738),
    .A1(net496),
    .S(_1493_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net3595),
    .A1(net491),
    .S(_1493_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(net2477),
    .A1(net484),
    .S(_1493_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net3028),
    .A1(net479),
    .S(_1493_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(net3356),
    .A1(net476),
    .S(_1493_),
    .X(_0152_));
 sky130_fd_sc_hd__and4_4 _4271_ (.A(net411),
    .B(net408),
    .C(net2454),
    .D(net503),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(net3395),
    .A1(net499),
    .S(_1494_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(net3542),
    .A1(net491),
    .S(_1494_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4274_ (.A0(net2948),
    .A1(net487),
    .S(_1494_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(net2458),
    .A1(net483),
    .S(_1494_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(net3281),
    .A1(net476),
    .S(_1494_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_8 _4277_ (.A(net3805),
    .B(net608),
    .Y(_1495_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(_1495_),
    .B(net3476),
    .Y(_1496_));
 sky130_fd_sc_hd__o21ai_1 _4279_ (.A1(_1495_),
    .A2(_1368_),
    .B1(_1496_),
    .Y(_0158_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(_1297_),
    .A1(net3405),
    .S(_1495_),
    .X(_0159_));
 sky130_fd_sc_hd__nand2_1 _4281_ (.A(_1495_),
    .B(net3413),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_1 _4282_ (.A1(_1495_),
    .A2(_1231_),
    .B1(_1497_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _4283_ (.A(_1495_),
    .B(net3451),
    .Y(_1498_));
 sky130_fd_sc_hd__o21ai_1 _4284_ (.A1(_1495_),
    .A2(_1171_),
    .B1(_1498_),
    .Y(_0161_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_1495_),
    .B(net3548),
    .Y(_1499_));
 sky130_fd_sc_hd__o21ai_2 _4286_ (.A1(_1495_),
    .A2(clknet_1_0__leaf__1111_),
    .B1(_1499_),
    .Y(_0162_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(_1022_),
    .A1(net3408),
    .S(_1495_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(_0988_),
    .A1(net3386),
    .S(_1495_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_0953_),
    .A1(net3432),
    .S(_1495_),
    .X(_0165_));
 sky130_fd_sc_hd__nand2_8 _4290_ (.A(net3808),
    .B(net608),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(_1500_),
    .B(net3500),
    .Y(_1501_));
 sky130_fd_sc_hd__o21ai_1 _4292_ (.A1(_1500_),
    .A2(_1368_),
    .B1(_1501_),
    .Y(_0166_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_1297_),
    .A1(net3424),
    .S(_1500_),
    .X(_0167_));
 sky130_fd_sc_hd__nand2_1 _4294_ (.A(_1500_),
    .B(net3439),
    .Y(_1502_));
 sky130_fd_sc_hd__o21ai_1 _4295_ (.A1(_1500_),
    .A2(_1231_),
    .B1(_1502_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _4296_ (.A(_1500_),
    .B(net3461),
    .Y(_1503_));
 sky130_fd_sc_hd__o21ai_1 _4297_ (.A1(_1500_),
    .A2(_1171_),
    .B1(_1503_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_1500_),
    .B(net3494),
    .Y(_1504_));
 sky130_fd_sc_hd__o21ai_2 _4299_ (.A1(_1500_),
    .A2(clknet_1_0__leaf__1111_),
    .B1(_1504_),
    .Y(_0170_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(_1022_),
    .A1(net3471),
    .S(_1500_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(_0988_),
    .A1(net3506),
    .S(_1500_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(_0953_),
    .A1(net3524),
    .S(_1500_),
    .X(_0173_));
 sky130_fd_sc_hd__and3_2 _4303_ (.A(net378),
    .B(net370),
    .C(net501),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(net3780),
    .A1(net495),
    .S(_1505_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(net3092),
    .A1(net489),
    .S(_1505_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(net2511),
    .A1(net484),
    .S(_1505_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(net3082),
    .A1(net479),
    .S(_1505_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(net3678),
    .A1(net474),
    .S(_1505_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_8 _4309_ (.A(net3809),
    .B(net607),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_1506_),
    .B(net3442),
    .Y(_1507_));
 sky130_fd_sc_hd__o21ai_1 _4311_ (.A1(_1506_),
    .A2(_1368_),
    .B1(_1507_),
    .Y(_0179_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(_1297_),
    .A1(net3419),
    .S(_1506_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_1506_),
    .B(net3410),
    .Y(_1508_));
 sky130_fd_sc_hd__o21ai_1 _4314_ (.A1(_1506_),
    .A2(_1231_),
    .B1(_1508_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_1506_),
    .B(net3473),
    .Y(_1509_));
 sky130_fd_sc_hd__o21ai_1 _4316_ (.A1(_1506_),
    .A2(_1171_),
    .B1(_1509_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_1506_),
    .B(net3535),
    .Y(_1510_));
 sky130_fd_sc_hd__o21ai_2 _4318_ (.A1(_1506_),
    .A2(clknet_1_0__leaf__1111_),
    .B1(_1510_),
    .Y(_0183_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(_1022_),
    .A1(net3429),
    .S(_1506_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(_0988_),
    .A1(net3391),
    .S(_1506_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(_0953_),
    .A1(net3486),
    .S(_1506_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_4 _4322_ (.A(_1024_),
    .B(net502),
    .Y(_1511_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(net496),
    .A1(net3785),
    .S(_1511_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(net489),
    .A1(net3136),
    .S(_1511_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(net484),
    .A1(net2635),
    .S(_1511_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(net479),
    .A1(net3014),
    .S(_1511_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(net474),
    .A1(net3614),
    .S(_1511_),
    .X(_0191_));
 sky130_fd_sc_hd__and4_4 _4328_ (.A(net413),
    .B(net409),
    .C(net378),
    .D(net501),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(net3723),
    .A1(net496),
    .S(_1512_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(net3117),
    .A1(net489),
    .S(_1512_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(net2277),
    .A1(net485),
    .S(_1512_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(net2950),
    .A1(net479),
    .S(_1512_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(net3668),
    .A1(net474),
    .S(_1512_),
    .X(_0196_));
 sky130_fd_sc_hd__and4_4 _4334_ (.A(net420),
    .B(net411),
    .C(net2454),
    .D(net671),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(net3771),
    .A1(net496),
    .S(_1513_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(net3631),
    .A1(net491),
    .S(_1513_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(net1094),
    .A1(net484),
    .S(_1513_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(net2599),
    .A1(net483),
    .S(_1513_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _4339_ (.A0(net3351),
    .A1(net476),
    .S(_1513_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_4 _4340_ (.A(_1031_),
    .B(net502),
    .Y(_1514_));
 sky130_fd_sc_hd__mux2_1 _4341_ (.A0(net496),
    .A1(net3711),
    .S(_1514_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(net667),
    .A1(net2463),
    .S(_1514_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(net484),
    .A1(net2613),
    .S(_1514_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(net479),
    .A1(net3016),
    .S(_1514_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(net474),
    .A1(net3562),
    .S(_1514_),
    .X(_0206_));
 sky130_fd_sc_hd__and4_4 _4346_ (.A(net415),
    .B(net410),
    .C(net378),
    .D(net501),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(net3731),
    .A1(net495),
    .S(_1515_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4348_ (.A0(net3148),
    .A1(net489),
    .S(_1515_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(net2622),
    .A1(net484),
    .S(_1515_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(net3056),
    .A1(net479),
    .S(_1515_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(net3648),
    .A1(net474),
    .S(_1515_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_2 _4352_ (.A(net2454),
    .B(net375),
    .C(net503),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(net3404),
    .A1(net499),
    .S(_1516_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(net3558),
    .A1(net491),
    .S(_1516_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _4355_ (.A0(net2992),
    .A1(net487),
    .S(_1516_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(net2597),
    .A1(net483),
    .S(_1516_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4357_ (.A0(net3294),
    .A1(net476),
    .S(_1516_),
    .X(_0216_));
 sky130_fd_sc_hd__and4_4 _4358_ (.A(net391),
    .B(net411),
    .C(net408),
    .D(net503),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(net3446),
    .A1(net499),
    .S(_1517_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(net3644),
    .A1(net491),
    .S(_1517_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _4361_ (.A0(net2999),
    .A1(net487),
    .S(_1517_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(net2578),
    .A1(net483),
    .S(_1517_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4363_ (.A0(net3292),
    .A1(net476),
    .S(_1517_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_2 _4364_ (.A(net390),
    .B(net370),
    .C(net502),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(net3727),
    .A1(net496),
    .S(_1518_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(net2982),
    .A1(net489),
    .S(_1518_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _4367_ (.A0(net2473),
    .A1(net484),
    .S(_1518_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(net2593),
    .A1(net480),
    .S(_1518_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _4369_ (.A0(net3673),
    .A1(net474),
    .S(_1518_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_4 _4370_ (.A(_1034_),
    .B(net503),
    .Y(_1519_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(net499),
    .A1(net3457),
    .S(_1519_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(net493),
    .A1(net3010),
    .S(_1519_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(net487),
    .A1(net3087),
    .S(_1519_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _4374_ (.A0(net483),
    .A1(net2643),
    .S(_1519_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _4375_ (.A0(net478),
    .A1(net2780),
    .S(_1519_),
    .X(_0231_));
 sky130_fd_sc_hd__and4_4 _4376_ (.A(net413),
    .B(net356),
    .C(net409),
    .D(net503),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _4377_ (.A0(net3497),
    .A1(net499),
    .S(_1520_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(net3646),
    .A1(net491),
    .S(_1520_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(net3100),
    .A1(net487),
    .S(_1520_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(net2611),
    .A1(net483),
    .S(_1520_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(net3390),
    .A1(net476),
    .S(_1520_),
    .X(_0236_));
 sky130_fd_sc_hd__nand4_4 _4382_ (.A(net420),
    .B(net358),
    .C(net409),
    .D(net503),
    .Y(_1521_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(net496),
    .A1(net3766),
    .S(_1521_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _4384_ (.A0(net491),
    .A1(net3551),
    .S(_1521_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(net485),
    .A1(net2361),
    .S(_1521_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(net480),
    .A1(net2436),
    .S(_1521_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _4387_ (.A0(net476),
    .A1(net3348),
    .S(_1521_),
    .X(_0241_));
 sky130_fd_sc_hd__nand4_4 _4388_ (.A(net680),
    .B(net409),
    .C(net2092),
    .D(net501),
    .Y(_1522_));
 sky130_fd_sc_hd__mux2_1 _4389_ (.A0(net496),
    .A1(net3328),
    .S(_1522_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(net491),
    .A1(net3340),
    .S(_1522_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _4391_ (.A0(net485),
    .A1(net980),
    .S(_1522_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(net480),
    .A1(net2367),
    .S(_1522_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(net474),
    .A1(net3324),
    .S(_1522_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_4 _4394_ (.A(_1040_),
    .B(net502),
    .Y(_1523_));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(net496),
    .A1(net3761),
    .S(_1523_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _4396_ (.A0(net667),
    .A1(net2393),
    .S(_1523_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(net485),
    .A1(net2218),
    .S(_1523_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _4398_ (.A0(net479),
    .A1(net2960),
    .S(_1523_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _4399_ (.A0(net474),
    .A1(net3566),
    .S(_1523_),
    .X(_0251_));
 sky130_fd_sc_hd__and4_4 _4400_ (.A(net410),
    .B(net680),
    .C(net2092),
    .D(net501),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(net3694),
    .A1(net496),
    .S(_1524_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _4402_ (.A0(net3682),
    .A1(net491),
    .S(_1524_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _4403_ (.A0(net2275),
    .A1(net485),
    .S(_1524_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(net2676),
    .A1(net480),
    .S(_1524_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(net3364),
    .A1(net476),
    .S(_1524_),
    .X(_0256_));
 sky130_fd_sc_hd__o31ai_2 _4406_ (.A1(net1869),
    .A2(net908),
    .A3(net67),
    .B1(_0932_),
    .Y(_1525_));
 sky130_fd_sc_hd__o211a_4 _4407_ (.A1(_0932_),
    .A2(_1472_),
    .B1(_1525_),
    .C1(net504),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(net2743),
    .A1(net498),
    .S(_0932_),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _4409_ (.A0(net3569),
    .A1(_1527_),
    .S(_1526_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(net3459),
    .A1(net492),
    .S(_0932_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _4411_ (.A0(net3639),
    .A1(_1528_),
    .S(_1526_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(net2144),
    .A1(net488),
    .S(_0932_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(net2706),
    .A1(_1529_),
    .S(_1526_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(net2241),
    .A1(net482),
    .S(_0932_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _4415_ (.A0(net2718),
    .A1(_1530_),
    .S(_1526_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _4416_ (.A0(net2783),
    .A1(net476),
    .S(_0932_),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _4417_ (.A0(net3577),
    .A1(_1531_),
    .S(_1526_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _4418_ (.A0(net2405),
    .A1(net473),
    .S(_0932_),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(net2755),
    .A1(_1532_),
    .S(_1526_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(net2627),
    .A1(net685),
    .S(_0932_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(net2812),
    .A1(_1533_),
    .S(_1526_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(net3023),
    .A1(net466),
    .S(_0932_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(net3276),
    .A1(_1534_),
    .S(_1526_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(\wbbd_state[1] ),
    .B(net3854),
    .Y(_1535_));
 sky130_fd_sc_hd__nor4b_2 _4425_ (.A(net3808),
    .B(net3809),
    .C(net3805),
    .D_N(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__nor3_2 _4426_ (.A(\wbbd_state[8] ),
    .B(\wbbd_state[9] ),
    .C(\wbbd_state[10] ),
    .Y(_1537_));
 sky130_fd_sc_hd__nor4_4 _4427_ (.A(net3876),
    .B(\wbbd_state[8] ),
    .C(\wbbd_state[9] ),
    .D(\wbbd_state[10] ),
    .Y(_1538_));
 sky130_fd_sc_hd__nand2b_4 _4428_ (.A_N(\wbbd_state[6] ),
    .B(net463),
    .Y(_1539_));
 sky130_fd_sc_hd__nand2b_1 _4429_ (.A_N(net3875),
    .B(net524),
    .Y(_1540_));
 sky130_fd_sc_hd__nand4b_1 _4430_ (.A_N(net3813),
    .B(_1536_),
    .C(_1538_),
    .D(_1540_),
    .Y(_0265_));
 sky130_fd_sc_hd__and3_4 _4431_ (.A(net388),
    .B(net380),
    .C(net504),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _4432_ (.A0(net3626),
    .A1(net498),
    .S(_1541_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(net3450),
    .A1(net492),
    .S(_1541_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _4434_ (.A0(net2181),
    .A1(net488),
    .S(_1541_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(net2262),
    .A1(net482),
    .S(_1541_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(net2709),
    .A1(net478),
    .S(_1541_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(net2109),
    .A1(net473),
    .S(_1541_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _4438_ (.A0(net2314),
    .A1(net685),
    .S(_1541_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(net2934),
    .A1(net466),
    .S(_1541_),
    .X(_0273_));
 sky130_fd_sc_hd__o311a_4 _4440_ (.A1(hkspi_disable),
    .A2(net908),
    .A3(net67),
    .B1(_0932_),
    .C1(net504),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(net2743),
    .A1(net1088),
    .S(_1542_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(net3459),
    .A1(net492),
    .S(_1542_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(net2144),
    .A1(net488),
    .S(_1542_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(net2241),
    .A1(net482),
    .S(_1542_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(net2783),
    .A1(net478),
    .S(_1542_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _4446_ (.A0(net2405),
    .A1(net473),
    .S(_1542_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(net2627),
    .A1(net685),
    .S(_1542_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(net3023),
    .A1(net466),
    .S(_1542_),
    .X(_0281_));
 sky130_fd_sc_hd__and4_2 _4449_ (.A(net391),
    .B(net413),
    .C(net2210),
    .D(net503),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _4450_ (.A0(net3423),
    .A1(net499),
    .S(_1543_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(net3554),
    .A1(net491),
    .S(_1543_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(net3098),
    .A1(net487),
    .S(_1543_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(net2670),
    .A1(net483),
    .S(_1543_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(net3383),
    .A1(net476),
    .S(_1543_),
    .X(_0286_));
 sky130_fd_sc_hd__and4_1 _4455_ (.A(net414),
    .B(net381),
    .C(net2210),
    .D(net671),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _4456_ (.A0(net3438),
    .A1(net499),
    .S(net780),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _4457_ (.A0(net3660),
    .A1(net491),
    .S(net780),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(net3045),
    .A1(net487),
    .S(net780),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(net2658),
    .A1(net483),
    .S(net780),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _4460_ (.A0(net2761),
    .A1(net478),
    .S(net780),
    .X(_0291_));
 sky130_fd_sc_hd__and4_4 _4461_ (.A(net391),
    .B(net420),
    .C(net411),
    .D(net503),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(net3527),
    .A1(net499),
    .S(_1545_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(net3612),
    .A1(net491),
    .S(_1545_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(net3037),
    .A1(net487),
    .S(_1545_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(net2574),
    .A1(net483),
    .S(_1545_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(net2751),
    .A1(net478),
    .S(_1545_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_4 _4467_ (.A(_1038_),
    .B(net503),
    .Y(_1546_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(net499),
    .A1(net3499),
    .S(_1546_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(net493),
    .A1(net3073),
    .S(_1546_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(net487),
    .A1(net3001),
    .S(_1546_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(net483),
    .A1(net2648),
    .S(_1546_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(net478),
    .A1(net2771),
    .S(_1546_),
    .X(_0301_));
 sky130_fd_sc_hd__and3_2 _4473_ (.A(net391),
    .B(net374),
    .C(net503),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(net3397),
    .A1(net499),
    .S(_1547_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(net3598),
    .A1(net491),
    .S(_1547_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(net3162),
    .A1(net487),
    .S(_1547_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(net2604),
    .A1(net483),
    .S(_1547_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(net3326),
    .A1(net476),
    .S(_1547_),
    .X(_0306_));
 sky130_fd_sc_hd__and3_2 _4479_ (.A(net381),
    .B(net371),
    .C(net503),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(net3428),
    .A1(net499),
    .S(_1548_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(net3112),
    .A1(net493),
    .S(_1548_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(net3041),
    .A1(net487),
    .S(_1548_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4483_ (.A0(net2673),
    .A1(net483),
    .S(_1548_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net3402),
    .A1(net476),
    .S(_1548_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_4 _4485_ (.A(_1042_),
    .B(net502),
    .Y(_1549_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(net495),
    .A1(net3753),
    .S(_1549_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(net489),
    .A1(net3144),
    .S(_1549_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(net484),
    .A1(net2651),
    .S(_1549_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(net479),
    .A1(net3043),
    .S(_1549_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(net474),
    .A1(net3680),
    .S(_1549_),
    .X(_0316_));
 sky130_fd_sc_hd__and4_4 _4491_ (.A(net412),
    .B(net381),
    .C(net408),
    .D(net503),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _4492_ (.A0(net3489),
    .A1(net499),
    .S(_1550_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(net3122),
    .A1(net493),
    .S(_1550_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(net3039),
    .A1(net487),
    .S(_1550_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(net2681),
    .A1(net483),
    .S(_1550_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(net3385),
    .A1(net476),
    .S(_1550_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_4 _4497_ (.A(_1050_),
    .B(net503),
    .Y(_1551_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(net499),
    .A1(net3491),
    .S(_1551_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(net493),
    .A1(net3131),
    .S(_1551_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(net487),
    .A1(net3061),
    .S(_1551_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _4501_ (.A0(net483),
    .A1(net2618),
    .S(_1551_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(net478),
    .A1(net2730),
    .S(_1551_),
    .X(_0326_));
 sky130_fd_sc_hd__and3_2 _4503_ (.A(net680),
    .B(net375),
    .C(net503),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(net3725),
    .A1(net496),
    .S(_1552_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(net3158),
    .A1(net489),
    .S(_1552_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(net2265),
    .A1(net485),
    .S(_1552_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(net2973),
    .A1(net479),
    .S(_1552_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(net3637),
    .A1(net474),
    .S(_1552_),
    .X(_0331_));
 sky130_fd_sc_hd__and4_4 _4509_ (.A(net357),
    .B(net410),
    .C(net2092),
    .D(net502),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(net3689),
    .A1(net496),
    .S(_1553_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(net3606),
    .A1(net491),
    .S(_1553_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(net2333),
    .A1(net485),
    .S(_1553_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(net2582),
    .A1(net483),
    .S(_1553_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(net3335),
    .A1(net476),
    .S(_1553_),
    .X(_0336_));
 sky130_fd_sc_hd__and4_4 _4515_ (.A(net416),
    .B(net411),
    .C(net354),
    .D(net503),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _4516_ (.A0(net3736),
    .A1(net496),
    .S(_1554_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _4517_ (.A0(net3587),
    .A1(net491),
    .S(_1554_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(net942),
    .A1(net485),
    .S(_1554_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(net2987),
    .A1(net479),
    .S(_1554_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(net3338),
    .A1(net476),
    .S(_1554_),
    .X(_0341_));
 sky130_fd_sc_hd__and3_2 _4521_ (.A(net358),
    .B(net371),
    .C(net503),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(net3399),
    .A1(net499),
    .S(_1555_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _4523_ (.A0(net3618),
    .A1(net491),
    .S(_1555_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(net3018),
    .A1(net487),
    .S(_1555_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(net2442),
    .A1(net483),
    .S(_1555_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(net3370),
    .A1(net476),
    .S(_1555_),
    .X(_0346_));
 sky130_fd_sc_hd__and3_4 _4527_ (.A(net680),
    .B(net374),
    .C(net501),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(net3764),
    .A1(net496),
    .S(_1556_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(net3164),
    .A1(net489),
    .S(_1556_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net2353),
    .A1(net485),
    .S(_1556_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(net2971),
    .A1(net479),
    .S(_1556_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net3153),
    .A1(net708),
    .S(_1556_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_4 _4533_ (.A(_1028_),
    .B(net503),
    .Y(_1557_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(net499),
    .A1(net3417),
    .S(_1557_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(net491),
    .A1(net3603),
    .S(_1557_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(net487),
    .A1(net3053),
    .S(_1557_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net483),
    .A1(net2608),
    .S(_1557_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(net476),
    .A1(net3353),
    .S(_1557_),
    .X(_0356_));
 sky130_fd_sc_hd__and4_1 _4539_ (.A(net660),
    .B(net410),
    .C(net680),
    .D(net502),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(net3775),
    .A1(net496),
    .S(net681),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _4541_ (.A0(net2001),
    .A1(net667),
    .S(net681),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(net2255),
    .A1(net485),
    .S(net681),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(net3012),
    .A1(net479),
    .S(net681),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _4544_ (.A0(net3635),
    .A1(net474),
    .S(net681),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_4 _4545_ (.A(_1046_),
    .B(net502),
    .Y(_1559_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(net496),
    .A1(net3715),
    .S(_1559_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(net491),
    .A1(net3600),
    .S(_1559_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _4548_ (.A0(net485),
    .A1(net2505),
    .S(_1559_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _4549_ (.A0(net480),
    .A1(net2557),
    .S(_1559_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(net476),
    .A1(net3314),
    .S(_1559_),
    .X(_0366_));
 sky130_fd_sc_hd__nand4_4 _4551_ (.A(net420),
    .B(net358),
    .C(net411),
    .D(net503),
    .Y(_1560_));
 sky130_fd_sc_hd__mux2_1 _4552_ (.A0(net499),
    .A1(net3517),
    .S(_1560_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(net493),
    .A1(net2996),
    .S(_1560_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _4554_ (.A0(net487),
    .A1(net2989),
    .S(_1560_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _4555_ (.A0(net483),
    .A1(net2655),
    .S(_1560_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(net476),
    .A1(net3345),
    .S(_1560_),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _4557_ (.A(net2066),
    .B(\wbbd_state[6] ),
    .Y(_1561_));
 sky130_fd_sc_hd__and4_2 _4558_ (.A(net112),
    .B(net111),
    .C(net114),
    .D(net113),
    .X(_1562_));
 sky130_fd_sc_hd__a21o_4 _4559_ (.A1(_1425_),
    .A2(_1426_),
    .B1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__nor3_4 _4560_ (.A(net112),
    .B(net114),
    .C(net113),
    .Y(_1564_));
 sky130_fd_sc_hd__and4_4 _4561_ (.A(net107),
    .B(net106),
    .C(net109),
    .D(net108),
    .X(_1565_));
 sky130_fd_sc_hd__nand4_4 _4562_ (.A(net107),
    .B(net106),
    .C(net109),
    .D(net108),
    .Y(_1566_));
 sky130_fd_sc_hd__nand4_4 _4563_ (.A(net103),
    .B(net102),
    .C(net105),
    .D(net104),
    .Y(_1567_));
 sky130_fd_sc_hd__nand4_4 _4564_ (.A(net130),
    .B(net129),
    .C(net101),
    .D(net100),
    .Y(_1568_));
 sky130_fd_sc_hd__nor2_8 _4565_ (.A(_1567_),
    .B(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__and2_4 _4566_ (.A(net612),
    .B(net614),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_8 _4567_ (.A(net612),
    .B(net614),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_4 _4568_ (.A(net610),
    .B(net611),
    .Y(_1572_));
 sky130_fd_sc_hd__and3_2 _4569_ (.A(net610),
    .B(net611),
    .C(net614),
    .X(_1573_));
 sky130_fd_sc_hd__nand3_4 _4570_ (.A(net610),
    .B(net612),
    .C(net614),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_8 _4571_ (.A(net616),
    .B(net618),
    .Y(_1575_));
 sky130_fd_sc_hd__and3_4 _4572_ (.A(net619),
    .B(net615),
    .C(net617),
    .X(_1576_));
 sky130_fd_sc_hd__nand3_4 _4573_ (.A(net619),
    .B(net615),
    .C(net617),
    .Y(_1577_));
 sky130_fd_sc_hd__and4_2 _4574_ (.A(net619),
    .B(net615),
    .C(net617),
    .D(net614),
    .X(_1578_));
 sky130_fd_sc_hd__nand4_4 _4575_ (.A(net621),
    .B(net616),
    .C(net618),
    .D(net614),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_2 _4576_ (.A(_1573_),
    .B(_1576_),
    .Y(_1580_));
 sky130_fd_sc_hd__nand3_4 _4577_ (.A(net610),
    .B(net609),
    .C(net612),
    .Y(_1581_));
 sky130_fd_sc_hd__nor2_8 _4578_ (.A(_1579_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__and4_4 _4579_ (.A(net610),
    .B(net609),
    .C(net612),
    .D(net614),
    .X(_1583_));
 sky130_fd_sc_hd__nand4_4 _4580_ (.A(net610),
    .B(net609),
    .C(net612),
    .D(net614),
    .Y(_1584_));
 sky130_fd_sc_hd__and4_4 _4581_ (.A(net621),
    .B(net562),
    .C(net616),
    .D(net618),
    .X(_1585_));
 sky130_fd_sc_hd__nand4_4 _4582_ (.A(net621),
    .B(net562),
    .C(net616),
    .D(net618),
    .Y(_1586_));
 sky130_fd_sc_hd__nor2_2 _4583_ (.A(_1584_),
    .B(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__nand4_4 _4584_ (.A(_1565_),
    .B(_1569_),
    .C(_1583_),
    .D(net558),
    .Y(_1588_));
 sky130_fd_sc_hd__nand4_2 _4585_ (.A(_1569_),
    .B(_1583_),
    .C(net558),
    .D(_0821_),
    .Y(_1589_));
 sky130_fd_sc_hd__nand4_4 _4586_ (.A(_1565_),
    .B(_1569_),
    .C(_1587_),
    .D(_0821_),
    .Y(_1590_));
 sky130_fd_sc_hd__a21boi_4 _4587_ (.A1(net111),
    .A2(_1588_),
    .B1_N(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__a2bb2o_4 _4588_ (.A1_N(_1566_),
    .A2_N(_1589_),
    .B1(_1588_),
    .B2(net111),
    .X(_1592_));
 sky130_fd_sc_hd__and2b_4 _4589_ (.A_N(net112),
    .B(net111),
    .X(_1593_));
 sky130_fd_sc_hd__and2b_4 _4590_ (.A_N(net111),
    .B(net112),
    .X(_1594_));
 sky130_fd_sc_hd__nor2_8 _4591_ (.A(_1593_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__o2111a_1 _4592_ (.A1(_1593_),
    .A2(_1594_),
    .B1(_1565_),
    .C1(_1569_),
    .D1(_1587_),
    .X(_1596_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_1588_),
    .B(net112),
    .Y(_1597_));
 sky130_fd_sc_hd__nor4_2 _4594_ (.A(net112),
    .B(net114),
    .C(net113),
    .D(_1591_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_8 _4595_ (.A(_1592_),
    .B(net559),
    .Y(_1599_));
 sky130_fd_sc_hd__and2b_2 _4596_ (.A_N(net621),
    .B(net562),
    .X(_1600_));
 sky130_fd_sc_hd__nand2b_4 _4597_ (.A_N(net620),
    .B(net561),
    .Y(_1601_));
 sky130_fd_sc_hd__and2b_4 _4598_ (.A_N(net617),
    .B(net615),
    .X(_1602_));
 sky130_fd_sc_hd__nand2b_4 _4599_ (.A_N(net617),
    .B(net615),
    .Y(_1603_));
 sky130_fd_sc_hd__nor2_8 _4600_ (.A(_1601_),
    .B(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__nand2_8 _4601_ (.A(net556),
    .B(_1602_),
    .Y(_1605_));
 sky130_fd_sc_hd__nor2_8 _4602_ (.A(net612),
    .B(net614),
    .Y(_1606_));
 sky130_fd_sc_hd__nor2_8 _4603_ (.A(net610),
    .B(net609),
    .Y(_1607_));
 sky130_fd_sc_hd__nor4_2 _4604_ (.A(net610),
    .B(net609),
    .C(net612),
    .D(net614),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_8 _4605_ (.A(_1606_),
    .B(_1607_),
    .Y(_1609_));
 sky130_fd_sc_hd__nor2_8 _4606_ (.A(net621),
    .B(net562),
    .Y(_1610_));
 sky130_fd_sc_hd__o211a_4 _4607_ (.A1(net621),
    .A2(net562),
    .B1(net616),
    .C1(net618),
    .X(_1611_));
 sky130_fd_sc_hd__o211ai_4 _4608_ (.A1(net621),
    .A2(net562),
    .B1(net616),
    .C1(net618),
    .Y(_1612_));
 sky130_fd_sc_hd__o2111ai_4 _4609_ (.A1(net621),
    .A2(net562),
    .B1(net616),
    .C1(net618),
    .D1(net614),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_2 _4610_ (.A(_1570_),
    .B(_1611_),
    .Y(_1614_));
 sky130_fd_sc_hd__o21bai_4 _4611_ (.A1(_0828_),
    .A2(_1612_),
    .B1_N(net612),
    .Y(_1615_));
 sky130_fd_sc_hd__o21ai_4 _4612_ (.A1(_1575_),
    .A2(_1610_),
    .B1(_0828_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_2 _4613_ (.A(_1613_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__a22oi_4 _4614_ (.A1(_1614_),
    .A2(_1615_),
    .B1(_1616_),
    .B2(_1613_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _4615_ (.A(_1573_),
    .B(_1611_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_2 _4616_ (.A(_1583_),
    .B(_1611_),
    .Y(_1620_));
 sky130_fd_sc_hd__o21bai_4 _4617_ (.A1(_1574_),
    .A2(net550),
    .B1_N(net609),
    .Y(_1621_));
 sky130_fd_sc_hd__o21bai_4 _4618_ (.A1(_1571_),
    .A2(net550),
    .B1_N(net610),
    .Y(_1622_));
 sky130_fd_sc_hd__o21ai_4 _4619_ (.A1(_1574_),
    .A2(net550),
    .B1(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a22oi_4 _4620_ (.A1(_1620_),
    .A2(_1621_),
    .B1(_1622_),
    .B2(_1619_),
    .Y(_1624_));
 sky130_fd_sc_hd__and2_4 _4621_ (.A(net429),
    .B(net428),
    .X(_1625_));
 sky130_fd_sc_hd__nand2_8 _4622_ (.A(net429),
    .B(_1624_),
    .Y(_1626_));
 sky130_fd_sc_hd__and3_1 _4623_ (.A(net363),
    .B(_1604_),
    .C(net552),
    .X(_1627_));
 sky130_fd_sc_hd__and3_4 _4624_ (.A(net619),
    .B(net561),
    .C(_1602_),
    .X(_1628_));
 sky130_fd_sc_hd__nand3_4 _4625_ (.A(net619),
    .B(net561),
    .C(_1602_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand2_4 _4626_ (.A(net614),
    .B(_1585_),
    .Y(_1630_));
 sky130_fd_sc_hd__o21bai_4 _4627_ (.A1(_1571_),
    .A2(net557),
    .B1_N(net610),
    .Y(_1631_));
 sky130_fd_sc_hd__nand3_2 _4628_ (.A(net562),
    .B(net610),
    .C(net612),
    .Y(_1632_));
 sky130_fd_sc_hd__o31a_4 _4629_ (.A1(_0828_),
    .A2(_1572_),
    .A3(net557),
    .B1(_1631_),
    .X(_1633_));
 sky130_fd_sc_hd__o21ai_4 _4630_ (.A1(_1574_),
    .A2(net557),
    .B1(_1631_),
    .Y(_1634_));
 sky130_fd_sc_hd__o21ai_2 _4631_ (.A1(_1574_),
    .A2(net557),
    .B1(net609),
    .Y(_1635_));
 sky130_fd_sc_hd__o31ai_4 _4632_ (.A1(net609),
    .A2(_1579_),
    .A3(_1632_),
    .B1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__nor2_4 _4633_ (.A(_1633_),
    .B(net427),
    .Y(_1637_));
 sky130_fd_sc_hd__a41o_4 _4634_ (.A1(net620),
    .A2(net561),
    .A3(net615),
    .A4(net617),
    .B1(net614),
    .X(_1638_));
 sky130_fd_sc_hd__a21boi_4 _4635_ (.A1(net561),
    .A2(_1578_),
    .B1_N(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__o21bai_4 _4636_ (.A1(_0828_),
    .A2(net557),
    .B1_N(net612),
    .Y(_1640_));
 sky130_fd_sc_hd__nor2_8 _4637_ (.A(net611),
    .B(_0828_),
    .Y(_1641_));
 sky130_fd_sc_hd__o21a_4 _4638_ (.A1(_1571_),
    .A2(net557),
    .B1(_1640_),
    .X(_1642_));
 sky130_fd_sc_hd__o21ai_4 _4639_ (.A1(_1571_),
    .A2(net557),
    .B1(_1640_),
    .Y(_1643_));
 sky130_fd_sc_hd__a21oi_4 _4640_ (.A1(_1630_),
    .A2(_1638_),
    .B1(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__nor4_2 _4641_ (.A(net427),
    .B(_1643_),
    .C(_1639_),
    .D(_1633_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand4_4 _4642_ (.A(_1565_),
    .B(_1569_),
    .C(_1583_),
    .D(_1611_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand4_1 _4643_ (.A(_1565_),
    .B(_1569_),
    .C(_1583_),
    .D(_1611_),
    .Y(_1647_));
 sky130_fd_sc_hd__a41oi_4 _4644_ (.A1(_1565_),
    .A2(_1569_),
    .A3(_1583_),
    .A4(_1611_),
    .B1(_0821_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand4_4 _4645_ (.A(_1569_),
    .B(_0821_),
    .C(_1565_),
    .D(_1611_),
    .Y(_1649_));
 sky130_fd_sc_hd__nor2_4 _4646_ (.A(_1584_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__a2bb2oi_2 _4647_ (.A1_N(_1584_),
    .A2_N(_1649_),
    .B1(_1647_),
    .B2(net111),
    .Y(_1651_));
 sky130_fd_sc_hd__nand2_4 _4648_ (.A(_1646_),
    .B(net112),
    .Y(_1652_));
 sky130_fd_sc_hd__nand4bb_4 _4649_ (.A_N(_1595_),
    .B_N(_1620_),
    .C(_1565_),
    .D(_1569_),
    .Y(_1653_));
 sky130_fd_sc_hd__o21a_4 _4650_ (.A1(_1595_),
    .A2(_1646_),
    .B1(_1652_),
    .X(_1654_));
 sky130_fd_sc_hd__o21ai_4 _4651_ (.A1(_1595_),
    .A2(_1646_),
    .B1(_1652_),
    .Y(_1655_));
 sky130_fd_sc_hd__o211a_4 _4652_ (.A1(_1646_),
    .A2(_1595_),
    .B1(_1563_),
    .C1(_1652_),
    .X(_1656_));
 sky130_fd_sc_hd__o21a_4 _4653_ (.A1(_1648_),
    .A2(_1650_),
    .B1(net560),
    .X(_1657_));
 sky130_fd_sc_hd__o21ai_4 _4654_ (.A1(_1648_),
    .A2(_1650_),
    .B1(net560),
    .Y(_1658_));
 sky130_fd_sc_hd__o311a_4 _4655_ (.A1(_1571_),
    .A2(_1575_),
    .A3(_1610_),
    .B1(_1615_),
    .C1(_1617_),
    .X(_1659_));
 sky130_fd_sc_hd__o211ai_4 _4656_ (.A1(_1571_),
    .A2(_1612_),
    .B1(_1615_),
    .C1(_1617_),
    .Y(_1660_));
 sky130_fd_sc_hd__and4_4 _4657_ (.A(_1624_),
    .B(_1617_),
    .C(_1615_),
    .D(_1614_),
    .X(_1661_));
 sky130_fd_sc_hd__and3_2 _4658_ (.A(net428),
    .B(_1657_),
    .C(_1659_),
    .X(_1662_));
 sky130_fd_sc_hd__nand2_2 _4659_ (.A(_1657_),
    .B(_1661_),
    .Y(_1663_));
 sky130_fd_sc_hd__a41oi_4 _4660_ (.A1(net619),
    .A2(net615),
    .A3(net617),
    .A4(net614),
    .B1(net611),
    .Y(_1664_));
 sky130_fd_sc_hd__a31o_4 _4661_ (.A1(net619),
    .A2(net615),
    .A3(net617),
    .B1(net614),
    .X(_1665_));
 sky130_fd_sc_hd__a21oi_4 _4662_ (.A1(_1665_),
    .A2(net611),
    .B1(_1664_),
    .Y(_1666_));
 sky130_fd_sc_hd__o21bai_4 _4663_ (.A1(_1571_),
    .A2(_1577_),
    .B1_N(net610),
    .Y(_1667_));
 sky130_fd_sc_hd__o21ai_4 _4664_ (.A1(_1572_),
    .A2(_1579_),
    .B1(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__and2b_4 _4665_ (.A_N(net609),
    .B(net610),
    .X(_1669_));
 sky130_fd_sc_hd__nand2b_4 _4666_ (.A_N(net609),
    .B(net610),
    .Y(_1670_));
 sky130_fd_sc_hd__nor3_2 _4667_ (.A(_1571_),
    .B(_1577_),
    .C(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__nand4_4 _4668_ (.A(net611),
    .B(net614),
    .C(_1576_),
    .D(_1669_),
    .Y(_1672_));
 sky130_fd_sc_hd__o21a_4 _4669_ (.A1(_1574_),
    .A2(_1577_),
    .B1(net609),
    .X(_1673_));
 sky130_fd_sc_hd__o21ai_4 _4670_ (.A1(_1572_),
    .A2(_1579_),
    .B1(net609),
    .Y(_1674_));
 sky130_fd_sc_hd__o311a_4 _4671_ (.A1(_1571_),
    .A2(_1577_),
    .A3(_1670_),
    .B1(_1674_),
    .C1(_1668_),
    .X(_1675_));
 sky130_fd_sc_hd__a211o_4 _4672_ (.A1(_1580_),
    .A2(_1667_),
    .B1(_1671_),
    .C1(_1673_),
    .X(_1676_));
 sky130_fd_sc_hd__nand3_2 _4673_ (.A(net111),
    .B(_1569_),
    .C(_1582_),
    .Y(_1677_));
 sky130_fd_sc_hd__nand4_4 _4674_ (.A(net111),
    .B(_1565_),
    .C(_1569_),
    .D(_1582_),
    .Y(_1678_));
 sky130_fd_sc_hd__nand3_2 _4675_ (.A(_1565_),
    .B(_1569_),
    .C(_1582_),
    .Y(_1679_));
 sky130_fd_sc_hd__a31o_2 _4676_ (.A1(_1565_),
    .A2(_1569_),
    .A3(_1582_),
    .B1(net111),
    .X(_1680_));
 sky130_fd_sc_hd__o2bb2ai_4 _4677_ (.A1_N(_0821_),
    .A2_N(_1679_),
    .B1(_1677_),
    .B2(_1566_),
    .Y(_1681_));
 sky130_fd_sc_hd__and3_4 _4678_ (.A(_1680_),
    .B(_1564_),
    .C(_1678_),
    .X(_1682_));
 sky130_fd_sc_hd__nand3_4 _4679_ (.A(_1680_),
    .B(_1564_),
    .C(_1678_),
    .Y(_1683_));
 sky130_fd_sc_hd__and3_1 _4680_ (.A(_1628_),
    .B(_1657_),
    .C(_1661_),
    .X(_1684_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_1628_),
    .B(_1662_),
    .Y(_1685_));
 sky130_fd_sc_hd__a21boi_4 _4682_ (.A1(_1588_),
    .A2(net111),
    .B1_N(_1563_),
    .Y(_1686_));
 sky130_fd_sc_hd__o21a_4 _4683_ (.A1(_1566_),
    .A2(_1589_),
    .B1(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__a21oi_4 _4684_ (.A1(net112),
    .A2(_1588_),
    .B1(_1596_),
    .Y(_1688_));
 sky130_fd_sc_hd__o21ai_4 _4685_ (.A1(_1588_),
    .A2(_1595_),
    .B1(_1597_),
    .Y(_1689_));
 sky130_fd_sc_hd__and3_4 _4686_ (.A(_1688_),
    .B(_1590_),
    .C(_1686_),
    .X(_1690_));
 sky130_fd_sc_hd__nand3_4 _4687_ (.A(_1688_),
    .B(_1590_),
    .C(_1686_),
    .Y(_1691_));
 sky130_fd_sc_hd__o21a_4 _4688_ (.A1(_1427_),
    .A2(_1562_),
    .B1(_1595_),
    .X(_1692_));
 sky130_fd_sc_hd__a21boi_4 _4689_ (.A1(_1678_),
    .A2(_1680_),
    .B1_N(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_8 _4690_ (.A(net400),
    .B(_1692_),
    .Y(_1694_));
 sky130_fd_sc_hd__and3_2 _4691_ (.A(net558),
    .B(_1681_),
    .C(_1692_),
    .X(_1695_));
 sky130_fd_sc_hd__nand3_4 _4692_ (.A(net558),
    .B(_1681_),
    .C(_1692_),
    .Y(_1696_));
 sky130_fd_sc_hd__a21oi_4 _4693_ (.A1(_1630_),
    .A2(_1638_),
    .B1(_1642_),
    .Y(_1697_));
 sky130_fd_sc_hd__nor4_4 _4694_ (.A(_1633_),
    .B(net427),
    .C(net460),
    .D(_1642_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_2 _4695_ (.A(_1637_),
    .B(_1697_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_1695_),
    .B(net396),
    .Y(_1700_));
 sky130_fd_sc_hd__and3_4 _4697_ (.A(net612),
    .B(_1669_),
    .C(_0828_),
    .X(_1701_));
 sky130_fd_sc_hd__nand3_4 _4698_ (.A(net612),
    .B(_1669_),
    .C(_0828_),
    .Y(_1702_));
 sky130_fd_sc_hd__nor3_4 _4699_ (.A(net620),
    .B(net561),
    .C(net615),
    .Y(_1703_));
 sky130_fd_sc_hd__nand2b_4 _4700_ (.A_N(net616),
    .B(net551),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_8 _4701_ (.A(net615),
    .B(net617),
    .Y(_1705_));
 sky130_fd_sc_hd__nor4_4 _4702_ (.A(net621),
    .B(net561),
    .C(net615),
    .D(net618),
    .Y(_1706_));
 sky130_fd_sc_hd__nand2_8 _4703_ (.A(net551),
    .B(_1705_),
    .Y(_1707_));
 sky130_fd_sc_hd__nor4_4 _4704_ (.A(net112),
    .B(net111),
    .C(net114),
    .D(net113),
    .Y(_1708_));
 sky130_fd_sc_hd__nand3b_1 _4705_ (.A_N(net112),
    .B(_1426_),
    .C(_0821_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_4 _4706_ (.A(net546),
    .B(net542),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_4 _4707_ (.A(_1701_),
    .B(net542),
    .Y(_1711_));
 sky130_fd_sc_hd__and3_4 _4708_ (.A(net615),
    .B(net617),
    .C(net551),
    .X(_1712_));
 sky130_fd_sc_hd__nand3_4 _4709_ (.A(net616),
    .B(net618),
    .C(_1610_),
    .Y(_1713_));
 sky130_fd_sc_hd__and3_2 _4710_ (.A(_1712_),
    .B(_0821_),
    .C(_1564_),
    .X(_1714_));
 sky130_fd_sc_hd__and2_2 _4711_ (.A(_1636_),
    .B(_1634_),
    .X(_1715_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(_1636_),
    .B(_1634_),
    .Y(_1716_));
 sky130_fd_sc_hd__a211o_2 _4713_ (.A1(_1630_),
    .A2(_1638_),
    .B1(_1642_),
    .C1(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__and2b_4 _4714_ (.A_N(net610),
    .B(net609),
    .X(_1718_));
 sky130_fd_sc_hd__nor4b_2 _4715_ (.A(net610),
    .B(net613),
    .C(net614),
    .D_N(net609),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_4 _4716_ (.A(_1606_),
    .B(_1718_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2_4 _4717_ (.A(net542),
    .B(net540),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _4718_ (.A(_1714_),
    .B(net539),
    .Y(_1722_));
 sky130_fd_sc_hd__and4bb_4 _4719_ (.A_N(net610),
    .B_N(net613),
    .C(net125),
    .D(net609),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_4 _4720_ (.A(_1641_),
    .B(_1718_),
    .Y(_1724_));
 sky130_fd_sc_hd__nor3_4 _4721_ (.A(net619),
    .B(net561),
    .C(_1603_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_8 _4722_ (.A(_1602_),
    .B(net551),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2_4 _4723_ (.A(net543),
    .B(net456),
    .Y(_1727_));
 sky130_fd_sc_hd__o21a_4 _4724_ (.A1(_1427_),
    .A2(_1562_),
    .B1(_1651_),
    .X(_1728_));
 sky130_fd_sc_hd__and4_1 _4725_ (.A(net401),
    .B(_1652_),
    .C(_1653_),
    .D(_1563_),
    .X(_1729_));
 sky130_fd_sc_hd__nand4_4 _4726_ (.A(net401),
    .B(_1652_),
    .C(_1653_),
    .D(_1563_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_4 _4727_ (.A(net542),
    .B(_1723_),
    .Y(_1731_));
 sky130_fd_sc_hd__and3_1 _4728_ (.A(net542),
    .B(_1723_),
    .C(net455),
    .X(_1732_));
 sky130_fd_sc_hd__and4b_2 _4729_ (.A_N(net611),
    .B(_1637_),
    .C(_1638_),
    .D(_1630_),
    .X(_1733_));
 sky130_fd_sc_hd__nand3b_4 _4730_ (.A_N(net611),
    .B(_1637_),
    .C(_1639_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_1687_),
    .B(_1689_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand4_4 _4732_ (.A(net558),
    .B(_1689_),
    .C(_1591_),
    .D(_1563_),
    .Y(_1736_));
 sky130_fd_sc_hd__and3_4 _4733_ (.A(_1630_),
    .B(_1638_),
    .C(net611),
    .X(_1737_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(net612),
    .B(net460),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_1715_),
    .B(_1737_),
    .Y(_1739_));
 sky130_fd_sc_hd__and3b_4 _4736_ (.A_N(net610),
    .B(net609),
    .C(net613),
    .X(_1740_));
 sky130_fd_sc_hd__nand2_4 _4737_ (.A(_1570_),
    .B(_1718_),
    .Y(_1741_));
 sky130_fd_sc_hd__o32a_1 _4738_ (.A1(_1710_),
    .A2(_1716_),
    .A3(_1738_),
    .B1(_1741_),
    .B2(_1727_),
    .X(_1742_));
 sky130_fd_sc_hd__o21a_1 _4739_ (.A1(_1734_),
    .A2(_1736_),
    .B1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__and4bb_4 _4740_ (.A_N(net127),
    .B_N(net125),
    .C(net613),
    .D(net609),
    .X(_1744_));
 sky130_fd_sc_hd__nand2_8 _4741_ (.A(_1740_),
    .B(_0828_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2b_4 _4742_ (.A_N(net615),
    .B(net617),
    .Y(_1746_));
 sky130_fd_sc_hd__nor3_2 _4743_ (.A(net620),
    .B(net561),
    .C(_1746_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_4 _4744_ (.A(net618),
    .B(_1703_),
    .Y(_1748_));
 sky130_fd_sc_hd__and3_1 _4745_ (.A(_1570_),
    .B(_1718_),
    .C(net453),
    .X(_1749_));
 sky130_fd_sc_hd__nand4_1 _4746_ (.A(_1591_),
    .B(_1688_),
    .C(_1749_),
    .D(_1563_),
    .Y(_1750_));
 sky130_fd_sc_hd__and4b_4 _4747_ (.A_N(net621),
    .B(net562),
    .C(net616),
    .D(net618),
    .X(_1751_));
 sky130_fd_sc_hd__nand3_4 _4748_ (.A(net616),
    .B(net618),
    .C(_1600_),
    .Y(_1752_));
 sky130_fd_sc_hd__a21oi_2 _4749_ (.A1(_0828_),
    .A2(_1612_),
    .B1(_1615_),
    .Y(_1753_));
 sky130_fd_sc_hd__and3_2 _4750_ (.A(_1606_),
    .B(_1607_),
    .C(_1751_),
    .X(_1754_));
 sky130_fd_sc_hd__a221oi_2 _4751_ (.A1(_1608_),
    .A2(_1628_),
    .B1(net455),
    .B2(_1744_),
    .C1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__o221a_1 _4752_ (.A1(_1710_),
    .A2(_1745_),
    .B1(_1755_),
    .B2(_1691_),
    .C1(_1750_),
    .X(_1756_));
 sky130_fd_sc_hd__and3_2 _4753_ (.A(_1644_),
    .B(_1634_),
    .C(_1636_),
    .X(_1757_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_1714_),
    .B(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand4_4 _4755_ (.A(_1591_),
    .B(_1688_),
    .C(net453),
    .D(_1563_),
    .Y(_1759_));
 sky130_fd_sc_hd__and3_1 _4756_ (.A(net558),
    .B(net555),
    .C(net542),
    .X(_1760_));
 sky130_fd_sc_hd__o22a_1 _4757_ (.A1(_1696_),
    .A2(_1734_),
    .B1(_1745_),
    .B2(_1759_),
    .X(_1761_));
 sky130_fd_sc_hd__and3_4 _4758_ (.A(_1628_),
    .B(_1681_),
    .C(_1692_),
    .X(_1762_));
 sky130_fd_sc_hd__nand2_8 _4759_ (.A(_1628_),
    .B(net397),
    .Y(_1763_));
 sky130_fd_sc_hd__nand4_1 _4760_ (.A(_1743_),
    .B(_1756_),
    .C(_1761_),
    .D(_1758_),
    .Y(_1764_));
 sky130_fd_sc_hd__nand3b_4 _4761_ (.A_N(net612),
    .B(net460),
    .C(_1715_),
    .Y(_1765_));
 sky130_fd_sc_hd__and4b_1 _4762_ (.A_N(net612),
    .B(net460),
    .C(_1714_),
    .D(_1715_),
    .X(_1766_));
 sky130_fd_sc_hd__nor3_1 _4763_ (.A(_1732_),
    .B(_1766_),
    .C(_1764_),
    .Y(_1767_));
 sky130_fd_sc_hd__o211ai_1 _4764_ (.A1(_1704_),
    .A2(_1731_),
    .B1(_1722_),
    .C1(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__and3_1 _4765_ (.A(net542),
    .B(net539),
    .C(net455),
    .X(_1769_));
 sky130_fd_sc_hd__nor2_1 _4766_ (.A(_1769_),
    .B(_1768_),
    .Y(_1770_));
 sky130_fd_sc_hd__nor2_8 _4767_ (.A(net128),
    .B(_1634_),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2b_1 _4768_ (.A_N(net609),
    .B(_1633_),
    .Y(_1772_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_1737_),
    .B(_1771_),
    .Y(_1773_));
 sky130_fd_sc_hd__nand4_1 _4770_ (.A(net543),
    .B(_1712_),
    .C(_1737_),
    .D(_1771_),
    .Y(_1774_));
 sky130_fd_sc_hd__o211ai_1 _4771_ (.A1(_1704_),
    .A2(_1721_),
    .B1(_1774_),
    .C1(_1770_),
    .Y(_1775_));
 sky130_fd_sc_hd__and3_4 _4772_ (.A(net612),
    .B(net125),
    .C(_1669_),
    .X(_1776_));
 sky130_fd_sc_hd__and3_2 _4773_ (.A(_1570_),
    .B(_1669_),
    .C(net542),
    .X(_1777_));
 sky130_fd_sc_hd__nand2_4 _4774_ (.A(net543),
    .B(_1776_),
    .Y(_1778_));
 sky130_fd_sc_hd__and3_1 _4775_ (.A(net543),
    .B(net455),
    .C(_1776_),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_1 _4776_ (.A(_1779_),
    .B(_1775_),
    .Y(_1780_));
 sky130_fd_sc_hd__a211o_1 _4777_ (.A1(_1630_),
    .A2(_1638_),
    .B1(_1643_),
    .C1(_1772_),
    .X(_1781_));
 sky130_fd_sc_hd__nand4_1 _4778_ (.A(_1644_),
    .B(net543),
    .C(_1712_),
    .D(_1771_),
    .Y(_1782_));
 sky130_fd_sc_hd__o211ai_1 _4779_ (.A1(_1704_),
    .A2(_1778_),
    .B1(_1782_),
    .C1(_1780_),
    .Y(_1783_));
 sky130_fd_sc_hd__and3_1 _4780_ (.A(_1701_),
    .B(net543),
    .C(net455),
    .X(_1784_));
 sky130_fd_sc_hd__nor2_1 _4781_ (.A(_1784_),
    .B(_1783_),
    .Y(_1785_));
 sky130_fd_sc_hd__and4b_1 _4782_ (.A_N(net612),
    .B(net460),
    .C(_1690_),
    .D(_1771_),
    .X(_1786_));
 sky130_fd_sc_hd__nand4b_4 _4783_ (.A_N(net612),
    .B(net460),
    .C(_1690_),
    .D(_1771_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_1 _4784_ (.A(_1712_),
    .B(_1786_),
    .Y(_1788_));
 sky130_fd_sc_hd__o211ai_1 _4785_ (.A1(_1704_),
    .A2(_1711_),
    .B1(_1788_),
    .C1(_1785_),
    .Y(_1789_));
 sky130_fd_sc_hd__and4bb_4 _4786_ (.A_N(net609),
    .B_N(net612),
    .C(net125),
    .D(net610),
    .X(_1790_));
 sky130_fd_sc_hd__nand2_1 _4787_ (.A(_1641_),
    .B(_1669_),
    .Y(_1791_));
 sky130_fd_sc_hd__and3_4 _4788_ (.A(_1790_),
    .B(_0821_),
    .C(net560),
    .X(_1792_));
 sky130_fd_sc_hd__nand2_2 _4789_ (.A(net543),
    .B(_1790_),
    .Y(_1793_));
 sky130_fd_sc_hd__and3_1 _4790_ (.A(net543),
    .B(net455),
    .C(_1790_),
    .X(_1794_));
 sky130_fd_sc_hd__nor2_1 _4791_ (.A(_1794_),
    .B(_1789_),
    .Y(_1795_));
 sky130_fd_sc_hd__o21ai_1 _4792_ (.A1(_1704_),
    .A2(_1793_),
    .B1(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_1697_),
    .B(_1771_),
    .Y(_1797_));
 sky130_fd_sc_hd__and3_1 _4794_ (.A(_1697_),
    .B(_1714_),
    .C(_1771_),
    .X(_1798_));
 sky130_fd_sc_hd__and4bb_4 _4795_ (.A_N(net609),
    .B_N(net611),
    .C(net610),
    .D(_0828_),
    .X(_1799_));
 sky130_fd_sc_hd__nand2_4 _4796_ (.A(_1606_),
    .B(_1669_),
    .Y(_1800_));
 sky130_fd_sc_hd__and3_1 _4797_ (.A(_1606_),
    .B(_1669_),
    .C(net542),
    .X(_1801_));
 sky130_fd_sc_hd__nand2_4 _4798_ (.A(net543),
    .B(_1799_),
    .Y(_1802_));
 sky130_fd_sc_hd__and3_1 _4799_ (.A(net543),
    .B(net456),
    .C(_1799_),
    .X(_1803_));
 sky130_fd_sc_hd__nor3_1 _4800_ (.A(_1798_),
    .B(_1803_),
    .C(_1796_),
    .Y(_1804_));
 sky130_fd_sc_hd__and3_2 _4801_ (.A(_1637_),
    .B(net460),
    .C(_1642_),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_1 _4802_ (.A(_1637_),
    .B(_1737_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _4803_ (.A(_1714_),
    .B(_1805_),
    .Y(_1807_));
 sky130_fd_sc_hd__o211ai_1 _4804_ (.A1(_1704_),
    .A2(_1802_),
    .B1(_1807_),
    .C1(_1804_),
    .Y(_1808_));
 sky130_fd_sc_hd__and3_4 _4805_ (.A(net611),
    .B(net614),
    .C(_1607_),
    .X(_1809_));
 sky130_fd_sc_hd__nand2_2 _4806_ (.A(_1570_),
    .B(_1607_),
    .Y(_1810_));
 sky130_fd_sc_hd__and3_1 _4807_ (.A(_1690_),
    .B(net456),
    .C(_1809_),
    .X(_1811_));
 sky130_fd_sc_hd__and3_1 _4808_ (.A(_1690_),
    .B(net454),
    .C(_1809_),
    .X(_1812_));
 sky130_fd_sc_hd__nor3_1 _4809_ (.A(_1811_),
    .B(_1812_),
    .C(_1808_),
    .Y(_1813_));
 sky130_fd_sc_hd__nand4_1 _4810_ (.A(_1687_),
    .B(_1688_),
    .C(net549),
    .D(_1809_),
    .Y(_1814_));
 sky130_fd_sc_hd__nand4_1 _4811_ (.A(_1645_),
    .B(_1687_),
    .C(_1688_),
    .D(_1712_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand3_1 _4812_ (.A(_1813_),
    .B(_1814_),
    .C(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__and3_4 _4813_ (.A(net611),
    .B(_1607_),
    .C(_0828_),
    .X(_1817_));
 sky130_fd_sc_hd__nand3_4 _4814_ (.A(net613),
    .B(_1607_),
    .C(_0828_),
    .Y(_1818_));
 sky130_fd_sc_hd__and3_1 _4815_ (.A(net543),
    .B(net456),
    .C(_1817_),
    .X(_1819_));
 sky130_fd_sc_hd__and3_1 _4816_ (.A(_1690_),
    .B(net454),
    .C(_1817_),
    .X(_1820_));
 sky130_fd_sc_hd__and3_1 _4817_ (.A(_1817_),
    .B(_0821_),
    .C(net560),
    .X(_1821_));
 sky130_fd_sc_hd__nor3_1 _4818_ (.A(_1819_),
    .B(_1820_),
    .C(_1816_),
    .Y(_1822_));
 sky130_fd_sc_hd__and3b_4 _4819_ (.A_N(net615),
    .B(net561),
    .C(net619),
    .X(_1823_));
 sky130_fd_sc_hd__and3_4 _4820_ (.A(net619),
    .B(net561),
    .C(_1705_),
    .X(_1824_));
 sky130_fd_sc_hd__nand3_4 _4821_ (.A(net619),
    .B(net561),
    .C(_1705_),
    .Y(_1825_));
 sky130_fd_sc_hd__nand4_4 _4822_ (.A(_1687_),
    .B(_1698_),
    .C(_1824_),
    .D(_1689_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand4_1 _4823_ (.A(_1592_),
    .B(_1805_),
    .C(net560),
    .D(net558),
    .Y(_1827_));
 sky130_fd_sc_hd__nand4_1 _4824_ (.A(_1822_),
    .B(_1826_),
    .C(_1827_),
    .D(_1700_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor4_2 _4825_ (.A(net112),
    .B(net114),
    .C(net113),
    .D(_0821_),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_8 _4826_ (.A(_1426_),
    .B(_1593_),
    .Y(_1830_));
 sky130_fd_sc_hd__and3_1 _4827_ (.A(_1426_),
    .B(_1593_),
    .C(_1817_),
    .X(_1831_));
 sky130_fd_sc_hd__nand2_1 _4828_ (.A(_1817_),
    .B(net451),
    .Y(_1832_));
 sky130_fd_sc_hd__and3_1 _4829_ (.A(_1751_),
    .B(_1817_),
    .C(net452),
    .X(_1833_));
 sky130_fd_sc_hd__nor3_1 _4830_ (.A(_1684_),
    .B(_1833_),
    .C(_1828_),
    .Y(_1834_));
 sky130_fd_sc_hd__nor4b_4 _4831_ (.A(net127),
    .B(net128),
    .C(net613),
    .D_N(net125),
    .Y(_1835_));
 sky130_fd_sc_hd__nand2_8 _4832_ (.A(_1607_),
    .B(_1641_),
    .Y(_1836_));
 sky130_fd_sc_hd__and3_1 _4833_ (.A(net559),
    .B(_1733_),
    .C(_1592_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_2 _4834_ (.A(net363),
    .B(_1733_),
    .Y(_1838_));
 sky130_fd_sc_hd__o32a_1 _4835_ (.A1(_1586_),
    .A2(_1599_),
    .A3(_1836_),
    .B1(_1838_),
    .B2(_1629_),
    .X(_1839_));
 sky130_fd_sc_hd__nand4_1 _4836_ (.A(net364),
    .B(_1607_),
    .C(_1641_),
    .D(_1751_),
    .Y(_1840_));
 sky130_fd_sc_hd__nand3_1 _4837_ (.A(_1834_),
    .B(_1839_),
    .C(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__and4_1 _4838_ (.A(net619),
    .B(net561),
    .C(net617),
    .D(_1837_),
    .X(_1842_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_1823_),
    .B(_1837_),
    .Y(_1843_));
 sky130_fd_sc_hd__and4b_4 _4840_ (.A_N(net615),
    .B(net617),
    .C(net619),
    .D(net561),
    .X(_1844_));
 sky130_fd_sc_hd__nor3_1 _4841_ (.A(_1627_),
    .B(_1842_),
    .C(_1841_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2b_4 _4842_ (.A_N(net616),
    .B(net556),
    .Y(_1846_));
 sky130_fd_sc_hd__nor2_8 _4843_ (.A(_1601_),
    .B(_1746_),
    .Y(_1847_));
 sky130_fd_sc_hd__nand3b_4 _4844_ (.A_N(net616),
    .B(net618),
    .C(net556),
    .Y(_1848_));
 sky130_fd_sc_hd__and3_1 _4845_ (.A(_1426_),
    .B(_1593_),
    .C(net552),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_4 _4846_ (.A(net552),
    .B(net449),
    .Y(_1850_));
 sky130_fd_sc_hd__and3_2 _4847_ (.A(net552),
    .B(net451),
    .C(_1847_),
    .X(_1851_));
 sky130_fd_sc_hd__a31oi_1 _4848_ (.A1(net362),
    .A2(net395),
    .A3(net535),
    .B1(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__and3_1 _4849_ (.A(_1682_),
    .B(net395),
    .C(_1824_),
    .X(_1853_));
 sky130_fd_sc_hd__nand4_4 _4850_ (.A(net559),
    .B(net396),
    .C(_1824_),
    .D(_1592_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand3_1 _4851_ (.A(_1845_),
    .B(_1852_),
    .C(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__o31a_4 _4852_ (.A1(_1586_),
    .A2(_1599_),
    .A3(_1699_),
    .B1(\wbbd_state[9] ),
    .X(_1856_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_1657_),
    .B(_1751_),
    .Y(_1857_));
 sky130_fd_sc_hd__o31a_2 _4854_ (.A1(_1626_),
    .A2(_1658_),
    .A3(_1752_),
    .B1(\wbbd_state[10] ),
    .X(_1858_));
 sky130_fd_sc_hd__o2111ai_4 _4855_ (.A1(_1648_),
    .A2(_1650_),
    .B1(_1656_),
    .C1(_1844_),
    .D1(_1625_),
    .Y(_1859_));
 sky130_fd_sc_hd__nor3b_2 _4856_ (.A(net561),
    .B(net615),
    .C_N(net619),
    .Y(_1860_));
 sky130_fd_sc_hd__and3b_4 _4857_ (.A_N(net561),
    .B(_1705_),
    .C(net619),
    .X(_1861_));
 sky130_fd_sc_hd__nand3b_4 _4858_ (.A_N(net561),
    .B(_1705_),
    .C(net619),
    .Y(_1862_));
 sky130_fd_sc_hd__and3_1 _4859_ (.A(_1661_),
    .B(net361),
    .C(_1861_),
    .X(_1863_));
 sky130_fd_sc_hd__nor2_4 _4860_ (.A(net128),
    .B(_1623_),
    .Y(_1864_));
 sky130_fd_sc_hd__and4_4 _4861_ (.A(_1580_),
    .B(_1667_),
    .C(_1672_),
    .D(_1674_),
    .X(_1865_));
 sky130_fd_sc_hd__a311o_2 _4862_ (.A1(net611),
    .A2(_1578_),
    .A3(_1669_),
    .B1(_1673_),
    .C1(_1668_),
    .X(_1866_));
 sky130_fd_sc_hd__o21a_4 _4863_ (.A1(net614),
    .A2(_1576_),
    .B1(_1664_),
    .X(_1867_));
 sky130_fd_sc_hd__and3_4 _4864_ (.A(net400),
    .B(_1692_),
    .C(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(net397),
    .B(_1867_),
    .Y(_1869_));
 sky130_fd_sc_hd__and3_1 _4866_ (.A(net448),
    .B(net394),
    .C(_1868_),
    .X(_1870_));
 sky130_fd_sc_hd__and3_2 _4867_ (.A(net429),
    .B(_1654_),
    .C(_1728_),
    .X(_1871_));
 sky130_fd_sc_hd__o311a_4 _4868_ (.A1(_1575_),
    .A2(_1584_),
    .A3(_1610_),
    .B1(_1621_),
    .C1(_1623_),
    .X(_1872_));
 sky130_fd_sc_hd__o211ai_4 _4869_ (.A1(_1584_),
    .A2(net550),
    .B1(_1621_),
    .C1(_1623_),
    .Y(_1873_));
 sky130_fd_sc_hd__and3_4 _4870_ (.A(net429),
    .B(net360),
    .C(_1872_),
    .X(_1874_));
 sky130_fd_sc_hd__and4bb_4 _4871_ (.A_N(net562),
    .B_N(net618),
    .C(net616),
    .D(net621),
    .X(_1875_));
 sky130_fd_sc_hd__nand3b_4 _4872_ (.A_N(net561),
    .B(_1602_),
    .C(net619),
    .Y(_1876_));
 sky130_fd_sc_hd__o22a_4 _4873_ (.A1(_1571_),
    .A2(_1577_),
    .B1(net611),
    .B2(_1665_),
    .X(_1877_));
 sky130_fd_sc_hd__a2bb2o_4 _4874_ (.A1_N(net611),
    .A2_N(_1665_),
    .B1(_1576_),
    .B2(_1570_),
    .X(_1878_));
 sky130_fd_sc_hd__and3_4 _4875_ (.A(net400),
    .B(_1692_),
    .C(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a22oi_4 _4876_ (.A1(_1580_),
    .A2(_1667_),
    .B1(_1672_),
    .B2(_1674_),
    .Y(_1880_));
 sky130_fd_sc_hd__nand2_4 _4877_ (.A(_1874_),
    .B(net532),
    .Y(_1881_));
 sky130_fd_sc_hd__nand4_1 _4878_ (.A(net360),
    .B(net426),
    .C(net448),
    .D(_1872_),
    .Y(_1882_));
 sky130_fd_sc_hd__and4bb_4 _4879_ (.A_N(net562),
    .B_N(net616),
    .C(net618),
    .D(net621),
    .X(_1883_));
 sky130_fd_sc_hd__nand2_4 _4880_ (.A(net617),
    .B(net534),
    .Y(_1884_));
 sky130_fd_sc_hd__and3_2 _4881_ (.A(_1654_),
    .B(_1728_),
    .C(_1883_),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(net399),
    .B(_1883_),
    .Y(_1886_));
 sky130_fd_sc_hd__and3_2 _4883_ (.A(_1868_),
    .B(_1880_),
    .C(_1883_),
    .X(_1887_));
 sky130_fd_sc_hd__nand4_2 _4884_ (.A(net360),
    .B(_1753_),
    .C(_1872_),
    .D(_1875_),
    .Y(_1888_));
 sky130_fd_sc_hd__and3_1 _4885_ (.A(_1604_),
    .B(_1654_),
    .C(_1728_),
    .X(_1889_));
 sky130_fd_sc_hd__nand2_2 _4886_ (.A(_1604_),
    .B(net360),
    .Y(_1890_));
 sky130_fd_sc_hd__and4b_4 _4887_ (.A_N(net562),
    .B(net616),
    .C(net121),
    .D(net621),
    .X(_1891_));
 sky130_fd_sc_hd__nand4b_4 _4888_ (.A_N(net561),
    .B(net615),
    .C(net617),
    .D(net619),
    .Y(_1892_));
 sky130_fd_sc_hd__nor2_2 _4889_ (.A(_1660_),
    .B(_1873_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand4_2 _4890_ (.A(net401),
    .B(_1656_),
    .C(net531),
    .D(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand4_1 _4891_ (.A(net401),
    .B(_1656_),
    .C(_1875_),
    .D(_1893_),
    .Y(_1895_));
 sky130_fd_sc_hd__and3_4 _4892_ (.A(_1616_),
    .B(net613),
    .C(_1613_),
    .X(_1896_));
 sky130_fd_sc_hd__nand2_1 _4893_ (.A(net397),
    .B(net531),
    .Y(_1897_));
 sky130_fd_sc_hd__nand4_1 _4894_ (.A(net399),
    .B(_1872_),
    .C(net531),
    .D(_1896_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand4_2 _4895_ (.A(_1654_),
    .B(_1563_),
    .C(net401),
    .D(_1754_),
    .Y(_1899_));
 sky130_fd_sc_hd__nand4_4 _4896_ (.A(_1625_),
    .B(_1628_),
    .C(net401),
    .D(_1656_),
    .Y(_1900_));
 sky130_fd_sc_hd__o31a_1 _4897_ (.A1(_1626_),
    .A2(_1629_),
    .A3(_1730_),
    .B1(_1899_),
    .X(_1901_));
 sky130_fd_sc_hd__nand4_4 _4898_ (.A(_1563_),
    .B(_1655_),
    .C(_1754_),
    .D(net401),
    .Y(_1902_));
 sky130_fd_sc_hd__o2111ai_2 _4899_ (.A1(_1571_),
    .A2(_1612_),
    .B1(_1615_),
    .C1(net533),
    .D1(_1872_),
    .Y(_1903_));
 sky130_fd_sc_hd__o311a_1 _4900_ (.A1(_1605_),
    .A2(_1626_),
    .A3(_1730_),
    .B1(_1899_),
    .C1(_1900_),
    .X(_1904_));
 sky130_fd_sc_hd__o2111a_1 _4901_ (.A1(_1730_),
    .A2(_1903_),
    .B1(_1902_),
    .C1(_1898_),
    .D1(_1895_),
    .X(_1905_));
 sky130_fd_sc_hd__nand4_1 _4902_ (.A(_1904_),
    .B(_1905_),
    .C(_1888_),
    .D(_1894_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand4_1 _4903_ (.A(net360),
    .B(_1872_),
    .C(net531),
    .D(_1896_),
    .Y(_1907_));
 sky130_fd_sc_hd__nor2_1 _4904_ (.A(_1887_),
    .B(_1906_),
    .Y(_1908_));
 sky130_fd_sc_hd__nand4_2 _4905_ (.A(net360),
    .B(net426),
    .C(_1872_),
    .D(net531),
    .Y(_1909_));
 sky130_fd_sc_hd__nand4_1 _4906_ (.A(_1908_),
    .B(_1909_),
    .C(_1881_),
    .D(_1882_),
    .Y(_1910_));
 sky130_fd_sc_hd__and3_1 _4907_ (.A(_1871_),
    .B(_1872_),
    .C(net531),
    .X(_1911_));
 sky130_fd_sc_hd__a211oi_1 _4908_ (.A1(net533),
    .A2(_1874_),
    .B1(_1911_),
    .C1(_1910_),
    .Y(_1912_));
 sky130_fd_sc_hd__and4_2 _4909_ (.A(_1613_),
    .B(net394),
    .C(_1616_),
    .D(net613),
    .X(_1913_));
 sky130_fd_sc_hd__and4b_2 _4910_ (.A_N(net561),
    .B(_1602_),
    .C(net394),
    .D(net619),
    .X(_1914_));
 sky130_fd_sc_hd__nand4_4 _4911_ (.A(net360),
    .B(net394),
    .C(net532),
    .D(_1896_),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(_1885_),
    .B(_1913_),
    .Y(_1916_));
 sky130_fd_sc_hd__nand3_1 _4913_ (.A(_1912_),
    .B(_1915_),
    .C(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__and4_1 _4914_ (.A(net360),
    .B(net448),
    .C(net394),
    .D(_1896_),
    .X(_1918_));
 sky130_fd_sc_hd__and3_1 _4915_ (.A(net360),
    .B(net531),
    .C(_1913_),
    .X(_1919_));
 sky130_fd_sc_hd__nor3_1 _4916_ (.A(_1918_),
    .B(_1919_),
    .C(_1917_),
    .Y(_1920_));
 sky130_fd_sc_hd__nand4_2 _4917_ (.A(_1659_),
    .B(net360),
    .C(net394),
    .D(_1875_),
    .Y(_1921_));
 sky130_fd_sc_hd__nand4_1 _4918_ (.A(_1659_),
    .B(net399),
    .C(net394),
    .D(_1883_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand3_1 _4919_ (.A(_1920_),
    .B(_1921_),
    .C(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__and4_1 _4920_ (.A(_1659_),
    .B(net360),
    .C(net448),
    .D(net394),
    .X(_1924_));
 sky130_fd_sc_hd__and4_1 _4921_ (.A(_1659_),
    .B(net399),
    .C(net394),
    .D(net531),
    .X(_1925_));
 sky130_fd_sc_hd__nor3_1 _4922_ (.A(_1924_),
    .B(_1925_),
    .C(_1923_),
    .Y(_1926_));
 sky130_fd_sc_hd__nand4_1 _4923_ (.A(net361),
    .B(net426),
    .C(net394),
    .D(_1875_),
    .Y(_1927_));
 sky130_fd_sc_hd__nand4_2 _4924_ (.A(net398),
    .B(net394),
    .C(_1867_),
    .D(_1883_),
    .Y(_1928_));
 sky130_fd_sc_hd__nand3_1 _4925_ (.A(_1926_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__and4_1 _4926_ (.A(net399),
    .B(net426),
    .C(net394),
    .D(net531),
    .X(_1930_));
 sky130_fd_sc_hd__nor3_1 _4927_ (.A(_1870_),
    .B(_1930_),
    .C(_1929_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_1871_),
    .B(_1914_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand3_1 _4929_ (.A(net394),
    .B(_1879_),
    .C(_1883_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand3_1 _4930_ (.A(_1931_),
    .B(_1932_),
    .C(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__and3_1 _4931_ (.A(net448),
    .B(_1864_),
    .C(_1871_),
    .X(_1935_));
 sky130_fd_sc_hd__and4_1 _4932_ (.A(net429),
    .B(net399),
    .C(_1864_),
    .D(_1891_),
    .X(_1936_));
 sky130_fd_sc_hd__and3_1 _4933_ (.A(_1864_),
    .B(_1871_),
    .C(net531),
    .X(_1937_));
 sky130_fd_sc_hd__nor3_1 _4934_ (.A(_1935_),
    .B(_1937_),
    .C(_1934_),
    .Y(_1938_));
 sky130_fd_sc_hd__and3_1 _4935_ (.A(net428),
    .B(net361),
    .C(_1896_),
    .X(_1939_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(net428),
    .B(_1896_),
    .Y(_1940_));
 sky130_fd_sc_hd__nand4_1 _4937_ (.A(net428),
    .B(net361),
    .C(_1875_),
    .D(_1896_),
    .Y(_1941_));
 sky130_fd_sc_hd__o211ai_1 _4938_ (.A1(_1886_),
    .A2(_1940_),
    .B1(_1941_),
    .C1(_1938_),
    .Y(_1942_));
 sky130_fd_sc_hd__and4_1 _4939_ (.A(net428),
    .B(net361),
    .C(net448),
    .D(_1896_),
    .X(_1943_));
 sky130_fd_sc_hd__and4_1 _4940_ (.A(net428),
    .B(net361),
    .C(_1891_),
    .D(_1896_),
    .X(_1944_));
 sky130_fd_sc_hd__nor3_1 _4941_ (.A(_1943_),
    .B(_1944_),
    .C(_1942_),
    .Y(_1945_));
 sky130_fd_sc_hd__nand4_1 _4942_ (.A(_1654_),
    .B(_1661_),
    .C(_1728_),
    .D(net532),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _4943_ (.A(_1661_),
    .B(_1885_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand3_1 _4944_ (.A(_1945_),
    .B(_1946_),
    .C(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nor2_8 _4945_ (.A(net121),
    .B(_1846_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_8 _4946_ (.A(net556),
    .B(_1705_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand4_4 _4947_ (.A(_1655_),
    .B(_1728_),
    .C(net429),
    .D(net428),
    .Y(_1951_));
 sky130_fd_sc_hd__and4_1 _4948_ (.A(_1625_),
    .B(_1655_),
    .C(_1728_),
    .D(_1949_),
    .X(_1952_));
 sky130_fd_sc_hd__nor3_1 _4949_ (.A(_1863_),
    .B(_1952_),
    .C(_1948_),
    .Y(_1953_));
 sky130_fd_sc_hd__nand4_1 _4950_ (.A(_1625_),
    .B(net401),
    .C(_1656_),
    .D(_1751_),
    .Y(_1954_));
 sky130_fd_sc_hd__o2111a_1 _4951_ (.A1(_1857_),
    .A2(_1940_),
    .B1(_1954_),
    .C1(_1685_),
    .D1(_1953_),
    .X(_1955_));
 sky130_fd_sc_hd__nand2_1 _4952_ (.A(_1604_),
    .B(_1662_),
    .Y(_1956_));
 sky130_fd_sc_hd__and3_4 _4953_ (.A(net428),
    .B(_1657_),
    .C(net426),
    .X(_1957_));
 sky130_fd_sc_hd__nand3_4 _4954_ (.A(net428),
    .B(_1657_),
    .C(net426),
    .Y(_1958_));
 sky130_fd_sc_hd__a32o_1 _4955_ (.A1(_1657_),
    .A2(_1661_),
    .A3(_1751_),
    .B1(_1957_),
    .B2(_1604_),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_2 _4956_ (.A(_1629_),
    .B(_1876_),
    .Y(_1960_));
 sky130_fd_sc_hd__a21oi_1 _4957_ (.A1(_1957_),
    .A2(_1960_),
    .B1(_1959_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand3_1 _4958_ (.A(_1955_),
    .B(_1956_),
    .C(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a32o_1 _4959_ (.A1(_1657_),
    .A2(_1661_),
    .A3(_1847_),
    .B1(_1957_),
    .B2(_1712_),
    .X(_1963_));
 sky130_fd_sc_hd__nor2_1 _4960_ (.A(_1846_),
    .B(_1958_),
    .Y(_1964_));
 sky130_fd_sc_hd__a211oi_1 _4961_ (.A1(net532),
    .A2(_1957_),
    .B1(_1964_),
    .C1(_1963_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(_1962_),
    .B(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__a21o_1 _4963_ (.A1(_1575_),
    .A2(_1746_),
    .B1(_1601_),
    .X(_1967_));
 sky130_fd_sc_hd__o211ai_4 _4964_ (.A1(_1967_),
    .A2(_1958_),
    .B1(_1859_),
    .C1(_1966_),
    .Y(_1968_));
 sky130_fd_sc_hd__a31o_1 _4965_ (.A1(_1625_),
    .A2(_1682_),
    .A3(_1824_),
    .B1(_1851_),
    .X(_1969_));
 sky130_fd_sc_hd__and3_1 _4966_ (.A(_1625_),
    .B(_1657_),
    .C(_1949_),
    .X(_1970_));
 sky130_fd_sc_hd__o31ai_4 _4967_ (.A1(_1970_),
    .A2(_1969_),
    .A3(_1968_),
    .B1(_1858_),
    .Y(_1971_));
 sky130_fd_sc_hd__o41a_1 _4968_ (.A1(_1877_),
    .A2(net530),
    .A3(_1676_),
    .A4(_1683_),
    .B1(\wbbd_state[8] ),
    .X(_1972_));
 sky130_fd_sc_hd__o41ai_4 _4969_ (.A1(_1877_),
    .A2(net530),
    .A3(_1676_),
    .A4(_1683_),
    .B1(\wbbd_state[8] ),
    .Y(_1973_));
 sky130_fd_sc_hd__and3_1 _4970_ (.A(_1657_),
    .B(_1661_),
    .C(net532),
    .X(_1974_));
 sky130_fd_sc_hd__o21a_4 _4971_ (.A1(_1575_),
    .A2(_1601_),
    .B1(_1713_),
    .X(_1975_));
 sky130_fd_sc_hd__o211a_2 _4972_ (.A1(_1712_),
    .A2(_1751_),
    .B1(_1817_),
    .C1(net449),
    .X(_1976_));
 sky130_fd_sc_hd__a211o_2 _4973_ (.A1(_1713_),
    .A2(_1752_),
    .B1(_1818_),
    .C1(_1830_),
    .X(_1977_));
 sky130_fd_sc_hd__and4_1 _4974_ (.A(_1666_),
    .B(_1668_),
    .C(_1672_),
    .D(_1674_),
    .X(_1978_));
 sky130_fd_sc_hd__a211o_1 _4975_ (.A1(net611),
    .A2(_1665_),
    .B1(_1664_),
    .C1(_1676_),
    .X(_1979_));
 sky130_fd_sc_hd__a211o_1 _4976_ (.A1(_1629_),
    .A2(_1876_),
    .B1(_1979_),
    .C1(_1830_),
    .X(_1980_));
 sky130_fd_sc_hd__and3_2 _4977_ (.A(_1687_),
    .B(_1688_),
    .C(_1824_),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_2 _4978_ (.A(_1690_),
    .B(_1824_),
    .Y(_1982_));
 sky130_fd_sc_hd__and3_2 _4979_ (.A(_1666_),
    .B(net400),
    .C(_1692_),
    .X(_1983_));
 sky130_fd_sc_hd__a211o_1 _4980_ (.A1(net611),
    .A2(_1665_),
    .B1(_1664_),
    .C1(_1694_),
    .X(_1984_));
 sky130_fd_sc_hd__and3_2 _4981_ (.A(_1675_),
    .B(_1824_),
    .C(_1983_),
    .X(_1985_));
 sky130_fd_sc_hd__nand4_2 _4982_ (.A(_1666_),
    .B(_1675_),
    .C(net398),
    .D(net535),
    .Y(_1986_));
 sky130_fd_sc_hd__and3_1 _4983_ (.A(net558),
    .B(net398),
    .C(_1817_),
    .X(_1987_));
 sky130_fd_sc_hd__and3_4 _4984_ (.A(_1665_),
    .B(net611),
    .C(_1579_),
    .X(_1988_));
 sky130_fd_sc_hd__and3_4 _4985_ (.A(net400),
    .B(_1692_),
    .C(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(net398),
    .B(_1988_),
    .Y(_1990_));
 sky130_fd_sc_hd__nand4_1 _4987_ (.A(_1675_),
    .B(net397),
    .C(_1824_),
    .D(_1988_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand4_1 _4988_ (.A(_1675_),
    .B(net397),
    .C(net535),
    .D(_1988_),
    .Y(_1992_));
 sky130_fd_sc_hd__and3_1 _4989_ (.A(_1824_),
    .B(net425),
    .C(_1879_),
    .X(_1993_));
 sky130_fd_sc_hd__nand4_1 _4990_ (.A(net397),
    .B(net535),
    .C(net425),
    .D(_1878_),
    .Y(_1994_));
 sky130_fd_sc_hd__nand4_1 _4991_ (.A(net397),
    .B(_1878_),
    .C(net425),
    .D(_1628_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand4_1 _4992_ (.A(net558),
    .B(net397),
    .C(net425),
    .D(_1867_),
    .Y(_1996_));
 sky130_fd_sc_hd__and3_1 _4993_ (.A(net535),
    .B(net425),
    .C(_1868_),
    .X(_1997_));
 sky130_fd_sc_hd__and3_1 _4994_ (.A(_1628_),
    .B(net425),
    .C(_1868_),
    .X(_1998_));
 sky130_fd_sc_hd__nand4_1 _4995_ (.A(_1666_),
    .B(net397),
    .C(_1824_),
    .D(net425),
    .Y(_1999_));
 sky130_fd_sc_hd__nand4_1 _4996_ (.A(_1666_),
    .B(net397),
    .C(net535),
    .D(net425),
    .Y(_2000_));
 sky130_fd_sc_hd__nand4_4 _4997_ (.A(_1628_),
    .B(_1693_),
    .C(_1737_),
    .D(_1771_),
    .Y(_2001_));
 sky130_fd_sc_hd__o211a_2 _4998_ (.A1(net459),
    .A2(_1673_),
    .B1(net558),
    .C1(_1668_),
    .X(_2002_));
 sky130_fd_sc_hd__and3_1 _4999_ (.A(net397),
    .B(_1878_),
    .C(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__and3_1 _5000_ (.A(_1824_),
    .B(_1879_),
    .C(_1880_),
    .X(_2004_));
 sky130_fd_sc_hd__o2111ai_4 _5001_ (.A1(net459),
    .A2(_1673_),
    .B1(_1668_),
    .C1(net535),
    .D1(_1879_),
    .Y(_2005_));
 sky130_fd_sc_hd__o2111ai_2 _5002_ (.A1(net459),
    .A2(_1673_),
    .B1(_1668_),
    .C1(_1879_),
    .D1(_1628_),
    .Y(_2006_));
 sky130_fd_sc_hd__a31o_1 _5003_ (.A1(_1565_),
    .A2(_1569_),
    .A3(_1582_),
    .B1(_1594_),
    .X(_2007_));
 sky130_fd_sc_hd__o2111ai_4 _5004_ (.A1(net112),
    .A2(_0821_),
    .B1(_1565_),
    .C1(_1569_),
    .D1(_1582_),
    .Y(_2008_));
 sky130_fd_sc_hd__nand3_4 _5005_ (.A(_1563_),
    .B(_2007_),
    .C(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__o31ai_1 _5006_ (.A1(_1609_),
    .A2(net530),
    .A3(_2009_),
    .B1(_1694_),
    .Y(_2010_));
 sky130_fd_sc_hd__nand2_2 _5007_ (.A(net552),
    .B(net532),
    .Y(_2011_));
 sky130_fd_sc_hd__o31a_1 _5008_ (.A1(_1712_),
    .A2(net532),
    .A3(net531),
    .B1(net552),
    .X(_2012_));
 sky130_fd_sc_hd__o211a_1 _5009_ (.A1(net459),
    .A2(_1673_),
    .B1(_1666_),
    .C1(_1668_),
    .X(_2013_));
 sky130_fd_sc_hd__o21a_1 _5010_ (.A1(_1666_),
    .A2(_1988_),
    .B1(net424),
    .X(_2014_));
 sky130_fd_sc_hd__nand4_1 _5011_ (.A(_2014_),
    .B(_1823_),
    .C(_1692_),
    .D(net400),
    .Y(_2015_));
 sky130_fd_sc_hd__nand3_2 _5012_ (.A(net400),
    .B(_1692_),
    .C(_2013_),
    .Y(_2016_));
 sky130_fd_sc_hd__and3_2 _5013_ (.A(_1628_),
    .B(net397),
    .C(_2013_),
    .X(_2017_));
 sky130_fd_sc_hd__nand4_2 _5014_ (.A(net400),
    .B(_1692_),
    .C(_1988_),
    .D(_2002_),
    .Y(_2018_));
 sky130_fd_sc_hd__a31o_1 _5015_ (.A1(net558),
    .A2(net424),
    .A3(_1989_),
    .B1(_2017_),
    .X(_2019_));
 sky130_fd_sc_hd__o211ai_1 _5016_ (.A1(_1629_),
    .A2(_2016_),
    .B1(_2018_),
    .C1(_2015_),
    .Y(_2020_));
 sky130_fd_sc_hd__a21oi_1 _5017_ (.A1(_2010_),
    .A2(_2012_),
    .B1(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_1983_),
    .B(_2002_),
    .Y(_2022_));
 sky130_fd_sc_hd__o2111ai_1 _5019_ (.A1(net459),
    .A2(_1673_),
    .B1(_1668_),
    .C1(_1868_),
    .D1(_1628_),
    .Y(_2023_));
 sky130_fd_sc_hd__o2111ai_2 _5020_ (.A1(net459),
    .A2(_1673_),
    .B1(_1668_),
    .C1(net535),
    .D1(_1868_),
    .Y(_2024_));
 sky130_fd_sc_hd__nand4_1 _5021_ (.A(_2021_),
    .B(_2022_),
    .C(_2023_),
    .D(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__and3_1 _5022_ (.A(_1824_),
    .B(_1868_),
    .C(_1880_),
    .X(_2026_));
 sky130_fd_sc_hd__nor2_1 _5023_ (.A(_2026_),
    .B(_2025_),
    .Y(_2027_));
 sky130_fd_sc_hd__o2111ai_4 _5024_ (.A1(net459),
    .A2(_1673_),
    .B1(_1668_),
    .C1(_1868_),
    .D1(net558),
    .Y(_2028_));
 sky130_fd_sc_hd__nand4_2 _5025_ (.A(_2027_),
    .B(_2028_),
    .C(_2005_),
    .D(_2006_),
    .Y(_2029_));
 sky130_fd_sc_hd__nor3_1 _5026_ (.A(_2003_),
    .B(_2004_),
    .C(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand4_1 _5027_ (.A(net397),
    .B(net535),
    .C(net425),
    .D(_1988_),
    .Y(_2031_));
 sky130_fd_sc_hd__nand3_1 _5028_ (.A(_2030_),
    .B(_2031_),
    .C(_2001_),
    .Y(_2032_));
 sky130_fd_sc_hd__and3_1 _5029_ (.A(_1824_),
    .B(net425),
    .C(_1989_),
    .X(_2033_));
 sky130_fd_sc_hd__and3_1 _5030_ (.A(net558),
    .B(net425),
    .C(_1989_),
    .X(_2034_));
 sky130_fd_sc_hd__nor3_1 _5031_ (.A(_2033_),
    .B(_2034_),
    .C(_2032_),
    .Y(_2035_));
 sky130_fd_sc_hd__a2111o_1 _5032_ (.A1(net611),
    .A2(_1665_),
    .B1(_1664_),
    .C1(_1866_),
    .D1(_1763_),
    .X(_2036_));
 sky130_fd_sc_hd__nand4_1 _5033_ (.A(_2035_),
    .B(_2036_),
    .C(_1999_),
    .D(_2000_),
    .Y(_2037_));
 sky130_fd_sc_hd__and3_1 _5034_ (.A(net558),
    .B(net425),
    .C(_1983_),
    .X(_2038_));
 sky130_fd_sc_hd__nor4_1 _5035_ (.A(_1997_),
    .B(_1998_),
    .C(_2038_),
    .D(_2037_),
    .Y(_2039_));
 sky130_fd_sc_hd__o311a_1 _5036_ (.A1(_1825_),
    .A2(_1866_),
    .A3(_1869_),
    .B1(_1996_),
    .C1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__nand3_1 _5037_ (.A(_2040_),
    .B(_1995_),
    .C(_1994_),
    .Y(_2041_));
 sky130_fd_sc_hd__and3_1 _5038_ (.A(net558),
    .B(net425),
    .C(_1879_),
    .X(_2042_));
 sky130_fd_sc_hd__nor3_1 _5039_ (.A(_1993_),
    .B(_2042_),
    .C(_2041_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand4_1 _5040_ (.A(_1628_),
    .B(_1675_),
    .C(net397),
    .D(_1988_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand4_1 _5041_ (.A(_2043_),
    .B(_2044_),
    .C(_1991_),
    .D(_1992_),
    .Y(_2045_));
 sky130_fd_sc_hd__nor2_1 _5042_ (.A(_1987_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__a2111o_1 _5043_ (.A1(net611),
    .A2(_1665_),
    .B1(_1676_),
    .C1(_1664_),
    .D1(_1763_),
    .X(_2047_));
 sky130_fd_sc_hd__nand3_1 _5044_ (.A(_2046_),
    .B(_2047_),
    .C(_1986_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand3_1 _5045_ (.A(_1675_),
    .B(net448),
    .C(_1878_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_1 _5046_ (.A(_2009_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__nor3_1 _5047_ (.A(_1985_),
    .B(_2050_),
    .C(_2048_),
    .Y(_2051_));
 sky130_fd_sc_hd__nand4_1 _5048_ (.A(_1675_),
    .B(net398),
    .C(_1878_),
    .D(net531),
    .Y(_2052_));
 sky130_fd_sc_hd__nand4_1 _5049_ (.A(_1675_),
    .B(_1682_),
    .C(net531),
    .D(_1988_),
    .Y(_2053_));
 sky130_fd_sc_hd__and3_1 _5050_ (.A(_1712_),
    .B(_1817_),
    .C(net450),
    .X(_2054_));
 sky130_fd_sc_hd__nand3_1 _5051_ (.A(_2051_),
    .B(_2052_),
    .C(_2053_),
    .Y(_2055_));
 sky130_fd_sc_hd__nor3_1 _5052_ (.A(_1974_),
    .B(_2054_),
    .C(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__and3_4 _5053_ (.A(_1675_),
    .B(_1682_),
    .C(_1867_),
    .X(_2057_));
 sky130_fd_sc_hd__a32oi_2 _5054_ (.A1(_1682_),
    .A2(net536),
    .A3(net531),
    .B1(_2057_),
    .B2(net532),
    .Y(_2058_));
 sky130_fd_sc_hd__nand4_1 _5055_ (.A(_1592_),
    .B(_1712_),
    .C(net537),
    .D(net559),
    .Y(_2059_));
 sky130_fd_sc_hd__nand3_1 _5056_ (.A(_2056_),
    .B(_2058_),
    .C(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5057_ (.A(net534),
    .B(_2057_),
    .Y(_2061_));
 sky130_fd_sc_hd__and4b_1 _5058_ (.A_N(net562),
    .B(net617),
    .C(_2057_),
    .D(net619),
    .X(_2062_));
 sky130_fd_sc_hd__and3_2 _5059_ (.A(net552),
    .B(_1725_),
    .C(net450),
    .X(_2063_));
 sky130_fd_sc_hd__nor3_1 _5060_ (.A(_2063_),
    .B(_2062_),
    .C(_2060_),
    .Y(_2064_));
 sky130_fd_sc_hd__and3_1 _5061_ (.A(net552),
    .B(net454),
    .C(net450),
    .X(_2065_));
 sky130_fd_sc_hd__o32a_1 _5062_ (.A1(_1609_),
    .A2(_1658_),
    .A3(_1884_),
    .B1(_1850_),
    .B2(_1748_),
    .X(_2066_));
 sky130_fd_sc_hd__nand4_1 _5063_ (.A(_1682_),
    .B(_1878_),
    .C(net448),
    .D(_1675_),
    .Y(_2067_));
 sky130_fd_sc_hd__nand3_1 _5064_ (.A(_2064_),
    .B(_2066_),
    .C(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__nand2_2 _5065_ (.A(net360),
    .B(_1847_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2_2 _5066_ (.A(_1792_),
    .B(_1847_),
    .Y(_2070_));
 sky130_fd_sc_hd__and3_1 _5067_ (.A(_1701_),
    .B(net542),
    .C(_1847_),
    .X(_2071_));
 sky130_fd_sc_hd__nand3_1 _5068_ (.A(_1701_),
    .B(net545),
    .C(_1847_),
    .Y(_2072_));
 sky130_fd_sc_hd__and3_4 _5069_ (.A(net556),
    .B(_1705_),
    .C(net542),
    .X(_2073_));
 sky130_fd_sc_hd__a22o_1 _5070_ (.A1(net546),
    .A2(_1835_),
    .B1(_1891_),
    .B2(net555),
    .X(_2074_));
 sky130_fd_sc_hd__nor4b_4 _5071_ (.A(net111),
    .B(net114),
    .C(net113),
    .D_N(net112),
    .Y(_2075_));
 sky130_fd_sc_hd__nand4_1 _5072_ (.A(net551),
    .B(_1705_),
    .C(_1835_),
    .D(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_8 _5073_ (.A(_1603_),
    .B(_1746_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand4_1 _5074_ (.A(_2077_),
    .B(_1740_),
    .C(net543),
    .D(net556),
    .Y(_2078_));
 sky130_fd_sc_hd__o311ai_1 _5075_ (.A1(_1609_),
    .A2(net458),
    .A3(_1713_),
    .B1(_2076_),
    .C1(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__a21oi_1 _5076_ (.A1(net542),
    .A2(_2074_),
    .B1(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_4 _5077_ (.A(net543),
    .B(_1744_),
    .Y(_2081_));
 sky130_fd_sc_hd__o32a_1 _5078_ (.A1(_1575_),
    .A2(_1601_),
    .A3(_1731_),
    .B1(_1950_),
    .B2(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__and3_1 _5079_ (.A(_1570_),
    .B(_1718_),
    .C(_1949_),
    .X(_2083_));
 sky130_fd_sc_hd__o32a_1 _5080_ (.A1(net457),
    .A2(_1741_),
    .A3(_1950_),
    .B1(_2081_),
    .B2(_1752_),
    .X(_2084_));
 sky130_fd_sc_hd__nand4_2 _5081_ (.A(_2077_),
    .B(_1723_),
    .C(net542),
    .D(net556),
    .Y(_2085_));
 sky130_fd_sc_hd__o221a_1 _5082_ (.A1(_1721_),
    .A2(_1752_),
    .B1(_1950_),
    .B2(_1731_),
    .C1(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__o32a_1 _5083_ (.A1(net458),
    .A2(_1724_),
    .A3(_1950_),
    .B1(_1752_),
    .B2(_1721_),
    .X(_2087_));
 sky130_fd_sc_hd__nand4_1 _5084_ (.A(_2080_),
    .B(_2082_),
    .C(_2084_),
    .D(_2086_),
    .Y(_2088_));
 sky130_fd_sc_hd__a31oi_1 _5085_ (.A1(_1604_),
    .A2(net543),
    .A3(net539),
    .B1(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_1751_),
    .B(_1777_),
    .Y(_2090_));
 sky130_fd_sc_hd__o211ai_1 _5087_ (.A1(_1721_),
    .A2(_1846_),
    .B1(_2090_),
    .C1(_2089_),
    .Y(_2091_));
 sky130_fd_sc_hd__a21oi_1 _5088_ (.A1(_1604_),
    .A2(_1777_),
    .B1(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand4_4 _5089_ (.A(_1701_),
    .B(_0821_),
    .C(_1564_),
    .D(_1751_),
    .Y(_2093_));
 sky130_fd_sc_hd__o211ai_1 _5090_ (.A1(_1778_),
    .A2(_1846_),
    .B1(_2093_),
    .C1(_2092_),
    .Y(_2094_));
 sky130_fd_sc_hd__and3_1 _5091_ (.A(net556),
    .B(_1602_),
    .C(_1701_),
    .X(_2095_));
 sky130_fd_sc_hd__a211oi_1 _5092_ (.A1(net542),
    .A2(_2095_),
    .B1(_2071_),
    .C1(_2094_),
    .Y(_2096_));
 sky130_fd_sc_hd__o21ai_1 _5093_ (.A1(_1711_),
    .A2(_1950_),
    .B1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_1751_),
    .B(_1792_),
    .Y(_2098_));
 sky130_fd_sc_hd__a31oi_1 _5095_ (.A1(net616),
    .A2(net556),
    .A3(_1792_),
    .B1(_2097_),
    .Y(_2099_));
 sky130_fd_sc_hd__nand2_1 _5096_ (.A(_1792_),
    .B(_1949_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand3_1 _5097_ (.A(_2099_),
    .B(_2100_),
    .C(_2070_),
    .Y(_2101_));
 sky130_fd_sc_hd__a31oi_2 _5098_ (.A1(net616),
    .A2(net556),
    .A3(_1801_),
    .B1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__o21ai_1 _5099_ (.A1(_1802_),
    .A2(_1846_),
    .B1(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__and3_1 _5100_ (.A(_1570_),
    .B(_1607_),
    .C(net543),
    .X(_2104_));
 sky130_fd_sc_hd__a31oi_2 _5101_ (.A1(net615),
    .A2(net556),
    .A3(_2104_),
    .B1(_2103_),
    .Y(_2105_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_1809_),
    .B(_2073_),
    .Y(_2106_));
 sky130_fd_sc_hd__o311ai_2 _5103_ (.A1(net457),
    .A2(_1810_),
    .A3(_1848_),
    .B1(_2106_),
    .C1(_2105_),
    .Y(_2107_));
 sky130_fd_sc_hd__a31oi_1 _5104_ (.A1(net615),
    .A2(net556),
    .A3(_1821_),
    .B1(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__and3_1 _5105_ (.A(net543),
    .B(_1817_),
    .C(_1847_),
    .X(_2109_));
 sky130_fd_sc_hd__o31ai_1 _5106_ (.A1(net457),
    .A2(_1818_),
    .A3(_1848_),
    .B1(_2108_),
    .Y(_2110_));
 sky130_fd_sc_hd__and3_1 _5107_ (.A(net552),
    .B(net548),
    .C(net543),
    .X(_2111_));
 sky130_fd_sc_hd__a31o_1 _5108_ (.A1(net552),
    .A2(_1747_),
    .A3(net529),
    .B1(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__and3_1 _5109_ (.A(net548),
    .B(_1809_),
    .C(net452),
    .X(_2113_));
 sky130_fd_sc_hd__and3_1 _5110_ (.A(_1703_),
    .B(_1809_),
    .C(net452),
    .X(_2114_));
 sky130_fd_sc_hd__nor3_1 _5111_ (.A(_2113_),
    .B(_2112_),
    .C(_2110_),
    .Y(_2115_));
 sky130_fd_sc_hd__o221a_1 _5112_ (.A1(_1832_),
    .A2(net530),
    .B1(_1977_),
    .B2(net562),
    .C1(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__and3_1 _5113_ (.A(_1712_),
    .B(net452),
    .C(net538),
    .X(_2117_));
 sky130_fd_sc_hd__a31o_1 _5114_ (.A1(net548),
    .A2(_1817_),
    .A3(net452),
    .B1(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__and3_2 _5115_ (.A(_1426_),
    .B(_1593_),
    .C(net538),
    .X(_2119_));
 sky130_fd_sc_hd__o32a_1 _5116_ (.A1(_1713_),
    .A2(_1830_),
    .A3(_1836_),
    .B1(_1832_),
    .B2(_1707_),
    .X(_2120_));
 sky130_fd_sc_hd__o311ai_4 _5117_ (.A1(_1830_),
    .A2(_1836_),
    .A3(net530),
    .B1(_2120_),
    .C1(_2116_),
    .Y(_2121_));
 sky130_fd_sc_hd__and3_1 _5118_ (.A(net548),
    .B(net451),
    .C(net537),
    .X(_2122_));
 sky130_fd_sc_hd__a211o_1 _5119_ (.A1(_1725_),
    .A2(_2119_),
    .B1(_2122_),
    .C1(_2121_),
    .X(_2123_));
 sky130_fd_sc_hd__a21oi_1 _5120_ (.A1(_1849_),
    .A2(net532),
    .B1(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__a211o_1 _5121_ (.A1(_1726_),
    .A2(_1884_),
    .B1(_1830_),
    .C1(_1609_),
    .X(_2125_));
 sky130_fd_sc_hd__nand3b_1 _5122_ (.A_N(_2065_),
    .B(_2124_),
    .C(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__o31a_1 _5123_ (.A1(_1609_),
    .A2(_1707_),
    .A3(_1830_),
    .B1(net463),
    .X(_2127_));
 sky130_fd_sc_hd__a21o_1 _5124_ (.A1(_2126_),
    .A2(_2127_),
    .B1(net461),
    .X(_2128_));
 sky130_fd_sc_hd__a221oi_2 _5125_ (.A1(_1855_),
    .A2(_1856_),
    .B1(_2068_),
    .B2(_1972_),
    .C1(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__a22oi_1 _5126_ (.A1(net463),
    .A2(_1561_),
    .B1(_2129_),
    .B2(_1971_),
    .Y(_0372_));
 sky130_fd_sc_hd__and3_1 _5127_ (.A(net363),
    .B(net402),
    .C(_1824_),
    .X(_2130_));
 sky130_fd_sc_hd__o211a_1 _5128_ (.A1(_1699_),
    .A2(_1736_),
    .B1(_1826_),
    .C1(_1700_),
    .X(_2131_));
 sky130_fd_sc_hd__a31o_1 _5129_ (.A1(_1690_),
    .A2(net456),
    .A3(_1817_),
    .B1(_1985_),
    .X(_2132_));
 sky130_fd_sc_hd__o22a_1 _5130_ (.A1(_1707_),
    .A2(_1711_),
    .B1(_1787_),
    .B2(_1629_),
    .X(_2133_));
 sky130_fd_sc_hd__o31a_1 _5131_ (.A1(_1707_),
    .A2(net458),
    .A3(_1720_),
    .B1(_2001_),
    .X(_2134_));
 sky130_fd_sc_hd__o22a_1 _5132_ (.A1(_1726_),
    .A2(_1731_),
    .B1(_1765_),
    .B2(_1982_),
    .X(_2135_));
 sky130_fd_sc_hd__a31o_1 _5133_ (.A1(net615),
    .A2(net618),
    .A3(net556),
    .B1(_1891_),
    .X(_2136_));
 sky130_fd_sc_hd__and3_1 _5134_ (.A(net555),
    .B(net542),
    .C(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__a22oi_2 _5135_ (.A1(net455),
    .A2(_1744_),
    .B1(_1757_),
    .B2(_1824_),
    .Y(_2138_));
 sky130_fd_sc_hd__o21ba_1 _5136_ (.A1(_1691_),
    .A2(_2138_),
    .B1_N(_2137_),
    .X(_2139_));
 sky130_fd_sc_hd__a211o_1 _5137_ (.A1(_1699_),
    .A2(_1739_),
    .B1(_1825_),
    .C1(_1691_),
    .X(_2140_));
 sky130_fd_sc_hd__nand4_1 _5138_ (.A(_1687_),
    .B(_1688_),
    .C(_1698_),
    .D(_1824_),
    .Y(_2141_));
 sky130_fd_sc_hd__and4b_1 _5139_ (.A_N(_2017_),
    .B(_2139_),
    .C(_2140_),
    .D(_1743_),
    .X(_2142_));
 sky130_fd_sc_hd__o32a_1 _5140_ (.A1(_1629_),
    .A2(_1691_),
    .A3(_1765_),
    .B1(_1745_),
    .B2(_1710_),
    .X(_2143_));
 sky130_fd_sc_hd__o221a_1 _5141_ (.A1(_1710_),
    .A2(_1745_),
    .B1(_1763_),
    .B2(_1765_),
    .C1(_2142_),
    .X(_2144_));
 sky130_fd_sc_hd__o32a_1 _5142_ (.A1(_1629_),
    .A2(_1694_),
    .A3(_1717_),
    .B1(_1724_),
    .B2(_1710_),
    .X(_2145_));
 sky130_fd_sc_hd__and3_1 _5143_ (.A(_2135_),
    .B(_2144_),
    .C(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__o32a_1 _5144_ (.A1(_1691_),
    .A2(_1717_),
    .A3(_1825_),
    .B1(_1727_),
    .B2(_1720_),
    .X(_2147_));
 sky130_fd_sc_hd__nand3_1 _5145_ (.A(_2134_),
    .B(_2146_),
    .C(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__a31o_1 _5146_ (.A1(_1737_),
    .A2(_1771_),
    .A3(_1981_),
    .B1(_1779_),
    .X(_2149_));
 sky130_fd_sc_hd__a32o_1 _5147_ (.A1(_1644_),
    .A2(_1762_),
    .A3(_1771_),
    .B1(_1777_),
    .B2(net546),
    .X(_2150_));
 sky130_fd_sc_hd__nor3_1 _5148_ (.A(_2148_),
    .B(_2149_),
    .C(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__o32a_1 _5149_ (.A1(_1691_),
    .A2(_1781_),
    .A3(_1825_),
    .B1(_1702_),
    .B2(_1727_),
    .X(_2152_));
 sky130_fd_sc_hd__and3_1 _5150_ (.A(_2133_),
    .B(_2151_),
    .C(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__o32a_1 _5151_ (.A1(net457),
    .A2(_1726_),
    .A3(_1791_),
    .B1(_1825_),
    .B2(_1787_),
    .X(_2154_));
 sky130_fd_sc_hd__a32oi_4 _5152_ (.A1(_1697_),
    .A2(_1762_),
    .A3(_1771_),
    .B1(_1792_),
    .B2(net547),
    .Y(_2155_));
 sky130_fd_sc_hd__and3_1 _5153_ (.A(_2153_),
    .B(_2154_),
    .C(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__o32a_1 _5154_ (.A1(_1691_),
    .A2(_1797_),
    .A3(_1825_),
    .B1(_1800_),
    .B2(_1727_),
    .X(_2157_));
 sky130_fd_sc_hd__o32a_1 _5155_ (.A1(_1629_),
    .A2(_1694_),
    .A3(_1806_),
    .B1(_1800_),
    .B2(_1710_),
    .X(_2158_));
 sky130_fd_sc_hd__nand3_1 _5156_ (.A(_2156_),
    .B(_2157_),
    .C(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__a32o_1 _5157_ (.A1(net543),
    .A2(net456),
    .A3(_1809_),
    .B1(_1981_),
    .B2(_1805_),
    .X(_2160_));
 sky130_fd_sc_hd__and3_1 _5158_ (.A(_1628_),
    .B(net402),
    .C(_1690_),
    .X(_2161_));
 sky130_fd_sc_hd__a31o_1 _5159_ (.A1(_1690_),
    .A2(net549),
    .A3(_1809_),
    .B1(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__nor4_1 _5160_ (.A(_2132_),
    .B(_2159_),
    .C(_2160_),
    .D(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__a211o_1 _5161_ (.A1(_1752_),
    .A2(net530),
    .B1(_1830_),
    .C1(_1818_),
    .X(_2164_));
 sky130_fd_sc_hd__a211o_1 _5162_ (.A1(_1752_),
    .A2(net530),
    .B1(_1830_),
    .C1(_1818_),
    .X(_2165_));
 sky130_fd_sc_hd__nand3_1 _5163_ (.A(_2131_),
    .B(_2163_),
    .C(_2164_),
    .Y(_2166_));
 sky130_fd_sc_hd__nor2_1 _5164_ (.A(_2130_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__o32a_2 _5165_ (.A1(_1599_),
    .A2(_1752_),
    .A3(_1836_),
    .B1(_1838_),
    .B2(_1713_),
    .X(_2168_));
 sky130_fd_sc_hd__a31oi_4 _5166_ (.A1(net362),
    .A2(net395),
    .A3(net535),
    .B1(_2063_),
    .Y(_2169_));
 sky130_fd_sc_hd__nand4_1 _5167_ (.A(_2167_),
    .B(_2168_),
    .C(_2169_),
    .D(_1843_),
    .Y(_2170_));
 sky130_fd_sc_hd__o31a_1 _5168_ (.A1(_1853_),
    .A2(_2065_),
    .A3(_2170_),
    .B1(_1856_),
    .X(_2171_));
 sky130_fd_sc_hd__o32a_1 _5169_ (.A1(_1676_),
    .A2(_1876_),
    .A3(_1984_),
    .B1(_1696_),
    .B2(_1818_),
    .X(_2172_));
 sky130_fd_sc_hd__a31o_1 _5170_ (.A1(_1675_),
    .A2(net532),
    .A3(_1989_),
    .B1(_2042_),
    .X(_2173_));
 sky130_fd_sc_hd__a32o_1 _5171_ (.A1(net558),
    .A2(_1865_),
    .A3(_1868_),
    .B1(_1879_),
    .B2(_1914_),
    .X(_2174_));
 sky130_fd_sc_hd__a22o_1 _5172_ (.A1(_1874_),
    .A2(net532),
    .B1(_2002_),
    .B2(_1868_),
    .X(_2175_));
 sky130_fd_sc_hd__o32a_1 _5173_ (.A1(_1609_),
    .A2(net530),
    .A3(_2009_),
    .B1(_2049_),
    .B2(_1694_),
    .X(_2176_));
 sky130_fd_sc_hd__a21oi_4 _5174_ (.A1(net617),
    .A2(_1823_),
    .B1(net448),
    .Y(_2177_));
 sky130_fd_sc_hd__a21o_1 _5175_ (.A1(_1876_),
    .A2(_2177_),
    .B1(_2016_),
    .X(_2178_));
 sky130_fd_sc_hd__o311a_1 _5176_ (.A1(_1609_),
    .A2(_1694_),
    .A3(_1975_),
    .B1(_2018_),
    .C1(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__o21ai_1 _5177_ (.A1(net535),
    .A2(net448),
    .B1(net424),
    .Y(_2180_));
 sky130_fd_sc_hd__o21a_1 _5178_ (.A1(net535),
    .A2(net448),
    .B1(_1880_),
    .X(_2181_));
 sky130_fd_sc_hd__o211ai_2 _5179_ (.A1(_2180_),
    .A2(_1990_),
    .B1(_2176_),
    .C1(_2179_),
    .Y(_2182_));
 sky130_fd_sc_hd__and3_1 _5180_ (.A(_1868_),
    .B(net532),
    .C(_1880_),
    .X(_2183_));
 sky130_fd_sc_hd__o211a_1 _5181_ (.A1(net535),
    .A2(net448),
    .B1(_1868_),
    .C1(_1880_),
    .X(_2184_));
 sky130_fd_sc_hd__a2111oi_1 _5182_ (.A1(_1983_),
    .A2(_2002_),
    .B1(_2183_),
    .C1(_2184_),
    .D1(_2182_),
    .Y(_2185_));
 sky130_fd_sc_hd__nand4_1 _5183_ (.A(net397),
    .B(_1878_),
    .C(net448),
    .D(_1675_),
    .Y(_2186_));
 sky130_fd_sc_hd__o31a_1 _5184_ (.A1(_1609_),
    .A2(net530),
    .A3(_2009_),
    .B1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__nand3_1 _5185_ (.A(_2185_),
    .B(_2028_),
    .C(_1881_),
    .Y(_2188_));
 sky130_fd_sc_hd__a31o_1 _5186_ (.A1(net425),
    .A2(net532),
    .A3(_1989_),
    .B1(_2003_),
    .X(_2189_));
 sky130_fd_sc_hd__a211o_1 _5187_ (.A1(_2181_),
    .A2(_1879_),
    .B1(_2189_),
    .C1(_2188_),
    .X(_2190_));
 sky130_fd_sc_hd__o21a_1 _5188_ (.A1(net535),
    .A2(net448),
    .B1(_1865_),
    .X(_2191_));
 sky130_fd_sc_hd__a31o_1 _5189_ (.A1(net394),
    .A2(net532),
    .A3(_1983_),
    .B1(_2034_),
    .X(_2192_));
 sky130_fd_sc_hd__a211o_1 _5190_ (.A1(_1989_),
    .A2(_2191_),
    .B1(_2192_),
    .C1(_2190_),
    .X(_2193_));
 sky130_fd_sc_hd__a31o_1 _5191_ (.A1(net394),
    .A2(_1868_),
    .A3(net532),
    .B1(_2038_),
    .X(_2194_));
 sky130_fd_sc_hd__a211o_1 _5192_ (.A1(_1983_),
    .A2(_2191_),
    .B1(_2193_),
    .C1(_2194_),
    .X(_2195_));
 sky130_fd_sc_hd__a311o_1 _5193_ (.A1(net397),
    .A2(_1867_),
    .A3(_2191_),
    .B1(_2195_),
    .C1(_2174_),
    .X(_2196_));
 sky130_fd_sc_hd__a311oi_2 _5194_ (.A1(net397),
    .A2(_2191_),
    .A3(_1878_),
    .B1(_2173_),
    .C1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__o311a_1 _5195_ (.A1(_1676_),
    .A2(_2177_),
    .A3(_1990_),
    .B1(_2172_),
    .C1(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__o311a_1 _5196_ (.A1(_1676_),
    .A2(_1862_),
    .A3(_1984_),
    .B1(_1986_),
    .C1(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__a2111o_1 _5197_ (.A1(_1862_),
    .A2(net530),
    .B1(_1877_),
    .C1(_1676_),
    .D1(_2009_),
    .X(_2200_));
 sky130_fd_sc_hd__o311a_1 _5198_ (.A1(_1676_),
    .A2(_1897_),
    .A3(_1877_),
    .B1(_2200_),
    .C1(_2199_),
    .X(_2201_));
 sky130_fd_sc_hd__nand4b_2 _5199_ (.A_N(net617),
    .B(_1682_),
    .C(net534),
    .D(_1978_),
    .Y(_2202_));
 sky130_fd_sc_hd__and3_1 _5200_ (.A(_2201_),
    .B(_2202_),
    .C(_1977_),
    .X(_2203_));
 sky130_fd_sc_hd__a32oi_2 _5201_ (.A1(_1682_),
    .A2(_1712_),
    .A3(net536),
    .B1(_2057_),
    .B2(_1628_),
    .Y(_2204_));
 sky130_fd_sc_hd__and3_1 _5202_ (.A(_2203_),
    .B(_2204_),
    .C(_2061_),
    .X(_2205_));
 sky130_fd_sc_hd__nand4_1 _5203_ (.A(_1682_),
    .B(_1878_),
    .C(net535),
    .D(_1675_),
    .Y(_2206_));
 sky130_fd_sc_hd__o31a_1 _5204_ (.A1(_1609_),
    .A2(_1683_),
    .A3(_1884_),
    .B1(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__a31o_1 _5205_ (.A1(net362),
    .A2(net552),
    .A3(net454),
    .B1(_1973_),
    .X(_2208_));
 sky130_fd_sc_hd__a21oi_1 _5206_ (.A1(_2205_),
    .A2(_2207_),
    .B1(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__a21o_1 _5207_ (.A1(_1629_),
    .A2(_1713_),
    .B1(_1663_),
    .X(_2210_));
 sky130_fd_sc_hd__o31ai_1 _5208_ (.A1(net458),
    .A2(_1800_),
    .A3(_1950_),
    .B1(_1933_),
    .Y(_2211_));
 sky130_fd_sc_hd__o2bb2a_1 _5209_ (.A1_N(_1885_),
    .A2_N(_1913_),
    .B1(_1950_),
    .B2(_1778_),
    .X(_2212_));
 sky130_fd_sc_hd__o31a_1 _5210_ (.A1(_1605_),
    .A2(_1720_),
    .A3(_1730_),
    .B1(_1909_),
    .X(_2213_));
 sky130_fd_sc_hd__o21ai_1 _5211_ (.A1(_1720_),
    .A2(_1890_),
    .B1(_1909_),
    .Y(_2214_));
 sky130_fd_sc_hd__a31o_1 _5212_ (.A1(net545),
    .A2(_1723_),
    .A3(_1949_),
    .B1(_1887_),
    .X(_2215_));
 sky130_fd_sc_hd__and4_1 _5213_ (.A(_1659_),
    .B(net360),
    .C(_1872_),
    .D(_1883_),
    .X(_2216_));
 sky130_fd_sc_hd__o31a_1 _5214_ (.A1(_1626_),
    .A2(_1730_),
    .A3(_1950_),
    .B1(_1902_),
    .X(_2217_));
 sky130_fd_sc_hd__o31a_1 _5215_ (.A1(_1626_),
    .A2(_1713_),
    .A3(_1730_),
    .B1(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__and3_2 _5216_ (.A(_1880_),
    .B(_1883_),
    .C(_1988_),
    .X(_2219_));
 sky130_fd_sc_hd__a31o_1 _5217_ (.A1(_1872_),
    .A2(_1883_),
    .A3(_1896_),
    .B1(_2083_),
    .X(_2220_));
 sky130_fd_sc_hd__o21ai_1 _5218_ (.A1(_2083_),
    .A2(_2219_),
    .B1(net360),
    .Y(_2221_));
 sky130_fd_sc_hd__o2111ai_2 _5219_ (.A1(_1745_),
    .A2(_1890_),
    .B1(_1900_),
    .C1(_1907_),
    .D1(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__a32o_1 _5220_ (.A1(_1659_),
    .A2(_1872_),
    .A3(_1883_),
    .B1(_1949_),
    .B2(_1744_),
    .X(_2223_));
 sky130_fd_sc_hd__a21oi_1 _5221_ (.A1(net360),
    .A2(_2223_),
    .B1(_2222_),
    .Y(_2224_));
 sky130_fd_sc_hd__nand4_1 _5222_ (.A(_1604_),
    .B(net401),
    .C(_1656_),
    .D(_1723_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand4_1 _5223_ (.A(_2218_),
    .B(_2224_),
    .C(_2225_),
    .D(_1894_),
    .Y(_2226_));
 sky130_fd_sc_hd__nor3_1 _5224_ (.A(_2214_),
    .B(_2215_),
    .C(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a32oi_2 _5225_ (.A1(_1871_),
    .A2(_1872_),
    .A3(_1883_),
    .B1(_2073_),
    .B2(net541),
    .Y(_2228_));
 sky130_fd_sc_hd__a32o_1 _5226_ (.A1(_1871_),
    .A2(_1872_),
    .A3(_1883_),
    .B1(_2073_),
    .B2(net541),
    .X(_2229_));
 sky130_fd_sc_hd__a21oi_2 _5227_ (.A1(_1776_),
    .A2(_1889_),
    .B1(_1911_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand4_1 _5228_ (.A(_2212_),
    .B(_2227_),
    .C(_2228_),
    .D(_2230_),
    .Y(_2231_));
 sky130_fd_sc_hd__a31o_1 _5229_ (.A1(_1604_),
    .A2(_1701_),
    .A3(net360),
    .B1(_1919_),
    .X(_2232_));
 sky130_fd_sc_hd__a32o_1 _5230_ (.A1(_1659_),
    .A2(net394),
    .A3(_1885_),
    .B1(_2073_),
    .B2(_1701_),
    .X(_2233_));
 sky130_fd_sc_hd__nor3_1 _5231_ (.A(_2231_),
    .B(_2232_),
    .C(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__a21oi_1 _5232_ (.A1(_1790_),
    .A2(_1889_),
    .B1(_1925_),
    .Y(_2235_));
 sky130_fd_sc_hd__a32o_1 _5233_ (.A1(net426),
    .A2(net394),
    .A3(_1885_),
    .B1(_2073_),
    .B2(_1790_),
    .X(_2236_));
 sky130_fd_sc_hd__a32oi_1 _5234_ (.A1(net394),
    .A2(_1868_),
    .A3(_1883_),
    .B1(_2073_),
    .B2(_1790_),
    .Y(_2237_));
 sky130_fd_sc_hd__and3_1 _5235_ (.A(_2234_),
    .B(_2235_),
    .C(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__a21oi_1 _5236_ (.A1(_1799_),
    .A2(_1889_),
    .B1(_1930_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand3b_1 _5237_ (.A_N(_2211_),
    .B(_2238_),
    .C(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__a31o_1 _5238_ (.A1(_1604_),
    .A2(net361),
    .A3(_1809_),
    .B1(_1936_),
    .X(_2241_));
 sky130_fd_sc_hd__a311o_1 _5239_ (.A1(_1604_),
    .A2(net361),
    .A3(_1809_),
    .B1(_1937_),
    .C1(_2240_),
    .X(_2242_));
 sky130_fd_sc_hd__a22o_1 _5240_ (.A1(net556),
    .A2(_1705_),
    .B1(net533),
    .B2(net618),
    .X(_2243_));
 sky130_fd_sc_hd__a21o_1 _5241_ (.A1(_1939_),
    .A2(_2243_),
    .B1(_2242_),
    .X(_2244_));
 sky130_fd_sc_hd__a31o_1 _5242_ (.A1(_1604_),
    .A2(_1661_),
    .A3(net361),
    .B1(_1944_),
    .X(_2245_));
 sky130_fd_sc_hd__and3_1 _5243_ (.A(_1661_),
    .B(net361),
    .C(_2243_),
    .X(_2246_));
 sky130_fd_sc_hd__nor3_1 _5244_ (.A(_2246_),
    .B(_2245_),
    .C(_2244_),
    .Y(_2247_));
 sky130_fd_sc_hd__o22a_1 _5245_ (.A1(_1575_),
    .A2(_1601_),
    .B1(net618),
    .B2(_1846_),
    .X(_2248_));
 sky130_fd_sc_hd__o32a_1 _5246_ (.A1(_1626_),
    .A2(_1730_),
    .A3(_1752_),
    .B1(_1951_),
    .B2(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__and3_1 _5247_ (.A(_2210_),
    .B(_2247_),
    .C(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__and3_1 _5248_ (.A(_1657_),
    .B(_1661_),
    .C(_1949_),
    .X(_2251_));
 sky130_fd_sc_hd__o21ai_1 _5249_ (.A1(_1663_),
    .A2(_1950_),
    .B1(_2250_),
    .Y(_2252_));
 sky130_fd_sc_hd__a31o_1 _5250_ (.A1(net620),
    .A2(_1602_),
    .A3(_1957_),
    .B1(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__a31o_1 _5251_ (.A1(_1625_),
    .A2(_1682_),
    .A3(_1883_),
    .B1(_1851_),
    .X(_2254_));
 sky130_fd_sc_hd__nor3_1 _5252_ (.A(_2254_),
    .B(_1964_),
    .C(_2253_),
    .Y(_2255_));
 sky130_fd_sc_hd__a31oi_1 _5253_ (.A1(net552),
    .A2(_1703_),
    .A3(net529),
    .B1(_2111_),
    .Y(_2256_));
 sky130_fd_sc_hd__o22a_1 _5254_ (.A1(_1711_),
    .A2(_1713_),
    .B1(_1778_),
    .B2(_1950_),
    .X(_2257_));
 sky130_fd_sc_hd__o31a_4 _5255_ (.A1(net620),
    .A2(net562),
    .A3(_1746_),
    .B1(_1605_),
    .X(_2258_));
 sky130_fd_sc_hd__a211o_1 _5256_ (.A1(_1605_),
    .A2(_1748_),
    .B1(_1720_),
    .C1(net458),
    .X(_2259_));
 sky130_fd_sc_hd__a2bb2o_1 _5257_ (.A1_N(_2258_),
    .A2_N(_2081_),
    .B1(net539),
    .B2(_1714_),
    .X(_2260_));
 sky130_fd_sc_hd__a31o_1 _5258_ (.A1(net542),
    .A2(_1723_),
    .A3(net453),
    .B1(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__o31a_1 _5259_ (.A1(_1609_),
    .A2(net458),
    .A3(_1748_),
    .B1(_2076_),
    .X(_2262_));
 sky130_fd_sc_hd__nand4_1 _5260_ (.A(_1606_),
    .B(_1607_),
    .C(net542),
    .D(net531),
    .Y(_2263_));
 sky130_fd_sc_hd__o221a_1 _5261_ (.A1(_1713_),
    .A2(_1731_),
    .B1(_1950_),
    .B2(_2081_),
    .C1(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__o32a_1 _5262_ (.A1(net458),
    .A2(_1741_),
    .A3(_2258_),
    .B1(_2081_),
    .B2(_1713_),
    .X(_2265_));
 sky130_fd_sc_hd__a31o_1 _5263_ (.A1(_1604_),
    .A2(net542),
    .A3(_1723_),
    .B1(_1760_),
    .X(_2266_));
 sky130_fd_sc_hd__a31oi_2 _5264_ (.A1(net125),
    .A2(_1718_),
    .A3(_2073_),
    .B1(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand4_1 _5265_ (.A(_2262_),
    .B(_2264_),
    .C(_2265_),
    .D(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__nor3b_1 _5266_ (.A(_2261_),
    .B(_2268_),
    .C_N(_2259_),
    .Y(_2269_));
 sky130_fd_sc_hd__o2bb2a_1 _5267_ (.A1_N(_1714_),
    .A2_N(_1776_),
    .B1(_1950_),
    .B2(_1721_),
    .X(_2270_));
 sky130_fd_sc_hd__o211a_1 _5268_ (.A1(_2258_),
    .A2(_1778_),
    .B1(_2270_),
    .C1(_2269_),
    .X(_2271_));
 sky130_fd_sc_hd__o311a_1 _5269_ (.A1(_1702_),
    .A2(_2258_),
    .A3(net457),
    .B1(_2257_),
    .C1(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__o32a_1 _5270_ (.A1(_1702_),
    .A2(net457),
    .A3(_1950_),
    .B1(_1793_),
    .B2(_1713_),
    .X(_2273_));
 sky130_fd_sc_hd__o211a_1 _5271_ (.A1(_2258_),
    .A2(_1793_),
    .B1(_2273_),
    .C1(_2272_),
    .X(_2274_));
 sky130_fd_sc_hd__o221a_1 _5272_ (.A1(_1713_),
    .A2(_1802_),
    .B1(_1950_),
    .B2(_1793_),
    .C1(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__o32a_1 _5273_ (.A1(net457),
    .A2(_1713_),
    .A3(_1810_),
    .B1(_1950_),
    .B2(_1802_),
    .X(_2276_));
 sky130_fd_sc_hd__o211a_1 _5274_ (.A1(_2258_),
    .A2(_1802_),
    .B1(_2276_),
    .C1(_2275_),
    .X(_2277_));
 sky130_fd_sc_hd__o31a_1 _5275_ (.A1(net457),
    .A2(_1810_),
    .A3(_2258_),
    .B1(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__o31a_1 _5276_ (.A1(net457),
    .A2(_1713_),
    .A3(_1818_),
    .B1(_2106_),
    .X(_2279_));
 sky130_fd_sc_hd__o211a_1 _5277_ (.A1(_1604_),
    .A2(_1747_),
    .B1(_1817_),
    .C1(net543),
    .X(_2280_));
 sky130_fd_sc_hd__and4b_1 _5278_ (.A_N(_2280_),
    .B(_2279_),
    .C(_2278_),
    .D(_2256_),
    .X(_2281_));
 sky130_fd_sc_hd__o21ai_1 _5279_ (.A1(_1577_),
    .A2(_1832_),
    .B1(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__a31o_1 _5280_ (.A1(net364),
    .A2(net454),
    .A3(_1817_),
    .B1(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__a31o_1 _5281_ (.A1(net364),
    .A2(net538),
    .A3(_2136_),
    .B1(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__and4_1 _5282_ (.A(net617),
    .B(_1703_),
    .C(net450),
    .D(net538),
    .X(_2285_));
 sky130_fd_sc_hd__a21oi_1 _5283_ (.A1(_1725_),
    .A2(_2119_),
    .B1(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__a31o_1 _5284_ (.A1(net551),
    .A2(_2077_),
    .A3(_2119_),
    .B1(_2284_),
    .X(_2287_));
 sky130_fd_sc_hd__a31o_1 _5285_ (.A1(net554),
    .A2(_1725_),
    .A3(net451),
    .B1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__a31o_1 _5286_ (.A1(_1604_),
    .A2(net552),
    .A3(_1682_),
    .B1(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__o21ai_2 _5287_ (.A1(net454),
    .A2(_1847_),
    .B1(_1849_),
    .Y(_2290_));
 sky130_fd_sc_hd__o31ai_2 _5288_ (.A1(_1851_),
    .A2(_2065_),
    .A3(_2289_),
    .B1(_2127_),
    .Y(_2291_));
 sky130_fd_sc_hd__a211o_1 _5289_ (.A1(_1862_),
    .A2(_1950_),
    .B1(_1626_),
    .C1(_1658_),
    .X(_2292_));
 sky130_fd_sc_hd__a21bo_1 _5290_ (.A1(_2255_),
    .A2(_2292_),
    .B1_N(_1858_),
    .X(_2293_));
 sky130_fd_sc_hd__a2111o_1 _5291_ (.A1(_1825_),
    .A2(_1862_),
    .B1(_1676_),
    .C1(_1877_),
    .D1(_1683_),
    .X(_2294_));
 sky130_fd_sc_hd__o2111ai_2 _5292_ (.A1(_1973_),
    .A2(_2294_),
    .B1(_2291_),
    .C1(_1539_),
    .D1(_2293_),
    .Y(_2295_));
 sky130_fd_sc_hd__o32a_1 _5293_ (.A1(_2171_),
    .A2(_2209_),
    .A3(_2295_),
    .B1(_1539_),
    .B2(net2206),
    .X(_0373_));
 sky130_fd_sc_hd__nand3_1 _5294_ (.A(_1856_),
    .B(_2290_),
    .C(_1854_),
    .Y(_2296_));
 sky130_fd_sc_hd__nand4_2 _5295_ (.A(_1592_),
    .B(net402),
    .C(net535),
    .D(net559),
    .Y(_2297_));
 sky130_fd_sc_hd__o221a_1 _5296_ (.A1(_1724_),
    .A2(_1759_),
    .B1(_1765_),
    .B2(_1696_),
    .C1(_2135_),
    .X(_2298_));
 sky130_fd_sc_hd__nand2_1 _5297_ (.A(_1695_),
    .B(_1757_),
    .Y(_2299_));
 sky130_fd_sc_hd__a211o_1 _5298_ (.A1(_1586_),
    .A2(_1825_),
    .B1(_1739_),
    .C1(_1691_),
    .X(_2300_));
 sky130_fd_sc_hd__o311a_1 _5299_ (.A1(net458),
    .A2(_1726_),
    .A3(_1741_),
    .B1(_1750_),
    .C1(_2300_),
    .X(_2301_));
 sky130_fd_sc_hd__a211o_1 _5300_ (.A1(_1629_),
    .A2(_1713_),
    .B1(_1691_),
    .C1(_1609_),
    .X(_2302_));
 sky130_fd_sc_hd__o311a_1 _5301_ (.A1(net557),
    .A2(_1734_),
    .A3(_1735_),
    .B1(_2141_),
    .C1(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__o221a_1 _5302_ (.A1(_1745_),
    .A2(_1759_),
    .B1(_1691_),
    .B2(_2138_),
    .C1(_2299_),
    .X(_2304_));
 sky130_fd_sc_hd__and4_1 _5303_ (.A(_2298_),
    .B(_2301_),
    .C(_2303_),
    .D(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__o32a_1 _5304_ (.A1(_1571_),
    .A2(_1696_),
    .A3(_1716_),
    .B1(_1720_),
    .B2(_1759_),
    .X(_2306_));
 sky130_fd_sc_hd__o221a_1 _5305_ (.A1(_1720_),
    .A2(_1727_),
    .B1(_1982_),
    .B2(_1717_),
    .C1(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_2305_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__a32o_1 _5307_ (.A1(_1695_),
    .A2(_1737_),
    .A3(_1771_),
    .B1(_1777_),
    .B2(net453),
    .X(_2309_));
 sky130_fd_sc_hd__nor3_1 _5308_ (.A(_2149_),
    .B(_2308_),
    .C(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__o221a_1 _5309_ (.A1(_1702_),
    .A2(_1759_),
    .B1(_1781_),
    .B2(_1696_),
    .C1(_2152_),
    .X(_2311_));
 sky130_fd_sc_hd__o221a_1 _5310_ (.A1(_1586_),
    .A2(_1787_),
    .B1(_1793_),
    .B2(_1748_),
    .C1(_2154_),
    .X(_2312_));
 sky130_fd_sc_hd__and3_1 _5311_ (.A(_2310_),
    .B(_2311_),
    .C(_2312_),
    .X(_2313_));
 sky130_fd_sc_hd__o32a_1 _5312_ (.A1(_1571_),
    .A2(_1696_),
    .A3(_1772_),
    .B1(_1800_),
    .B2(_1759_),
    .X(_2314_));
 sky130_fd_sc_hd__o221a_1 _5313_ (.A1(_1727_),
    .A2(_1800_),
    .B1(_1982_),
    .B2(_1797_),
    .C1(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(_2313_),
    .B(_2315_),
    .Y(_2316_));
 sky130_fd_sc_hd__a311o_1 _5315_ (.A1(net558),
    .A2(_1690_),
    .A3(_1805_),
    .B1(_1812_),
    .C1(_2160_),
    .X(_2317_));
 sky130_fd_sc_hd__o32a_1 _5316_ (.A1(_1609_),
    .A2(_1629_),
    .A3(_1735_),
    .B1(_1759_),
    .B2(_1818_),
    .X(_2318_));
 sky130_fd_sc_hd__nor4b_1 _5317_ (.A(_2132_),
    .B(_2316_),
    .C(_2317_),
    .D_N(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__a211o_1 _5318_ (.A1(_1586_),
    .A2(_1825_),
    .B1(_1806_),
    .C1(_1599_),
    .X(_2320_));
 sky130_fd_sc_hd__and3_1 _5319_ (.A(_2319_),
    .B(_2320_),
    .C(_2165_),
    .X(_2321_));
 sky130_fd_sc_hd__o2111a_1 _5320_ (.A1(_1629_),
    .A2(_1838_),
    .B1(_2168_),
    .C1(_2297_),
    .D1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__o32a_1 _5321_ (.A1(_1599_),
    .A2(_1605_),
    .A3(_1626_),
    .B1(_1850_),
    .B2(_1876_),
    .X(_2323_));
 sky130_fd_sc_hd__a31oi_2 _5322_ (.A1(_2169_),
    .A2(_2322_),
    .A3(_2323_),
    .B1(_2296_),
    .Y(_2324_));
 sky130_fd_sc_hd__o2111a_1 _5323_ (.A1(net448),
    .A2(net531),
    .B1(_1988_),
    .C1(_1682_),
    .D1(_1675_),
    .X(_2325_));
 sky130_fd_sc_hd__nor2_1 _5324_ (.A(_1976_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__o2bb2a_1 _5325_ (.A1_N(net402),
    .A2_N(_1981_),
    .B1(_2009_),
    .B2(_2011_),
    .X(_2327_));
 sky130_fd_sc_hd__o31a_1 _5326_ (.A1(_1676_),
    .A2(_1984_),
    .A3(_2177_),
    .B1(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__a211o_4 _5327_ (.A1(net620),
    .A2(_1705_),
    .B1(net535),
    .C1(net531),
    .X(_2329_));
 sky130_fd_sc_hd__and3_2 _5328_ (.A(net400),
    .B(_1692_),
    .C(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__o311a_2 _5329_ (.A1(_1823_),
    .A2(net448),
    .A3(net531),
    .B1(_1865_),
    .C1(net397),
    .X(_2331_));
 sky130_fd_sc_hd__o221a_1 _5330_ (.A1(_1609_),
    .A2(_1763_),
    .B1(_2011_),
    .B2(_1694_),
    .C1(_2176_),
    .X(_2332_));
 sky130_fd_sc_hd__o221ai_4 _5331_ (.A1(_1609_),
    .A2(_1763_),
    .B1(_2011_),
    .B2(_1694_),
    .C1(_2187_),
    .Y(_2333_));
 sky130_fd_sc_hd__a31o_1 _5332_ (.A1(net398),
    .A2(_2014_),
    .A3(_2329_),
    .B1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__a31o_1 _5333_ (.A1(_1867_),
    .A2(net424),
    .A3(_2330_),
    .B1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__a31o_1 _5334_ (.A1(_1878_),
    .A2(net424),
    .A3(_2330_),
    .B1(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__a31o_1 _5335_ (.A1(net425),
    .A2(_1989_),
    .A3(_2329_),
    .B1(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__a31o_1 _5336_ (.A1(_1666_),
    .A2(net425),
    .A3(_2330_),
    .B1(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__a31o_1 _5337_ (.A1(net425),
    .A2(_1867_),
    .A3(_2330_),
    .B1(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__a21oi_1 _5338_ (.A1(_1878_),
    .A2(_2331_),
    .B1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__nand4_2 _5339_ (.A(net398),
    .B(_2329_),
    .C(_1988_),
    .D(_1675_),
    .Y(_2341_));
 sky130_fd_sc_hd__nand4_1 _5340_ (.A(_2341_),
    .B(_2340_),
    .C(_2328_),
    .D(_2326_),
    .Y(_2342_));
 sky130_fd_sc_hd__a21bo_2 _5341_ (.A1(net532),
    .A2(_2057_),
    .B1_N(_2204_),
    .X(_2343_));
 sky130_fd_sc_hd__and3_2 _5342_ (.A(_1682_),
    .B(_1883_),
    .C(_1978_),
    .X(_2344_));
 sky130_fd_sc_hd__nor3_1 _5343_ (.A(_2344_),
    .B(_2343_),
    .C(_2342_),
    .Y(_2345_));
 sky130_fd_sc_hd__o31a_1 _5344_ (.A1(net620),
    .A2(_1603_),
    .A3(_1850_),
    .B1(_2207_),
    .X(_2346_));
 sky130_fd_sc_hd__a21oi_1 _5345_ (.A1(_2345_),
    .A2(_2346_),
    .B1(_1973_),
    .Y(_2347_));
 sky130_fd_sc_hd__o211a_4 _5346_ (.A1(_1751_),
    .A2(net448),
    .B1(_1654_),
    .C1(_1728_),
    .X(_2348_));
 sky130_fd_sc_hd__a31o_1 _5347_ (.A1(net429),
    .A2(_1864_),
    .A3(_2348_),
    .B1(_2211_),
    .X(_2349_));
 sky130_fd_sc_hd__o2111a_1 _5348_ (.A1(_1751_),
    .A2(net448),
    .B1(_1872_),
    .C1(net426),
    .D1(net360),
    .X(_2350_));
 sky130_fd_sc_hd__nor2_1 _5349_ (.A(_2215_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__o211a_1 _5350_ (.A1(_1751_),
    .A2(net448),
    .B1(_1893_),
    .C1(net361),
    .X(_2352_));
 sky130_fd_sc_hd__a211o_1 _5351_ (.A1(_1605_),
    .A2(_1876_),
    .B1(_1730_),
    .C1(_1626_),
    .X(_2353_));
 sky130_fd_sc_hd__a32oi_4 _5352_ (.A1(_1872_),
    .A2(_1896_),
    .A3(_2348_),
    .B1(_2220_),
    .B2(net360),
    .Y(_2354_));
 sky130_fd_sc_hd__o311a_1 _5353_ (.A1(_1626_),
    .A2(_1730_),
    .A3(_1950_),
    .B1(_1902_),
    .C1(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__a311oi_4 _5354_ (.A1(net360),
    .A2(_1744_),
    .A3(_1949_),
    .B1(_2216_),
    .C1(_2352_),
    .Y(_2356_));
 sky130_fd_sc_hd__and4_1 _5355_ (.A(_2351_),
    .B(_2353_),
    .C(_2355_),
    .D(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__o21ai_1 _5356_ (.A1(_1751_),
    .A2(net448),
    .B1(_1874_),
    .Y(_2358_));
 sky130_fd_sc_hd__a32o_1 _5357_ (.A1(net429),
    .A2(_1872_),
    .A3(_2348_),
    .B1(_2073_),
    .B2(net541),
    .X(_2359_));
 sky130_fd_sc_hd__a31oi_1 _5358_ (.A1(_1872_),
    .A2(_1879_),
    .A3(_1883_),
    .B1(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__a21boi_1 _5359_ (.A1(_1913_),
    .A2(_2348_),
    .B1_N(_2212_),
    .Y(_2361_));
 sky130_fd_sc_hd__a31oi_2 _5360_ (.A1(_1659_),
    .A2(net394),
    .A3(_2348_),
    .B1(_2233_),
    .Y(_2362_));
 sky130_fd_sc_hd__and4_1 _5361_ (.A(_2357_),
    .B(_2360_),
    .C(_2361_),
    .D(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__a31oi_2 _5362_ (.A1(net426),
    .A2(net394),
    .A3(_2348_),
    .B1(_2236_),
    .Y(_2364_));
 sky130_fd_sc_hd__nand3b_1 _5363_ (.A_N(_2349_),
    .B(_2363_),
    .C(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__o31a_1 _5364_ (.A1(_1751_),
    .A2(net533),
    .A3(_1949_),
    .B1(_1939_),
    .X(_2366_));
 sky130_fd_sc_hd__o21bai_2 _5365_ (.A1(_1605_),
    .A2(_1951_),
    .B1_N(_1863_),
    .Y(_2367_));
 sky130_fd_sc_hd__a31o_1 _5366_ (.A1(_1661_),
    .A2(net361),
    .A3(_2243_),
    .B1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__nor4_2 _5367_ (.A(_2366_),
    .B(_2246_),
    .C(_2365_),
    .D(_2367_),
    .Y(_2369_));
 sky130_fd_sc_hd__o31a_2 _5368_ (.A1(_1658_),
    .A2(_1940_),
    .A3(_2248_),
    .B1(_2210_),
    .X(_2370_));
 sky130_fd_sc_hd__a31o_1 _5369_ (.A1(_1605_),
    .A2(_1629_),
    .A3(_1876_),
    .B1(_1958_),
    .X(_2371_));
 sky130_fd_sc_hd__o2111ai_4 _5370_ (.A1(_1663_),
    .A2(_1848_),
    .B1(_2371_),
    .C1(_2370_),
    .D1(_2369_),
    .Y(_2372_));
 sky130_fd_sc_hd__o211a_1 _5371_ (.A1(_1725_),
    .A2(_1844_),
    .B1(_1625_),
    .C1(_1657_),
    .X(_2373_));
 sky130_fd_sc_hd__o31a_1 _5372_ (.A1(_2254_),
    .A2(_2372_),
    .A3(_2373_),
    .B1(_1858_),
    .X(_2374_));
 sky130_fd_sc_hd__a31o_1 _5373_ (.A1(_1748_),
    .A2(_1848_),
    .A3(_1884_),
    .B1(_1850_),
    .X(_2375_));
 sky130_fd_sc_hd__o211a_1 _5374_ (.A1(_1707_),
    .A2(_1850_),
    .B1(net463),
    .C1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__a31o_1 _5375_ (.A1(_1707_),
    .A2(_2258_),
    .A3(_1848_),
    .B1(_1711_),
    .X(_2377_));
 sky130_fd_sc_hd__a31o_1 _5376_ (.A1(_1707_),
    .A2(_1848_),
    .A3(_2258_),
    .B1(_1778_),
    .X(_2378_));
 sky130_fd_sc_hd__a31o_1 _5377_ (.A1(_2258_),
    .A2(_1848_),
    .A3(_1707_),
    .B1(_1721_),
    .X(_2379_));
 sky130_fd_sc_hd__a211o_1 _5378_ (.A1(_1707_),
    .A2(_1848_),
    .B1(_1745_),
    .C1(net458),
    .X(_2380_));
 sky130_fd_sc_hd__a211o_1 _5379_ (.A1(_1707_),
    .A2(_1848_),
    .B1(_1741_),
    .C1(net457),
    .X(_2381_));
 sky130_fd_sc_hd__a311o_1 _5380_ (.A1(_2258_),
    .A2(_1848_),
    .A3(_1707_),
    .B1(_1741_),
    .C1(net458),
    .X(_2382_));
 sky130_fd_sc_hd__o31a_1 _5381_ (.A1(_1704_),
    .A2(net458),
    .A3(_1724_),
    .B1(_2085_),
    .X(_2383_));
 sky130_fd_sc_hd__o311a_1 _5382_ (.A1(_1609_),
    .A2(net457),
    .A3(_1975_),
    .B1(_2262_),
    .C1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__o2111a_1 _5383_ (.A1(_2081_),
    .A2(_2258_),
    .B1(_2380_),
    .C1(_2382_),
    .D1(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__and3_1 _5384_ (.A(_2385_),
    .B(_2378_),
    .C(_2379_),
    .X(_2386_));
 sky130_fd_sc_hd__o41a_1 _5385_ (.A1(_1604_),
    .A2(_1706_),
    .A3(net453),
    .A4(_1847_),
    .B1(_1777_),
    .X(_2387_));
 sky130_fd_sc_hd__a211o_1 _5386_ (.A1(_1707_),
    .A2(_1848_),
    .B1(_1720_),
    .C1(net457),
    .X(_2388_));
 sky130_fd_sc_hd__and4b_1 _5387_ (.A_N(net616),
    .B(_1610_),
    .C(net543),
    .D(_1723_),
    .X(_2389_));
 sky130_fd_sc_hd__a41oi_4 _5388_ (.A1(net556),
    .A2(net542),
    .A3(_1723_),
    .A4(_2077_),
    .B1(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__a31o_1 _5389_ (.A1(_1605_),
    .A2(_1704_),
    .A3(_1848_),
    .B1(_1793_),
    .X(_2391_));
 sky130_fd_sc_hd__and3_1 _5390_ (.A(_2386_),
    .B(_2391_),
    .C(_2377_),
    .X(_2392_));
 sky130_fd_sc_hd__a41o_1 _5391_ (.A1(_1605_),
    .A2(_1707_),
    .A3(_1748_),
    .A4(_1848_),
    .B1(_1802_),
    .X(_2393_));
 sky130_fd_sc_hd__a311o_1 _5392_ (.A1(_2258_),
    .A2(_1848_),
    .A3(_1707_),
    .B1(_1810_),
    .C1(net457),
    .X(_2394_));
 sky130_fd_sc_hd__o41a_1 _5393_ (.A1(_1604_),
    .A2(_1706_),
    .A3(net453),
    .A4(_1847_),
    .B1(_2104_),
    .X(_2395_));
 sky130_fd_sc_hd__nand3_1 _5394_ (.A(_2392_),
    .B(_2393_),
    .C(_2394_),
    .Y(_2396_));
 sky130_fd_sc_hd__a31o_1 _5395_ (.A1(net554),
    .A2(_1712_),
    .A3(net529),
    .B1(_2280_),
    .X(_2397_));
 sky130_fd_sc_hd__a211o_1 _5396_ (.A1(_1821_),
    .A2(_1847_),
    .B1(_2396_),
    .C1(_2397_),
    .X(_2398_));
 sky130_fd_sc_hd__a211o_1 _5397_ (.A1(_1576_),
    .A2(_1831_),
    .B1(_2114_),
    .C1(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__a311o_1 _5398_ (.A1(_1713_),
    .A2(_1752_),
    .A3(net530),
    .B1(_1836_),
    .C1(_1830_),
    .X(_2400_));
 sky130_fd_sc_hd__nand4_1 _5399_ (.A(_1602_),
    .B(net551),
    .C(_1817_),
    .D(net450),
    .Y(_2401_));
 sky130_fd_sc_hd__nand3b_1 _5400_ (.A_N(_2399_),
    .B(_2400_),
    .C(_2401_),
    .Y(_2402_));
 sky130_fd_sc_hd__a31o_1 _5401_ (.A1(net364),
    .A2(_1602_),
    .A3(net553),
    .B1(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__a211o_1 _5402_ (.A1(_2376_),
    .A2(_2403_),
    .B1(net461),
    .C1(_2374_),
    .X(_2404_));
 sky130_fd_sc_hd__o32a_1 _5403_ (.A1(_2404_),
    .A2(_2347_),
    .A3(_2324_),
    .B1(net2295),
    .B2(_1539_),
    .X(_0374_));
 sky130_fd_sc_hd__nand4_1 _5404_ (.A(_1690_),
    .B(_1715_),
    .C(_1737_),
    .D(_1844_),
    .Y(_2405_));
 sky130_fd_sc_hd__and4bb_1 _5405_ (.A_N(_1760_),
    .B_N(_2137_),
    .C(_2405_),
    .D(_2303_),
    .X(_2406_));
 sky130_fd_sc_hd__a21oi_2 _5406_ (.A1(net618),
    .A2(_1823_),
    .B1(_1712_),
    .Y(_2407_));
 sky130_fd_sc_hd__a31o_1 _5407_ (.A1(net616),
    .A2(net121),
    .A3(net551),
    .B1(_1844_),
    .X(_2408_));
 sky130_fd_sc_hd__o21ai_2 _5408_ (.A1(_1712_),
    .A2(net535),
    .B1(_1690_),
    .Y(_2409_));
 sky130_fd_sc_hd__o311a_1 _5409_ (.A1(_1691_),
    .A2(_2407_),
    .A3(_1765_),
    .B1(_2143_),
    .C1(_2304_),
    .X(_2410_));
 sky130_fd_sc_hd__and3_1 _5410_ (.A(_1690_),
    .B(_1771_),
    .C(_2408_),
    .X(_2411_));
 sky130_fd_sc_hd__o211a_1 _5411_ (.A1(_2409_),
    .A2(_1773_),
    .B1(_2134_),
    .C1(_2307_),
    .X(_2412_));
 sky130_fd_sc_hd__o211a_1 _5412_ (.A1(_2407_),
    .A2(_1787_),
    .B1(_2133_),
    .C1(_2311_),
    .X(_2413_));
 sky130_fd_sc_hd__and4_1 _5413_ (.A(_2406_),
    .B(_2410_),
    .C(_2412_),
    .D(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__o2111ai_2 _5414_ (.A1(_1712_),
    .A2(net535),
    .B1(_1737_),
    .C1(_1637_),
    .D1(_1690_),
    .Y(_2415_));
 sky130_fd_sc_hd__o221a_1 _5415_ (.A1(_1710_),
    .A2(_1800_),
    .B1(_1806_),
    .B2(_1763_),
    .C1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__and3_1 _5416_ (.A(_2315_),
    .B(_2414_),
    .C(_2416_),
    .X(_2417_));
 sky130_fd_sc_hd__o21ba_1 _5417_ (.A1(_1699_),
    .A2(_1736_),
    .B1_N(_2132_),
    .X(_2418_));
 sky130_fd_sc_hd__and3_1 _5418_ (.A(_2418_),
    .B(_1826_),
    .C(_2318_),
    .X(_2419_));
 sky130_fd_sc_hd__and3_1 _5419_ (.A(_2210_),
    .B(_2417_),
    .C(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__o311a_1 _5420_ (.A1(_1599_),
    .A2(_1629_),
    .A3(_1734_),
    .B1(_2168_),
    .C1(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__o32a_1 _5421_ (.A1(_1599_),
    .A2(_1609_),
    .A3(_1629_),
    .B1(_1838_),
    .B2(_1586_),
    .X(_2422_));
 sky130_fd_sc_hd__and4_1 _5422_ (.A(_2421_),
    .B(_2422_),
    .C(_1843_),
    .D(_2297_),
    .X(_2423_));
 sky130_fd_sc_hd__and2_1 _5423_ (.A(_2200_),
    .B(_2328_),
    .X(_2424_));
 sky130_fd_sc_hd__o22a_1 _5424_ (.A1(_1629_),
    .A2(_1691_),
    .B1(_1730_),
    .B2(_1884_),
    .X(_2425_));
 sky130_fd_sc_hd__a31o_2 _5425_ (.A1(net617),
    .A2(net398),
    .A3(net534),
    .B1(_1762_),
    .X(_2426_));
 sky130_fd_sc_hd__o211a_1 _5426_ (.A1(_1628_),
    .A2(_1883_),
    .B1(net425),
    .C1(net397),
    .X(_2427_));
 sky130_fd_sc_hd__a31o_1 _5427_ (.A1(_1865_),
    .A2(_1988_),
    .A3(_2426_),
    .B1(_2189_),
    .X(_2428_));
 sky130_fd_sc_hd__a31o_1 _5428_ (.A1(_1878_),
    .A2(net424),
    .A3(_2330_),
    .B1(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__o31a_1 _5429_ (.A1(_1712_),
    .A2(_1751_),
    .A3(net531),
    .B1(net552),
    .X(_2430_));
 sky130_fd_sc_hd__o21ai_1 _5430_ (.A1(_2430_),
    .A2(_2219_),
    .B1(net398),
    .Y(_2431_));
 sky130_fd_sc_hd__o211a_1 _5431_ (.A1(_1883_),
    .A2(_1960_),
    .B1(_1868_),
    .C1(net424),
    .X(_2432_));
 sky130_fd_sc_hd__a31o_1 _5432_ (.A1(_1577_),
    .A2(_1825_),
    .A3(_2177_),
    .B1(_2016_),
    .X(_2433_));
 sky130_fd_sc_hd__nand3b_1 _5433_ (.A_N(_2333_),
    .B(_2431_),
    .C(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__a221o_1 _5434_ (.A1(_1666_),
    .A2(_2331_),
    .B1(_2427_),
    .B2(_1867_),
    .C1(_2194_),
    .X(_2435_));
 sky130_fd_sc_hd__nor4_1 _5435_ (.A(_2432_),
    .B(_2434_),
    .C(_2435_),
    .D(_2429_),
    .Y(_2436_));
 sky130_fd_sc_hd__a31o_1 _5436_ (.A1(_1675_),
    .A2(_1988_),
    .A3(_2426_),
    .B1(_2173_),
    .X(_2437_));
 sky130_fd_sc_hd__a21oi_2 _5437_ (.A1(_1878_),
    .A2(_2331_),
    .B1(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__and4_1 _5438_ (.A(_2436_),
    .B(_1980_),
    .C(_2424_),
    .D(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__a32o_1 _5439_ (.A1(net552),
    .A2(_1682_),
    .A3(net532),
    .B1(net531),
    .B2(_2057_),
    .X(_2440_));
 sky130_fd_sc_hd__a21oi_1 _5440_ (.A1(net534),
    .A2(_2057_),
    .B1(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__and4bb_1 _5441_ (.A_N(_2343_),
    .B_N(_2344_),
    .C(_2439_),
    .D(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__a31o_1 _5442_ (.A1(net552),
    .A2(_1682_),
    .A3(_1883_),
    .B1(_2208_),
    .X(_2443_));
 sky130_fd_sc_hd__a21o_1 _5443_ (.A1(_1605_),
    .A2(_1876_),
    .B1(_1663_),
    .X(_2444_));
 sky130_fd_sc_hd__and4_1 _5444_ (.A(_2362_),
    .B(_2070_),
    .C(_1927_),
    .D(_2235_),
    .X(_2445_));
 sky130_fd_sc_hd__o211a_1 _5445_ (.A1(_1604_),
    .A2(_1847_),
    .B1(net360),
    .C1(_1723_),
    .X(_2446_));
 sky130_fd_sc_hd__o2111a_1 _5446_ (.A1(_1741_),
    .A2(_2069_),
    .B1(_2353_),
    .C1(_2218_),
    .D1(_1901_),
    .X(_2447_));
 sky130_fd_sc_hd__o41a_1 _5447_ (.A1(_1660_),
    .A2(_1730_),
    .A3(_1873_),
    .A4(_1892_),
    .B1(_2356_),
    .X(_2448_));
 sky130_fd_sc_hd__and4b_1 _5448_ (.A_N(_2446_),
    .B(_2447_),
    .C(_2448_),
    .D(_1888_),
    .X(_2449_));
 sky130_fd_sc_hd__o311a_1 _5449_ (.A1(_1571_),
    .A2(_1670_),
    .A3(_2069_),
    .B1(_1915_),
    .C1(_2230_),
    .X(_2450_));
 sky130_fd_sc_hd__and3b_1 _5450_ (.A_N(_2229_),
    .B(_2358_),
    .C(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__o311a_1 _5451_ (.A1(net458),
    .A2(_1724_),
    .A3(_1848_),
    .B1(_1888_),
    .C1(_2225_),
    .X(_2452_));
 sky130_fd_sc_hd__and3_1 _5452_ (.A(_2445_),
    .B(_2449_),
    .C(_2451_),
    .X(_2453_));
 sky130_fd_sc_hd__and3_1 _5453_ (.A(net361),
    .B(_1809_),
    .C(_1847_),
    .X(_2454_));
 sky130_fd_sc_hd__a2111o_1 _5454_ (.A1(net532),
    .A2(_1939_),
    .B1(_2241_),
    .C1(_2454_),
    .D1(_2349_),
    .X(_2455_));
 sky130_fd_sc_hd__o21ba_1 _5455_ (.A1(_1951_),
    .A2(_2248_),
    .B1_N(_2368_),
    .X(_2456_));
 sky130_fd_sc_hd__and4b_1 _5456_ (.A_N(_2455_),
    .B(_2444_),
    .C(_2453_),
    .D(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(_2457_),
    .B(_2371_),
    .Y(_2458_));
 sky130_fd_sc_hd__a31o_1 _5458_ (.A1(net552),
    .A2(_1657_),
    .A3(_1751_),
    .B1(_1964_),
    .X(_2459_));
 sky130_fd_sc_hd__a31o_1 _5459_ (.A1(_1604_),
    .A2(net552),
    .A3(_1657_),
    .B1(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__a211o_1 _5460_ (.A1(_1662_),
    .A2(_1847_),
    .B1(_2458_),
    .C1(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__and2b_1 _5461_ (.A_N(_1969_),
    .B(_2292_),
    .X(_2462_));
 sky130_fd_sc_hd__o311a_2 _5462_ (.A1(_1626_),
    .A2(_1658_),
    .A3(_1884_),
    .B1(_2462_),
    .C1(_1858_),
    .X(_2463_));
 sky130_fd_sc_hd__o2bb2a_1 _5463_ (.A1_N(_2463_),
    .A2_N(_2461_),
    .B1(_2443_),
    .B2(_2442_),
    .X(_2464_));
 sky130_fd_sc_hd__o21ai_1 _5464_ (.A1(_2296_),
    .A2(_2423_),
    .B1(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__a31o_1 _5465_ (.A1(_1605_),
    .A2(_1704_),
    .A3(_1848_),
    .B1(_2081_),
    .X(_2466_));
 sky130_fd_sc_hd__a211o_1 _5466_ (.A1(_1713_),
    .A2(_1726_),
    .B1(_1724_),
    .C1(net457),
    .X(_2467_));
 sky130_fd_sc_hd__and3_1 _5467_ (.A(_2082_),
    .B(_2466_),
    .C(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__a32o_1 _5468_ (.A1(_1570_),
    .A2(_1718_),
    .A3(net455),
    .B1(net558),
    .B2(net555),
    .X(_2469_));
 sky130_fd_sc_hd__o21ai_1 _5469_ (.A1(_2074_),
    .A2(_2469_),
    .B1(net542),
    .Y(_2470_));
 sky130_fd_sc_hd__o311a_1 _5470_ (.A1(_1609_),
    .A2(net457),
    .A3(_1975_),
    .B1(_2262_),
    .C1(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__o31a_2 _5471_ (.A1(net620),
    .A2(net562),
    .A3(_1603_),
    .B1(_1752_),
    .X(_2472_));
 sky130_fd_sc_hd__o2111a_1 _5472_ (.A1(_1778_),
    .A2(_2472_),
    .B1(_2388_),
    .C1(_2259_),
    .D1(_2270_),
    .X(_2473_));
 sky130_fd_sc_hd__and4b_1 _5473_ (.A_N(_1794_),
    .B(_2273_),
    .C(_2377_),
    .D(_2098_),
    .X(_2474_));
 sky130_fd_sc_hd__nand4_1 _5474_ (.A(_2468_),
    .B(_2471_),
    .C(_2473_),
    .D(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__a211o_1 _5475_ (.A1(_1726_),
    .A2(_1752_),
    .B1(_1810_),
    .C1(net457),
    .X(_2476_));
 sky130_fd_sc_hd__nand3_1 _5476_ (.A(_2276_),
    .B(_2393_),
    .C(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__a311o_1 _5477_ (.A1(net552),
    .A2(_1703_),
    .A3(net529),
    .B1(_2109_),
    .C1(_2397_),
    .X(_2478_));
 sky130_fd_sc_hd__nor3_1 _5478_ (.A(_2475_),
    .B(_2477_),
    .C(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__o31a_1 _5479_ (.A1(_1683_),
    .A2(_1818_),
    .A3(_1975_),
    .B1(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__o32a_1 _5480_ (.A1(_1707_),
    .A2(_1830_),
    .A3(_1836_),
    .B1(_1850_),
    .B2(_1713_),
    .X(_2481_));
 sky130_fd_sc_hd__and3_1 _5481_ (.A(_2286_),
    .B(_2401_),
    .C(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__nand3_1 _5482_ (.A(_2400_),
    .B(_2480_),
    .C(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__o311a_1 _5483_ (.A1(_1603_),
    .A2(_1609_),
    .A3(_1830_),
    .B1(_2376_),
    .C1(\wbbd_state[6] ),
    .X(_2484_));
 sky130_fd_sc_hd__a221o_1 _5484_ (.A1(net2087),
    .A2(net461),
    .B1(_2483_),
    .B2(_2484_),
    .C1(_2465_),
    .X(_0375_));
 sky130_fd_sc_hd__o211a_1 _5485_ (.A1(_2409_),
    .A2(_1717_),
    .B1(_2145_),
    .C1(_2298_),
    .X(_2485_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_2410_),
    .B(_2485_),
    .Y(_2486_));
 sky130_fd_sc_hd__o41a_1 _5487_ (.A1(net460),
    .A2(_1642_),
    .A3(_1772_),
    .A4(_2409_),
    .B1(_2155_),
    .X(_2487_));
 sky130_fd_sc_hd__nand3_1 _5488_ (.A(_2312_),
    .B(_2413_),
    .C(_2487_),
    .Y(_2488_));
 sky130_fd_sc_hd__a31o_1 _5489_ (.A1(net558),
    .A2(net363),
    .A3(net537),
    .B1(_2130_),
    .X(_2489_));
 sky130_fd_sc_hd__a211oi_2 _5490_ (.A1(_1628_),
    .A2(_1662_),
    .B1(_2054_),
    .C1(_2489_),
    .Y(_2490_));
 sky130_fd_sc_hd__and4_1 _5491_ (.A(_2419_),
    .B(_2320_),
    .C(_2165_),
    .D(_1700_),
    .X(_2491_));
 sky130_fd_sc_hd__and4bb_1 _5492_ (.A_N(_2486_),
    .B_N(_2488_),
    .C(_2490_),
    .D(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__o31ai_1 _5493_ (.A1(_1599_),
    .A2(_1836_),
    .A3(net530),
    .B1(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__o32a_1 _5494_ (.A1(_1599_),
    .A2(_1605_),
    .A3(_1609_),
    .B1(_1838_),
    .B2(_1586_),
    .X(_2494_));
 sky130_fd_sc_hd__a211o_1 _5495_ (.A1(_1629_),
    .A2(_1876_),
    .B1(_1599_),
    .C1(_1609_),
    .X(_2495_));
 sky130_fd_sc_hd__and3_1 _5496_ (.A(_1843_),
    .B(_2169_),
    .C(_2494_),
    .X(_2496_));
 sky130_fd_sc_hd__a31o_1 _5497_ (.A1(_1878_),
    .A2(net424),
    .A3(_2426_),
    .B1(_2175_),
    .X(_2497_));
 sky130_fd_sc_hd__a31o_1 _5498_ (.A1(_1867_),
    .A2(net424),
    .A3(_2330_),
    .B1(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__nor3b_1 _5499_ (.A(_2432_),
    .B(_2498_),
    .C_N(_2433_),
    .Y(_2499_));
 sky130_fd_sc_hd__a221o_1 _5500_ (.A1(_1867_),
    .A2(_2331_),
    .B1(_2427_),
    .B2(_1878_),
    .C1(_2174_),
    .X(_2500_));
 sky130_fd_sc_hd__nor2_1 _5501_ (.A(_2435_),
    .B(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hd__o311a_1 _5502_ (.A1(_1683_),
    .A2(_1836_),
    .A3(net530),
    .B1(_1980_),
    .C1(_2202_),
    .X(_2502_));
 sky130_fd_sc_hd__o311a_1 _5503_ (.A1(_1676_),
    .A2(_1877_),
    .A3(_1897_),
    .B1(_2326_),
    .C1(_2424_),
    .X(_2503_));
 sky130_fd_sc_hd__nand4_1 _5504_ (.A(_2499_),
    .B(_2501_),
    .C(_2502_),
    .D(_2503_),
    .Y(_2504_));
 sky130_fd_sc_hd__a31o_1 _5505_ (.A1(_1682_),
    .A2(_1751_),
    .A3(net536),
    .B1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__and4b_2 _5506_ (.A_N(_2208_),
    .B(_2294_),
    .C(_2346_),
    .D(_2441_),
    .X(_2506_));
 sky130_fd_sc_hd__o2111a_1 _5507_ (.A1(_1720_),
    .A2(_2069_),
    .B1(_2213_),
    .C1(_1881_),
    .D1(_2351_),
    .X(_2507_));
 sky130_fd_sc_hd__and3_2 _5508_ (.A(_2448_),
    .B(_2452_),
    .C(_2507_),
    .X(_2508_));
 sky130_fd_sc_hd__o311a_1 _5509_ (.A1(_1730_),
    .A2(_1800_),
    .A3(_1848_),
    .B1(_1932_),
    .C1(_2239_),
    .X(_2509_));
 sky130_fd_sc_hd__and3_1 _5510_ (.A(_2364_),
    .B(_2445_),
    .C(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__o311a_1 _5511_ (.A1(_1601_),
    .A2(_1663_),
    .A3(_2077_),
    .B1(_2444_),
    .C1(_2249_),
    .X(_2511_));
 sky130_fd_sc_hd__nand4_1 _5512_ (.A(_2370_),
    .B(_2508_),
    .C(_2510_),
    .D(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__a211o_1 _5513_ (.A1(_1712_),
    .A2(_1957_),
    .B1(_2368_),
    .C1(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__a22o_1 _5514_ (.A1(_2463_),
    .A2(_2513_),
    .B1(_2505_),
    .B2(_2506_),
    .X(_2514_));
 sky130_fd_sc_hd__a41o_1 _5515_ (.A1(_1854_),
    .A2(_1856_),
    .A3(_2290_),
    .A4(_2493_),
    .B1(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__o32a_1 _5516_ (.A1(net457),
    .A2(_1791_),
    .A3(_1950_),
    .B1(_1802_),
    .B2(_1713_),
    .X(_2516_));
 sky130_fd_sc_hd__o31a_1 _5517_ (.A1(net457),
    .A2(_1800_),
    .A3(_2472_),
    .B1(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__and3_1 _5518_ (.A(_2474_),
    .B(_2517_),
    .C(_2391_),
    .X(_2518_));
 sky130_fd_sc_hd__o211a_1 _5519_ (.A1(_1721_),
    .A2(_1726_),
    .B1(_2087_),
    .C1(_1722_),
    .X(_2519_));
 sky130_fd_sc_hd__nand3_1 _5520_ (.A(_2390_),
    .B(_2468_),
    .C(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__nand4_2 _5521_ (.A(_2390_),
    .B(_2468_),
    .C(_2518_),
    .D(_2519_),
    .Y(_2521_));
 sky130_fd_sc_hd__a211o_1 _5522_ (.A1(_1576_),
    .A2(_1831_),
    .B1(_2111_),
    .C1(_2114_),
    .X(_2522_));
 sky130_fd_sc_hd__a31o_1 _5523_ (.A1(_1703_),
    .A2(_1817_),
    .A3(net452),
    .B1(_1976_),
    .X(_2523_));
 sky130_fd_sc_hd__a311o_1 _5524_ (.A1(net552),
    .A2(_1703_),
    .A3(net529),
    .B1(_2522_),
    .C1(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__a2111o_1 _5525_ (.A1(_1821_),
    .A2(_1847_),
    .B1(_2397_),
    .C1(_2521_),
    .D1(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__a31o_1 _5526_ (.A1(net558),
    .A2(net449),
    .A3(net537),
    .B1(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__a221o_1 _5527_ (.A1(net2111),
    .A2(net461),
    .B1(_2484_),
    .B2(_2526_),
    .C1(_2515_),
    .X(_0376_));
 sky130_fd_sc_hd__o311a_1 _5528_ (.A1(_1599_),
    .A2(_1836_),
    .A3(net530),
    .B1(_2297_),
    .C1(_1856_),
    .X(_2527_));
 sky130_fd_sc_hd__and4_1 _5529_ (.A(_2168_),
    .B(_2495_),
    .C(_2496_),
    .D(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__o2111a_1 _5530_ (.A1(_1629_),
    .A2(_1838_),
    .B1(_1854_),
    .C1(_2164_),
    .D1(_2290_),
    .X(_2529_));
 sky130_fd_sc_hd__and4_1 _5531_ (.A(_2318_),
    .B(_2320_),
    .C(_1700_),
    .D(_1826_),
    .X(_2530_));
 sky130_fd_sc_hd__and4_1 _5532_ (.A(_2418_),
    .B(_2490_),
    .C(_2529_),
    .D(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__nand2_1 _5533_ (.A(_2528_),
    .B(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__a311oi_1 _5534_ (.A1(_1645_),
    .A2(_2408_),
    .A3(_1690_),
    .B1(_2162_),
    .C1(_2317_),
    .Y(_2533_));
 sky130_fd_sc_hd__and3_1 _5535_ (.A(_2315_),
    .B(_2416_),
    .C(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__o211ai_1 _5536_ (.A1(_1628_),
    .A2(net535),
    .B1(_1757_),
    .C1(_1690_),
    .Y(_2535_));
 sky130_fd_sc_hd__o211a_1 _5537_ (.A1(_1710_),
    .A2(_1739_),
    .B1(_1758_),
    .C1(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__and3_1 _5538_ (.A(_2301_),
    .B(_2406_),
    .C(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__and3b_1 _5539_ (.A_N(_2488_),
    .B(_2534_),
    .C(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__a2111oi_1 _5540_ (.A1(_1957_),
    .A2(_1960_),
    .B1(_2251_),
    .C1(_2373_),
    .D1(_1963_),
    .Y(_2539_));
 sky130_fd_sc_hd__and4bb_1 _5541_ (.A_N(_1959_),
    .B_N(_2460_),
    .C(_2539_),
    .D(_2444_),
    .X(_2540_));
 sky130_fd_sc_hd__o311a_1 _5542_ (.A1(_1626_),
    .A2(_1730_),
    .A3(_1752_),
    .B1(_2370_),
    .C1(_2463_),
    .X(_2541_));
 sky130_fd_sc_hd__and3_1 _5543_ (.A(_2456_),
    .B(_2540_),
    .C(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__o211a_1 _5544_ (.A1(_1847_),
    .A2(net532),
    .B1(_1661_),
    .C1(net361),
    .X(_2543_));
 sky130_fd_sc_hd__nor4_1 _5545_ (.A(_2245_),
    .B(_2366_),
    .C(_2455_),
    .D(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__o211a_1 _5546_ (.A1(_1745_),
    .A2(_1890_),
    .B1(_1895_),
    .C1(_1898_),
    .X(_2545_));
 sky130_fd_sc_hd__o2111a_2 _5547_ (.A1(_1745_),
    .A2(_2069_),
    .B1(_2354_),
    .C1(_2447_),
    .D1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__nand3_1 _5548_ (.A(_2510_),
    .B(_2544_),
    .C(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hd__a311oi_4 _5549_ (.A1(_1682_),
    .A2(_1751_),
    .A3(net536),
    .B1(_2344_),
    .C1(_2343_),
    .Y(_2548_));
 sky130_fd_sc_hd__nand4_2 _5550_ (.A(_2502_),
    .B(_2503_),
    .C(_2506_),
    .D(_2548_),
    .Y(_2549_));
 sky130_fd_sc_hd__o2111a_1 _5551_ (.A1(_1979_),
    .A2(_2425_),
    .B1(_2341_),
    .C1(_2172_),
    .D1(_2438_),
    .X(_2550_));
 sky130_fd_sc_hd__o211a_1 _5552_ (.A1(net532),
    .A2(_1883_),
    .B1(_2013_),
    .C1(net397),
    .X(_2551_));
 sky130_fd_sc_hd__a311oi_1 _5553_ (.A1(net424),
    .A2(_1988_),
    .A3(_2330_),
    .B1(_2551_),
    .C1(_2019_),
    .Y(_2552_));
 sky130_fd_sc_hd__and3_1 _5554_ (.A(_2332_),
    .B(_2431_),
    .C(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a31o_1 _5555_ (.A1(_2501_),
    .A2(_2550_),
    .A3(_2553_),
    .B1(_2549_),
    .X(_2554_));
 sky130_fd_sc_hd__o21ai_1 _5556_ (.A1(_2532_),
    .A2(_2538_),
    .B1(_2554_),
    .Y(_2555_));
 sky130_fd_sc_hd__a21o_1 _5557_ (.A1(_2542_),
    .A2(_2547_),
    .B1(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__a221o_1 _5558_ (.A1(net454),
    .A2(_1831_),
    .B1(_2119_),
    .B2(_1611_),
    .C1(_1976_),
    .X(_2557_));
 sky130_fd_sc_hd__nor4_1 _5559_ (.A(_2118_),
    .B(_2478_),
    .C(_2522_),
    .D(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__and3_1 _5560_ (.A(_2482_),
    .B(_2484_),
    .C(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__o31a_1 _5561_ (.A1(net457),
    .A2(_1818_),
    .A3(_2472_),
    .B1(_2279_),
    .X(_2560_));
 sky130_fd_sc_hd__nand4bb_1 _5562_ (.A_N(_2395_),
    .B_N(_2477_),
    .C(_2518_),
    .D(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__o311a_1 _5563_ (.A1(net457),
    .A2(_1726_),
    .A3(_1745_),
    .B1(_2084_),
    .C1(_2381_),
    .X(_2562_));
 sky130_fd_sc_hd__nand3_2 _5564_ (.A(_2265_),
    .B(_2471_),
    .C(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__o21a_1 _5565_ (.A1(_2561_),
    .A2(_2563_),
    .B1(_2559_),
    .X(_2564_));
 sky130_fd_sc_hd__a211o_1 _5566_ (.A1(net3856),
    .A2(net462),
    .B1(_2564_),
    .C1(_2556_),
    .X(_0377_));
 sky130_fd_sc_hd__a2111oi_1 _5567_ (.A1(_1644_),
    .A2(_2411_),
    .B1(_2309_),
    .C1(_2150_),
    .D1(_2149_),
    .Y(_2565_));
 sky130_fd_sc_hd__and3_1 _5568_ (.A(_2412_),
    .B(_2537_),
    .C(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__and3_1 _5569_ (.A(_2410_),
    .B(_2485_),
    .C(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__a31o_1 _5570_ (.A1(_1666_),
    .A2(net425),
    .A3(_2426_),
    .B1(_2192_),
    .X(_2568_));
 sky130_fd_sc_hd__a311oi_2 _5571_ (.A1(net425),
    .A2(_2329_),
    .A3(_1989_),
    .B1(_2568_),
    .C1(_2429_),
    .Y(_2569_));
 sky130_fd_sc_hd__and3_1 _5572_ (.A(_2499_),
    .B(_2553_),
    .C(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__and4b_1 _5573_ (.A_N(_2232_),
    .B(_2361_),
    .C(_1921_),
    .D(_2072_),
    .X(_2571_));
 sky130_fd_sc_hd__and2_1 _5574_ (.A(_2451_),
    .B(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__nand3_2 _5575_ (.A(_2508_),
    .B(_2546_),
    .C(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__o2bb2a_1 _5576_ (.A1_N(_2542_),
    .A2_N(_2573_),
    .B1(_2549_),
    .B2(_2570_),
    .X(_2574_));
 sky130_fd_sc_hd__o21ai_1 _5577_ (.A1(_2532_),
    .A2(_2567_),
    .B1(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__o2111ai_2 _5578_ (.A1(_1711_),
    .A2(_1726_),
    .B1(_2093_),
    .C1(_2257_),
    .D1(_2473_),
    .Y(_2576_));
 sky130_fd_sc_hd__o41a_2 _5579_ (.A1(_2387_),
    .A2(_2520_),
    .A3(_2563_),
    .A4(_2576_),
    .B1(_2559_),
    .X(_2577_));
 sky130_fd_sc_hd__a211o_1 _5580_ (.A1(net3864),
    .A2(net461),
    .B1(_2577_),
    .C1(_2575_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_4 _5581_ (.A(_1052_),
    .B(net502),
    .Y(_2578_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(net496),
    .A1(net3729),
    .S(_2578_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net491),
    .A1(net3560),
    .S(_2578_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _5584_ (.A0(net485),
    .A1(net2408),
    .S(_2578_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(net480),
    .A1(net2566),
    .S(_2578_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(net476),
    .A1(net3333),
    .S(_2578_),
    .X(_0383_));
 sky130_fd_sc_hd__and4_1 _5587_ (.A(net660),
    .B(net417),
    .C(net386),
    .D(net501),
    .X(_2579_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net3750),
    .A1(net495),
    .S(_2579_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(net3119),
    .A1(net489),
    .S(_2579_),
    .X(_0393_));
 sky130_fd_sc_hd__and4_4 _5590_ (.A(net419),
    .B(net2092),
    .C(net372),
    .D(net501),
    .X(_2580_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net3653),
    .A1(net495),
    .S(_2580_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(net3107),
    .A1(net489),
    .S(_2580_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net2545),
    .A1(net484),
    .S(_2580_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(net3133),
    .A1(net479),
    .S(_2580_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(net3641),
    .A1(net474),
    .S(_2580_),
    .X(_0398_));
 sky130_fd_sc_hd__and4_4 _5596_ (.A(net410),
    .B(net2092),
    .C(net372),
    .D(net501),
    .X(_2581_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net3675),
    .A1(net495),
    .S(_2581_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(net3155),
    .A1(net489),
    .S(_2581_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net2536),
    .A1(net484),
    .S(_2581_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(net3058),
    .A1(net479),
    .S(_2581_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net3650),
    .A1(net474),
    .S(_2581_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _5602_ (.A0(net2311),
    .A1(net472),
    .S(_2581_),
    .X(_0404_));
 sky130_fd_sc_hd__and3_4 _5603_ (.A(net385),
    .B(net376),
    .C(net501),
    .X(_2582_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(net3793),
    .A1(net495),
    .S(_2582_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(net3063),
    .A1(net489),
    .S(_2582_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(net2632),
    .A1(net484),
    .S(_2582_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _5607_ (.A0(net3102),
    .A1(net479),
    .S(_2582_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(net3656),
    .A1(net474),
    .S(_2582_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _5609_ (.A0(net2272),
    .A1(net472),
    .S(_2582_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(net3226),
    .A1(net468),
    .S(_2582_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(net2712),
    .A1(net465),
    .S(_2582_),
    .X(_0412_));
 sky130_fd_sc_hd__and4_1 _5612_ (.A(net660),
    .B(net385),
    .C(net410),
    .D(net501),
    .X(_2583_));
 sky130_fd_sc_hd__mux2_1 _5613_ (.A0(net3782),
    .A1(net495),
    .S(_2583_),
    .X(_0413_));
 sky130_fd_sc_hd__and3_2 _5614_ (.A(net383),
    .B(net756),
    .C(net671),
    .X(_2584_));
 sky130_fd_sc_hd__mux2_1 _5615_ (.A0(net3322),
    .A1(net497),
    .S(net2043),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(net2874),
    .A1(net490),
    .S(net2043),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _5617_ (.A0(net799),
    .A1(net486),
    .S(net2043),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _5618_ (.A0(net2560),
    .A1(net480),
    .S(net2043),
    .X(_0417_));
 sky130_fd_sc_hd__and3_1 _5619_ (.A(net906),
    .B(net374),
    .C(net501),
    .X(_2585_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(net3696),
    .A1(net495),
    .S(_2585_),
    .X(_0418_));
 sky130_fd_sc_hd__a31o_1 _5621_ (.A1(net660),
    .A2(net419),
    .A3(net906),
    .B1(net3564),
    .X(_2586_));
 sky130_fd_sc_hd__o211a_1 _5622_ (.A1(_1306_),
    .A2(net495),
    .B1(net1867),
    .C1(net501),
    .X(_0419_));
 sky130_fd_sc_hd__and3_4 _5623_ (.A(net372),
    .B(net370),
    .C(net501),
    .X(_2587_));
 sky130_fd_sc_hd__mux2_1 _5624_ (.A0(net3662),
    .A1(net474),
    .S(_2587_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _5625_ (.A0(net3089),
    .A1(net479),
    .S(_2587_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _5626_ (.A0(net2667),
    .A1(net484),
    .S(_2587_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net2336),
    .A1(net472),
    .S(_2587_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _5628_ (.A0(net3255),
    .A1(net468),
    .S(_2587_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _5629_ (.A0(net3077),
    .A1(net489),
    .S(_2587_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(net3755),
    .A1(net495),
    .S(_0959_),
    .X(_2588_));
 sky130_fd_sc_hd__and2_1 _5631_ (.A(net501),
    .B(net1930),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _5632_ (.A(net380),
    .B(net375),
    .C(net504),
    .X(_2589_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(net3623),
    .A1(net498),
    .S(_2589_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_2 _5634_ (.A(_1049_),
    .B(net504),
    .Y(_2590_));
 sky130_fd_sc_hd__mux2_1 _5635_ (.A0(net488),
    .A1(net2184),
    .S(_2590_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(net478),
    .A1(net2703),
    .S(_2590_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _5637_ (.A0(net492),
    .A1(net3514),
    .S(_2590_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _5638_ (.A0(net482),
    .A1(net2516),
    .S(_2590_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(net1088),
    .A1(net2746),
    .S(_2590_),
    .X(_0432_));
 sky130_fd_sc_hd__and4_1 _5640_ (.A(net417),
    .B(net415),
    .C(net372),
    .D(net501),
    .X(_2591_));
 sky130_fd_sc_hd__mux2_1 _5641_ (.A0(net3670),
    .A1(net495),
    .S(_2591_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _5642_ (.A0(net3186),
    .A1(net489),
    .S(_2591_),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_8 _5643_ (.A(_1016_),
    .B(net504),
    .Y(_2592_));
 sky130_fd_sc_hd__mux2_1 _5644_ (.A0(net495),
    .A1(net3687),
    .S(_2592_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(net489),
    .A1(net3051),
    .S(_2592_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _5646_ (.A0(net488),
    .A1(net2803),
    .S(_2592_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _5647_ (.A0(net479),
    .A1(net3110),
    .S(_2592_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(net477),
    .A1(net3258),
    .S(_2592_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _5649_ (.A0(net473),
    .A1(net2080),
    .S(_2592_),
    .X(_0440_));
 sky130_fd_sc_hd__o311ai_4 _5650_ (.A1(hkspi_disable),
    .A2(net908),
    .A3(net67),
    .B1(_0935_),
    .C1(net671),
    .Y(_2593_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(net497),
    .A1(net3373),
    .S(net351),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _5652_ (.A0(net490),
    .A1(net2918),
    .S(net351),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(net486),
    .A1(net2055),
    .S(_2593_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(net480),
    .A1(net2460),
    .S(net352),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(net708),
    .A1(net3173),
    .S(net352),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _5656_ (.A0(net472),
    .A1(net2355),
    .S(net352),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(net468),
    .A1(net3170),
    .S(net351),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _5658_ (.A0(net465),
    .A1(net2807),
    .S(net351),
    .X(_0448_));
 sky130_fd_sc_hd__and3_4 _5659_ (.A(net383),
    .B(net373),
    .C(net502),
    .X(_2594_));
 sky130_fd_sc_hd__mux2_1 _5660_ (.A0(net3359),
    .A1(net497),
    .S(_2594_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(net2963),
    .A1(net490),
    .S(_2594_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(net2147),
    .A1(net486),
    .S(_2594_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(net2485),
    .A1(net480),
    .S(_2594_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(net2975),
    .A1(net708),
    .S(_2594_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(net2928),
    .A1(net471),
    .S(_2594_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _5666_ (.A0(net3198),
    .A1(net468),
    .S(_2594_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _5667_ (.A0(net2843),
    .A1(net465),
    .S(_2594_),
    .X(_0456_));
 sky130_fd_sc_hd__nand2_8 _5668_ (.A(net2093),
    .B(net502),
    .Y(_2595_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(net497),
    .A1(net3436),
    .S(_2595_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(net490),
    .A1(net3094),
    .S(_2595_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(net486),
    .A1(net821),
    .S(net2094),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(net480),
    .A1(net2396),
    .S(net2094),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _5673_ (.A0(net708),
    .A1(net2906),
    .S(net2094),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(net471),
    .A1(net2805),
    .S(net2094),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(net468),
    .A1(net3049),
    .S(net2094),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(net465),
    .A1(net2810),
    .S(net2094),
    .X(_0464_));
 sky130_fd_sc_hd__and3_4 _5677_ (.A(net636),
    .B(net377),
    .C(net671),
    .X(_2596_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(net3381),
    .A1(net497),
    .S(_2596_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _5679_ (.A0(net2869),
    .A1(net490),
    .S(_2596_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _5680_ (.A0(net2063),
    .A1(net486),
    .S(_2596_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(net2340),
    .A1(net480),
    .S(_2596_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _5682_ (.A0(net3142),
    .A1(net708),
    .S(_2596_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _5683_ (.A0(net2969),
    .A1(net471),
    .S(_2596_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(net3218),
    .A1(net468),
    .S(_2596_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(net2827),
    .A1(net465),
    .S(_2596_),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_8 _5686_ (.A(_0895_),
    .B(net671),
    .Y(_2597_));
 sky130_fd_sc_hd__mux2_1 _5687_ (.A0(net497),
    .A1(net3366),
    .S(_2597_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(net490),
    .A1(net2952),
    .S(_2597_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(net486),
    .A1(net2076),
    .S(_2597_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _5690_ (.A0(net480),
    .A1(net2389),
    .S(_2597_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(net708),
    .A1(net2958),
    .S(_2597_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _5692_ (.A0(net471),
    .A1(net3008),
    .S(_2597_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(net468),
    .A1(net3178),
    .S(_2597_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(net465),
    .A1(net2833),
    .S(_2597_),
    .X(_0480_));
 sky130_fd_sc_hd__and3_4 _5695_ (.A(net387),
    .B(net377),
    .C(net502),
    .X(_2598_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(net3216),
    .A1(net497),
    .S(_2598_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(net2879),
    .A1(net490),
    .S(_2598_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(net2221),
    .A1(net486),
    .S(_2598_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(net2424),
    .A1(net480),
    .S(_2598_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(net3075),
    .A1(net708),
    .S(_2598_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(net3066),
    .A1(net471),
    .S(_2598_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(net3211),
    .A1(net468),
    .S(_2598_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _5703_ (.A0(net2799),
    .A1(net465),
    .S(_2598_),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_8 _5704_ (.A(_0939_),
    .B(net502),
    .Y(_2599_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(net497),
    .A1(net3362),
    .S(_2599_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(net490),
    .A1(net2946),
    .S(_2599_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(net486),
    .A1(net2523),
    .S(_2599_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(net480),
    .A1(net2678),
    .S(_2599_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(net708),
    .A1(net2956),
    .S(_2599_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(net471),
    .A1(net2923),
    .S(_2599_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(net469),
    .A1(net3250),
    .S(_2599_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(net465),
    .A1(net2853),
    .S(_2599_),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_8 _5713_ (.A(_0944_),
    .B(net671),
    .Y(_2600_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(net496),
    .A1(net3658),
    .S(_2600_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _5715_ (.A0(net490),
    .A1(net2881),
    .S(_2600_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(net486),
    .A1(net2047),
    .S(_2600_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(net480),
    .A1(net2246),
    .S(_2600_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(net474),
    .A1(net3580),
    .S(_2600_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(net471),
    .A1(net2839),
    .S(_2600_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(net468),
    .A1(net3189),
    .S(_2600_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(net465),
    .A1(net2801),
    .S(_2600_),
    .X(_0504_));
 sky130_fd_sc_hd__and4_4 _5722_ (.A(net417),
    .B(net416),
    .C(net377),
    .D(net502),
    .X(_2601_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(net3342),
    .A1(net497),
    .S(_2601_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(net1210),
    .A1(net490),
    .S(_2601_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(net2059),
    .A1(net486),
    .S(_2601_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(net2427),
    .A1(net481),
    .S(_2601_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net2984),
    .A1(net708),
    .S(_2601_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(net2317),
    .A1(net472),
    .S(_2601_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(net3235),
    .A1(net468),
    .S(_2601_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(net2887),
    .A1(net466),
    .S(_2601_),
    .X(_0512_));
 sky130_fd_sc_hd__and3_4 _5731_ (.A(net383),
    .B(net377),
    .C(net671),
    .X(_2602_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(net3789),
    .A1(net495),
    .S(_2602_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _5733_ (.A0(net2864),
    .A1(net490),
    .S(_2602_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(net2646),
    .A1(net484),
    .S(_2602_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5735_ (.A0(net2006),
    .A1(net2027),
    .S(_2602_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(net2911),
    .A1(net708),
    .S(_2602_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _5737_ (.A0(net3047),
    .A1(net471),
    .S(_2602_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(net3140),
    .A1(net468),
    .S(_2602_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(net2823),
    .A1(net465),
    .S(_2602_),
    .X(_0520_));
 sky130_fd_sc_hd__and3_4 _5740_ (.A(net392),
    .B(net404),
    .C(net504),
    .X(_2603_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(net3769),
    .A1(net498),
    .S(_2603_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _5742_ (.A0(net3616),
    .A1(net492),
    .S(_2603_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(net2198),
    .A1(net486),
    .S(_2603_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(net2526),
    .A1(net481),
    .S(_2603_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(net2734),
    .A1(net478),
    .S(_2603_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(net3184),
    .A1(net471),
    .S(_2603_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(net3240),
    .A1(net469),
    .S(_2603_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5748_ (.A0(net2885),
    .A1(net466),
    .S(_2603_),
    .X(_0528_));
 sky130_fd_sc_hd__and3_4 _5749_ (.A(net390),
    .B(net636),
    .C(net502),
    .X(_2604_));
 sky130_fd_sc_hd__mux2_1 _5750_ (.A0(net3368),
    .A1(net497),
    .S(_2604_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(net3146),
    .A1(net490),
    .S(_2604_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5752_ (.A0(net2585),
    .A1(net484),
    .S(_2604_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(net2268),
    .A1(net480),
    .S(_2604_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _5754_ (.A0(net3621),
    .A1(net474),
    .S(_2604_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5755_ (.A0(net2980),
    .A1(net471),
    .S(_2604_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(net3068),
    .A1(net468),
    .S(_2604_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _5757_ (.A0(net2795),
    .A1(net465),
    .S(_2604_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_8 _5758_ (.A(_0901_),
    .B(net672),
    .Y(_2605_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(net498),
    .A1(net3589),
    .S(_2605_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(net667),
    .A1(net2377),
    .S(_2605_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _5761_ (.A0(net486),
    .A1(net2321),
    .S(_2605_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(net481),
    .A1(net2330),
    .S(_2605_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(net477),
    .A1(net3290),
    .S(_2605_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(net471),
    .A1(net3080),
    .S(_2605_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(net468),
    .A1(net3245),
    .S(_2605_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(net465),
    .A1(net2815),
    .S(_2605_),
    .X(_0544_));
 sky130_fd_sc_hd__and3_4 _5767_ (.A(net392),
    .B(_0867_),
    .C(net504),
    .X(_2606_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net3701),
    .A1(net498),
    .S(_2606_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _5769_ (.A0(net3556),
    .A1(net492),
    .S(_2606_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(net2214),
    .A1(net488),
    .S(_2606_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(net2519),
    .A1(net481),
    .S(_2606_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(net3266),
    .A1(net477),
    .S(_2606_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _5773_ (.A0(net3006),
    .A1(net471),
    .S(_2606_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(net3260),
    .A1(net469),
    .S(_2606_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(net2234),
    .A1(net641),
    .S(_2606_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_0938_),
    .B(net672),
    .Y(_2607_));
 sky130_fd_sc_hd__mux2_1 _5777_ (.A0(net498),
    .A1(net3703),
    .S(net673),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(net667),
    .A1(net2369),
    .S(net673),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(net486),
    .A1(net2224),
    .S(net673),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(net481),
    .A1(net2281),
    .S(net673),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(net477),
    .A1(net3264),
    .S(net673),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(net471),
    .A1(net2954),
    .S(net673),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(net469),
    .A1(net3191),
    .S(net673),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(net466),
    .A1(net2898),
    .S(net673),
    .X(_0560_));
 sky130_fd_sc_hd__and3_4 _5785_ (.A(net392),
    .B(net388),
    .C(net504),
    .X(_2608_));
 sky130_fd_sc_hd__mux2_1 _5786_ (.A0(net1191),
    .A1(net1088),
    .S(_2608_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(net2013),
    .A1(net493),
    .S(_2608_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _5788_ (.A0(net3071),
    .A1(net487),
    .S(_2608_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(net2398),
    .A1(net481),
    .S(_2608_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _5790_ (.A0(net2767),
    .A1(net478),
    .S(_2608_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(net3021),
    .A1(net471),
    .S(_2608_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(net3207),
    .A1(net469),
    .S(_2608_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(net2872),
    .A1(net466),
    .S(_2608_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_8 _5794_ (.A(_0865_),
    .B(net671),
    .Y(_2609_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(net497),
    .A1(net3534),
    .S(_2609_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(net490),
    .A1(net3129),
    .S(_2609_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(net486),
    .A1(net2413),
    .S(_2609_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _5798_ (.A0(net481),
    .A1(net2563),
    .S(_2609_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _5799_ (.A0(net477),
    .A1(net3288),
    .S(_2609_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _5800_ (.A0(net471),
    .A1(net2876),
    .S(_2609_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(net469),
    .A1(net3166),
    .S(_2609_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _5802_ (.A0(net465),
    .A1(net2861),
    .S(_2609_),
    .X(_0576_));
 sky130_fd_sc_hd__and3_4 _5803_ (.A(net390),
    .B(net383),
    .C(net502),
    .X(_2610_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(net3797),
    .A1(net495),
    .S(_2610_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _5805_ (.A0(net3138),
    .A1(net489),
    .S(_2610_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _5806_ (.A0(net2589),
    .A1(net484),
    .S(_2610_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(net2481),
    .A1(net480),
    .S(_2610_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(net3026),
    .A1(net708),
    .S(_2610_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(net2921),
    .A1(net471),
    .S(_2610_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(net3238),
    .A1(net468),
    .S(_2610_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(net2916),
    .A1(net465),
    .S(_2610_),
    .X(_0584_));
 sky130_fd_sc_hd__and3_4 _5812_ (.A(net358),
    .B(net404),
    .C(net505),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5813_ (.A0(net3482),
    .A1(net499),
    .S(_2611_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(net3220),
    .A1(net490),
    .S(_2611_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _5815_ (.A0(net2615),
    .A1(net485),
    .S(_2611_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(net2533),
    .A1(net481),
    .S(_2611_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _5817_ (.A0(net3305),
    .A1(net477),
    .S(_2611_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _5818_ (.A0(net2966),
    .A1(net471),
    .S(_2611_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(net3150),
    .A1(net469),
    .S(_2611_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _5820_ (.A0(net2913),
    .A1(net465),
    .S(_2611_),
    .X(_0592_));
 sky130_fd_sc_hd__and3_4 _5821_ (.A(net358),
    .B(net636),
    .C(net505),
    .X(_2612_));
 sky130_fd_sc_hd__mux2_1 _5822_ (.A0(net3744),
    .A1(net498),
    .S(_2612_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _5823_ (.A0(net3213),
    .A1(net490),
    .S(_2612_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _5824_ (.A0(net2502),
    .A1(net486),
    .S(_2612_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(net2640),
    .A1(net481),
    .S(_2612_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _5826_ (.A0(net3317),
    .A1(net477),
    .S(_2612_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(net2173),
    .A1(net472),
    .S(_2612_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(net3230),
    .A1(net469),
    .S(_2612_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _5829_ (.A0(net2908),
    .A1(net466),
    .S(_2612_),
    .X(_0600_));
 sky130_fd_sc_hd__and4_4 _5830_ (.A(net646),
    .B(net358),
    .C(net414),
    .D(net504),
    .X(_2613_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(net3741),
    .A1(net498),
    .S(_2613_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(net3546),
    .A1(net492),
    .S(_2613_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(net2439),
    .A1(net486),
    .S(_2613_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _5834_ (.A0(net2624),
    .A1(net481),
    .S(_2613_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(net3330),
    .A1(net477),
    .S(_2613_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(net2305),
    .A1(net473),
    .S(_2613_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(net3204),
    .A1(net469),
    .S(_2613_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(net2158),
    .A1(net641),
    .S(_2613_),
    .X(_0608_));
 sky130_fd_sc_hd__and3_4 _5839_ (.A(net358),
    .B(_0867_),
    .C(net504),
    .X(_2614_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(net3454),
    .A1(net499),
    .S(_2614_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(net3628),
    .A1(net492),
    .S(_2614_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _5842_ (.A0(net3031),
    .A1(net487),
    .S(_2614_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(net2291),
    .A1(net482),
    .S(_2614_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(net2727),
    .A1(net478),
    .S(_2614_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(net2124),
    .A1(net473),
    .S(_2614_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(net2496),
    .A1(net685),
    .S(_2614_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _5847_ (.A0(net651),
    .A1(net641),
    .S(_2614_),
    .X(_0616_));
 sky130_fd_sc_hd__nand2_8 _5848_ (.A(_0861_),
    .B(net672),
    .Y(_2615_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(net1088),
    .A1(net2684),
    .S(_2615_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(net492),
    .A1(net3283),
    .S(_2615_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(net488),
    .A1(net2508),
    .S(_2615_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(net483),
    .A1(net2568),
    .S(_2615_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(net478),
    .A1(net2774),
    .S(_2615_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(net473),
    .A1(net2191),
    .S(_2615_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _5855_ (.A0(net685),
    .A1(net2493),
    .S(_2615_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(net466),
    .A1(net2903),
    .S(_2615_),
    .X(_0624_));
 sky130_fd_sc_hd__nand2_8 _5857_ (.A(_0913_),
    .B(net671),
    .Y(_2616_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(net498),
    .A1(net3699),
    .S(_2616_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(net667),
    .A1(net2499),
    .S(_2616_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(net486),
    .A1(net2431),
    .S(_2616_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(net481),
    .A1(net2467),
    .S(_2616_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(net477),
    .A1(net3279),
    .S(_2616_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(net472),
    .A1(net2308),
    .S(_2616_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(net469),
    .A1(net3182),
    .S(_2616_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(net466),
    .A1(net2856),
    .S(_2616_),
    .X(_0632_));
 sky130_fd_sc_hd__and4_4 _5866_ (.A(net646),
    .B(net358),
    .C(net416),
    .D(net504),
    .X(_2617_));
 sky130_fd_sc_hd__mux2_1 _5867_ (.A0(net3574),
    .A1(net498),
    .S(_2617_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(net3509),
    .A1(net492),
    .S(_2617_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(net2470),
    .A1(net488),
    .S(_2617_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(net2364),
    .A1(net482),
    .S(_2617_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(net3299),
    .A1(net477),
    .S(_2617_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(net2105),
    .A1(net473),
    .S(_2617_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(net2380),
    .A1(net685),
    .S(_2617_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(net2836),
    .A1(net466),
    .S(_2617_),
    .X(_0640_));
 sky130_fd_sc_hd__and3_4 _5875_ (.A(net359),
    .B(net383),
    .C(net502),
    .X(_2618_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(net3777),
    .A1(net498),
    .S(_2618_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(net2895),
    .A1(net490),
    .S(_2618_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(net2051),
    .A1(net486),
    .S(_2618_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _5879_ (.A0(net2551),
    .A1(net481),
    .S(_2618_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(net3296),
    .A1(net477),
    .S(_2618_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _5881_ (.A0(net3195),
    .A1(net471),
    .S(_2618_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(net3242),
    .A1(net468),
    .S(_2618_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _5883_ (.A0(net3003),
    .A1(net465),
    .S(_2618_),
    .X(_0648_));
 sky130_fd_sc_hd__and3_4 _5884_ (.A(net356),
    .B(net404),
    .C(net504),
    .X(_2619_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(net2738),
    .A1(net1088),
    .S(net2116),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _5886_ (.A0(net3228),
    .A1(net492),
    .S(net2116),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _5887_ (.A0(net837),
    .A1(net488),
    .S(net2116),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(net2244),
    .A1(net482),
    .S(net2116),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(net3320),
    .A1(net477),
    .S(net2116),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _5890_ (.A0(net2205),
    .A1(net473),
    .S(net2116),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _5891_ (.A0(net2375),
    .A1(net685),
    .S(net2116),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(net2891),
    .A1(net466),
    .S(net2116),
    .X(_0656_));
 sky130_fd_sc_hd__nand2_8 _5893_ (.A(net2071),
    .B(net502),
    .Y(_2620_));
 sky130_fd_sc_hd__mux2_1 _5894_ (.A0(net498),
    .A1(net3718),
    .S(net2072),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _5895_ (.A0(net492),
    .A1(net3512),
    .S(net2072),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(net486),
    .A1(net2491),
    .S(net2072),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(net481),
    .A1(net2422),
    .S(net2072),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _5898_ (.A0(net478),
    .A1(net720),
    .S(net2072),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _5899_ (.A0(net473),
    .A1(net811),
    .S(net2072),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _5900_ (.A0(net469),
    .A1(net3160),
    .S(net2072),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(net466),
    .A1(net2825),
    .S(net2072),
    .X(_0664_));
 sky130_fd_sc_hd__nand2_8 _5902_ (.A(_0880_),
    .B(net502),
    .Y(_2621_));
 sky130_fd_sc_hd__mux2_1 _5903_ (.A0(net497),
    .A1(net3505),
    .S(_2621_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(net490),
    .A1(net3572),
    .S(_2621_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _5905_ (.A0(net484),
    .A1(net2231),
    .S(_2621_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(net481),
    .A1(net2195),
    .S(_2621_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _5907_ (.A0(net708),
    .A1(net2941),
    .S(_2621_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(net473),
    .A1(net2128),
    .S(_2621_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _5909_ (.A0(net468),
    .A1(net3180),
    .S(_2621_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(net466),
    .A1(net2866),
    .S(_2621_),
    .X(_0672_));
 sky130_fd_sc_hd__and3_4 _5911_ (.A(_0867_),
    .B(net356),
    .C(net504),
    .X(_2622_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(net2841),
    .A1(net1088),
    .S(_2622_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _5913_ (.A0(net3585),
    .A1(net492),
    .S(_2622_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _5914_ (.A0(net2978),
    .A1(net487),
    .S(_2622_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _5915_ (.A0(net2252),
    .A1(net482),
    .S(_2622_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(net2749),
    .A1(net478),
    .S(_2622_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _5917_ (.A0(net2177),
    .A1(net473),
    .S(_2622_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _5918_ (.A0(net700),
    .A1(net685),
    .S(_2622_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _5919_ (.A0(net2926),
    .A1(net466),
    .S(_2622_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_8 _5920_ (.A(_0933_),
    .B(net504),
    .Y(_2623_));
 sky130_fd_sc_hd__mux2_1 _5921_ (.A0(net498),
    .A1(net3582),
    .S(_2623_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _5922_ (.A0(net492),
    .A1(net3223),
    .S(_2623_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _5923_ (.A0(net488),
    .A1(net2140),
    .S(_2623_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _5924_ (.A0(net482),
    .A1(net2166),
    .S(_2623_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(net477),
    .A1(net3233),
    .S(_2623_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(net473),
    .A1(net2084),
    .S(_2623_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _5927_ (.A0(net685),
    .A1(net2324),
    .S(_2623_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _5928_ (.A0(net466),
    .A1(net2820),
    .S(_2623_),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_8 _5929_ (.A(_0921_),
    .B(net504),
    .Y(_2624_));
 sky130_fd_sc_hd__mux2_1 _5930_ (.A0(net1088),
    .A1(net2818),
    .S(_2624_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(net492),
    .A1(net3503),
    .S(_2624_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _5932_ (.A0(net488),
    .A1(net2465),
    .S(_2624_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _5933_ (.A0(net482),
    .A1(net2489),
    .S(_2624_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _5934_ (.A0(net477),
    .A1(net3286),
    .S(_2624_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(net473),
    .A1(net2188),
    .S(_2624_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _5936_ (.A0(net685),
    .A1(net2434),
    .S(_2624_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(net641),
    .A1(net2134),
    .S(_2624_),
    .X(_0696_));
 sky130_fd_sc_hd__and4_1 _5938_ (.A(net646),
    .B(net416),
    .C(net356),
    .D(net504),
    .X(_2625_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(net3707),
    .A1(net498),
    .S(net647),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _5940_ (.A0(net2690),
    .A1(net493),
    .S(net647),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(net2327),
    .A1(net488),
    .S(net647),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(net2227),
    .A1(net482),
    .S(net647),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(net2700),
    .A1(net478),
    .S(net647),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(net2154),
    .A1(net473),
    .S(net647),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(net2358),
    .A1(net685),
    .S(net647),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _5946_ (.A0(net2120),
    .A1(net641),
    .S(net647),
    .X(_0704_));
 sky130_fd_sc_hd__and3_4 _5947_ (.A(net383),
    .B(net355),
    .C(net671),
    .X(_2626_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(net3787),
    .A1(net495),
    .S(_2626_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _5949_ (.A0(net2859),
    .A1(net490),
    .S(_2626_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(net2630),
    .A1(net484),
    .S(_2626_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _5951_ (.A0(net2448),
    .A1(net480),
    .S(_2626_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _5952_ (.A0(net2893),
    .A1(net708),
    .S(_2626_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _5953_ (.A0(net2994),
    .A1(net471),
    .S(_2626_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(net3193),
    .A1(net468),
    .S(_2626_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _5955_ (.A0(net2883),
    .A1(net465),
    .S(_2626_),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _5956_ (.A(net382),
    .B(net405),
    .C(net672),
    .X(_2627_));
 sky130_fd_sc_hd__mux2_1 _5957_ (.A0(net3720),
    .A1(net498),
    .S(net757),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _5958_ (.A0(net3529),
    .A1(net492),
    .S(net757),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _5959_ (.A0(net2162),
    .A1(net488),
    .S(net757),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _5960_ (.A0(net2386),
    .A1(net481),
    .S(net757),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _5961_ (.A0(net3268),
    .A1(net477),
    .S(net757),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(net2258),
    .A1(net473),
    .S(net757),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _5963_ (.A0(net2530),
    .A1(net685),
    .S(net757),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(net2931),
    .A1(net466),
    .S(net757),
    .X(_0720_));
 sky130_fd_sc_hd__and3_1 _5965_ (.A(net382),
    .B(net636),
    .C(net505),
    .X(_2628_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(net3733),
    .A1(net498),
    .S(net637),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _5967_ (.A0(net3034),
    .A1(net490),
    .S(net637),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(net2037),
    .A1(net2033),
    .S(net637),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(net2419),
    .A1(net481),
    .S(net637),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _5970_ (.A0(net3273),
    .A1(net477),
    .S(net637),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(net2238),
    .A1(net473),
    .S(net637),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _5972_ (.A0(net3201),
    .A1(net469),
    .S(net637),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _5973_ (.A0(net2151),
    .A1(net641),
    .S(net637),
    .X(_0728_));
 sky130_fd_sc_hd__nand2_8 _5974_ (.A(net696),
    .B(net504),
    .Y(_2629_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(net498),
    .A1(net3773),
    .S(_2629_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _5976_ (.A0(net492),
    .A1(net3532),
    .S(_2629_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(net488),
    .A1(net2410),
    .S(_2629_),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _5978_ (.A0(net481),
    .A1(net2372),
    .S(_2629_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _5979_ (.A0(net478),
    .A1(net2764),
    .S(_2629_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _5980_ (.A0(net473),
    .A1(net2137),
    .S(_2629_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _5981_ (.A0(net685),
    .A1(net2416),
    .S(_2629_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _5982_ (.A0(net641),
    .A1(net2131),
    .S(_2629_),
    .X(_0736_));
 sky130_fd_sc_hd__and3_4 _5983_ (.A(net387),
    .B(net380),
    .C(net672),
    .X(_2630_));
 sky130_fd_sc_hd__mux2_1 _5984_ (.A0(net3709),
    .A1(net498),
    .S(_2630_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _5985_ (.A0(net3544),
    .A1(net492),
    .S(_2630_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _5986_ (.A0(net2445),
    .A1(net488),
    .S(_2630_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _5987_ (.A0(net2402),
    .A1(net481),
    .S(_2630_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _5988_ (.A0(net3262),
    .A1(net477),
    .S(_2630_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _5989_ (.A0(net2302),
    .A1(net473),
    .S(_2630_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _5990_ (.A0(net2539),
    .A1(net685),
    .S(_2630_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _5991_ (.A0(net2901),
    .A1(net466),
    .S(_2630_),
    .X(_0744_));
 sky130_fd_sc_hd__and4_4 _5992_ (.A(net660),
    .B(net646),
    .C(net380),
    .D(net504),
    .X(_2631_));
 sky130_fd_sc_hd__mux2_1 _5993_ (.A0(net3713),
    .A1(net498),
    .S(net661),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _5994_ (.A0(net2383),
    .A1(net667),
    .S(net661),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _5995_ (.A0(net1994),
    .A1(net2033),
    .S(_2631_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _5996_ (.A0(net2343),
    .A1(net482),
    .S(net661),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _5997_ (.A0(net3271),
    .A1(net477),
    .S(net661),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _5998_ (.A0(net2170),
    .A1(net473),
    .S(net661),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _5999_ (.A0(net3176),
    .A1(net469),
    .S(net661),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _6000_ (.A0(net2202),
    .A1(net641),
    .S(net661),
    .X(_0752_));
 sky130_fd_sc_hd__o21bai_1 _6001_ (.A1(\xfer_state[3] ),
    .A2(\xfer_state[0] ),
    .B1_N(_1437_),
    .Y(_2632_));
 sky130_fd_sc_hd__a32o_1 _6002_ (.A1(_0823_),
    .A2(\xfer_state[0] ),
    .A3(serial_xfer),
    .B1(_2632_),
    .B2(net3877),
    .X(_0753_));
 sky130_fd_sc_hd__o31ai_4 _6003_ (.A1(\xfer_state[3] ),
    .A2(net527),
    .A3(net526),
    .B1(_1447_),
    .Y(_2633_));
 sky130_fd_sc_hd__a211o_1 _6004_ (.A1(net527),
    .A2(_1443_),
    .B1(\xfer_state[3] ),
    .C1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__nor2_1 _6005_ (.A(\xfer_count[0] ),
    .B(_2633_),
    .Y(_2635_));
 sky130_fd_sc_hd__and2_1 _6006_ (.A(_2633_),
    .B(\xfer_count[0] ),
    .X(_2636_));
 sky130_fd_sc_hd__o311a_1 _6007_ (.A1(\xfer_state[3] ),
    .A2(net527),
    .A3(net526),
    .B1(\xfer_count[0] ),
    .C1(_1447_),
    .X(_2637_));
 sky130_fd_sc_hd__o21a_1 _6008_ (.A1(_2635_),
    .A2(_2636_),
    .B1(_2634_),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _6009_ (.A(\xfer_state[3] ),
    .B(net527),
    .Y(_2638_));
 sky130_fd_sc_hd__nand2_1 _6010_ (.A(\xfer_count[1] ),
    .B(\xfer_count[0] ),
    .Y(_2639_));
 sky130_fd_sc_hd__o22a_1 _6011_ (.A1(\xfer_count[1] ),
    .A2(\xfer_count[0] ),
    .B1(\xfer_state[3] ),
    .B2(net527),
    .X(_2640_));
 sky130_fd_sc_hd__a32o_1 _6012_ (.A1(_1447_),
    .A2(_2639_),
    .A3(_2640_),
    .B1(_2633_),
    .B2(net3889),
    .X(_0755_));
 sky130_fd_sc_hd__nand3_1 _6013_ (.A(\xfer_count[1] ),
    .B(\xfer_count[2] ),
    .C(_2637_),
    .Y(_2641_));
 sky130_fd_sc_hd__a21o_1 _6014_ (.A1(\xfer_count[1] ),
    .A2(_2637_),
    .B1(\xfer_count[2] ),
    .X(_2642_));
 sky130_fd_sc_hd__and3_1 _6015_ (.A(_2634_),
    .B(_2641_),
    .C(_2642_),
    .X(_0756_));
 sky130_fd_sc_hd__a31o_1 _6016_ (.A1(\xfer_count[1] ),
    .A2(\xfer_count[2] ),
    .A3(_2637_),
    .B1(\xfer_count[3] ),
    .X(_2643_));
 sky130_fd_sc_hd__nand4_1 _6017_ (.A(\xfer_count[1] ),
    .B(\xfer_count[2] ),
    .C(\xfer_count[3] ),
    .D(_2637_),
    .Y(_2644_));
 sky130_fd_sc_hd__and3_1 _6018_ (.A(_2634_),
    .B(_2643_),
    .C(_2644_),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_8 _6019_ (.A(net526),
    .B(\xfer_state[0] ),
    .Y(_2645_));
 sky130_fd_sc_hd__mux2_1 _6020_ (.A0(net526),
    .A1(_2645_),
    .S(net3901),
    .X(_0758_));
 sky130_fd_sc_hd__and2b_4 _6021_ (.A_N(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2646_));
 sky130_fd_sc_hd__and2b_4 _6022_ (.A_N(\pad_count_1[0] ),
    .B(\pad_count_1[1] ),
    .X(_2647_));
 sky130_fd_sc_hd__nor2_4 _6023_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .Y(_2648_));
 sky130_fd_sc_hd__and2_4 _6024_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .X(_2649_));
 sky130_fd_sc_hd__o21ai_1 _6025_ (.A1(net447),
    .A2(net446),
    .B1(net526),
    .Y(_2650_));
 sky130_fd_sc_hd__o31a_1 _6026_ (.A1(net526),
    .A2(\xfer_state[0] ),
    .A3(\pad_count_1[1] ),
    .B1(_2650_),
    .X(_0759_));
 sky130_fd_sc_hd__o21a_1 _6027_ (.A1(\pad_count_1[1] ),
    .A2(\pad_count_1[0] ),
    .B1(net522),
    .X(_2651_));
 sky130_fd_sc_hd__nor3_1 _6028_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .C(net522),
    .Y(_2652_));
 sky130_fd_sc_hd__o21a_1 _6029_ (.A1(_2651_),
    .A2(_2652_),
    .B1(net526),
    .X(_2653_));
 sky130_fd_sc_hd__a21o_1 _6030_ (.A1(net522),
    .A2(_2645_),
    .B1(_2653_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_4 _6031_ (.A(net520),
    .B(net444),
    .Y(_2654_));
 sky130_fd_sc_hd__nor2_8 _6032_ (.A(net522),
    .B(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__o221a_1 _6033_ (.A1(net520),
    .A2(_2652_),
    .B1(net522),
    .B2(_2654_),
    .C1(net526),
    .X(_2656_));
 sky130_fd_sc_hd__a21o_1 _6034_ (.A1(net520),
    .A2(_2645_),
    .B1(_2656_),
    .X(_0761_));
 sky130_fd_sc_hd__nor2_8 _6035_ (.A(net520),
    .B(net522),
    .Y(_2657_));
 sky130_fd_sc_hd__nand3_4 _6036_ (.A(net444),
    .B(net442),
    .C(net510),
    .Y(_2658_));
 sky130_fd_sc_hd__a21o_1 _6037_ (.A1(_2658_),
    .A2(net526),
    .B1(_2645_),
    .X(_2659_));
 sky130_fd_sc_hd__o211a_1 _6038_ (.A1(net526),
    .A2(\xfer_state[0] ),
    .B1(net444),
    .C1(net442),
    .X(_2660_));
 sky130_fd_sc_hd__o21ai_1 _6039_ (.A1(net510),
    .A2(_2660_),
    .B1(_2659_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor3_1 _6040_ (.A(\pad_count_2[0] ),
    .B(net526),
    .C(\xfer_state[0] ),
    .Y(_2661_));
 sky130_fd_sc_hd__a21oi_1 _6041_ (.A1(\pad_count_2[0] ),
    .A2(net526),
    .B1(_2661_),
    .Y(_0763_));
 sky130_fd_sc_hd__and2_4 _6042_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2662_));
 sky130_fd_sc_hd__nor2_8 _6043_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .Y(_2663_));
 sky130_fd_sc_hd__and2b_4 _6044_ (.A_N(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .X(_2664_));
 sky130_fd_sc_hd__o21ai_1 _6045_ (.A1(_2662_),
    .A2(net441),
    .B1(net526),
    .Y(_2665_));
 sky130_fd_sc_hd__o31a_1 _6046_ (.A1(\pad_count_2[1] ),
    .A2(net526),
    .A3(\xfer_state[0] ),
    .B1(_2665_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(net515),
    .B(_2662_),
    .Y(_2666_));
 sky130_fd_sc_hd__a21o_1 _6048_ (.A1(\pad_count_2[1] ),
    .A2(\pad_count_2[0] ),
    .B1(net515),
    .X(_2667_));
 sky130_fd_sc_hd__a32o_1 _6049_ (.A1(_2666_),
    .A2(_2667_),
    .A3(net526),
    .B1(_2645_),
    .B2(net515),
    .X(_0765_));
 sky130_fd_sc_hd__nand4_4 _6050_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .C(net514),
    .D(net515),
    .Y(_2668_));
 sky130_fd_sc_hd__nand4_1 _6051_ (.A(net514),
    .B(net515),
    .C(net526),
    .D(_2662_),
    .Y(_2669_));
 sky130_fd_sc_hd__a31o_1 _6052_ (.A1(\pad_count_2[1] ),
    .A2(\pad_count_2[0] ),
    .A3(net515),
    .B1(net514),
    .X(_2670_));
 sky130_fd_sc_hd__a32o_1 _6053_ (.A1(_2670_),
    .A2(net526),
    .A3(_2668_),
    .B1(_2645_),
    .B2(net514),
    .X(_0766_));
 sky130_fd_sc_hd__a211o_1 _6054_ (.A1(_2668_),
    .A2(net526),
    .B1(\pad_count_2[4] ),
    .C1(_2645_),
    .X(_2671_));
 sky130_fd_sc_hd__a21bo_1 _6055_ (.A1(net3900),
    .A2(_2669_),
    .B1_N(_2671_),
    .X(_0767_));
 sky130_fd_sc_hd__and2b_4 _6056_ (.A_N(\pad_count_2[5] ),
    .B(\pad_count_2[4] ),
    .X(_2672_));
 sky130_fd_sc_hd__and3_4 _6057_ (.A(\pad_count_2[1] ),
    .B(\pad_count_2[0] ),
    .C(net439),
    .X(_2673_));
 sky130_fd_sc_hd__and3_4 _6058_ (.A(net514),
    .B(net515),
    .C(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__a211o_1 _6059_ (.A1(_2668_),
    .A2(\pad_count_2[5] ),
    .B1(_1439_),
    .C1(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__a22o_1 _6060_ (.A1(net3897),
    .A2(_2645_),
    .B1(_2675_),
    .B2(net526),
    .X(_0768_));
 sky130_fd_sc_hd__a211o_1 _6061_ (.A1(\xfer_count[1] ),
    .A2(\xfer_count[0] ),
    .B1(\xfer_count[2] ),
    .C1(\xfer_count[3] ),
    .X(_2676_));
 sky130_fd_sc_hd__a22o_1 _6062_ (.A1(_2638_),
    .A2(_2645_),
    .B1(_2676_),
    .B2(\xfer_state[3] ),
    .X(_2677_));
 sky130_fd_sc_hd__a211o_1 _6063_ (.A1(\xfer_state[3] ),
    .A2(_2676_),
    .B1(net513),
    .C1(net301),
    .X(_2678_));
 sky130_fd_sc_hd__a21bo_1 _6064_ (.A1(net3853),
    .A2(_2677_),
    .B1_N(_2678_),
    .X(_0769_));
 sky130_fd_sc_hd__nor3_1 _6065_ (.A(\xfer_count[2] ),
    .B(\xfer_count[3] ),
    .C(_0823_),
    .Y(_2679_));
 sky130_fd_sc_hd__a32o_1 _6066_ (.A1(_0822_),
    .A2(\xfer_count[0] ),
    .A3(_2679_),
    .B1(_2677_),
    .B2(net3869),
    .X(_0770_));
 sky130_fd_sc_hd__and2_4 _6067_ (.A(_0824_),
    .B(\xfer_state[2] ),
    .X(_2680_));
 sky130_fd_sc_hd__a21oi_4 _6068_ (.A1(net527),
    .A2(net301),
    .B1(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__a21o_1 _6069_ (.A1(net528),
    .A2(net301),
    .B1(_2680_),
    .X(_2682_));
 sky130_fd_sc_hd__and4bb_4 _6070_ (.A_N(net516),
    .B_N(net523),
    .C(net444),
    .D(net521),
    .X(_2683_));
 sky130_fd_sc_hd__and3b_1 _6071_ (.A_N(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .C(net442),
    .X(_2684_));
 sky130_fd_sc_hd__and3_4 _6072_ (.A(net518),
    .B(_2646_),
    .C(net443),
    .X(_2685_));
 sky130_fd_sc_hd__and3_4 _6073_ (.A(net520),
    .B(net522),
    .C(net447),
    .X(_2686_));
 sky130_fd_sc_hd__and3b_4 _6074_ (.A_N(\pad_count_1[0] ),
    .B(net442),
    .C(\pad_count_1[1] ),
    .X(_2687_));
 sky130_fd_sc_hd__and3_4 _6075_ (.A(net517),
    .B(net446),
    .C(net442),
    .X(_2688_));
 sky130_fd_sc_hd__a32o_1 _6076_ (.A1(\gpio_configure[29][0] ),
    .A2(net518),
    .A3(net423),
    .B1(_2688_),
    .B2(\gpio_configure[18][0] ),
    .X(_2689_));
 sky130_fd_sc_hd__a221o_1 _6077_ (.A1(\gpio_configure[8][0] ),
    .A2(_2683_),
    .B1(_2685_),
    .B2(\gpio_configure[17][0] ),
    .C1(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__and2b_4 _6078_ (.A_N(net520),
    .B(net522),
    .X(_2691_));
 sky130_fd_sc_hd__and4bb_4 _6079_ (.A_N(\pad_count_1[0] ),
    .B_N(net520),
    .C(net522),
    .D(\pad_count_1[1] ),
    .X(_2692_));
 sky130_fd_sc_hd__and3_4 _6080_ (.A(net519),
    .B(net446),
    .C(net438),
    .X(_2693_));
 sky130_fd_sc_hd__and4bb_4 _6081_ (.A_N(\pad_count_1[1] ),
    .B_N(net520),
    .C(net522),
    .D(\pad_count_1[0] ),
    .X(_2694_));
 sky130_fd_sc_hd__and3_4 _6082_ (.A(net447),
    .B(net438),
    .C(net510),
    .X(_2695_));
 sky130_fd_sc_hd__a32o_1 _6083_ (.A1(\gpio_configure[22][0] ),
    .A2(net519),
    .A3(_2692_),
    .B1(_2695_),
    .B2(\gpio_configure[5][0] ),
    .X(_2696_));
 sky130_fd_sc_hd__and4b_4 _6084_ (.A_N(net522),
    .B(net520),
    .C(\pad_count_1[0] ),
    .D(\pad_count_1[1] ),
    .X(_2697_));
 sky130_fd_sc_hd__and4b_4 _6085_ (.A_N(net523),
    .B(_2649_),
    .C(net516),
    .D(net521),
    .X(_2698_));
 sky130_fd_sc_hd__and3_2 _6086_ (.A(\pad_count_1[1] ),
    .B(\pad_count_1[0] ),
    .C(net437),
    .X(_2699_));
 sky130_fd_sc_hd__and3_4 _6087_ (.A(net518),
    .B(_2649_),
    .C(net437),
    .X(_2700_));
 sky130_fd_sc_hd__a221o_1 _6088_ (.A1(\gpio_configure[27][0] ),
    .A2(_2698_),
    .B1(_2700_),
    .B2(\gpio_configure[23][0] ),
    .C1(_2696_),
    .X(_2701_));
 sky130_fd_sc_hd__and3_4 _6089_ (.A(net520),
    .B(net522),
    .C(net444),
    .X(_2702_));
 sky130_fd_sc_hd__and4_4 _6090_ (.A(net520),
    .B(net523),
    .C(net444),
    .D(net510),
    .X(_2703_));
 sky130_fd_sc_hd__and3_4 _6091_ (.A(net521),
    .B(net523),
    .C(_2649_),
    .X(_2704_));
 sky130_fd_sc_hd__and4_4 _6092_ (.A(net517),
    .B(net520),
    .C(net523),
    .D(_2649_),
    .X(_2705_));
 sky130_fd_sc_hd__and4bb_4 _6093_ (.A_N(\pad_count_1[0] ),
    .B_N(net522),
    .C(net520),
    .D(\pad_count_1[1] ),
    .X(_2706_));
 sky130_fd_sc_hd__and4_4 _6094_ (.A(net519),
    .B(net521),
    .C(net523),
    .D(net444),
    .X(_2707_));
 sky130_fd_sc_hd__a32o_1 _6095_ (.A1(\gpio_configure[26][0] ),
    .A2(net518),
    .A3(net436),
    .B1(_2707_),
    .B2(\gpio_configure[28][0] ),
    .X(_2708_));
 sky130_fd_sc_hd__a221o_1 _6096_ (.A1(\gpio_configure[12][0] ),
    .A2(_2703_),
    .B1(_2705_),
    .B2(\gpio_configure[31][0] ),
    .C1(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__and3_4 _6097_ (.A(net518),
    .B(net445),
    .C(net437),
    .X(_2710_));
 sky130_fd_sc_hd__a32o_1 _6098_ (.A1(\gpio_configure[16][0] ),
    .A2(net445),
    .A3(net443),
    .B1(_2710_),
    .B2(\gpio_configure[20][0] ),
    .X(_2711_));
 sky130_fd_sc_hd__and4bb_4 _6099_ (.A_N(net516),
    .B_N(net522),
    .C(net447),
    .D(net520),
    .X(_2712_));
 sky130_fd_sc_hd__and4b_4 _6100_ (.A_N(net522),
    .B(net444),
    .C(net516),
    .D(net520),
    .X(_2713_));
 sky130_fd_sc_hd__a221o_1 _6101_ (.A1(\gpio_configure[9][0] ),
    .A2(_2712_),
    .B1(_2713_),
    .B2(\gpio_configure[24][0] ),
    .C1(_2711_),
    .X(_2714_));
 sky130_fd_sc_hd__nor4_1 _6102_ (.A(_2690_),
    .B(_2701_),
    .C(_2709_),
    .D(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__a32o_1 _6103_ (.A1(\gpio_configure[7][0] ),
    .A2(_2649_),
    .A3(net437),
    .B1(net436),
    .B2(\gpio_configure[10][0] ),
    .X(_2716_));
 sky130_fd_sc_hd__a221o_1 _6104_ (.A1(\gpio_configure[6][0] ),
    .A2(_2692_),
    .B1(_2704_),
    .B2(\gpio_configure[15][0] ),
    .C1(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__a32o_1 _6105_ (.A1(\gpio_configure[3][0] ),
    .A2(_2649_),
    .A3(net442),
    .B1(_2684_),
    .B2(\gpio_configure[1][0] ),
    .X(_2718_));
 sky130_fd_sc_hd__and3_4 _6106_ (.A(net520),
    .B(net522),
    .C(net446),
    .X(_2719_));
 sky130_fd_sc_hd__a32o_1 _6107_ (.A1(\gpio_configure[2][0] ),
    .A2(net446),
    .A3(net442),
    .B1(net422),
    .B2(\gpio_configure[14][0] ),
    .X(_2720_));
 sky130_fd_sc_hd__o31a_1 _6108_ (.A1(_2717_),
    .A2(_2718_),
    .A3(_2720_),
    .B1(net510),
    .X(_2721_));
 sky130_fd_sc_hd__and4_1 _6109_ (.A(net521),
    .B(net523),
    .C(net447),
    .D(net511),
    .X(_2722_));
 sky130_fd_sc_hd__and3_4 _6110_ (.A(net518),
    .B(_2649_),
    .C(net443),
    .X(_2723_));
 sky130_fd_sc_hd__and4bb_4 _6111_ (.A_N(net517),
    .B_N(net522),
    .C(_2649_),
    .D(net520),
    .X(_2724_));
 sky130_fd_sc_hd__and4b_4 _6112_ (.A_N(net523),
    .B(net447),
    .C(net517),
    .D(net521),
    .X(_2725_));
 sky130_fd_sc_hd__a32o_1 _6113_ (.A1(\gpio_configure[11][0] ),
    .A2(net511),
    .A3(_2697_),
    .B1(_2725_),
    .B2(\gpio_configure[25][0] ),
    .X(_2726_));
 sky130_fd_sc_hd__a221o_1 _6114_ (.A1(\gpio_configure[13][0] ),
    .A2(_2722_),
    .B1(_2723_),
    .B2(\gpio_configure[19][0] ),
    .C1(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__a32o_1 _6115_ (.A1(\gpio_configure[21][0] ),
    .A2(net447),
    .A3(net437),
    .B1(net422),
    .B2(\gpio_configure[30][0] ),
    .X(_2728_));
 sky130_fd_sc_hd__and3_4 _6116_ (.A(net438),
    .B(net512),
    .C(net444),
    .X(_2729_));
 sky130_fd_sc_hd__a32o_1 _6117_ (.A1(net512),
    .A2(net445),
    .A3(net443),
    .B1(_2729_),
    .B2(\gpio_configure[4][0] ),
    .X(_2730_));
 sky130_fd_sc_hd__a2111oi_1 _6118_ (.A1(net518),
    .A2(_2728_),
    .B1(_2730_),
    .C1(_2727_),
    .D1(_2721_),
    .Y(_2731_));
 sky130_fd_sc_hd__and4_4 _6119_ (.A(net520),
    .B(net523),
    .C(_2649_),
    .D(net510),
    .X(_2732_));
 sky130_fd_sc_hd__and3_4 _6120_ (.A(_2649_),
    .B(net437),
    .C(net510),
    .X(_2733_));
 sky130_fd_sc_hd__and3_4 _6121_ (.A(_2649_),
    .B(net442),
    .C(net510),
    .X(_2734_));
 sky130_fd_sc_hd__nand2_4 _6122_ (.A(net350),
    .B(net349),
    .Y(_2735_));
 sky130_fd_sc_hd__o211a_1 _6123_ (.A1(\gpio_configure[0][0] ),
    .A2(_2658_),
    .B1(net513),
    .C1(\xfer_state[2] ),
    .X(_2736_));
 sky130_fd_sc_hd__a22o_1 _6124_ (.A1(net3842),
    .A2(net353),
    .B1(_2735_),
    .B2(_2736_),
    .X(_0771_));
 sky130_fd_sc_hd__a32o_1 _6125_ (.A1(\gpio_configure[23][1] ),
    .A2(net519),
    .A3(_2699_),
    .B1(_2712_),
    .B2(\gpio_configure[9][1] ),
    .X(_2737_));
 sky130_fd_sc_hd__a221o_1 _6126_ (.A1(\gpio_configure[31][1] ),
    .A2(_2705_),
    .B1(_2725_),
    .B2(\gpio_configure[25][1] ),
    .C1(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__a32o_1 _6127_ (.A1(\gpio_configure[27][1] ),
    .A2(net519),
    .A3(_2697_),
    .B1(_2733_),
    .B2(\gpio_configure[7][1] ),
    .X(_2739_));
 sky130_fd_sc_hd__a221o_1 _6128_ (.A1(\gpio_configure[18][1] ),
    .A2(_2688_),
    .B1(_2734_),
    .B2(\gpio_configure[3][1] ),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__a32o_1 _6129_ (.A1(\gpio_configure[21][1] ),
    .A2(net447),
    .A3(net438),
    .B1(net422),
    .B2(\gpio_configure[30][1] ),
    .X(_2741_));
 sky130_fd_sc_hd__a221o_1 _6130_ (.A1(\gpio_configure[24][1] ),
    .A2(_2655_),
    .B1(net436),
    .B2(\gpio_configure[26][1] ),
    .C1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__o211a_1 _6131_ (.A1(\gpio_configure[16][1] ),
    .A2(net510),
    .B1(net444),
    .C1(net442),
    .X(_2743_));
 sky130_fd_sc_hd__a221o_1 _6132_ (.A1(\gpio_configure[5][1] ),
    .A2(_2695_),
    .B1(_2707_),
    .B2(\gpio_configure[28][1] ),
    .C1(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__a2111o_4 _6133_ (.A1(net519),
    .A2(_2742_),
    .B1(_2744_),
    .C1(_2738_),
    .D1(_2740_),
    .X(_2745_));
 sky130_fd_sc_hd__a22o_1 _6134_ (.A1(\gpio_configure[10][1] ),
    .A2(net436),
    .B1(net422),
    .B2(\gpio_configure[14][1] ),
    .X(_2746_));
 sky130_fd_sc_hd__a221o_1 _6135_ (.A1(\gpio_configure[8][1] ),
    .A2(_2655_),
    .B1(net423),
    .B2(\gpio_configure[13][1] ),
    .C1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__and3_1 _6136_ (.A(\gpio_configure[2][1] ),
    .B(net446),
    .C(net442),
    .X(_2748_));
 sky130_fd_sc_hd__a32o_1 _6137_ (.A1(\gpio_configure[1][1] ),
    .A2(net447),
    .A3(net442),
    .B1(_2692_),
    .B2(\gpio_configure[6][1] ),
    .X(_2749_));
 sky130_fd_sc_hd__a2111o_1 _6138_ (.A1(\gpio_configure[11][1] ),
    .A2(_2697_),
    .B1(_2748_),
    .C1(_2749_),
    .D1(_2747_),
    .X(_2750_));
 sky130_fd_sc_hd__a32o_1 _6139_ (.A1(\gpio_configure[15][1] ),
    .A2(_2704_),
    .A3(net512),
    .B1(\gpio_configure[4][1] ),
    .B2(_2729_),
    .X(_2751_));
 sky130_fd_sc_hd__a221o_1 _6140_ (.A1(\gpio_configure[17][1] ),
    .A2(_2685_),
    .B1(_2710_),
    .B2(\gpio_configure[20][1] ),
    .C1(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__a32o_1 _6141_ (.A1(\gpio_configure[29][1] ),
    .A2(net519),
    .A3(net423),
    .B1(_2723_),
    .B2(\gpio_configure[19][1] ),
    .X(_2753_));
 sky130_fd_sc_hd__a221o_1 _6142_ (.A1(\gpio_configure[22][1] ),
    .A2(_2693_),
    .B1(_2703_),
    .B2(\gpio_configure[12][1] ),
    .C1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__a211o_2 _6143_ (.A1(net512),
    .A2(_2750_),
    .B1(_2752_),
    .C1(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__and3_1 _6144_ (.A(net447),
    .B(net443),
    .C(net511),
    .X(_2756_));
 sky130_fd_sc_hd__o221ai_4 _6145_ (.A1(_2658_),
    .A2(\gpio_configure[0][1] ),
    .B1(_2755_),
    .B2(_2745_),
    .C1(net513),
    .Y(_2757_));
 sky130_fd_sc_hd__o2bb2a_1 _6146_ (.A1_N(net528),
    .A2_N(\serial_data_staging_1[0] ),
    .B1(_1446_),
    .B2(_2680_),
    .X(_2758_));
 sky130_fd_sc_hd__o2bb2a_1 _6147_ (.A1_N(_2758_),
    .A2_N(_2757_),
    .B1(_2682_),
    .B2(net3843),
    .X(_0772_));
 sky130_fd_sc_hd__a32o_1 _6148_ (.A1(\gpio_configure[26][2] ),
    .A2(net517),
    .A3(net436),
    .B1(_2729_),
    .B2(\gpio_configure[4][2] ),
    .X(_2759_));
 sky130_fd_sc_hd__a221o_1 _6149_ (.A1(\gpio_configure[31][2] ),
    .A2(_2705_),
    .B1(_2733_),
    .B2(\gpio_configure[7][2] ),
    .C1(_2759_),
    .X(_2760_));
 sky130_fd_sc_hd__a32o_4 _6150_ (.A1(\gpio_configure[29][2] ),
    .A2(\pad_count_1[4] ),
    .A3(net423),
    .B1(_2700_),
    .B2(\gpio_configure[23][2] ),
    .X(_2761_));
 sky130_fd_sc_hd__o211a_1 _6151_ (.A1(\gpio_configure[16][2] ),
    .A2(net510),
    .B1(net444),
    .C1(net442),
    .X(_2762_));
 sky130_fd_sc_hd__a2111o_1 _6152_ (.A1(\gpio_configure[25][2] ),
    .A2(_2725_),
    .B1(_2762_),
    .C1(_2761_),
    .D1(_2760_),
    .X(_2763_));
 sky130_fd_sc_hd__a32o_1 _6153_ (.A1(\gpio_configure[22][2] ),
    .A2(net517),
    .A3(_2692_),
    .B1(_2732_),
    .B2(\gpio_configure[15][2] ),
    .X(_2764_));
 sky130_fd_sc_hd__a221oi_2 _6154_ (.A1(\gpio_configure[9][2] ),
    .A2(_2712_),
    .B1(_2723_),
    .B2(\gpio_configure[19][2] ),
    .C1(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__a32o_1 _6155_ (.A1(\gpio_configure[5][2] ),
    .A2(net512),
    .A3(_2694_),
    .B1(_2688_),
    .B2(\gpio_configure[18][2] ),
    .X(_2766_));
 sky130_fd_sc_hd__a221oi_1 _6156_ (.A1(\gpio_configure[11][2] ),
    .A2(_2724_),
    .B1(_2734_),
    .B2(\gpio_configure[3][2] ),
    .C1(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__nand3b_1 _6157_ (.A_N(_2763_),
    .B(_2765_),
    .C(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__a22o_1 _6158_ (.A1(\gpio_configure[12][2] ),
    .A2(_2702_),
    .B1(net422),
    .B2(\gpio_configure[14][2] ),
    .X(_2769_));
 sky130_fd_sc_hd__a41o_1 _6159_ (.A1(\gpio_configure[13][2] ),
    .A2(net521),
    .A3(net522),
    .A4(net447),
    .B1(net517),
    .X(_2770_));
 sky130_fd_sc_hd__a221o_1 _6160_ (.A1(\gpio_configure[2][2] ),
    .A2(_2687_),
    .B1(_2692_),
    .B2(\gpio_configure[6][2] ),
    .C1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__a211o_1 _6161_ (.A1(\gpio_configure[10][2] ),
    .A2(net436),
    .B1(_2769_),
    .C1(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__a41o_1 _6162_ (.A1(\gpio_configure[30][2] ),
    .A2(net521),
    .A3(net523),
    .A4(net446),
    .B1(net511),
    .X(_2773_));
 sky130_fd_sc_hd__a221o_2 _6163_ (.A1(\gpio_configure[21][2] ),
    .A2(_2694_),
    .B1(_2702_),
    .B2(\gpio_configure[28][2] ),
    .C1(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__a32o_1 _6164_ (.A1(net510),
    .A2(_2684_),
    .A3(\gpio_configure[1][2] ),
    .B1(_2710_),
    .B2(\gpio_configure[20][2] ),
    .X(_2775_));
 sky130_fd_sc_hd__a32o_1 _6165_ (.A1(\gpio_configure[27][2] ),
    .A2(net516),
    .A3(_2697_),
    .B1(_2713_),
    .B2(\gpio_configure[24][2] ),
    .X(_2776_));
 sky130_fd_sc_hd__a221o_1 _6166_ (.A1(\gpio_configure[8][2] ),
    .A2(_2683_),
    .B1(_2685_),
    .B2(\gpio_configure[17][2] ),
    .C1(_2776_),
    .X(_2777_));
 sky130_fd_sc_hd__a211o_1 _6167_ (.A1(_2772_),
    .A2(_2774_),
    .B1(_2775_),
    .C1(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__o221a_1 _6168_ (.A1(_2658_),
    .A2(\gpio_configure[0][2] ),
    .B1(_2778_),
    .B2(_2768_),
    .C1(net513),
    .X(_2779_));
 sky130_fd_sc_hd__a211o_1 _6169_ (.A1(net528),
    .A2(net3843),
    .B1(net353),
    .C1(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__o31a_1 _6170_ (.A1(net3852),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_2780_),
    .X(_0773_));
 sky130_fd_sc_hd__a32o_1 _6171_ (.A1(\gpio_configure[2][3] ),
    .A2(net446),
    .A3(net443),
    .B1(_2692_),
    .B2(\gpio_configure[6][3] ),
    .X(_2781_));
 sky130_fd_sc_hd__a221o_1 _6172_ (.A1(\gpio_configure[10][3] ),
    .A2(net436),
    .B1(net422),
    .B2(\gpio_configure[14][3] ),
    .C1(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__o211a_1 _6173_ (.A1(\gpio_configure[16][3] ),
    .A2(net511),
    .B1(net445),
    .C1(net443),
    .X(_2783_));
 sky130_fd_sc_hd__a31o_1 _6174_ (.A1(\gpio_configure[12][3] ),
    .A2(_2702_),
    .A3(net511),
    .B1(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__a221o_1 _6175_ (.A1(\gpio_configure[5][3] ),
    .A2(_2695_),
    .B1(_2712_),
    .B2(\gpio_configure[9][3] ),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a32o_1 _6176_ (.A1(\gpio_configure[11][3] ),
    .A2(net511),
    .A3(_2697_),
    .B1(_2683_),
    .B2(\gpio_configure[8][3] ),
    .X(_2786_));
 sky130_fd_sc_hd__a221o_1 _6177_ (.A1(\gpio_configure[4][3] ),
    .A2(_2729_),
    .B1(_2732_),
    .B2(\gpio_configure[15][3] ),
    .C1(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__a211o_4 _6178_ (.A1(net512),
    .A2(_2782_),
    .B1(_2785_),
    .C1(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__a32o_1 _6179_ (.A1(\gpio_configure[21][3] ),
    .A2(net447),
    .A3(net438),
    .B1(net423),
    .B2(\gpio_configure[29][3] ),
    .X(_2789_));
 sky130_fd_sc_hd__a32o_1 _6180_ (.A1(\gpio_configure[23][3] ),
    .A2(_2649_),
    .A3(net438),
    .B1(net422),
    .B2(\gpio_configure[30][3] ),
    .X(_2790_));
 sky130_fd_sc_hd__a211o_1 _6181_ (.A1(\gpio_configure[31][3] ),
    .A2(_2704_),
    .B1(_2789_),
    .C1(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__a32o_1 _6182_ (.A1(\gpio_configure[18][3] ),
    .A2(net519),
    .A3(_2687_),
    .B1(_2733_),
    .B2(\gpio_configure[7][3] ),
    .X(_2792_));
 sky130_fd_sc_hd__a221o_1 _6183_ (.A1(\gpio_configure[13][3] ),
    .A2(_2722_),
    .B1(_2723_),
    .B2(\gpio_configure[19][3] ),
    .C1(_2792_),
    .X(_2793_));
 sky130_fd_sc_hd__a221o_1 _6184_ (.A1(\gpio_configure[17][3] ),
    .A2(_2685_),
    .B1(_2756_),
    .B2(\gpio_configure[1][3] ),
    .C1(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__a32o_1 _6185_ (.A1(\gpio_configure[22][3] ),
    .A2(net519),
    .A3(_2692_),
    .B1(_2707_),
    .B2(\gpio_configure[28][3] ),
    .X(_2795_));
 sky130_fd_sc_hd__a221o_1 _6186_ (.A1(\gpio_configure[27][3] ),
    .A2(_2698_),
    .B1(_2725_),
    .B2(\gpio_configure[25][3] ),
    .C1(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__a32o_1 _6187_ (.A1(\gpio_configure[26][3] ),
    .A2(net519),
    .A3(_2706_),
    .B1(_2713_),
    .B2(\gpio_configure[24][3] ),
    .X(_2797_));
 sky130_fd_sc_hd__a221o_1 _6188_ (.A1(\gpio_configure[20][3] ),
    .A2(_2710_),
    .B1(_2734_),
    .B2(\gpio_configure[3][3] ),
    .C1(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__a2111o_4 _6189_ (.A1(_2791_),
    .A2(net519),
    .B1(_2796_),
    .C1(_2794_),
    .D1(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__o221a_1 _6190_ (.A1(\gpio_configure[0][3] ),
    .A2(_2658_),
    .B1(_2788_),
    .B2(_2799_),
    .C1(net513),
    .X(_2800_));
 sky130_fd_sc_hd__a211o_1 _6191_ (.A1(net528),
    .A2(\serial_data_staging_1[2] ),
    .B1(net353),
    .C1(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__o31a_1 _6192_ (.A1(net3831),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_2801_),
    .X(_0774_));
 sky130_fd_sc_hd__a32o_1 _6193_ (.A1(\gpio_configure[26][4] ),
    .A2(net519),
    .A3(_2706_),
    .B1(_2723_),
    .B2(\gpio_configure[19][4] ),
    .X(_2802_));
 sky130_fd_sc_hd__a221o_1 _6194_ (.A1(\gpio_configure[5][4] ),
    .A2(_2695_),
    .B1(_2733_),
    .B2(\gpio_configure[7][4] ),
    .C1(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__a32o_1 _6195_ (.A1(\gpio_configure[27][4] ),
    .A2(net519),
    .A3(_2697_),
    .B1(_2729_),
    .B2(\gpio_configure[4][4] ),
    .X(_2804_));
 sky130_fd_sc_hd__a221o_1 _6196_ (.A1(\gpio_configure[20][4] ),
    .A2(_2710_),
    .B1(_2734_),
    .B2(\gpio_configure[3][4] ),
    .C1(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__o211a_1 _6197_ (.A1(\gpio_configure[16][4] ),
    .A2(net511),
    .B1(net444),
    .C1(net443),
    .X(_2806_));
 sky130_fd_sc_hd__a32o_1 _6198_ (.A1(net511),
    .A2(_2702_),
    .A3(\gpio_configure[12][4] ),
    .B1(_2732_),
    .B2(\gpio_configure[15][4] ),
    .X(_2807_));
 sky130_fd_sc_hd__a2111o_2 _6199_ (.A1(\gpio_configure[25][4] ),
    .A2(_2725_),
    .B1(_2806_),
    .C1(_2807_),
    .D1(_2805_),
    .X(_2808_));
 sky130_fd_sc_hd__a32o_1 _6200_ (.A1(\gpio_configure[23][4] ),
    .A2(_2649_),
    .A3(net437),
    .B1(net423),
    .B2(\gpio_configure[29][4] ),
    .X(_2809_));
 sky130_fd_sc_hd__a32o_1 _6201_ (.A1(\gpio_configure[21][4] ),
    .A2(net447),
    .A3(net438),
    .B1(_2702_),
    .B2(\gpio_configure[28][4] ),
    .X(_2810_));
 sky130_fd_sc_hd__a211o_1 _6202_ (.A1(\gpio_configure[30][4] ),
    .A2(net422),
    .B1(_2809_),
    .C1(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__a32o_1 _6203_ (.A1(\gpio_configure[6][4] ),
    .A2(_2647_),
    .A3(net438),
    .B1(_2697_),
    .B2(\gpio_configure[11][4] ),
    .X(_2812_));
 sky130_fd_sc_hd__a221o_1 _6204_ (.A1(\gpio_configure[10][4] ),
    .A2(_2706_),
    .B1(_2719_),
    .B2(\gpio_configure[14][4] ),
    .C1(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__a32o_1 _6205_ (.A1(\gpio_configure[1][4] ),
    .A2(_2646_),
    .A3(net443),
    .B1(_2655_),
    .B2(\gpio_configure[8][4] ),
    .X(_2814_));
 sky130_fd_sc_hd__a32o_1 _6206_ (.A1(\gpio_configure[2][4] ),
    .A2(_2647_),
    .A3(_2657_),
    .B1(_2686_),
    .B2(\gpio_configure[13][4] ),
    .X(_2815_));
 sky130_fd_sc_hd__o31a_1 _6207_ (.A1(_2813_),
    .A2(_2814_),
    .A3(_2815_),
    .B1(net512),
    .X(_2816_));
 sky130_fd_sc_hd__a32o_1 _6208_ (.A1(\gpio_configure[18][4] ),
    .A2(net518),
    .A3(_2687_),
    .B1(_2713_),
    .B2(\gpio_configure[24][4] ),
    .X(_2817_));
 sky130_fd_sc_hd__a221o_1 _6209_ (.A1(\gpio_configure[22][4] ),
    .A2(_2693_),
    .B1(_2705_),
    .B2(\gpio_configure[31][4] ),
    .C1(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__a221o_1 _6210_ (.A1(\gpio_configure[17][4] ),
    .A2(_2685_),
    .B1(_2712_),
    .B2(\gpio_configure[9][4] ),
    .C1(_2818_),
    .X(_2819_));
 sky130_fd_sc_hd__a211o_1 _6211_ (.A1(net519),
    .A2(_2811_),
    .B1(_2816_),
    .C1(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__nor3_4 _6212_ (.A(_2803_),
    .B(_2808_),
    .C(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__o21ai_1 _6213_ (.A1(\gpio_configure[0][4] ),
    .A2(_2658_),
    .B1(net513),
    .Y(_2822_));
 sky130_fd_sc_hd__a2bb2o_1 _6214_ (.A1_N(_2822_),
    .A2_N(_2821_),
    .B1(\serial_data_staging_1[3] ),
    .B2(net528),
    .X(_2823_));
 sky130_fd_sc_hd__mux2_1 _6215_ (.A0(_2823_),
    .A1(net3823),
    .S(_2681_),
    .X(_0775_));
 sky130_fd_sc_hd__a32o_1 _6216_ (.A1(\gpio_configure[26][5] ),
    .A2(net519),
    .A3(net436),
    .B1(_2710_),
    .B2(\gpio_configure[20][5] ),
    .X(_2824_));
 sky130_fd_sc_hd__a221o_1 _6217_ (.A1(\gpio_configure[22][5] ),
    .A2(_2693_),
    .B1(_2698_),
    .B2(\gpio_configure[27][5] ),
    .C1(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__o211a_1 _6218_ (.A1(\gpio_configure[16][5] ),
    .A2(net510),
    .B1(net444),
    .C1(net442),
    .X(_2826_));
 sky130_fd_sc_hd__a32o_1 _6219_ (.A1(\gpio_configure[29][5] ),
    .A2(net516),
    .A3(net423),
    .B1(_2685_),
    .B2(\gpio_configure[17][5] ),
    .X(_2827_));
 sky130_fd_sc_hd__a2111o_1 _6220_ (.A1(\gpio_configure[8][5] ),
    .A2(_2683_),
    .B1(_2826_),
    .C1(_2827_),
    .D1(_2825_),
    .X(_2828_));
 sky130_fd_sc_hd__a32o_1 _6221_ (.A1(\gpio_configure[5][5] ),
    .A2(net512),
    .A3(_2694_),
    .B1(_2703_),
    .B2(\gpio_configure[12][5] ),
    .X(_2829_));
 sky130_fd_sc_hd__a32o_1 _6222_ (.A1(\gpio_configure[18][5] ),
    .A2(net519),
    .A3(_2687_),
    .B1(_2707_),
    .B2(\gpio_configure[28][5] ),
    .X(_2830_));
 sky130_fd_sc_hd__a221o_1 _6223_ (.A1(\gpio_configure[31][5] ),
    .A2(_2705_),
    .B1(_2725_),
    .B2(\gpio_configure[25][5] ),
    .C1(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__a2111o_2 _6224_ (.A1(\gpio_configure[23][5] ),
    .A2(_2700_),
    .B1(_2828_),
    .C1(_2829_),
    .D1(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__a32o_1 _6225_ (.A1(\gpio_configure[1][5] ),
    .A2(net447),
    .A3(net442),
    .B1(net436),
    .B2(\gpio_configure[10][5] ),
    .X(_2833_));
 sky130_fd_sc_hd__a221o_1 _6226_ (.A1(\gpio_configure[2][5] ),
    .A2(_2687_),
    .B1(net422),
    .B2(\gpio_configure[14][5] ),
    .C1(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__a32o_1 _6227_ (.A1(\gpio_configure[6][5] ),
    .A2(net446),
    .A3(net438),
    .B1(_2697_),
    .B2(\gpio_configure[11][5] ),
    .X(_2835_));
 sky130_fd_sc_hd__a2111o_1 _6228_ (.A1(\gpio_configure[13][5] ),
    .A2(net423),
    .B1(net516),
    .C1(_2835_),
    .D1(_2834_),
    .X(_2836_));
 sky130_fd_sc_hd__a41o_1 _6229_ (.A1(\gpio_configure[30][5] ),
    .A2(net521),
    .A3(net523),
    .A4(net446),
    .B1(net510),
    .X(_2837_));
 sky130_fd_sc_hd__a221o_1 _6230_ (.A1(\gpio_configure[24][5] ),
    .A2(_2655_),
    .B1(_2694_),
    .B2(\gpio_configure[21][5] ),
    .C1(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__a32o_1 _6231_ (.A1(\gpio_configure[15][5] ),
    .A2(_2704_),
    .A3(net512),
    .B1(\gpio_configure[9][5] ),
    .B2(_2712_),
    .X(_2839_));
 sky130_fd_sc_hd__a22o_1 _6232_ (.A1(\gpio_configure[19][5] ),
    .A2(_2723_),
    .B1(_2729_),
    .B2(\gpio_configure[4][5] ),
    .X(_2840_));
 sky130_fd_sc_hd__a221o_1 _6233_ (.A1(\gpio_configure[7][5] ),
    .A2(_2733_),
    .B1(_2734_),
    .B2(\gpio_configure[3][5] ),
    .C1(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__a211o_1 _6234_ (.A1(_2836_),
    .A2(_2838_),
    .B1(_2839_),
    .C1(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__o21a_1 _6235_ (.A1(\gpio_configure[0][5] ),
    .A2(_2658_),
    .B1(net513),
    .X(_2843_));
 sky130_fd_sc_hd__o21a_1 _6236_ (.A1(_2832_),
    .A2(_2842_),
    .B1(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__a211o_1 _6237_ (.A1(net528),
    .A2(net3823),
    .B1(net353),
    .C1(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__o31a_1 _6238_ (.A1(net3844),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_2845_),
    .X(_0776_));
 sky130_fd_sc_hd__a22o_1 _6239_ (.A1(\gpio_configure[11][6] ),
    .A2(_2697_),
    .B1(_2706_),
    .B2(\gpio_configure[10][6] ),
    .X(_2846_));
 sky130_fd_sc_hd__a31o_1 _6240_ (.A1(\gpio_configure[6][6] ),
    .A2(net446),
    .A3(net438),
    .B1(net517),
    .X(_2847_));
 sky130_fd_sc_hd__a32o_1 _6241_ (.A1(\gpio_configure[1][6] ),
    .A2(net447),
    .A3(net442),
    .B1(_2687_),
    .B2(\gpio_configure[2][6] ),
    .X(_2848_));
 sky130_fd_sc_hd__a221o_1 _6242_ (.A1(\gpio_configure[13][6] ),
    .A2(net423),
    .B1(net422),
    .B2(\gpio_configure[14][6] ),
    .C1(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__a2111o_1 _6243_ (.A1(\gpio_configure[12][6] ),
    .A2(_2702_),
    .B1(_2846_),
    .C1(_2847_),
    .D1(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__a41o_1 _6244_ (.A1(\gpio_configure[30][6] ),
    .A2(net521),
    .A3(net523),
    .A4(net446),
    .B1(net511),
    .X(_2851_));
 sky130_fd_sc_hd__a221o_1 _6245_ (.A1(\gpio_configure[24][6] ),
    .A2(_2655_),
    .B1(_2694_),
    .B2(\gpio_configure[21][6] ),
    .C1(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__a32o_1 _6246_ (.A1(\gpio_configure[29][6] ),
    .A2(net516),
    .A3(_2686_),
    .B1(_2698_),
    .B2(\gpio_configure[27][6] ),
    .X(_2853_));
 sky130_fd_sc_hd__a221o_1 _6247_ (.A1(\gpio_configure[4][6] ),
    .A2(_2729_),
    .B1(_2734_),
    .B2(\gpio_configure[3][6] ),
    .C1(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__a32o_1 _6248_ (.A1(\gpio_configure[18][6] ),
    .A2(net517),
    .A3(_2687_),
    .B1(_2733_),
    .B2(\gpio_configure[7][6] ),
    .X(_2855_));
 sky130_fd_sc_hd__a221o_1 _6249_ (.A1(\gpio_configure[17][6] ),
    .A2(_2685_),
    .B1(_2712_),
    .B2(\gpio_configure[9][6] ),
    .C1(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a32o_1 _6250_ (.A1(\gpio_configure[26][6] ),
    .A2(net517),
    .A3(net436),
    .B1(_2710_),
    .B2(\gpio_configure[20][6] ),
    .X(_2857_));
 sky130_fd_sc_hd__a221o_1 _6251_ (.A1(\gpio_configure[8][6] ),
    .A2(_2683_),
    .B1(_2725_),
    .B2(\gpio_configure[25][6] ),
    .C1(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__o211a_1 _6252_ (.A1(\gpio_configure[16][6] ),
    .A2(net512),
    .B1(net444),
    .C1(net443),
    .X(_2859_));
 sky130_fd_sc_hd__a32o_1 _6253_ (.A1(\gpio_configure[22][6] ),
    .A2(net517),
    .A3(_2692_),
    .B1(_2707_),
    .B2(\gpio_configure[28][6] ),
    .X(_2860_));
 sky130_fd_sc_hd__a32o_1 _6254_ (.A1(\gpio_configure[15][6] ),
    .A2(_2704_),
    .A3(net512),
    .B1(\gpio_configure[23][6] ),
    .B2(_2700_),
    .X(_2861_));
 sky130_fd_sc_hd__a221o_1 _6255_ (.A1(\gpio_configure[5][6] ),
    .A2(_2695_),
    .B1(_2723_),
    .B2(\gpio_configure[19][6] ),
    .C1(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__a2111o_1 _6256_ (.A1(\gpio_configure[31][6] ),
    .A2(_2705_),
    .B1(_2859_),
    .C1(_2860_),
    .D1(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__nor4_1 _6257_ (.A(_2854_),
    .B(_2856_),
    .C(_2858_),
    .D(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__a21bo_2 _6258_ (.A1(_2850_),
    .A2(_2852_),
    .B1_N(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__o21a_1 _6259_ (.A1(\gpio_configure[0][6] ),
    .A2(_2658_),
    .B1(_0824_),
    .X(_2866_));
 sky130_fd_sc_hd__a221o_1 _6260_ (.A1(net528),
    .A2(net3844),
    .B1(_2865_),
    .B2(_2866_),
    .C1(net353),
    .X(_2867_));
 sky130_fd_sc_hd__o31a_1 _6261_ (.A1(net3866),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_2867_),
    .X(_0777_));
 sky130_fd_sc_hd__a22o_1 _6262_ (.A1(\gpio_configure[12][7] ),
    .A2(_2702_),
    .B1(_2706_),
    .B2(\gpio_configure[10][7] ),
    .X(_2868_));
 sky130_fd_sc_hd__a31o_1 _6263_ (.A1(\gpio_configure[4][7] ),
    .A2(net444),
    .A3(net438),
    .B1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__a32o_1 _6264_ (.A1(\gpio_configure[1][7] ),
    .A2(net447),
    .A3(net443),
    .B1(_2687_),
    .B2(\gpio_configure[2][7] ),
    .X(_2870_));
 sky130_fd_sc_hd__a221o_1 _6265_ (.A1(\gpio_configure[13][7] ),
    .A2(_2686_),
    .B1(_2692_),
    .B2(\gpio_configure[6][7] ),
    .C1(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__a2111o_1 _6266_ (.A1(\gpio_configure[14][7] ),
    .A2(net422),
    .B1(net519),
    .C1(_2871_),
    .D1(_2869_),
    .X(_2872_));
 sky130_fd_sc_hd__a32o_1 _6267_ (.A1(\gpio_configure[21][7] ),
    .A2(net447),
    .A3(net438),
    .B1(net422),
    .B2(\gpio_configure[30][7] ),
    .X(_2873_));
 sky130_fd_sc_hd__a211o_1 _6268_ (.A1(\gpio_configure[24][7] ),
    .A2(_2655_),
    .B1(_2873_),
    .C1(net512),
    .X(_2874_));
 sky130_fd_sc_hd__a32o_1 _6269_ (.A1(\gpio_configure[31][7] ),
    .A2(net519),
    .A3(_2704_),
    .B1(_2734_),
    .B2(\gpio_configure[3][7] ),
    .X(_2875_));
 sky130_fd_sc_hd__o211a_1 _6270_ (.A1(\gpio_configure[16][7] ),
    .A2(net512),
    .B1(net444),
    .C1(net443),
    .X(_2876_));
 sky130_fd_sc_hd__a32o_1 _6271_ (.A1(\gpio_configure[18][7] ),
    .A2(\pad_count_1[4] ),
    .A3(_2687_),
    .B1(_2733_),
    .B2(\gpio_configure[7][7] ),
    .X(_2877_));
 sky130_fd_sc_hd__a221o_1 _6272_ (.A1(\gpio_configure[9][7] ),
    .A2(_2712_),
    .B1(_2725_),
    .B2(\gpio_configure[25][7] ),
    .C1(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__a2111o_1 _6273_ (.A1(\gpio_configure[22][7] ),
    .A2(_2693_),
    .B1(_2875_),
    .C1(_2876_),
    .D1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a32o_1 _6274_ (.A1(\gpio_configure[29][7] ),
    .A2(net519),
    .A3(net423),
    .B1(_2698_),
    .B2(\gpio_configure[27][7] ),
    .X(_2880_));
 sky130_fd_sc_hd__a221o_1 _6275_ (.A1(\gpio_configure[23][7] ),
    .A2(_2700_),
    .B1(_2707_),
    .B2(\gpio_configure[28][7] ),
    .C1(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__a32o_1 _6276_ (.A1(\gpio_configure[26][7] ),
    .A2(net519),
    .A3(_2706_),
    .B1(_2732_),
    .B2(\gpio_configure[15][7] ),
    .X(_2882_));
 sky130_fd_sc_hd__a221o_1 _6277_ (.A1(\gpio_configure[17][7] ),
    .A2(_2685_),
    .B1(_2710_),
    .B2(\gpio_configure[20][7] ),
    .C1(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__a32o_1 _6278_ (.A1(\gpio_configure[11][7] ),
    .A2(net512),
    .A3(_2697_),
    .B1(_2723_),
    .B2(\gpio_configure[19][7] ),
    .X(_2884_));
 sky130_fd_sc_hd__a221o_1 _6279_ (.A1(\gpio_configure[8][7] ),
    .A2(_2683_),
    .B1(_2695_),
    .B2(\gpio_configure[5][7] ),
    .C1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__nor4_1 _6280_ (.A(_2879_),
    .B(_2881_),
    .C(_2883_),
    .D(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__a21bo_4 _6281_ (.A1(_2872_),
    .A2(_2874_),
    .B1_N(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__o21a_1 _6282_ (.A1(\gpio_configure[0][7] ),
    .A2(_2658_),
    .B1(net513),
    .X(_2888_));
 sky130_fd_sc_hd__a22o_1 _6283_ (.A1(net528),
    .A2(\serial_data_staging_1[6] ),
    .B1(_2887_),
    .B2(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__mux2_1 _6284_ (.A0(_2889_),
    .A1(net3868),
    .S(net353),
    .X(_0778_));
 sky130_fd_sc_hd__a32o_1 _6285_ (.A1(\gpio_configure[4][8] ),
    .A2(net444),
    .A3(net437),
    .B1(net436),
    .B2(\gpio_configure[10][8] ),
    .X(_2890_));
 sky130_fd_sc_hd__a31o_1 _6286_ (.A1(\gpio_configure[6][8] ),
    .A2(net446),
    .A3(net437),
    .B1(net516),
    .X(_2891_));
 sky130_fd_sc_hd__a32o_1 _6287_ (.A1(\gpio_configure[1][8] ),
    .A2(net447),
    .A3(net442),
    .B1(net422),
    .B2(\gpio_configure[14][8] ),
    .X(_2892_));
 sky130_fd_sc_hd__a221o_1 _6288_ (.A1(\gpio_configure[13][8] ),
    .A2(net423),
    .B1(_2687_),
    .B2(\gpio_configure[2][8] ),
    .C1(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__a2111o_1 _6289_ (.A1(\gpio_configure[12][8] ),
    .A2(_2702_),
    .B1(_2890_),
    .C1(_2891_),
    .D1(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a41o_1 _6290_ (.A1(\gpio_configure[30][8] ),
    .A2(net520),
    .A3(net522),
    .A4(net446),
    .B1(net510),
    .X(_2895_));
 sky130_fd_sc_hd__a221o_1 _6291_ (.A1(\gpio_configure[24][8] ),
    .A2(_2655_),
    .B1(_2694_),
    .B2(\gpio_configure[21][8] ),
    .C1(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__a32o_1 _6292_ (.A1(\gpio_configure[22][8] ),
    .A2(net516),
    .A3(_2692_),
    .B1(_2707_),
    .B2(\gpio_configure[28][8] ),
    .X(_2897_));
 sky130_fd_sc_hd__a221o_1 _6293_ (.A1(\gpio_configure[8][8] ),
    .A2(_2683_),
    .B1(_2700_),
    .B2(\gpio_configure[23][8] ),
    .C1(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__a32o_1 _6294_ (.A1(\gpio_configure[7][8] ),
    .A2(_2699_),
    .A3(net510),
    .B1(\gpio_configure[3][8] ),
    .B2(_2734_),
    .X(_2899_));
 sky130_fd_sc_hd__o211a_1 _6295_ (.A1(\gpio_configure[16][8] ),
    .A2(net510),
    .B1(net444),
    .C1(net442),
    .X(_2900_));
 sky130_fd_sc_hd__a2111o_1 _6296_ (.A1(\gpio_configure[31][8] ),
    .A2(_2705_),
    .B1(_2900_),
    .C1(_2899_),
    .D1(_2898_),
    .X(_2901_));
 sky130_fd_sc_hd__a32o_1 _6297_ (.A1(\gpio_configure[26][8] ),
    .A2(net516),
    .A3(net436),
    .B1(_2732_),
    .B2(\gpio_configure[15][8] ),
    .X(_2902_));
 sky130_fd_sc_hd__a221o_1 _6298_ (.A1(\gpio_configure[19][8] ),
    .A2(_2723_),
    .B1(_2725_),
    .B2(\gpio_configure[25][8] ),
    .C1(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__a32o_1 _6299_ (.A1(\gpio_configure[27][8] ),
    .A2(net516),
    .A3(_2697_),
    .B1(_2710_),
    .B2(\gpio_configure[20][8] ),
    .X(_2904_));
 sky130_fd_sc_hd__a221o_1 _6300_ (.A1(\gpio_configure[5][8] ),
    .A2(_2695_),
    .B1(_2724_),
    .B2(\gpio_configure[11][8] ),
    .C1(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__a32o_1 _6301_ (.A1(\gpio_configure[29][8] ),
    .A2(net516),
    .A3(net423),
    .B1(_2685_),
    .B2(\gpio_configure[17][8] ),
    .X(_2906_));
 sky130_fd_sc_hd__a221o_1 _6302_ (.A1(\gpio_configure[18][8] ),
    .A2(_2688_),
    .B1(_2712_),
    .B2(\gpio_configure[9][8] ),
    .C1(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__nor4_1 _6303_ (.A(_2901_),
    .B(_2903_),
    .C(_2905_),
    .D(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__a21bo_1 _6304_ (.A1(_2894_),
    .A2(_2896_),
    .B1_N(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__o21a_1 _6305_ (.A1(\gpio_configure[0][8] ),
    .A2(_2658_),
    .B1(net513),
    .X(_2910_));
 sky130_fd_sc_hd__a22o_1 _6306_ (.A1(net527),
    .A2(\serial_data_staging_1[7] ),
    .B1(_2909_),
    .B2(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__mux2_1 _6307_ (.A0(_2911_),
    .A1(net3819),
    .S(net353),
    .X(_0779_));
 sky130_fd_sc_hd__a32o_1 _6308_ (.A1(\gpio_configure[4][9] ),
    .A2(net445),
    .A3(net437),
    .B1(net436),
    .B2(\gpio_configure[10][9] ),
    .X(_2912_));
 sky130_fd_sc_hd__a31o_1 _6309_ (.A1(\gpio_configure[6][9] ),
    .A2(net446),
    .A3(net437),
    .B1(net518),
    .X(_2913_));
 sky130_fd_sc_hd__a32o_1 _6310_ (.A1(\gpio_configure[1][9] ),
    .A2(_2646_),
    .A3(net443),
    .B1(net422),
    .B2(\gpio_configure[14][9] ),
    .X(_2914_));
 sky130_fd_sc_hd__a221o_1 _6311_ (.A1(\gpio_configure[13][9] ),
    .A2(net423),
    .B1(_2687_),
    .B2(\gpio_configure[2][9] ),
    .C1(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__a2111o_1 _6312_ (.A1(\gpio_configure[12][9] ),
    .A2(_2702_),
    .B1(_2912_),
    .C1(_2913_),
    .D1(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__a32o_1 _6313_ (.A1(\gpio_configure[21][9] ),
    .A2(_2646_),
    .A3(net437),
    .B1(net422),
    .B2(\gpio_configure[30][9] ),
    .X(_2917_));
 sky130_fd_sc_hd__a211o_1 _6314_ (.A1(\gpio_configure[24][9] ),
    .A2(_2655_),
    .B1(_2917_),
    .C1(net511),
    .X(_2918_));
 sky130_fd_sc_hd__a32o_1 _6315_ (.A1(\gpio_configure[27][9] ),
    .A2(net518),
    .A3(_2697_),
    .B1(_2688_),
    .B2(\gpio_configure[18][9] ),
    .X(_2919_));
 sky130_fd_sc_hd__a221o_1 _6316_ (.A1(\gpio_configure[25][9] ),
    .A2(_2725_),
    .B1(_2734_),
    .B2(\gpio_configure[3][9] ),
    .C1(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__and3_1 _6317_ (.A(\gpio_configure[29][9] ),
    .B(\pad_count_1[4] ),
    .C(net423),
    .X(_2921_));
 sky130_fd_sc_hd__a32o_1 _6318_ (.A1(\gpio_configure[26][9] ),
    .A2(net518),
    .A3(net436),
    .B1(_2705_),
    .B2(\gpio_configure[31][9] ),
    .X(_2922_));
 sky130_fd_sc_hd__a2111o_1 _6319_ (.A1(\gpio_configure[20][9] ),
    .A2(_2710_),
    .B1(_2921_),
    .C1(_2922_),
    .D1(_2920_),
    .X(_2923_));
 sky130_fd_sc_hd__a32o_1 _6320_ (.A1(\gpio_configure[11][9] ),
    .A2(net511),
    .A3(_2697_),
    .B1(_2685_),
    .B2(\gpio_configure[17][9] ),
    .X(_2924_));
 sky130_fd_sc_hd__a221o_1 _6321_ (.A1(\gpio_configure[8][9] ),
    .A2(_2683_),
    .B1(_2723_),
    .B2(\gpio_configure[19][9] ),
    .C1(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__o211a_1 _6322_ (.A1(\gpio_configure[16][9] ),
    .A2(net511),
    .B1(net445),
    .C1(net443),
    .X(_2926_));
 sky130_fd_sc_hd__a31o_1 _6323_ (.A1(\gpio_configure[15][9] ),
    .A2(_2704_),
    .A3(net511),
    .B1(_2926_),
    .X(_2927_));
 sky130_fd_sc_hd__a221o_1 _6324_ (.A1(\gpio_configure[5][9] ),
    .A2(_2695_),
    .B1(_2707_),
    .B2(\gpio_configure[28][9] ),
    .C1(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__a32o_1 _6325_ (.A1(\gpio_configure[22][9] ),
    .A2(net518),
    .A3(_2692_),
    .B1(_2712_),
    .B2(\gpio_configure[9][9] ),
    .X(_2929_));
 sky130_fd_sc_hd__a221o_1 _6326_ (.A1(\gpio_configure[23][9] ),
    .A2(_2700_),
    .B1(_2733_),
    .B2(\gpio_configure[7][9] ),
    .C1(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__nor4_1 _6327_ (.A(_2923_),
    .B(_2925_),
    .C(_2928_),
    .D(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__a21bo_4 _6328_ (.A1(_2916_),
    .A2(_2918_),
    .B1_N(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__o21a_1 _6329_ (.A1(\gpio_configure[0][9] ),
    .A2(_2658_),
    .B1(net513),
    .X(_2933_));
 sky130_fd_sc_hd__a22o_1 _6330_ (.A1(net527),
    .A2(net3819),
    .B1(_2932_),
    .B2(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__mux2_1 _6331_ (.A0(_2934_),
    .A1(net3841),
    .S(net353),
    .X(_0780_));
 sky130_fd_sc_hd__and3_1 _6332_ (.A(\gpio_configure[26][10] ),
    .B(net516),
    .C(net436),
    .X(_2935_));
 sky130_fd_sc_hd__a32o_1 _6333_ (.A1(\gpio_configure[21][10] ),
    .A2(net447),
    .A3(net437),
    .B1(net422),
    .B2(\gpio_configure[30][10] ),
    .X(_2936_));
 sky130_fd_sc_hd__o211a_1 _6334_ (.A1(\gpio_configure[16][10] ),
    .A2(net510),
    .B1(net444),
    .C1(net442),
    .X(_2937_));
 sky130_fd_sc_hd__a32o_1 _6335_ (.A1(\gpio_configure[4][10] ),
    .A2(net444),
    .A3(net437),
    .B1(net423),
    .B2(\gpio_configure[13][10] ),
    .X(_2938_));
 sky130_fd_sc_hd__a32o_1 _6336_ (.A1(\gpio_configure[2][10] ),
    .A2(net446),
    .A3(net442),
    .B1(net436),
    .B2(\gpio_configure[10][10] ),
    .X(_2939_));
 sky130_fd_sc_hd__a32o_1 _6337_ (.A1(\gpio_configure[1][10] ),
    .A2(net447),
    .A3(net442),
    .B1(net422),
    .B2(\gpio_configure[14][10] ),
    .X(_2940_));
 sky130_fd_sc_hd__a31o_1 _6338_ (.A1(\gpio_configure[6][10] ),
    .A2(net446),
    .A3(net437),
    .B1(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__o31a_1 _6339_ (.A1(_2938_),
    .A2(_2939_),
    .A3(_2941_),
    .B1(net510),
    .X(_2942_));
 sky130_fd_sc_hd__a221o_1 _6340_ (.A1(\gpio_configure[31][10] ),
    .A2(_2705_),
    .B1(_2732_),
    .B2(\gpio_configure[15][10] ),
    .C1(_2937_),
    .X(_2943_));
 sky130_fd_sc_hd__a211o_1 _6341_ (.A1(net516),
    .A2(_2936_),
    .B1(_2943_),
    .C1(_2942_),
    .X(_2944_));
 sky130_fd_sc_hd__a32o_1 _6342_ (.A1(\gpio_configure[27][10] ),
    .A2(net516),
    .A3(_2697_),
    .B1(_2734_),
    .B2(\gpio_configure[3][10] ),
    .X(_2945_));
 sky130_fd_sc_hd__a31o_1 _6343_ (.A1(\gpio_configure[7][10] ),
    .A2(net510),
    .A3(_2699_),
    .B1(_2945_),
    .X(_2946_));
 sky130_fd_sc_hd__a32o_1 _6344_ (.A1(\gpio_configure[11][10] ),
    .A2(net510),
    .A3(_2697_),
    .B1(_2725_),
    .B2(\gpio_configure[25][10] ),
    .X(_2947_));
 sky130_fd_sc_hd__a32o_1 _6345_ (.A1(\gpio_configure[29][10] ),
    .A2(net516),
    .A3(net423),
    .B1(_2723_),
    .B2(\gpio_configure[19][10] ),
    .X(_2948_));
 sky130_fd_sc_hd__a221o_1 _6346_ (.A1(\gpio_configure[5][10] ),
    .A2(_2695_),
    .B1(_2710_),
    .B2(\gpio_configure[20][10] ),
    .C1(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__a211o_1 _6347_ (.A1(\gpio_configure[23][10] ),
    .A2(_2700_),
    .B1(_2947_),
    .C1(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__a32o_1 _6348_ (.A1(\gpio_configure[28][10] ),
    .A2(net516),
    .A3(_2702_),
    .B1(_2713_),
    .B2(\gpio_configure[24][10] ),
    .X(_2951_));
 sky130_fd_sc_hd__a221o_1 _6349_ (.A1(\gpio_configure[8][10] ),
    .A2(_2683_),
    .B1(_2703_),
    .B2(\gpio_configure[12][10] ),
    .C1(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__a32o_1 _6350_ (.A1(\gpio_configure[22][10] ),
    .A2(net516),
    .A3(_2692_),
    .B1(_2685_),
    .B2(\gpio_configure[17][10] ),
    .X(_2953_));
 sky130_fd_sc_hd__a2111o_1 _6351_ (.A1(\gpio_configure[18][10] ),
    .A2(_2688_),
    .B1(_2953_),
    .C1(_2935_),
    .D1(_2952_),
    .X(_2954_));
 sky130_fd_sc_hd__a2111o_1 _6352_ (.A1(\gpio_configure[9][10] ),
    .A2(_2712_),
    .B1(_2946_),
    .C1(_2950_),
    .D1(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__o221a_1 _6353_ (.A1(\gpio_configure[0][10] ),
    .A2(_2658_),
    .B1(_2944_),
    .B2(_2955_),
    .C1(net513),
    .X(_2956_));
 sky130_fd_sc_hd__a211o_1 _6354_ (.A1(net527),
    .A2(\serial_data_staging_1[9] ),
    .B1(net353),
    .C1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__o31a_1 _6355_ (.A1(net3839),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_2957_),
    .X(_0781_));
 sky130_fd_sc_hd__a32o_1 _6356_ (.A1(\gpio_configure[26][11] ),
    .A2(net518),
    .A3(net436),
    .B1(_2688_),
    .B2(\gpio_configure[18][11] ),
    .X(_2958_));
 sky130_fd_sc_hd__a221o_1 _6357_ (.A1(\gpio_configure[27][11] ),
    .A2(_2698_),
    .B1(_2732_),
    .B2(\gpio_configure[15][11] ),
    .C1(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__a32o_1 _6358_ (.A1(\gpio_configure[22][11] ),
    .A2(net518),
    .A3(_2692_),
    .B1(_2733_),
    .B2(\gpio_configure[7][11] ),
    .X(_2960_));
 sky130_fd_sc_hd__a221oi_4 _6359_ (.A1(\gpio_configure[17][11] ),
    .A2(_2685_),
    .B1(_2712_),
    .B2(\gpio_configure[9][11] ),
    .C1(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__a32o_1 _6360_ (.A1(\gpio_configure[5][11] ),
    .A2(net511),
    .A3(_2694_),
    .B1(_2710_),
    .B2(\gpio_configure[20][11] ),
    .X(_2962_));
 sky130_fd_sc_hd__a221oi_4 _6361_ (.A1(\gpio_configure[11][11] ),
    .A2(_2724_),
    .B1(_2734_),
    .B2(\gpio_configure[3][11] ),
    .C1(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__nand3b_4 _6362_ (.A_N(_2959_),
    .B(_2961_),
    .C(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__a32o_1 _6363_ (.A1(\gpio_configure[23][11] ),
    .A2(_2649_),
    .A3(net437),
    .B1(net423),
    .B2(\gpio_configure[29][11] ),
    .X(_2965_));
 sky130_fd_sc_hd__a221o_1 _6364_ (.A1(\gpio_configure[28][11] ),
    .A2(_2702_),
    .B1(net422),
    .B2(\gpio_configure[30][11] ),
    .C1(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__a31o_1 _6365_ (.A1(\gpio_configure[21][11] ),
    .A2(_2646_),
    .A3(net437),
    .B1(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__a32o_1 _6366_ (.A1(\gpio_configure[1][11] ),
    .A2(_2646_),
    .A3(net443),
    .B1(_2692_),
    .B2(\gpio_configure[6][11] ),
    .X(_2968_));
 sky130_fd_sc_hd__a221o_1 _6367_ (.A1(\gpio_configure[13][11] ),
    .A2(net423),
    .B1(net436),
    .B2(\gpio_configure[10][11] ),
    .C1(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__a32o_1 _6368_ (.A1(\gpio_configure[2][11] ),
    .A2(net446),
    .A3(net443),
    .B1(_2655_),
    .B2(\gpio_configure[8][11] ),
    .X(_2970_));
 sky130_fd_sc_hd__a32o_1 _6369_ (.A1(\gpio_configure[4][11] ),
    .A2(net445),
    .A3(net437),
    .B1(net422),
    .B2(\gpio_configure[14][11] ),
    .X(_2971_));
 sky130_fd_sc_hd__o31a_1 _6370_ (.A1(_2969_),
    .A2(_2970_),
    .A3(_2971_),
    .B1(net511),
    .X(_2972_));
 sky130_fd_sc_hd__a32o_1 _6371_ (.A1(\gpio_configure[12][11] ),
    .A2(_2702_),
    .A3(net511),
    .B1(\gpio_configure[24][11] ),
    .B2(_2713_),
    .X(_2973_));
 sky130_fd_sc_hd__a32o_1 _6372_ (.A1(\gpio_configure[31][11] ),
    .A2(net518),
    .A3(_2704_),
    .B1(_2723_),
    .B2(\gpio_configure[19][11] ),
    .X(_2974_));
 sky130_fd_sc_hd__o211a_1 _6373_ (.A1(\gpio_configure[16][11] ),
    .A2(net511),
    .B1(net445),
    .C1(net443),
    .X(_2975_));
 sky130_fd_sc_hd__a2111o_1 _6374_ (.A1(\gpio_configure[25][11] ),
    .A2(_2725_),
    .B1(_2973_),
    .C1(_2975_),
    .D1(_2974_),
    .X(_2976_));
 sky130_fd_sc_hd__a211o_2 _6375_ (.A1(net518),
    .A2(_2967_),
    .B1(_2972_),
    .C1(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__o221ai_4 _6376_ (.A1(\gpio_configure[0][11] ),
    .A2(_2658_),
    .B1(_2964_),
    .B2(_2977_),
    .C1(net513),
    .Y(_2978_));
 sky130_fd_sc_hd__o2bb2a_1 _6377_ (.A1_N(net527),
    .A2_N(\serial_data_staging_1[10] ),
    .B1(_1446_),
    .B2(_2680_),
    .X(_2979_));
 sky130_fd_sc_hd__o2bb2a_1 _6378_ (.A1_N(_2979_),
    .A2_N(_2978_),
    .B1(_2682_),
    .B2(net3862),
    .X(_0782_));
 sky130_fd_sc_hd__a32o_1 _6379_ (.A1(\gpio_configure[6][12] ),
    .A2(net446),
    .A3(net437),
    .B1(net422),
    .B2(\gpio_configure[14][12] ),
    .X(_2980_));
 sky130_fd_sc_hd__a31o_1 _6380_ (.A1(\gpio_configure[4][12] ),
    .A2(net445),
    .A3(net437),
    .B1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__a32o_1 _6381_ (.A1(\gpio_configure[1][12] ),
    .A2(_2646_),
    .A3(net443),
    .B1(net436),
    .B2(\gpio_configure[10][12] ),
    .X(_2982_));
 sky130_fd_sc_hd__a221o_1 _6382_ (.A1(\gpio_configure[13][12] ),
    .A2(net423),
    .B1(_2702_),
    .B2(\gpio_configure[12][12] ),
    .C1(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__a2111o_1 _6383_ (.A1(\gpio_configure[2][12] ),
    .A2(_2687_),
    .B1(net518),
    .C1(_2983_),
    .D1(_2981_),
    .X(_2984_));
 sky130_fd_sc_hd__a41o_1 _6384_ (.A1(\gpio_configure[30][12] ),
    .A2(net520),
    .A3(net522),
    .A4(net446),
    .B1(net511),
    .X(_2985_));
 sky130_fd_sc_hd__a221o_1 _6385_ (.A1(\gpio_configure[24][12] ),
    .A2(_2655_),
    .B1(_2694_),
    .B2(\gpio_configure[21][12] ),
    .C1(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__a22o_1 _6386_ (.A1(\gpio_configure[25][12] ),
    .A2(_2725_),
    .B1(_2734_),
    .B2(\gpio_configure[3][12] ),
    .X(_2987_));
 sky130_fd_sc_hd__o211a_1 _6387_ (.A1(\gpio_configure[16][12] ),
    .A2(net511),
    .B1(net445),
    .C1(net443),
    .X(_2988_));
 sky130_fd_sc_hd__a32o_1 _6388_ (.A1(\gpio_configure[27][12] ),
    .A2(net518),
    .A3(_2697_),
    .B1(_2695_),
    .B2(\gpio_configure[5][12] ),
    .X(_2989_));
 sky130_fd_sc_hd__a221o_1 _6389_ (.A1(\gpio_configure[9][12] ),
    .A2(_2712_),
    .B1(_2724_),
    .B2(\gpio_configure[11][12] ),
    .C1(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__a2111o_1 _6390_ (.A1(\gpio_configure[7][12] ),
    .A2(_2733_),
    .B1(_2987_),
    .C1(_2988_),
    .D1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__a32o_1 _6391_ (.A1(\gpio_configure[26][12] ),
    .A2(net518),
    .A3(net436),
    .B1(_2688_),
    .B2(\gpio_configure[18][12] ),
    .X(_2992_));
 sky130_fd_sc_hd__a221o_1 _6392_ (.A1(\gpio_configure[20][12] ),
    .A2(_2710_),
    .B1(_2723_),
    .B2(\gpio_configure[19][12] ),
    .C1(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__a32o_1 _6393_ (.A1(\gpio_configure[28][12] ),
    .A2(net518),
    .A3(_2702_),
    .B1(_2705_),
    .B2(\gpio_configure[31][12] ),
    .X(_2994_));
 sky130_fd_sc_hd__a221o_1 _6394_ (.A1(\gpio_configure[23][12] ),
    .A2(_2700_),
    .B1(_2732_),
    .B2(\gpio_configure[15][12] ),
    .C1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__a32o_1 _6395_ (.A1(\gpio_configure[29][12] ),
    .A2(\pad_count_1[4] ),
    .A3(net423),
    .B1(_2685_),
    .B2(\gpio_configure[17][12] ),
    .X(_2996_));
 sky130_fd_sc_hd__a221o_1 _6396_ (.A1(\gpio_configure[8][12] ),
    .A2(_2683_),
    .B1(_2693_),
    .B2(\gpio_configure[22][12] ),
    .C1(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__nor4_1 _6397_ (.A(_2991_),
    .B(_2993_),
    .C(_2995_),
    .D(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__a21bo_4 _6398_ (.A1(_2984_),
    .A2(_2986_),
    .B1_N(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__o21a_1 _6399_ (.A1(\gpio_configure[0][12] ),
    .A2(_2658_),
    .B1(net513),
    .X(_3000_));
 sky130_fd_sc_hd__a22o_1 _6400_ (.A1(net527),
    .A2(\serial_data_staging_1[11] ),
    .B1(_2999_),
    .B2(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__mux2_1 _6401_ (.A0(_3001_),
    .A1(net3858),
    .S(net353),
    .X(_0783_));
 sky130_fd_sc_hd__nor2_8 _6402_ (.A(net514),
    .B(net515),
    .Y(_3002_));
 sky130_fd_sc_hd__and3_4 _6403_ (.A(_1438_),
    .B(_1439_),
    .C(net435),
    .X(_3003_));
 sky130_fd_sc_hd__nor2_8 _6404_ (.A(\pad_count_2[4] ),
    .B(\pad_count_2[5] ),
    .Y(_3004_));
 sky130_fd_sc_hd__and4_4 _6405_ (.A(net514),
    .B(\pad_count_2[2] ),
    .C(net441),
    .D(net432),
    .X(_3005_));
 sky130_fd_sc_hd__and4bb_4 _6406_ (.A_N(\pad_count_2[1] ),
    .B_N(\pad_count_2[4] ),
    .C(\pad_count_2[5] ),
    .D(_1440_),
    .X(_3006_));
 sky130_fd_sc_hd__and3_4 _6407_ (.A(_1439_),
    .B(net441),
    .C(net435),
    .X(_3007_));
 sky130_fd_sc_hd__nor4_4 _6408_ (.A(_3003_),
    .B(_3005_),
    .C(_3006_),
    .D(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__and4_4 _6409_ (.A(net514),
    .B(net515),
    .C(_2662_),
    .D(net432),
    .X(_3009_));
 sky130_fd_sc_hd__and3_1 _6410_ (.A(\pad_count_2[1] ),
    .B(_1440_),
    .C(net432),
    .X(_3010_));
 sky130_fd_sc_hd__a2111oi_1 _6411_ (.A1(_2664_),
    .A2(net432),
    .B1(_3009_),
    .C1(_3010_),
    .D1(net439),
    .Y(_3011_));
 sky130_fd_sc_hd__and3_4 _6412_ (.A(_1438_),
    .B(net435),
    .C(net432),
    .X(_3012_));
 sky130_fd_sc_hd__and3_4 _6413_ (.A(_2662_),
    .B(net435),
    .C(net433),
    .X(_3013_));
 sky130_fd_sc_hd__and4_4 _6414_ (.A(net514),
    .B(net515),
    .C(_1438_),
    .D(net432),
    .X(_3014_));
 sky130_fd_sc_hd__and3_4 _6415_ (.A(_1439_),
    .B(_2664_),
    .C(net435),
    .X(_3015_));
 sky130_fd_sc_hd__and4bb_1 _6416_ (.A_N(net515),
    .B_N(_2664_),
    .C(net432),
    .D(net514),
    .X(_3016_));
 sky130_fd_sc_hd__and3_4 _6417_ (.A(_1439_),
    .B(_2662_),
    .C(net435),
    .X(_3017_));
 sky130_fd_sc_hd__and3_4 _6418_ (.A(_1440_),
    .B(_2663_),
    .C(net434),
    .X(_3018_));
 sky130_fd_sc_hd__nor4_1 _6419_ (.A(_3015_),
    .B(_3016_),
    .C(_3017_),
    .D(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__nor4b_4 _6420_ (.A(_3012_),
    .B(_3013_),
    .C(_3014_),
    .D_N(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__and3_4 _6421_ (.A(_1440_),
    .B(_2664_),
    .C(net432),
    .X(_3021_));
 sky130_fd_sc_hd__and3_4 _6422_ (.A(_2664_),
    .B(net435),
    .C(net434),
    .X(_3022_));
 sky130_fd_sc_hd__and3_4 _6423_ (.A(_1438_),
    .B(_1440_),
    .C(net432),
    .X(_3023_));
 sky130_fd_sc_hd__and3_4 _6424_ (.A(_1439_),
    .B(_1440_),
    .C(_2663_),
    .X(_3024_));
 sky130_fd_sc_hd__and3_4 _6425_ (.A(_1440_),
    .B(_2662_),
    .C(net434),
    .X(_3025_));
 sky130_fd_sc_hd__and3_4 _6426_ (.A(net514),
    .B(net515),
    .C(_2664_),
    .X(_3026_));
 sky130_fd_sc_hd__and3_4 _6427_ (.A(_1439_),
    .B(_1440_),
    .C(_2664_),
    .X(_3027_));
 sky130_fd_sc_hd__and4bb_4 _6428_ (.A_N(\pad_count_2[1] ),
    .B_N(net515),
    .C(net514),
    .D(\pad_count_2[0] ),
    .X(_3028_));
 sky130_fd_sc_hd__and4b_4 _6429_ (.A_N(net515),
    .B(net514),
    .C(\pad_count_2[0] ),
    .D(\pad_count_2[1] ),
    .X(_3029_));
 sky130_fd_sc_hd__and3_4 _6430_ (.A(_3008_),
    .B(net393),
    .C(_3020_),
    .X(_3030_));
 sky130_fd_sc_hd__nand3_4 _6431_ (.A(_3008_),
    .B(net393),
    .C(_3020_),
    .Y(_3031_));
 sky130_fd_sc_hd__a22o_1 _6432_ (.A1(\gpio_configure[31][0] ),
    .A2(_2674_),
    .B1(_3024_),
    .B2(\gpio_configure[36][0] ),
    .X(_3032_));
 sky130_fd_sc_hd__and4bb_4 _6433_ (.A_N(net514),
    .B_N(\pad_count_2[5] ),
    .C(\pad_count_2[4] ),
    .D(net515),
    .X(_3033_));
 sky130_fd_sc_hd__and3_4 _6434_ (.A(_1440_),
    .B(_2662_),
    .C(net439),
    .X(_3034_));
 sky130_fd_sc_hd__and4_4 _6435_ (.A(net514),
    .B(net515),
    .C(_2664_),
    .D(net439),
    .X(_3035_));
 sky130_fd_sc_hd__a22o_1 _6436_ (.A1(\gpio_configure[5][0] ),
    .A2(_3021_),
    .B1(_3035_),
    .B2(\gpio_configure[29][0] ),
    .X(_3036_));
 sky130_fd_sc_hd__a221o_1 _6437_ (.A1(\gpio_configure[34][0] ),
    .A2(_3003_),
    .B1(_3034_),
    .B2(\gpio_configure[23][0] ),
    .C1(_3036_),
    .X(_3037_));
 sky130_fd_sc_hd__a22o_1 _6438_ (.A1(\gpio_configure[14][0] ),
    .A2(_3014_),
    .B1(_3015_),
    .B2(\gpio_configure[33][0] ),
    .X(_3038_));
 sky130_fd_sc_hd__a211o_1 _6439_ (.A1(\gpio_configure[15][0] ),
    .A2(_3009_),
    .B1(_3037_),
    .C1(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__a2111oi_4 _6440_ (.A1(\gpio_configure[37][0] ),
    .A2(_3027_),
    .B1(_3032_),
    .C1(_3039_),
    .D1(_3030_),
    .Y(_3040_));
 sky130_fd_sc_hd__and4bb_4 _6441_ (.A_N(net515),
    .B_N(\pad_count_2[5] ),
    .C(\pad_count_2[4] ),
    .D(net514),
    .X(_3041_));
 sky130_fd_sc_hd__a32o_1 _6442_ (.A1(\gpio_configure[27][0] ),
    .A2(net439),
    .A3(net431),
    .B1(_3022_),
    .B2(\gpio_configure[1][0] ),
    .X(_3042_));
 sky130_fd_sc_hd__and3_4 _6443_ (.A(_1440_),
    .B(_2664_),
    .C(net440),
    .X(_3043_));
 sky130_fd_sc_hd__a32o_1 _6444_ (.A1(\gpio_configure[21][0] ),
    .A2(_2664_),
    .A3(net430),
    .B1(_3023_),
    .B2(\gpio_configure[6][0] ),
    .X(_3044_));
 sky130_fd_sc_hd__a221o_1 _6445_ (.A1(\gpio_configure[32][0] ),
    .A2(_3007_),
    .B1(_3012_),
    .B2(\gpio_configure[2][0] ),
    .C1(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__and4_4 _6446_ (.A(net514),
    .B(\pad_count_2[2] ),
    .C(_1438_),
    .D(net439),
    .X(_3046_));
 sky130_fd_sc_hd__and3_4 _6447_ (.A(_1440_),
    .B(net441),
    .C(net440),
    .X(_3047_));
 sky130_fd_sc_hd__a32o_1 _6448_ (.A1(\gpio_configure[20][0] ),
    .A2(_2663_),
    .A3(net430),
    .B1(_3046_),
    .B2(\gpio_configure[30][0] ),
    .X(_3048_));
 sky130_fd_sc_hd__a221o_1 _6449_ (.A1(\gpio_configure[4][0] ),
    .A2(_3018_),
    .B1(_3025_),
    .B2(\gpio_configure[7][0] ),
    .C1(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__a2111o_1 _6450_ (.A1(\gpio_configure[35][0] ),
    .A2(_3017_),
    .B1(_3042_),
    .C1(_3045_),
    .D1(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__and4b_4 _6451_ (.A_N(\pad_count_2[2] ),
    .B(_2664_),
    .C(net439),
    .D(\pad_count_2[3] ),
    .X(_3051_));
 sky130_fd_sc_hd__and4b_4 _6452_ (.A_N(\pad_count_2[2] ),
    .B(net441),
    .C(net432),
    .D(\pad_count_2[3] ),
    .X(_3052_));
 sky130_fd_sc_hd__a32o_1 _6453_ (.A1(\gpio_configure[25][0] ),
    .A2(net440),
    .A3(_3028_),
    .B1(_3052_),
    .B2(\gpio_configure[8][0] ),
    .X(_3053_));
 sky130_fd_sc_hd__and4b_4 _6454_ (.A_N(\pad_count_2[2] ),
    .B(_1438_),
    .C(net439),
    .D(\pad_count_2[3] ),
    .X(_3054_));
 sky130_fd_sc_hd__and3_4 _6455_ (.A(_1438_),
    .B(_1440_),
    .C(net439),
    .X(_3055_));
 sky130_fd_sc_hd__a221o_1 _6456_ (.A1(\gpio_configure[26][0] ),
    .A2(_3054_),
    .B1(_3055_),
    .B2(\gpio_configure[22][0] ),
    .C1(_3053_),
    .X(_3056_));
 sky130_fd_sc_hd__and4b_4 _6457_ (.A_N(\pad_count_2[2] ),
    .B(net441),
    .C(net439),
    .D(\pad_count_2[3] ),
    .X(_3057_));
 sky130_fd_sc_hd__a32o_1 _6458_ (.A1(\gpio_configure[19][0] ),
    .A2(_2673_),
    .A3(_3002_),
    .B1(_3057_),
    .B2(\gpio_configure[24][0] ),
    .X(_3058_));
 sky130_fd_sc_hd__and3_1 _6459_ (.A(\gpio_configure[9][0] ),
    .B(net434),
    .C(_3028_),
    .X(_3059_));
 sky130_fd_sc_hd__and4_4 _6460_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .C(_2664_),
    .D(net432),
    .X(_3060_));
 sky130_fd_sc_hd__a2111o_2 _6461_ (.A1(\gpio_configure[13][0] ),
    .A2(_3060_),
    .B1(_3059_),
    .C1(_3058_),
    .D1(_3056_),
    .X(_3061_));
 sky130_fd_sc_hd__and4b_4 _6462_ (.A_N(net515),
    .B(_1438_),
    .C(net432),
    .D(net514),
    .X(_3062_));
 sky130_fd_sc_hd__and3_4 _6463_ (.A(_1438_),
    .B(net439),
    .C(net435),
    .X(_3063_));
 sky130_fd_sc_hd__a22o_1 _6464_ (.A1(\gpio_configure[12][0] ),
    .A2(_3005_),
    .B1(_3063_),
    .B2(\gpio_configure[18][0] ),
    .X(_3064_));
 sky130_fd_sc_hd__a221o_1 _6465_ (.A1(\gpio_configure[3][0] ),
    .A2(_3013_),
    .B1(_3062_),
    .B2(\gpio_configure[10][0] ),
    .C1(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__and4_4 _6466_ (.A(\pad_count_2[3] ),
    .B(\pad_count_2[2] ),
    .C(net441),
    .D(net439),
    .X(_3066_));
 sky130_fd_sc_hd__and3_4 _6467_ (.A(_2664_),
    .B(net439),
    .C(net435),
    .X(_3067_));
 sky130_fd_sc_hd__and3_4 _6468_ (.A(net441),
    .B(net439),
    .C(net435),
    .X(_3068_));
 sky130_fd_sc_hd__a32o_1 _6469_ (.A1(\gpio_configure[11][0] ),
    .A2(net434),
    .A3(_3029_),
    .B1(_3068_),
    .B2(\gpio_configure[16][0] ),
    .X(_3069_));
 sky130_fd_sc_hd__a221o_1 _6470_ (.A1(\gpio_configure[28][0] ),
    .A2(_3066_),
    .B1(_3067_),
    .B2(\gpio_configure[17][0] ),
    .C1(_3069_),
    .X(_3070_));
 sky130_fd_sc_hd__nor4_2 _6471_ (.A(_3050_),
    .B(_3061_),
    .C(_3065_),
    .D(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__o2bb2a_1 _6472_ (.A1_N(net348),
    .A2_N(_3071_),
    .B1(\gpio_configure[0][0] ),
    .B2(_3031_),
    .X(_3072_));
 sky130_fd_sc_hd__a32o_1 _6473_ (.A1(_3072_),
    .A2(net513),
    .A3(\xfer_state[2] ),
    .B1(net353),
    .B2(net3837),
    .X(_0784_));
 sky130_fd_sc_hd__a32o_1 _6474_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][1] ),
    .A3(_3006_),
    .B1(_2674_),
    .B2(\gpio_configure[31][1] ),
    .X(_3073_));
 sky130_fd_sc_hd__a32o_1 _6475_ (.A1(\gpio_configure[21][1] ),
    .A2(_2664_),
    .A3(_3033_),
    .B1(_3005_),
    .B2(\gpio_configure[12][1] ),
    .X(_3074_));
 sky130_fd_sc_hd__a221o_1 _6476_ (.A1(\gpio_configure[30][1] ),
    .A2(_3046_),
    .B1(_3047_),
    .B2(\gpio_configure[20][1] ),
    .C1(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__a22o_1 _6477_ (.A1(\gpio_configure[29][1] ),
    .A2(_3035_),
    .B1(_3066_),
    .B2(\gpio_configure[28][1] ),
    .X(_3076_));
 sky130_fd_sc_hd__a211o_1 _6478_ (.A1(\gpio_configure[15][1] ),
    .A2(_3009_),
    .B1(_3075_),
    .C1(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__a2111o_1 _6479_ (.A1(\gpio_configure[36][1] ),
    .A2(_3024_),
    .B1(_3073_),
    .C1(_3077_),
    .D1(_3030_),
    .X(_3078_));
 sky130_fd_sc_hd__a32o_1 _6480_ (.A1(\gpio_configure[19][1] ),
    .A2(_2673_),
    .A3(_3002_),
    .B1(_3021_),
    .B2(\gpio_configure[5][1] ),
    .X(_3079_));
 sky130_fd_sc_hd__a32o_1 _6481_ (.A1(\gpio_configure[22][1] ),
    .A2(_1438_),
    .A3(_3033_),
    .B1(_3025_),
    .B2(\gpio_configure[7][1] ),
    .X(_3080_));
 sky130_fd_sc_hd__a221o_2 _6482_ (.A1(\gpio_configure[14][1] ),
    .A2(_3014_),
    .B1(_3015_),
    .B2(\gpio_configure[33][1] ),
    .C1(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__a32o_1 _6483_ (.A1(\gpio_configure[9][1] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3062_),
    .B2(\gpio_configure[10][1] ),
    .X(_3082_));
 sky130_fd_sc_hd__a221o_1 _6484_ (.A1(\gpio_configure[3][1] ),
    .A2(_3013_),
    .B1(_3054_),
    .B2(\gpio_configure[26][1] ),
    .C1(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__a2111oi_4 _6485_ (.A1(\gpio_configure[25][1] ),
    .A2(_3051_),
    .B1(_3079_),
    .C1(_3081_),
    .D1(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__a32o_1 _6486_ (.A1(\gpio_configure[11][1] ),
    .A2(net433),
    .A3(net431),
    .B1(_3022_),
    .B2(\gpio_configure[1][1] ),
    .X(_3085_));
 sky130_fd_sc_hd__a221o_1 _6487_ (.A1(\gpio_configure[2][1] ),
    .A2(_3012_),
    .B1(_3067_),
    .B2(\gpio_configure[17][1] ),
    .C1(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__a32o_1 _6488_ (.A1(\gpio_configure[24][1] ),
    .A2(net441),
    .A3(_3041_),
    .B1(_3023_),
    .B2(\gpio_configure[6][1] ),
    .X(_3087_));
 sky130_fd_sc_hd__a221o_1 _6489_ (.A1(\gpio_configure[34][1] ),
    .A2(_3003_),
    .B1(_3007_),
    .B2(\gpio_configure[32][1] ),
    .C1(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__a32o_1 _6490_ (.A1(\gpio_configure[27][1] ),
    .A2(net440),
    .A3(_3029_),
    .B1(_3017_),
    .B2(\gpio_configure[35][1] ),
    .X(_3089_));
 sky130_fd_sc_hd__a221o_1 _6491_ (.A1(\gpio_configure[23][1] ),
    .A2(_3034_),
    .B1(_3060_),
    .B2(\gpio_configure[13][1] ),
    .C1(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__a22o_1 _6492_ (.A1(\gpio_configure[4][1] ),
    .A2(_3018_),
    .B1(_3052_),
    .B2(\gpio_configure[8][1] ),
    .X(_3091_));
 sky130_fd_sc_hd__a221o_1 _6493_ (.A1(\gpio_configure[18][1] ),
    .A2(_3063_),
    .B1(_3068_),
    .B2(\gpio_configure[16][1] ),
    .C1(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__nor4_2 _6494_ (.A(_3086_),
    .B(_3088_),
    .C(_3090_),
    .D(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__nand3b_4 _6495_ (.A_N(_3078_),
    .B(_3084_),
    .C(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__o21a_1 _6496_ (.A1(\gpio_configure[0][1] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3095_));
 sky130_fd_sc_hd__a22o_1 _6497_ (.A1(net528),
    .A2(\serial_data_staging_2[0] ),
    .B1(_3094_),
    .B2(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__mux2_1 _6498_ (.A0(_3096_),
    .A1(net3817),
    .S(net353),
    .X(_0785_));
 sky130_fd_sc_hd__a32o_1 _6499_ (.A1(\gpio_configure[26][2] ),
    .A2(_1438_),
    .A3(_3041_),
    .B1(_3025_),
    .B2(\gpio_configure[7][2] ),
    .X(_3097_));
 sky130_fd_sc_hd__a32o_1 _6500_ (.A1(\gpio_configure[11][2] ),
    .A2(net432),
    .A3(net431),
    .B1(_3057_),
    .B2(\gpio_configure[24][2] ),
    .X(_3098_));
 sky130_fd_sc_hd__a221o_1 _6501_ (.A1(\gpio_configure[31][2] ),
    .A2(_2674_),
    .B1(_3022_),
    .B2(\gpio_configure[1][2] ),
    .C1(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__a221o_1 _6502_ (.A1(\gpio_configure[15][2] ),
    .A2(_3009_),
    .B1(_3013_),
    .B2(\gpio_configure[3][2] ),
    .C1(_3097_),
    .X(_3100_));
 sky130_fd_sc_hd__a32o_1 _6503_ (.A1(\gpio_configure[9][2] ),
    .A2(net433),
    .A3(_3028_),
    .B1(_3005_),
    .B2(\gpio_configure[12][2] ),
    .X(_3101_));
 sky130_fd_sc_hd__a32o_1 _6504_ (.A1(\gpio_configure[13][2] ),
    .A2(net433),
    .A3(_3026_),
    .B1(_3051_),
    .B2(\gpio_configure[25][2] ),
    .X(_3102_));
 sky130_fd_sc_hd__a221o_1 _6505_ (.A1(\gpio_configure[2][2] ),
    .A2(_3012_),
    .B1(_3021_),
    .B2(\gpio_configure[5][2] ),
    .C1(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__a211o_1 _6506_ (.A1(\gpio_configure[6][2] ),
    .A2(_3023_),
    .B1(_3101_),
    .C1(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__a32o_1 _6507_ (.A1(\gpio_configure[19][2] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3003_),
    .B2(\gpio_configure[34][2] ),
    .X(_3105_));
 sky130_fd_sc_hd__a31o_1 _6508_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][2] ),
    .A3(_3006_),
    .B1(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__a221o_1 _6509_ (.A1(\gpio_configure[4][2] ),
    .A2(_3018_),
    .B1(_3024_),
    .B2(\gpio_configure[36][2] ),
    .C1(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__a41o_1 _6510_ (.A1(\gpio_configure[32][2] ),
    .A2(_1439_),
    .A3(net441),
    .A4(net435),
    .B1(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__a2111o_1 _6511_ (.A1(\gpio_configure[10][2] ),
    .A2(_3062_),
    .B1(_3100_),
    .C1(_3104_),
    .D1(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__a22o_1 _6512_ (.A1(\gpio_configure[29][2] ),
    .A2(_3035_),
    .B1(_3046_),
    .B2(\gpio_configure[30][2] ),
    .X(_3110_));
 sky130_fd_sc_hd__a32o_1 _6513_ (.A1(\gpio_configure[23][2] ),
    .A2(_2662_),
    .A3(net430),
    .B1(_3066_),
    .B2(\gpio_configure[28][2] ),
    .X(_3111_));
 sky130_fd_sc_hd__a31o_1 _6514_ (.A1(\gpio_configure[20][2] ),
    .A2(_2663_),
    .A3(net430),
    .B1(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__a221o_1 _6515_ (.A1(\gpio_configure[35][2] ),
    .A2(_3017_),
    .B1(_3043_),
    .B2(\gpio_configure[21][2] ),
    .C1(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__a211o_4 _6516_ (.A1(\gpio_configure[33][2] ),
    .A2(_3015_),
    .B1(_3110_),
    .C1(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__a32o_1 _6517_ (.A1(\gpio_configure[27][2] ),
    .A2(net439),
    .A3(net431),
    .B1(_3052_),
    .B2(\gpio_configure[8][2] ),
    .X(_3115_));
 sky130_fd_sc_hd__a221o_1 _6518_ (.A1(\gpio_configure[14][2] ),
    .A2(_3014_),
    .B1(_3067_),
    .B2(\gpio_configure[17][2] ),
    .C1(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__a221o_1 _6519_ (.A1(\gpio_configure[22][2] ),
    .A2(_3055_),
    .B1(_3063_),
    .B2(\gpio_configure[18][2] ),
    .C1(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__a2111o_1 _6520_ (.A1(\gpio_configure[16][2] ),
    .A2(_3068_),
    .B1(_3030_),
    .C1(_3117_),
    .D1(_3114_),
    .X(_3118_));
 sky130_fd_sc_hd__o32a_1 _6521_ (.A1(_3099_),
    .A2(_3109_),
    .A3(_3118_),
    .B1(_3031_),
    .B2(\gpio_configure[0][2] ),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _6522_ (.A0(_3119_),
    .A1(net3817),
    .S(net528),
    .X(_3120_));
 sky130_fd_sc_hd__mux2_1 _6523_ (.A0(_3120_),
    .A1(net3829),
    .S(_2681_),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _6524_ (.A1(\gpio_configure[31][3] ),
    .A2(_2674_),
    .B1(_3009_),
    .B2(\gpio_configure[15][3] ),
    .X(_3121_));
 sky130_fd_sc_hd__a32o_1 _6525_ (.A1(\gpio_configure[27][3] ),
    .A2(net440),
    .A3(_3029_),
    .B1(_3067_),
    .B2(\gpio_configure[17][3] ),
    .X(_3122_));
 sky130_fd_sc_hd__a221o_1 _6526_ (.A1(\gpio_configure[35][3] ),
    .A2(_3017_),
    .B1(_3066_),
    .B2(\gpio_configure[28][3] ),
    .C1(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__a32o_1 _6527_ (.A1(\gpio_configure[11][3] ),
    .A2(net434),
    .A3(net431),
    .B1(_3055_),
    .B2(\gpio_configure[22][3] ),
    .X(_3124_));
 sky130_fd_sc_hd__a211o_1 _6528_ (.A1(\gpio_configure[36][3] ),
    .A2(_3024_),
    .B1(_3123_),
    .C1(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__a2111o_1 _6529_ (.A1(\gpio_configure[37][3] ),
    .A2(_3027_),
    .B1(_3121_),
    .C1(_3125_),
    .D1(_3030_),
    .X(_3126_));
 sky130_fd_sc_hd__a22o_1 _6530_ (.A1(\gpio_configure[34][3] ),
    .A2(_3003_),
    .B1(_3063_),
    .B2(\gpio_configure[18][3] ),
    .X(_3127_));
 sky130_fd_sc_hd__a32o_1 _6531_ (.A1(\gpio_configure[19][3] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3047_),
    .B2(\gpio_configure[20][3] ),
    .X(_3128_));
 sky130_fd_sc_hd__a221o_2 _6532_ (.A1(\gpio_configure[1][3] ),
    .A2(_3022_),
    .B1(_3043_),
    .B2(\gpio_configure[21][3] ),
    .C1(_3128_),
    .X(_3129_));
 sky130_fd_sc_hd__a32o_1 _6533_ (.A1(\gpio_configure[9][3] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3051_),
    .B2(\gpio_configure[25][3] ),
    .X(_3130_));
 sky130_fd_sc_hd__a221o_1 _6534_ (.A1(\gpio_configure[32][3] ),
    .A2(_3007_),
    .B1(_3025_),
    .B2(\gpio_configure[7][3] ),
    .C1(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__a2111oi_4 _6535_ (.A1(\gpio_configure[2][3] ),
    .A2(_3012_),
    .B1(_3127_),
    .C1(_3129_),
    .D1(_3131_),
    .Y(_3132_));
 sky130_fd_sc_hd__a32o_1 _6536_ (.A1(\gpio_configure[23][3] ),
    .A2(_2662_),
    .A3(_3033_),
    .B1(_3046_),
    .B2(\gpio_configure[30][3] ),
    .X(_3133_));
 sky130_fd_sc_hd__a221o_1 _6537_ (.A1(\gpio_configure[10][3] ),
    .A2(_3062_),
    .B1(_3068_),
    .B2(\gpio_configure[16][3] ),
    .C1(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__a32o_1 _6538_ (.A1(\gpio_configure[6][3] ),
    .A2(_1441_),
    .A3(net434),
    .B1(_3013_),
    .B2(\gpio_configure[3][3] ),
    .X(_3135_));
 sky130_fd_sc_hd__a221o_1 _6539_ (.A1(\gpio_configure[33][3] ),
    .A2(_3015_),
    .B1(_3035_),
    .B2(\gpio_configure[29][3] ),
    .C1(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__a22o_1 _6540_ (.A1(\gpio_configure[12][3] ),
    .A2(_3005_),
    .B1(_3060_),
    .B2(\gpio_configure[13][3] ),
    .X(_3137_));
 sky130_fd_sc_hd__a221o_1 _6541_ (.A1(\gpio_configure[14][3] ),
    .A2(_3014_),
    .B1(_3021_),
    .B2(\gpio_configure[5][3] ),
    .C1(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__a32o_1 _6542_ (.A1(\gpio_configure[24][3] ),
    .A2(_2663_),
    .A3(_3041_),
    .B1(_3052_),
    .B2(\gpio_configure[8][3] ),
    .X(_3139_));
 sky130_fd_sc_hd__a221o_1 _6543_ (.A1(\gpio_configure[4][3] ),
    .A2(_3018_),
    .B1(_3054_),
    .B2(\gpio_configure[26][3] ),
    .C1(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__nor4_2 _6544_ (.A(_3134_),
    .B(_3136_),
    .C(_3138_),
    .D(_3140_),
    .Y(_3141_));
 sky130_fd_sc_hd__nand3b_4 _6545_ (.A_N(_3126_),
    .B(_3132_),
    .C(_3141_),
    .Y(_3142_));
 sky130_fd_sc_hd__o21a_1 _6546_ (.A1(\gpio_configure[0][3] ),
    .A2(_3031_),
    .B1(_0824_),
    .X(_3143_));
 sky130_fd_sc_hd__a22o_1 _6547_ (.A1(net528),
    .A2(\serial_data_staging_2[2] ),
    .B1(_3142_),
    .B2(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__mux2_1 _6548_ (.A0(_3144_),
    .A1(net3826),
    .S(_2681_),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _6549_ (.A1(\gpio_configure[36][4] ),
    .A2(_3024_),
    .B1(_3027_),
    .B2(\gpio_configure[37][4] ),
    .X(_3145_));
 sky130_fd_sc_hd__a32o_1 _6550_ (.A1(\gpio_configure[21][4] ),
    .A2(_2664_),
    .A3(net430),
    .B1(_3046_),
    .B2(\gpio_configure[30][4] ),
    .X(_3146_));
 sky130_fd_sc_hd__a221o_1 _6551_ (.A1(\gpio_configure[6][4] ),
    .A2(_3023_),
    .B1(_3052_),
    .B2(\gpio_configure[8][4] ),
    .C1(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__a22o_1 _6552_ (.A1(\gpio_configure[18][4] ),
    .A2(_3063_),
    .B1(_3067_),
    .B2(\gpio_configure[17][4] ),
    .X(_3148_));
 sky130_fd_sc_hd__a211o_1 _6553_ (.A1(\gpio_configure[31][4] ),
    .A2(_2674_),
    .B1(_3147_),
    .C1(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__a2111o_1 _6554_ (.A1(\gpio_configure[15][4] ),
    .A2(_3009_),
    .B1(_3145_),
    .C1(_3149_),
    .D1(_3030_),
    .X(_3150_));
 sky130_fd_sc_hd__a32o_1 _6555_ (.A1(\gpio_configure[19][4] ),
    .A2(_2673_),
    .A3(_3002_),
    .B1(_3060_),
    .B2(\gpio_configure[13][4] ),
    .X(_3151_));
 sky130_fd_sc_hd__a32o_1 _6556_ (.A1(\gpio_configure[9][4] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3014_),
    .B2(\gpio_configure[14][4] ),
    .X(_3152_));
 sky130_fd_sc_hd__a221o_1 _6557_ (.A1(\gpio_configure[35][4] ),
    .A2(_3017_),
    .B1(_3034_),
    .B2(\gpio_configure[23][4] ),
    .C1(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__a32o_1 _6558_ (.A1(\gpio_configure[20][4] ),
    .A2(_2663_),
    .A3(net430),
    .B1(_3066_),
    .B2(\gpio_configure[28][4] ),
    .X(_3154_));
 sky130_fd_sc_hd__a221o_1 _6559_ (.A1(\gpio_configure[5][4] ),
    .A2(_3021_),
    .B1(_3062_),
    .B2(\gpio_configure[10][4] ),
    .C1(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__a2111oi_4 _6560_ (.A1(\gpio_configure[12][4] ),
    .A2(_3005_),
    .B1(_3151_),
    .C1(_3153_),
    .D1(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__a32o_1 _6561_ (.A1(\gpio_configure[11][4] ),
    .A2(net434),
    .A3(_3029_),
    .B1(_3068_),
    .B2(\gpio_configure[16][4] ),
    .X(_3157_));
 sky130_fd_sc_hd__a221o_1 _6562_ (.A1(\gpio_configure[4][4] ),
    .A2(_3018_),
    .B1(_3051_),
    .B2(\gpio_configure[25][4] ),
    .C1(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__a32o_1 _6563_ (.A1(\gpio_configure[24][4] ),
    .A2(_2663_),
    .A3(_3041_),
    .B1(_3025_),
    .B2(\gpio_configure[7][4] ),
    .X(_3159_));
 sky130_fd_sc_hd__a221o_1 _6564_ (.A1(\gpio_configure[2][4] ),
    .A2(_3012_),
    .B1(_3054_),
    .B2(\gpio_configure[26][4] ),
    .C1(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__a22o_1 _6565_ (.A1(\gpio_configure[3][4] ),
    .A2(_3013_),
    .B1(_3022_),
    .B2(\gpio_configure[1][4] ),
    .X(_3161_));
 sky130_fd_sc_hd__a221o_1 _6566_ (.A1(\gpio_configure[34][4] ),
    .A2(_3003_),
    .B1(_3007_),
    .B2(\gpio_configure[32][4] ),
    .C1(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__a32o_1 _6567_ (.A1(\gpio_configure[27][4] ),
    .A2(net440),
    .A3(_3029_),
    .B1(_3055_),
    .B2(\gpio_configure[22][4] ),
    .X(_3163_));
 sky130_fd_sc_hd__a221o_1 _6568_ (.A1(\gpio_configure[33][4] ),
    .A2(_3015_),
    .B1(_3035_),
    .B2(\gpio_configure[29][4] ),
    .C1(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__nor4_2 _6569_ (.A(_3158_),
    .B(_3160_),
    .C(_3162_),
    .D(_3164_),
    .Y(_3165_));
 sky130_fd_sc_hd__nand3b_4 _6570_ (.A_N(_3150_),
    .B(_3156_),
    .C(_3165_),
    .Y(_3166_));
 sky130_fd_sc_hd__o21a_1 _6571_ (.A1(\gpio_configure[0][4] ),
    .A2(_3031_),
    .B1(_0824_),
    .X(_3167_));
 sky130_fd_sc_hd__a22o_1 _6572_ (.A1(net528),
    .A2(net3826),
    .B1(_3166_),
    .B2(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_1 _6573_ (.A0(_3168_),
    .A1(net3833),
    .S(_2681_),
    .X(_0788_));
 sky130_fd_sc_hd__and3_1 _6574_ (.A(\gpio_configure[20][5] ),
    .B(net441),
    .C(_3033_),
    .X(_3169_));
 sky130_fd_sc_hd__a32o_1 _6575_ (.A1(\gpio_configure[9][5] ),
    .A2(net433),
    .A3(_3028_),
    .B1(_3062_),
    .B2(\gpio_configure[10][5] ),
    .X(_3170_));
 sky130_fd_sc_hd__a221o_1 _6576_ (.A1(\gpio_configure[12][5] ),
    .A2(_3005_),
    .B1(_3023_),
    .B2(\gpio_configure[6][5] ),
    .C1(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__a32o_1 _6577_ (.A1(\gpio_configure[25][5] ),
    .A2(net440),
    .A3(_3028_),
    .B1(_3021_),
    .B2(\gpio_configure[5][5] ),
    .X(_3172_));
 sky130_fd_sc_hd__a31o_1 _6578_ (.A1(\gpio_configure[13][5] ),
    .A2(net433),
    .A3(_3026_),
    .B1(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__a32o_1 _6579_ (.A1(\gpio_configure[11][5] ),
    .A2(net433),
    .A3(net431),
    .B1(_2674_),
    .B2(\gpio_configure[31][5] ),
    .X(_3174_));
 sky130_fd_sc_hd__a221o_1 _6580_ (.A1(\gpio_configure[1][5] ),
    .A2(_3022_),
    .B1(_3057_),
    .B2(\gpio_configure[24][5] ),
    .C1(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__a221o_1 _6581_ (.A1(\gpio_configure[7][5] ),
    .A2(_3025_),
    .B1(_3054_),
    .B2(\gpio_configure[26][5] ),
    .C1(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__a221o_1 _6582_ (.A1(\gpio_configure[15][5] ),
    .A2(_3009_),
    .B1(_3013_),
    .B2(\gpio_configure[3][5] ),
    .C1(_3176_),
    .X(_3177_));
 sky130_fd_sc_hd__a32o_1 _6583_ (.A1(\gpio_configure[19][5] ),
    .A2(_2673_),
    .A3(_3002_),
    .B1(_3003_),
    .B2(\gpio_configure[34][5] ),
    .X(_3178_));
 sky130_fd_sc_hd__a31o_1 _6584_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][5] ),
    .A3(_3006_),
    .B1(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__a221o_4 _6585_ (.A1(\gpio_configure[4][5] ),
    .A2(_3018_),
    .B1(_3024_),
    .B2(\gpio_configure[36][5] ),
    .C1(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__a211o_1 _6586_ (.A1(\gpio_configure[32][5] ),
    .A2(_3007_),
    .B1(_3177_),
    .C1(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__a2111o_1 _6587_ (.A1(\gpio_configure[2][5] ),
    .A2(_3012_),
    .B1(_3171_),
    .C1(_3173_),
    .D1(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__a32o_1 _6588_ (.A1(\gpio_configure[22][5] ),
    .A2(_1438_),
    .A3(net430),
    .B1(_3063_),
    .B2(\gpio_configure[18][5] ),
    .X(_3183_));
 sky130_fd_sc_hd__a32o_1 _6589_ (.A1(\gpio_configure[27][5] ),
    .A2(net439),
    .A3(net431),
    .B1(_3068_),
    .B2(\gpio_configure[16][5] ),
    .X(_3184_));
 sky130_fd_sc_hd__a221o_1 _6590_ (.A1(\gpio_configure[8][5] ),
    .A2(_3052_),
    .B1(_3067_),
    .B2(\gpio_configure[17][5] ),
    .C1(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__a221o_1 _6591_ (.A1(\gpio_configure[21][5] ),
    .A2(_3043_),
    .B1(_3046_),
    .B2(\gpio_configure[30][5] ),
    .C1(_3169_),
    .X(_3186_));
 sky130_fd_sc_hd__a32o_1 _6592_ (.A1(\gpio_configure[23][5] ),
    .A2(_2662_),
    .A3(_3033_),
    .B1(_3066_),
    .B2(\gpio_configure[28][5] ),
    .X(_3187_));
 sky130_fd_sc_hd__a221o_1 _6593_ (.A1(\gpio_configure[33][5] ),
    .A2(_3015_),
    .B1(_3017_),
    .B2(\gpio_configure[35][5] ),
    .C1(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__a211o_4 _6594_ (.A1(\gpio_configure[29][5] ),
    .A2(_3035_),
    .B1(_3186_),
    .C1(_3188_),
    .X(_3189_));
 sky130_fd_sc_hd__a2111o_1 _6595_ (.A1(\gpio_configure[14][5] ),
    .A2(_3014_),
    .B1(_3183_),
    .C1(_3185_),
    .D1(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__o21a_1 _6596_ (.A1(\gpio_configure[0][5] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3191_));
 sky130_fd_sc_hd__o31a_1 _6597_ (.A1(_3190_),
    .A2(_3030_),
    .A3(_3182_),
    .B1(_3191_),
    .X(_3192_));
 sky130_fd_sc_hd__a211o_1 _6598_ (.A1(net528),
    .A2(net3833),
    .B1(net353),
    .C1(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__o31a_1 _6599_ (.A1(net3863),
    .A2(_1446_),
    .A3(_2680_),
    .B1(_3193_),
    .X(_0789_));
 sky130_fd_sc_hd__and3_1 _6600_ (.A(\gpio_configure[27][6] ),
    .B(net439),
    .C(net431),
    .X(_3194_));
 sky130_fd_sc_hd__a22o_1 _6601_ (.A1(\gpio_configure[29][6] ),
    .A2(_3035_),
    .B1(_3046_),
    .B2(\gpio_configure[30][6] ),
    .X(_3195_));
 sky130_fd_sc_hd__a22o_1 _6602_ (.A1(\gpio_configure[8][6] ),
    .A2(_3052_),
    .B1(_3063_),
    .B2(\gpio_configure[18][6] ),
    .X(_3196_));
 sky130_fd_sc_hd__a32o_1 _6603_ (.A1(\gpio_configure[24][6] ),
    .A2(net441),
    .A3(_3041_),
    .B1(_2674_),
    .B2(\gpio_configure[31][6] ),
    .X(_3197_));
 sky130_fd_sc_hd__a31o_1 _6604_ (.A1(\gpio_configure[11][6] ),
    .A2(net433),
    .A3(net431),
    .B1(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__a32o_1 _6605_ (.A1(\gpio_configure[26][6] ),
    .A2(_1438_),
    .A3(_3041_),
    .B1(_3009_),
    .B2(\gpio_configure[15][6] ),
    .X(_3199_));
 sky130_fd_sc_hd__a221o_1 _6606_ (.A1(\gpio_configure[3][6] ),
    .A2(_3013_),
    .B1(_3025_),
    .B2(\gpio_configure[7][6] ),
    .C1(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__a32o_1 _6607_ (.A1(\gpio_configure[9][6] ),
    .A2(net433),
    .A3(_3028_),
    .B1(_3005_),
    .B2(\gpio_configure[12][6] ),
    .X(_3201_));
 sky130_fd_sc_hd__a32o_1 _6608_ (.A1(\gpio_configure[13][6] ),
    .A2(net433),
    .A3(_3026_),
    .B1(_3051_),
    .B2(\gpio_configure[25][6] ),
    .X(_3202_));
 sky130_fd_sc_hd__a221o_1 _6609_ (.A1(\gpio_configure[2][6] ),
    .A2(_3012_),
    .B1(_3021_),
    .B2(\gpio_configure[5][6] ),
    .C1(_3202_),
    .X(_3203_));
 sky130_fd_sc_hd__a211o_1 _6610_ (.A1(\gpio_configure[10][6] ),
    .A2(_3062_),
    .B1(_3201_),
    .C1(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__a32o_1 _6611_ (.A1(\gpio_configure[19][6] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3003_),
    .B2(\gpio_configure[34][6] ),
    .X(_3205_));
 sky130_fd_sc_hd__a31o_1 _6612_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][6] ),
    .A3(_3006_),
    .B1(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__a221o_1 _6613_ (.A1(\gpio_configure[4][6] ),
    .A2(_3018_),
    .B1(_3024_),
    .B2(\gpio_configure[36][6] ),
    .C1(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__a41o_1 _6614_ (.A1(\gpio_configure[32][6] ),
    .A2(_1439_),
    .A3(net441),
    .A4(net435),
    .B1(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__a2111o_1 _6615_ (.A1(\gpio_configure[6][6] ),
    .A2(_3023_),
    .B1(_3200_),
    .C1(_3204_),
    .D1(_3208_),
    .X(_3209_));
 sky130_fd_sc_hd__a32o_1 _6616_ (.A1(\gpio_configure[20][6] ),
    .A2(net441),
    .A3(net430),
    .B1(_3043_),
    .B2(\gpio_configure[21][6] ),
    .X(_3210_));
 sky130_fd_sc_hd__a221o_1 _6617_ (.A1(\gpio_configure[35][6] ),
    .A2(_3017_),
    .B1(_3066_),
    .B2(\gpio_configure[28][6] ),
    .C1(_3195_),
    .X(_3211_));
 sky130_fd_sc_hd__a221o_1 _6618_ (.A1(\gpio_configure[33][6] ),
    .A2(_3015_),
    .B1(_3055_),
    .B2(\gpio_configure[22][6] ),
    .C1(_3196_),
    .X(_3212_));
 sky130_fd_sc_hd__a221o_1 _6619_ (.A1(\gpio_configure[14][6] ),
    .A2(_3014_),
    .B1(_3067_),
    .B2(\gpio_configure[17][6] ),
    .C1(_3194_),
    .X(_3213_));
 sky130_fd_sc_hd__a2111o_1 _6620_ (.A1(\gpio_configure[16][6] ),
    .A2(_3068_),
    .B1(_3212_),
    .C1(_3213_),
    .D1(_3030_),
    .X(_3214_));
 sky130_fd_sc_hd__a2111o_1 _6621_ (.A1(\gpio_configure[23][6] ),
    .A2(_3034_),
    .B1(_3210_),
    .C1(_3211_),
    .D1(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__a2111o_2 _6622_ (.A1(\gpio_configure[1][6] ),
    .A2(_3022_),
    .B1(_3198_),
    .C1(_3209_),
    .D1(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__o21a_1 _6623_ (.A1(\gpio_configure[0][6] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3217_));
 sky130_fd_sc_hd__a22o_1 _6624_ (.A1(net528),
    .A2(\serial_data_staging_2[5] ),
    .B1(_3216_),
    .B2(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__mux2_1 _6625_ (.A0(_3218_),
    .A1(net3835),
    .S(net353),
    .X(_0790_));
 sky130_fd_sc_hd__a22o_1 _6626_ (.A1(\gpio_configure[31][7] ),
    .A2(_2674_),
    .B1(_3009_),
    .B2(\gpio_configure[15][7] ),
    .X(_3219_));
 sky130_fd_sc_hd__a32o_1 _6627_ (.A1(\gpio_configure[9][7] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3005_),
    .B2(\gpio_configure[12][7] ),
    .X(_3220_));
 sky130_fd_sc_hd__a221o_1 _6628_ (.A1(\gpio_configure[3][7] ),
    .A2(_3013_),
    .B1(_3063_),
    .B2(\gpio_configure[18][7] ),
    .C1(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__a22o_1 _6629_ (.A1(\gpio_configure[32][7] ),
    .A2(_3007_),
    .B1(_3035_),
    .B2(\gpio_configure[29][7] ),
    .X(_3222_));
 sky130_fd_sc_hd__a211o_1 _6630_ (.A1(\gpio_configure[36][7] ),
    .A2(_3024_),
    .B1(_3221_),
    .C1(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__a2111oi_4 _6631_ (.A1(\gpio_configure[37][7] ),
    .A2(_3027_),
    .B1(_3219_),
    .C1(_3223_),
    .D1(_3030_),
    .Y(_3224_));
 sky130_fd_sc_hd__a22o_1 _6632_ (.A1(\gpio_configure[34][7] ),
    .A2(_3003_),
    .B1(_3018_),
    .B2(\gpio_configure[4][7] ),
    .X(_3225_));
 sky130_fd_sc_hd__a32o_1 _6633_ (.A1(\gpio_configure[11][7] ),
    .A2(_3004_),
    .A3(net431),
    .B1(_3022_),
    .B2(\gpio_configure[1][7] ),
    .X(_3226_));
 sky130_fd_sc_hd__a221o_1 _6634_ (.A1(\gpio_configure[6][7] ),
    .A2(_3023_),
    .B1(_3054_),
    .B2(\gpio_configure[26][7] ),
    .C1(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__a22o_1 _6635_ (.A1(\gpio_configure[7][7] ),
    .A2(_3025_),
    .B1(_3060_),
    .B2(\gpio_configure[13][7] ),
    .X(_3228_));
 sky130_fd_sc_hd__a221o_1 _6636_ (.A1(\gpio_configure[30][7] ),
    .A2(_3046_),
    .B1(_3066_),
    .B2(\gpio_configure[28][7] ),
    .C1(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__a2111o_1 _6637_ (.A1(\gpio_configure[2][7] ),
    .A2(_3012_),
    .B1(_3225_),
    .C1(_3227_),
    .D1(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__a32o_1 _6638_ (.A1(\gpio_configure[24][7] ),
    .A2(_2663_),
    .A3(_3041_),
    .B1(_3043_),
    .B2(\gpio_configure[21][7] ),
    .X(_3231_));
 sky130_fd_sc_hd__a221o_1 _6639_ (.A1(\gpio_configure[8][7] ),
    .A2(_3052_),
    .B1(_3068_),
    .B2(\gpio_configure[16][7] ),
    .C1(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__a32o_1 _6640_ (.A1(\gpio_configure[20][7] ),
    .A2(_2663_),
    .A3(net430),
    .B1(_3034_),
    .B2(\gpio_configure[23][7] ),
    .X(_3233_));
 sky130_fd_sc_hd__a221o_1 _6641_ (.A1(\gpio_configure[5][7] ),
    .A2(_3021_),
    .B1(_3062_),
    .B2(\gpio_configure[10][7] ),
    .C1(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__a32o_1 _6642_ (.A1(\gpio_configure[25][7] ),
    .A2(net440),
    .A3(_3028_),
    .B1(_3017_),
    .B2(\gpio_configure[35][7] ),
    .X(_3235_));
 sky130_fd_sc_hd__a221o_1 _6643_ (.A1(\gpio_configure[33][7] ),
    .A2(_3015_),
    .B1(_3067_),
    .B2(\gpio_configure[17][7] ),
    .C1(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__a32o_1 _6644_ (.A1(\gpio_configure[27][7] ),
    .A2(net440),
    .A3(_3029_),
    .B1(_3014_),
    .B2(\gpio_configure[14][7] ),
    .X(_3237_));
 sky130_fd_sc_hd__and3_1 _6645_ (.A(\gpio_configure[19][7] ),
    .B(_2673_),
    .C(_3002_),
    .X(_3238_));
 sky130_fd_sc_hd__a2111o_1 _6646_ (.A1(\gpio_configure[22][7] ),
    .A2(_3055_),
    .B1(_3238_),
    .C1(_3237_),
    .D1(_3236_),
    .X(_3239_));
 sky130_fd_sc_hd__nor4_1 _6647_ (.A(_3230_),
    .B(_3232_),
    .C(_3234_),
    .D(_3239_),
    .Y(_3240_));
 sky130_fd_sc_hd__o2bb2a_1 _6648_ (.A1_N(_3224_),
    .A2_N(net347),
    .B1(\gpio_configure[0][7] ),
    .B2(_3031_),
    .X(_3241_));
 sky130_fd_sc_hd__mux2_1 _6649_ (.A0(_3241_),
    .A1(net3835),
    .S(net528),
    .X(_3242_));
 sky130_fd_sc_hd__mux2_1 _6650_ (.A0(_3242_),
    .A1(net3850),
    .S(net353),
    .X(_0791_));
 sky130_fd_sc_hd__and3_1 _6651_ (.A(\gpio_configure[11][8] ),
    .B(net432),
    .C(net431),
    .X(_3243_));
 sky130_fd_sc_hd__a22o_1 _6652_ (.A1(\gpio_configure[35][8] ),
    .A2(_3017_),
    .B1(_3046_),
    .B2(\gpio_configure[30][8] ),
    .X(_3244_));
 sky130_fd_sc_hd__a221o_1 _6653_ (.A1(\gpio_configure[29][8] ),
    .A2(_3035_),
    .B1(_3043_),
    .B2(\gpio_configure[21][8] ),
    .C1(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__a221o_1 _6654_ (.A1(\gpio_configure[23][8] ),
    .A2(_3034_),
    .B1(_3066_),
    .B2(\gpio_configure[28][8] ),
    .C1(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__a32o_1 _6655_ (.A1(\gpio_configure[26][8] ),
    .A2(_1438_),
    .A3(_3041_),
    .B1(_3025_),
    .B2(\gpio_configure[7][8] ),
    .X(_3247_));
 sky130_fd_sc_hd__a221o_1 _6656_ (.A1(\gpio_configure[31][8] ),
    .A2(_2674_),
    .B1(_3057_),
    .B2(\gpio_configure[24][8] ),
    .C1(_3243_),
    .X(_3248_));
 sky130_fd_sc_hd__a221o_1 _6657_ (.A1(\gpio_configure[15][8] ),
    .A2(_3009_),
    .B1(_3013_),
    .B2(\gpio_configure[3][8] ),
    .C1(_3247_),
    .X(_3249_));
 sky130_fd_sc_hd__a32o_1 _6658_ (.A1(\gpio_configure[9][8] ),
    .A2(net432),
    .A3(_3028_),
    .B1(_3005_),
    .B2(\gpio_configure[12][8] ),
    .X(_3250_));
 sky130_fd_sc_hd__a221o_1 _6659_ (.A1(\gpio_configure[6][8] ),
    .A2(_3023_),
    .B1(_3062_),
    .B2(\gpio_configure[10][8] ),
    .C1(_3250_),
    .X(_3251_));
 sky130_fd_sc_hd__a31o_1 _6660_ (.A1(\gpio_configure[13][8] ),
    .A2(net432),
    .A3(_3026_),
    .B1(_3251_),
    .X(_3252_));
 sky130_fd_sc_hd__a221o_1 _6661_ (.A1(\gpio_configure[2][8] ),
    .A2(_3012_),
    .B1(_3021_),
    .B2(\gpio_configure[5][8] ),
    .C1(_3252_),
    .X(_3253_));
 sky130_fd_sc_hd__a31o_1 _6662_ (.A1(\gpio_configure[25][8] ),
    .A2(net440),
    .A3(_3028_),
    .B1(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__a32o_1 _6663_ (.A1(\gpio_configure[19][8] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3003_),
    .B2(\gpio_configure[34][8] ),
    .X(_3255_));
 sky130_fd_sc_hd__a31o_1 _6664_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][8] ),
    .A3(_3006_),
    .B1(_3255_),
    .X(_3256_));
 sky130_fd_sc_hd__a221o_4 _6665_ (.A1(\gpio_configure[4][8] ),
    .A2(_3018_),
    .B1(_3024_),
    .B2(\gpio_configure[36][8] ),
    .C1(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__a2111o_1 _6666_ (.A1(\gpio_configure[32][8] ),
    .A2(_3007_),
    .B1(_3249_),
    .C1(_3254_),
    .D1(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__a32o_1 _6667_ (.A1(\gpio_configure[22][8] ),
    .A2(_1438_),
    .A3(net430),
    .B1(_3063_),
    .B2(\gpio_configure[18][8] ),
    .X(_3259_));
 sky130_fd_sc_hd__a32o_1 _6668_ (.A1(\gpio_configure[27][8] ),
    .A2(net439),
    .A3(net431),
    .B1(_3052_),
    .B2(\gpio_configure[8][8] ),
    .X(_3260_));
 sky130_fd_sc_hd__a221o_1 _6669_ (.A1(\gpio_configure[14][8] ),
    .A2(_3014_),
    .B1(_3067_),
    .B2(\gpio_configure[17][8] ),
    .C1(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__a211o_1 _6670_ (.A1(\gpio_configure[16][8] ),
    .A2(_3068_),
    .B1(_3259_),
    .C1(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__a211o_1 _6671_ (.A1(\gpio_configure[33][8] ),
    .A2(_3015_),
    .B1(_3262_),
    .C1(_3030_),
    .X(_3263_));
 sky130_fd_sc_hd__a2111o_1 _6672_ (.A1(\gpio_configure[1][8] ),
    .A2(_3022_),
    .B1(_3248_),
    .C1(_3258_),
    .D1(_3263_),
    .X(_3264_));
 sky130_fd_sc_hd__a311o_2 _6673_ (.A1(\gpio_configure[20][8] ),
    .A2(net441),
    .A3(net430),
    .B1(_3246_),
    .C1(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__o21a_1 _6674_ (.A1(\gpio_configure[0][8] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3266_));
 sky130_fd_sc_hd__a22o_1 _6675_ (.A1(net528),
    .A2(net3850),
    .B1(_3265_),
    .B2(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(_3267_),
    .A1(net3851),
    .S(net353),
    .X(_0792_));
 sky130_fd_sc_hd__a22o_1 _6677_ (.A1(\gpio_configure[31][9] ),
    .A2(_2674_),
    .B1(_3009_),
    .B2(\gpio_configure[15][9] ),
    .X(_3268_));
 sky130_fd_sc_hd__a32o_1 _6678_ (.A1(\gpio_configure[11][9] ),
    .A2(net434),
    .A3(net431),
    .B1(_3023_),
    .B2(\gpio_configure[6][9] ),
    .X(_3269_));
 sky130_fd_sc_hd__a221o_1 _6679_ (.A1(\gpio_configure[34][9] ),
    .A2(_3003_),
    .B1(_3051_),
    .B2(\gpio_configure[25][9] ),
    .C1(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__a32o_1 _6680_ (.A1(\gpio_configure[23][9] ),
    .A2(_2662_),
    .A3(net430),
    .B1(_3063_),
    .B2(\gpio_configure[18][9] ),
    .X(_3271_));
 sky130_fd_sc_hd__a211o_1 _6681_ (.A1(\gpio_configure[37][9] ),
    .A2(_3027_),
    .B1(_3270_),
    .C1(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__a2111o_1 _6682_ (.A1(\gpio_configure[36][9] ),
    .A2(_3024_),
    .B1(_3268_),
    .C1(_3272_),
    .D1(_3030_),
    .X(_3273_));
 sky130_fd_sc_hd__a32o_1 _6683_ (.A1(\gpio_configure[27][9] ),
    .A2(net440),
    .A3(net431),
    .B1(_3047_),
    .B2(\gpio_configure[20][9] ),
    .X(_3274_));
 sky130_fd_sc_hd__a32o_1 _6684_ (.A1(\gpio_configure[9][9] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3060_),
    .B2(\gpio_configure[13][9] ),
    .X(_3275_));
 sky130_fd_sc_hd__a221o_2 _6685_ (.A1(\gpio_configure[12][9] ),
    .A2(_3005_),
    .B1(_3062_),
    .B2(\gpio_configure[10][9] ),
    .C1(_3275_),
    .X(_3276_));
 sky130_fd_sc_hd__a32o_1 _6686_ (.A1(\gpio_configure[19][9] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3025_),
    .B2(\gpio_configure[7][9] ),
    .X(_3277_));
 sky130_fd_sc_hd__a221o_2 _6687_ (.A1(\gpio_configure[2][9] ),
    .A2(_3012_),
    .B1(_3057_),
    .B2(\gpio_configure[24][9] ),
    .C1(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__a2111oi_4 _6688_ (.A1(\gpio_configure[17][9] ),
    .A2(_3067_),
    .B1(_3274_),
    .C1(_3276_),
    .D1(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__a32o_1 _6689_ (.A1(\gpio_configure[22][9] ),
    .A2(_1438_),
    .A3(net430),
    .B1(_3007_),
    .B2(\gpio_configure[32][9] ),
    .X(_3280_));
 sky130_fd_sc_hd__a221o_1 _6690_ (.A1(\gpio_configure[21][9] ),
    .A2(_3043_),
    .B1(_3068_),
    .B2(\gpio_configure[16][9] ),
    .C1(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__a22o_1 _6691_ (.A1(\gpio_configure[4][9] ),
    .A2(_3018_),
    .B1(_3021_),
    .B2(\gpio_configure[5][9] ),
    .X(_3282_));
 sky130_fd_sc_hd__a221o_1 _6692_ (.A1(\gpio_configure[14][9] ),
    .A2(_3014_),
    .B1(_3015_),
    .B2(\gpio_configure[33][9] ),
    .C1(_3282_),
    .X(_3283_));
 sky130_fd_sc_hd__a32o_1 _6693_ (.A1(\gpio_configure[26][9] ),
    .A2(_1438_),
    .A3(_3041_),
    .B1(_3066_),
    .B2(\gpio_configure[28][9] ),
    .X(_3284_));
 sky130_fd_sc_hd__a221o_1 _6694_ (.A1(\gpio_configure[29][9] ),
    .A2(_3035_),
    .B1(_3052_),
    .B2(\gpio_configure[8][9] ),
    .C1(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__a22o_1 _6695_ (.A1(\gpio_configure[35][9] ),
    .A2(_3017_),
    .B1(_3046_),
    .B2(\gpio_configure[30][9] ),
    .X(_3286_));
 sky130_fd_sc_hd__a221o_1 _6696_ (.A1(\gpio_configure[3][9] ),
    .A2(_3013_),
    .B1(_3022_),
    .B2(\gpio_configure[1][9] ),
    .C1(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__nor4_2 _6697_ (.A(_3281_),
    .B(_3283_),
    .C(_3285_),
    .D(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__nand3b_4 _6698_ (.A_N(_3273_),
    .B(_3279_),
    .C(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__o21a_1 _6699_ (.A1(\gpio_configure[0][9] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3290_));
 sky130_fd_sc_hd__a22o_1 _6700_ (.A1(net528),
    .A2(\serial_data_staging_2[8] ),
    .B1(_3289_),
    .B2(_3290_),
    .X(_3291_));
 sky130_fd_sc_hd__mux2_1 _6701_ (.A0(_3291_),
    .A1(net3814),
    .S(net353),
    .X(_0793_));
 sky130_fd_sc_hd__and3_1 _6702_ (.A(\gpio_configure[19][10] ),
    .B(_2673_),
    .C(net435),
    .X(_3292_));
 sky130_fd_sc_hd__a32o_1 _6703_ (.A1(\gpio_configure[25][10] ),
    .A2(net439),
    .A3(_3028_),
    .B1(_3021_),
    .B2(\gpio_configure[5][10] ),
    .X(_3293_));
 sky130_fd_sc_hd__a31o_1 _6704_ (.A1(\gpio_configure[13][10] ),
    .A2(net432),
    .A3(_3026_),
    .B1(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__a32o_1 _6705_ (.A1(\gpio_configure[9][10] ),
    .A2(net432),
    .A3(_3028_),
    .B1(_3005_),
    .B2(\gpio_configure[12][10] ),
    .X(_3295_));
 sky130_fd_sc_hd__a221o_1 _6706_ (.A1(\gpio_configure[6][10] ),
    .A2(_3023_),
    .B1(_3062_),
    .B2(\gpio_configure[10][10] ),
    .C1(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__a32o_1 _6707_ (.A1(\gpio_configure[24][10] ),
    .A2(net441),
    .A3(_3041_),
    .B1(_2674_),
    .B2(\gpio_configure[31][10] ),
    .X(_3297_));
 sky130_fd_sc_hd__a31o_1 _6708_ (.A1(\gpio_configure[11][10] ),
    .A2(net432),
    .A3(net431),
    .B1(_3297_),
    .X(_3298_));
 sky130_fd_sc_hd__a221o_1 _6709_ (.A1(\gpio_configure[15][10] ),
    .A2(_3009_),
    .B1(_3022_),
    .B2(\gpio_configure[1][10] ),
    .C1(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__a221o_1 _6710_ (.A1(\gpio_configure[7][10] ),
    .A2(_3025_),
    .B1(_3054_),
    .B2(\gpio_configure[26][10] ),
    .C1(_3299_),
    .X(_3300_));
 sky130_fd_sc_hd__a221o_2 _6711_ (.A1(\gpio_configure[34][10] ),
    .A2(_3003_),
    .B1(_3024_),
    .B2(\gpio_configure[36][10] ),
    .C1(_3292_),
    .X(_3301_));
 sky130_fd_sc_hd__a221o_4 _6712_ (.A1(\gpio_configure[32][10] ),
    .A2(_3007_),
    .B1(_3027_),
    .B2(\gpio_configure[37][10] ),
    .C1(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__a41o_1 _6713_ (.A1(\gpio_configure[4][10] ),
    .A2(_1440_),
    .A3(net441),
    .A4(net432),
    .B1(_3302_),
    .X(_3303_));
 sky130_fd_sc_hd__a2111o_1 _6714_ (.A1(\gpio_configure[3][10] ),
    .A2(_3013_),
    .B1(_3296_),
    .C1(_3300_),
    .D1(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__a211o_1 _6715_ (.A1(\gpio_configure[2][10] ),
    .A2(_3012_),
    .B1(_3294_),
    .C1(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__a32o_1 _6716_ (.A1(\gpio_configure[23][10] ),
    .A2(_2662_),
    .A3(net430),
    .B1(_3066_),
    .B2(\gpio_configure[28][10] ),
    .X(_3306_));
 sky130_fd_sc_hd__a221o_1 _6717_ (.A1(\gpio_configure[33][10] ),
    .A2(_3015_),
    .B1(_3017_),
    .B2(\gpio_configure[35][10] ),
    .C1(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__a32o_1 _6718_ (.A1(\gpio_configure[20][10] ),
    .A2(net441),
    .A3(net430),
    .B1(_3043_),
    .B2(\gpio_configure[21][10] ),
    .X(_3308_));
 sky130_fd_sc_hd__a221o_1 _6719_ (.A1(\gpio_configure[29][10] ),
    .A2(_3035_),
    .B1(_3046_),
    .B2(\gpio_configure[30][10] ),
    .C1(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__a32o_1 _6720_ (.A1(\gpio_configure[22][10] ),
    .A2(_1438_),
    .A3(net430),
    .B1(_3063_),
    .B2(\gpio_configure[18][10] ),
    .X(_3310_));
 sky130_fd_sc_hd__a32o_1 _6721_ (.A1(\gpio_configure[27][10] ),
    .A2(net439),
    .A3(net431),
    .B1(_3052_),
    .B2(\gpio_configure[8][10] ),
    .X(_3311_));
 sky130_fd_sc_hd__a221o_1 _6722_ (.A1(\gpio_configure[14][10] ),
    .A2(_3014_),
    .B1(_3067_),
    .B2(\gpio_configure[17][10] ),
    .C1(_3311_),
    .X(_3312_));
 sky130_fd_sc_hd__a2111o_1 _6723_ (.A1(\gpio_configure[16][10] ),
    .A2(_3068_),
    .B1(_3309_),
    .C1(_3310_),
    .D1(_3312_),
    .X(_3313_));
 sky130_fd_sc_hd__a31o_1 _6724_ (.A1(_3008_),
    .A2(net393),
    .A3(_3020_),
    .B1(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__o32a_1 _6725_ (.A1(_3305_),
    .A2(_3307_),
    .A3(_3314_),
    .B1(_3031_),
    .B2(\gpio_configure[0][10] ),
    .X(_3315_));
 sky130_fd_sc_hd__mux2_1 _6726_ (.A0(_3315_),
    .A1(net3814),
    .S(net527),
    .X(_3316_));
 sky130_fd_sc_hd__mux2_1 _6727_ (.A0(_3316_),
    .A1(net3825),
    .S(net353),
    .X(_0794_));
 sky130_fd_sc_hd__a32o_1 _6728_ (.A1(\pad_count_2[0] ),
    .A2(\gpio_configure[37][11] ),
    .A3(_3006_),
    .B1(_3009_),
    .B2(\gpio_configure[15][11] ),
    .X(_3317_));
 sky130_fd_sc_hd__a32o_1 _6729_ (.A1(\gpio_configure[6][11] ),
    .A2(_1441_),
    .A3(net434),
    .B1(_3022_),
    .B2(\gpio_configure[1][11] ),
    .X(_3318_));
 sky130_fd_sc_hd__a221o_1 _6730_ (.A1(\gpio_configure[34][11] ),
    .A2(_3003_),
    .B1(_3012_),
    .B2(\gpio_configure[2][11] ),
    .C1(_3318_),
    .X(_3319_));
 sky130_fd_sc_hd__a22o_1 _6731_ (.A1(\gpio_configure[4][11] ),
    .A2(_3018_),
    .B1(_3046_),
    .B2(\gpio_configure[30][11] ),
    .X(_3320_));
 sky130_fd_sc_hd__a211o_1 _6732_ (.A1(\gpio_configure[36][11] ),
    .A2(_3024_),
    .B1(_3319_),
    .C1(_3320_),
    .X(_3321_));
 sky130_fd_sc_hd__a2111oi_2 _6733_ (.A1(\gpio_configure[31][11] ),
    .A2(_2674_),
    .B1(_3317_),
    .C1(_3321_),
    .D1(_3030_),
    .Y(_3322_));
 sky130_fd_sc_hd__a32o_1 _6734_ (.A1(\gpio_configure[23][11] ),
    .A2(_2662_),
    .A3(net430),
    .B1(_3014_),
    .B2(\gpio_configure[14][11] ),
    .X(_3323_));
 sky130_fd_sc_hd__a32o_1 _6735_ (.A1(\gpio_configure[9][11] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3051_),
    .B2(\gpio_configure[25][11] ),
    .X(_3324_));
 sky130_fd_sc_hd__a221o_1 _6736_ (.A1(\gpio_configure[12][11] ),
    .A2(_3005_),
    .B1(_3060_),
    .B2(\gpio_configure[13][11] ),
    .C1(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__a22o_1 _6737_ (.A1(\gpio_configure[3][11] ),
    .A2(_3013_),
    .B1(_3062_),
    .B2(\gpio_configure[10][11] ),
    .X(_3326_));
 sky130_fd_sc_hd__a221o_1 _6738_ (.A1(\gpio_configure[7][11] ),
    .A2(_3025_),
    .B1(_3057_),
    .B2(\gpio_configure[24][11] ),
    .C1(_3326_),
    .X(_3327_));
 sky130_fd_sc_hd__a2111o_2 _6739_ (.A1(\gpio_configure[16][11] ),
    .A2(_3068_),
    .B1(_3323_),
    .C1(_3325_),
    .D1(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__a32o_1 _6740_ (.A1(\gpio_configure[27][11] ),
    .A2(net440),
    .A3(net431),
    .B1(_3035_),
    .B2(\gpio_configure[29][11] ),
    .X(_3329_));
 sky130_fd_sc_hd__a221o_1 _6741_ (.A1(\gpio_configure[33][11] ),
    .A2(_3015_),
    .B1(_3047_),
    .B2(\gpio_configure[20][11] ),
    .C1(_3329_),
    .X(_3330_));
 sky130_fd_sc_hd__a32o_1 _6742_ (.A1(\gpio_configure[26][11] ),
    .A2(_1438_),
    .A3(_3041_),
    .B1(_3043_),
    .B2(\gpio_configure[21][11] ),
    .X(_3331_));
 sky130_fd_sc_hd__a221o_1 _6743_ (.A1(\gpio_configure[32][11] ),
    .A2(_3007_),
    .B1(_3021_),
    .B2(\gpio_configure[5][11] ),
    .C1(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__a32o_1 _6744_ (.A1(\gpio_configure[22][11] ),
    .A2(_1438_),
    .A3(net430),
    .B1(_3017_),
    .B2(\gpio_configure[35][11] ),
    .X(_3333_));
 sky130_fd_sc_hd__a221o_1 _6745_ (.A1(\gpio_configure[28][11] ),
    .A2(_3066_),
    .B1(_3067_),
    .B2(\gpio_configure[17][11] ),
    .C1(_3333_),
    .X(_3334_));
 sky130_fd_sc_hd__a32o_1 _6746_ (.A1(\gpio_configure[11][11] ),
    .A2(net434),
    .A3(net431),
    .B1(_3063_),
    .B2(\gpio_configure[18][11] ),
    .X(_3335_));
 sky130_fd_sc_hd__and3_1 _6747_ (.A(\gpio_configure[19][11] ),
    .B(_2673_),
    .C(net435),
    .X(_3336_));
 sky130_fd_sc_hd__a2111o_1 _6748_ (.A1(\gpio_configure[8][11] ),
    .A2(_3052_),
    .B1(_3336_),
    .C1(_3335_),
    .D1(_3334_),
    .X(_3337_));
 sky130_fd_sc_hd__nor4_4 _6749_ (.A(_3328_),
    .B(_3330_),
    .C(_3332_),
    .D(_3337_),
    .Y(_3338_));
 sky130_fd_sc_hd__o2bb2a_1 _6750_ (.A1_N(net346),
    .A2_N(_3338_),
    .B1(\gpio_configure[0][11] ),
    .B2(_3031_),
    .X(_3339_));
 sky130_fd_sc_hd__mux2_1 _6751_ (.A0(_3339_),
    .A1(net3825),
    .S(net527),
    .X(_3340_));
 sky130_fd_sc_hd__mux2_1 _6752_ (.A0(_3340_),
    .A1(net3828),
    .S(net353),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _6753_ (.A1(\gpio_configure[36][12] ),
    .A2(_3024_),
    .B1(_3027_),
    .B2(\gpio_configure[37][12] ),
    .X(_3341_));
 sky130_fd_sc_hd__a32o_1 _6754_ (.A1(\gpio_configure[19][12] ),
    .A2(_2673_),
    .A3(net435),
    .B1(_3043_),
    .B2(\gpio_configure[21][12] ),
    .X(_3342_));
 sky130_fd_sc_hd__a221o_1 _6755_ (.A1(\gpio_configure[18][12] ),
    .A2(_3063_),
    .B1(_3066_),
    .B2(\gpio_configure[28][12] ),
    .C1(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__a32o_1 _6756_ (.A1(\gpio_configure[24][12] ),
    .A2(net441),
    .A3(_3041_),
    .B1(_3018_),
    .B2(\gpio_configure[4][12] ),
    .X(_3344_));
 sky130_fd_sc_hd__a211o_1 _6757_ (.A1(\gpio_configure[31][12] ),
    .A2(_2674_),
    .B1(_3343_),
    .C1(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__a2111o_1 _6758_ (.A1(\gpio_configure[15][12] ),
    .A2(_3009_),
    .B1(_3341_),
    .C1(_3345_),
    .D1(_3030_),
    .X(_3346_));
 sky130_fd_sc_hd__a32o_1 _6759_ (.A1(\gpio_configure[6][12] ),
    .A2(_1441_),
    .A3(net434),
    .B1(_3067_),
    .B2(\gpio_configure[17][12] ),
    .X(_3347_));
 sky130_fd_sc_hd__a32o_1 _6760_ (.A1(\gpio_configure[27][12] ),
    .A2(net440),
    .A3(net431),
    .B1(_3015_),
    .B2(\gpio_configure[33][12] ),
    .X(_3348_));
 sky130_fd_sc_hd__a221o_4 _6761_ (.A1(\gpio_configure[30][12] ),
    .A2(_3046_),
    .B1(_3052_),
    .B2(\gpio_configure[8][12] ),
    .C1(_3348_),
    .X(_3349_));
 sky130_fd_sc_hd__a32o_1 _6762_ (.A1(\gpio_configure[20][12] ),
    .A2(net441),
    .A3(net430),
    .B1(_3068_),
    .B2(\gpio_configure[16][12] ),
    .X(_3350_));
 sky130_fd_sc_hd__a221o_1 _6763_ (.A1(\gpio_configure[34][12] ),
    .A2(_3003_),
    .B1(_3035_),
    .B2(\gpio_configure[29][12] ),
    .C1(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__a2111oi_4 _6764_ (.A1(\gpio_configure[25][12] ),
    .A2(_3051_),
    .B1(_3347_),
    .C1(_3349_),
    .D1(_3351_),
    .Y(_3352_));
 sky130_fd_sc_hd__a22o_1 _6765_ (.A1(\gpio_configure[3][12] ),
    .A2(_3013_),
    .B1(_3060_),
    .B2(\gpio_configure[13][12] ),
    .X(_3353_));
 sky130_fd_sc_hd__a221o_1 _6766_ (.A1(\gpio_configure[32][12] ),
    .A2(_3007_),
    .B1(_3054_),
    .B2(\gpio_configure[26][12] ),
    .C1(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__a32o_1 _6767_ (.A1(\gpio_configure[9][12] ),
    .A2(net434),
    .A3(_3028_),
    .B1(_3062_),
    .B2(\gpio_configure[10][12] ),
    .X(_3355_));
 sky130_fd_sc_hd__a221o_1 _6768_ (.A1(\gpio_configure[12][12] ),
    .A2(_3005_),
    .B1(_3025_),
    .B2(\gpio_configure[7][12] ),
    .C1(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__a32o_1 _6769_ (.A1(\gpio_configure[11][12] ),
    .A2(net434),
    .A3(net431),
    .B1(_3021_),
    .B2(\gpio_configure[5][12] ),
    .X(_3357_));
 sky130_fd_sc_hd__a221o_1 _6770_ (.A1(\gpio_configure[14][12] ),
    .A2(_3014_),
    .B1(_3055_),
    .B2(\gpio_configure[22][12] ),
    .C1(_3357_),
    .X(_3358_));
 sky130_fd_sc_hd__a32o_1 _6771_ (.A1(\gpio_configure[23][12] ),
    .A2(_2662_),
    .A3(net430),
    .B1(_3017_),
    .B2(\gpio_configure[35][12] ),
    .X(_3359_));
 sky130_fd_sc_hd__a221o_1 _6772_ (.A1(\gpio_configure[2][12] ),
    .A2(_3012_),
    .B1(_3022_),
    .B2(\gpio_configure[1][12] ),
    .C1(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__nor4_2 _6773_ (.A(_3354_),
    .B(_3356_),
    .C(_3358_),
    .D(_3360_),
    .Y(_3361_));
 sky130_fd_sc_hd__nand3b_4 _6774_ (.A_N(_3346_),
    .B(_3352_),
    .C(_3361_),
    .Y(_3362_));
 sky130_fd_sc_hd__o21a_1 _6775_ (.A1(\gpio_configure[0][12] ),
    .A2(_3031_),
    .B1(net513),
    .X(_3363_));
 sky130_fd_sc_hd__a22o_1 _6776_ (.A1(net527),
    .A2(net3828),
    .B1(_3362_),
    .B2(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__mux2_1 _6777_ (.A0(_3364_),
    .A1(net3865),
    .S(net353),
    .X(_0796_));
 sky130_fd_sc_hd__o41ai_1 _6778_ (.A1(\wbbd_state[0] ),
    .A2(\wbbd_state[1] ),
    .A3(net3854),
    .A4(\wbbd_state[7] ),
    .B1(_1445_),
    .Y(_3365_));
 sky130_fd_sc_hd__a22o_1 _6779_ (.A1(net3810),
    .A2(_1445_),
    .B1(_3365_),
    .B2(net3883),
    .X(_0797_));
 sky130_fd_sc_hd__nand2_8 _6780_ (.A(\wbbd_state[1] ),
    .B(net608),
    .Y(_3366_));
 sky130_fd_sc_hd__nand2_1 _6781_ (.A(_3366_),
    .B(net3539),
    .Y(_3367_));
 sky130_fd_sc_hd__o21ai_1 _6782_ (.A1(_3366_),
    .A2(_1368_),
    .B1(_3367_),
    .Y(_0798_));
 sky130_fd_sc_hd__mux2_1 _6783_ (.A0(_1297_),
    .A1(net3519),
    .S(_3366_),
    .X(_0799_));
 sky130_fd_sc_hd__nand2_1 _6784_ (.A(_3366_),
    .B(net3447),
    .Y(_3368_));
 sky130_fd_sc_hd__o21ai_1 _6785_ (.A1(_3366_),
    .A2(_1231_),
    .B1(_3368_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _6786_ (.A(_3366_),
    .B(net3463),
    .Y(_3369_));
 sky130_fd_sc_hd__o21ai_1 _6787_ (.A1(_3366_),
    .A2(_1171_),
    .B1(_3369_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _6788_ (.A(_3366_),
    .B(net3704),
    .Y(_3370_));
 sky130_fd_sc_hd__o21ai_2 _6789_ (.A1(net3811),
    .A2(clknet_1_0__leaf__1111_),
    .B1(_3370_),
    .Y(_0802_));
 sky130_fd_sc_hd__mux2_1 _6790_ (.A0(_1022_),
    .A1(net3537),
    .S(_3366_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _6791_ (.A0(_0988_),
    .A1(net3492),
    .S(_3366_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _6792_ (.A0(_0953_),
    .A1(net3484),
    .S(_3366_),
    .X(_0805_));
 sky130_fd_sc_hd__a21bo_1 _6793_ (.A1(net170),
    .A2(net165),
    .B1_N(\wbbd_state[6] ),
    .X(_3371_));
 sky130_fd_sc_hd__nand2_1 _6794_ (.A(net168),
    .B(net170),
    .Y(_3372_));
 sky130_fd_sc_hd__nand2_1 _6795_ (.A(net170),
    .B(net167),
    .Y(_3373_));
 sky130_fd_sc_hd__a21bo_1 _6796_ (.A1(net170),
    .A2(net166),
    .B1_N(\wbbd_state[9] ),
    .X(_3374_));
 sky130_fd_sc_hd__a221o_1 _6797_ (.A1(\wbbd_state[10] ),
    .A2(_3372_),
    .B1(_3373_),
    .B2(\wbbd_state[8] ),
    .C1(_1538_),
    .X(_3375_));
 sky130_fd_sc_hd__nand3b_4 _6798_ (.A_N(_3375_),
    .B(_3374_),
    .C(_3371_),
    .Y(_3376_));
 sky130_fd_sc_hd__a22o_1 _6799_ (.A1(\wbbd_state[10] ),
    .A2(net148),
    .B1(net162),
    .B2(\wbbd_state[9] ),
    .X(_3377_));
 sky130_fd_sc_hd__a221o_1 _6800_ (.A1(\wbbd_state[8] ),
    .A2(net139),
    .B1(net132),
    .B2(_1537_),
    .C1(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__mux2_1 _6801_ (.A0(_3378_),
    .A1(net2660),
    .S(_3376_),
    .X(_0806_));
 sky130_fd_sc_hd__a22o_1 _6802_ (.A1(\wbbd_state[10] ),
    .A2(net149),
    .B1(net140),
    .B2(\wbbd_state[8] ),
    .X(_3379_));
 sky130_fd_sc_hd__a221o_1 _6803_ (.A1(\wbbd_state[9] ),
    .A2(net163),
    .B1(net143),
    .B2(_1537_),
    .C1(_3379_),
    .X(_3380_));
 sky130_fd_sc_hd__mux2_1 _6804_ (.A0(_3380_),
    .A1(net3845),
    .S(_3376_),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _6805_ (.A1(\wbbd_state[10] ),
    .A2(net150),
    .B1(net133),
    .B2(\wbbd_state[9] ),
    .X(_3381_));
 sky130_fd_sc_hd__a221o_1 _6806_ (.A1(\wbbd_state[8] ),
    .A2(net141),
    .B1(net154),
    .B2(net464),
    .C1(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__mux2_1 _6807_ (.A0(_3382_),
    .A1(net3821),
    .S(_3376_),
    .X(_0808_));
 sky130_fd_sc_hd__a22o_1 _6808_ (.A1(\wbbd_state[10] ),
    .A2(net151),
    .B1(net134),
    .B2(\wbbd_state[9] ),
    .X(_3383_));
 sky130_fd_sc_hd__a221o_1 _6809_ (.A1(\wbbd_state[8] ),
    .A2(net142),
    .B1(net157),
    .B2(net464),
    .C1(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__mux2_1 _6810_ (.A0(_3384_),
    .A1(net3867),
    .S(_3376_),
    .X(_0809_));
 sky130_fd_sc_hd__a22o_1 _6811_ (.A1(\wbbd_state[10] ),
    .A2(net152),
    .B1(net135),
    .B2(\wbbd_state[9] ),
    .X(_3385_));
 sky130_fd_sc_hd__a221o_1 _6812_ (.A1(\wbbd_state[8] ),
    .A2(net144),
    .B1(net158),
    .B2(net464),
    .C1(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__mux2_1 _6813_ (.A0(_3386_),
    .A1(net3822),
    .S(_3376_),
    .X(_0810_));
 sky130_fd_sc_hd__a22o_1 _6814_ (.A1(\wbbd_state[10] ),
    .A2(net153),
    .B1(net145),
    .B2(\wbbd_state[8] ),
    .X(_3387_));
 sky130_fd_sc_hd__a221o_1 _6815_ (.A1(\wbbd_state[9] ),
    .A2(net136),
    .B1(net159),
    .B2(net464),
    .C1(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__mux2_1 _6816_ (.A0(_3388_),
    .A1(net3857),
    .S(_3376_),
    .X(_0811_));
 sky130_fd_sc_hd__a22o_1 _6817_ (.A1(\wbbd_state[10] ),
    .A2(net155),
    .B1(net137),
    .B2(\wbbd_state[9] ),
    .X(_3389_));
 sky130_fd_sc_hd__a221o_1 _6818_ (.A1(\wbbd_state[8] ),
    .A2(net146),
    .B1(net160),
    .B2(net464),
    .C1(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__mux2_1 _6819_ (.A0(_3390_),
    .A1(net3816),
    .S(_3376_),
    .X(_0812_));
 sky130_fd_sc_hd__a22o_1 _6820_ (.A1(\wbbd_state[10] ),
    .A2(net156),
    .B1(net138),
    .B2(\wbbd_state[9] ),
    .X(_3391_));
 sky130_fd_sc_hd__a221o_1 _6821_ (.A1(\wbbd_state[8] ),
    .A2(net147),
    .B1(net161),
    .B2(net464),
    .C1(_3391_),
    .X(_3392_));
 sky130_fd_sc_hd__mux2_1 _6822_ (.A0(_3392_),
    .A1(net3830),
    .S(_3376_),
    .X(_0813_));
 sky130_fd_sc_hd__o41ai_2 _6823_ (.A1(net3875),
    .A2(net3813),
    .A3(net624),
    .A4(_1539_),
    .B1(_1536_),
    .Y(_0814_));
 sky130_fd_sc_hd__and3_1 _6824_ (.A(\wbbd_state[10] ),
    .B(net168),
    .C(net170),
    .X(_3393_));
 sky130_fd_sc_hd__a31o_1 _6825_ (.A1(\wbbd_state[9] ),
    .A2(net170),
    .A3(net166),
    .B1(_3393_),
    .X(_3394_));
 sky130_fd_sc_hd__a31o_1 _6826_ (.A1(\wbbd_state[8] ),
    .A2(net170),
    .A3(net167),
    .B1(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__nor2_1 _6827_ (.A(net3854),
    .B(net3893),
    .Y(_3396_));
 sky130_fd_sc_hd__o21a_1 _6828_ (.A1(net2039),
    .A2(\wbbd_state[6] ),
    .B1(_3371_),
    .X(_3397_));
 sky130_fd_sc_hd__a31o_1 _6829_ (.A1(net464),
    .A2(_3396_),
    .A3(_3397_),
    .B1(_3395_),
    .X(_0815_));
 sky130_fd_sc_hd__and2_1 _6830_ (.A(net570),
    .B(net367),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _6831_ (.A(net563),
    .B(net366),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _6832_ (.A(net563),
    .B(net366),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _6833_ (.A(net591),
    .B(net369),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _6834_ (.A(net592),
    .B(net369),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _6835_ (.A(net592),
    .B(net369),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _6836_ (.A(net592),
    .B(net369),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _6837_ (.A(net592),
    .B(net369),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _6838_ (.A(net592),
    .B(net369),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _6839_ (.A(net592),
    .B(net369),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _6840_ (.A(net570),
    .B(net367),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _6841_ (.A(net570),
    .B(net367),
    .X(_0032_));
 sky130_fd_sc_hd__and2_1 _6842_ (.A(net570),
    .B(net366),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _6843_ (.A(net570),
    .B(net367),
    .X(_0034_));
 sky130_fd_sc_hd__and2_1 _6844_ (.A(net563),
    .B(net366),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _6845_ (.A(net563),
    .B(net366),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _6846_ (.A(net563),
    .B(net366),
    .X(_0037_));
 sky130_fd_sc_hd__and2_1 _6847_ (.A(net563),
    .B(net366),
    .X(_0038_));
 sky130_fd_sc_hd__and2_1 _6848_ (.A(net563),
    .B(net366),
    .X(_0039_));
 sky130_fd_sc_hd__and2_1 _6849_ (.A(net563),
    .B(net366),
    .X(_0040_));
 sky130_fd_sc_hd__and2_1 _6850_ (.A(net570),
    .B(net367),
    .X(_0041_));
 sky130_fd_sc_hd__and2_1 _6851_ (.A(net570),
    .B(net368),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _6852_ (.A(net571),
    .B(net368),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _6853_ (.A(net571),
    .B(net368),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _6854_ (.A(net571),
    .B(net368),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _6855_ (.A(net571),
    .B(net368),
    .X(_0046_));
 sky130_fd_sc_hd__and2_1 _6856_ (.A(net570),
    .B(net368),
    .X(_0047_));
 sky130_fd_sc_hd__and2_1 _6857_ (.A(net570),
    .B(net366),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _6858_ (.A(net563),
    .B(net366),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _6859_ (.A(net563),
    .B(net366),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _6860_ (.A(net563),
    .B(net366),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _6861_ (.A(net570),
    .B(net366),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _6862_ (.A(net563),
    .B(net366),
    .X(_0053_));
 sky130_fd_sc_hd__and2_1 _6863_ (.A(net570),
    .B(net366),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _6864_ (.A(net563),
    .B(net366),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _6865_ (.A(net563),
    .B(net366),
    .X(_0056_));
 sky130_fd_sc_hd__and2_1 _6866_ (.A(net570),
    .B(net367),
    .X(_0057_));
 sky130_fd_sc_hd__and2_1 _6867_ (.A(net570),
    .B(net367),
    .X(_0058_));
 sky130_fd_sc_hd__and2_1 _6868_ (.A(net570),
    .B(net367),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _6869_ (.A(net570),
    .B(net366),
    .X(_0060_));
 sky130_fd_sc_hd__and2_1 _6870_ (.A(net571),
    .B(net368),
    .X(_0061_));
 sky130_fd_sc_hd__and2_1 _6871_ (.A(net571),
    .B(net368),
    .X(_0062_));
 sky130_fd_sc_hd__and2_1 _6872_ (.A(net570),
    .B(net368),
    .X(_0063_));
 sky130_fd_sc_hd__and2_1 _6873_ (.A(net570),
    .B(net367),
    .X(_0064_));
 sky130_fd_sc_hd__dfrtp_4 _6874_ (.CLK(clknet_leaf_14_csclk),
    .D(net1693),
    .RESET_B(net591),
    .Q(\gpio_configure[25][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6875_ (.CLK(clknet_leaf_19_csclk),
    .D(net1772),
    .RESET_B(net591),
    .Q(\gpio_configure[25][9] ));
 sky130_fd_sc_hd__dfstp_4 _6876_ (.CLK(clknet_leaf_14_csclk),
    .D(net1588),
    .SET_B(net591),
    .Q(\gpio_configure[25][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6877_ (.CLK(clknet_leaf_14_csclk),
    .D(net1091),
    .RESET_B(net591),
    .Q(\gpio_configure[25][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6878_ (.CLK(clknet_leaf_14_csclk),
    .D(net768),
    .RESET_B(net591),
    .Q(\gpio_configure[25][12] ));
 sky130_fd_sc_hd__dfrtn_1 _6879_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0070_),
    .RESET_B(_0019_),
    .Q(\hkspi.wrstb ));
 sky130_fd_sc_hd__dfrtp_2 _6880_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0071_),
    .RESET_B(_0020_),
    .Q(\hkspi.pre_pass_thru_user ));
 sky130_fd_sc_hd__dfstp_2 _6881_ (.CLK(net623),
    .D(_0018_),
    .SET_B(_0021_),
    .Q(\hkspi.sdoenb ));
 sky130_fd_sc_hd__dfrtp_4 _6882_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0072_),
    .RESET_B(_0023_),
    .Q(\hkspi.pre_pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_1 _6883_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0073_),
    .RESET_B(_0024_),
    .Q(\hkspi.odata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6884_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0074_),
    .RESET_B(_0025_),
    .Q(\hkspi.odata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6885_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0075_),
    .RESET_B(_0026_),
    .Q(\hkspi.odata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6886_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0076_),
    .RESET_B(_0027_),
    .Q(\hkspi.odata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6887_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0077_),
    .RESET_B(_0028_),
    .Q(\hkspi.odata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6888_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0078_),
    .RESET_B(_0029_),
    .Q(\hkspi.odata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6889_ (.CLK(clknet_2_3__leaf_mgmt_gpio_in[4]),
    .D(_0079_),
    .RESET_B(_0030_),
    .Q(\hkspi.odata[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6890_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0080_),
    .RESET_B(_0031_),
    .Q(\hkspi.fixed[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6891_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net3879),
    .RESET_B(_0032_),
    .Q(\hkspi.fixed[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6892_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0082_),
    .RESET_B(_0033_),
    .Q(\hkspi.fixed[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6893_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0083_),
    .RESET_B(_0034_),
    .Q(\hkspi.readmode ));
 sky130_fd_sc_hd__dfrtp_1 _6894_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0084_),
    .RESET_B(_0035_),
    .Q(\hkspi.writemode ));
 sky130_fd_sc_hd__dfrtp_4 _6895_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0085_),
    .RESET_B(_0036_),
    .Q(\hkspi.rdstb ));
 sky130_fd_sc_hd__dfrtp_4 _6896_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0086_),
    .RESET_B(_0037_),
    .Q(\hkspi.pass_thru_mgmt ));
 sky130_fd_sc_hd__dfrtp_4 _6897_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0087_),
    .RESET_B(_0038_),
    .Q(\hkspi.pass_thru_mgmt_delay ));
 sky130_fd_sc_hd__dfrtp_4 _6898_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0088_),
    .RESET_B(_0039_),
    .Q(\hkspi.pass_thru_user ));
 sky130_fd_sc_hd__dfrtp_4 _6899_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net3847),
    .RESET_B(_0040_),
    .Q(\hkspi.pass_thru_user_delay ));
 sky130_fd_sc_hd__dfrtp_4 _6900_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0090_),
    .RESET_B(_0041_),
    .Q(\hkspi.addr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6901_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0091_),
    .RESET_B(_0042_),
    .Q(\hkspi.addr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6902_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0092_),
    .RESET_B(_0043_),
    .Q(\hkspi.addr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6903_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0093_),
    .RESET_B(_0044_),
    .Q(\hkspi.addr[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6904_ (.CLK(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0094_),
    .RESET_B(_0045_),
    .Q(\hkspi.addr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6905_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0095_),
    .RESET_B(_0046_),
    .Q(\hkspi.addr[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6906_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0096_),
    .RESET_B(_0047_),
    .Q(\hkspi.addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6907_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0097_),
    .RESET_B(_0048_),
    .Q(\hkspi.addr[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6908_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0098_),
    .RESET_B(_0049_),
    .Q(\hkspi.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6909_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0099_),
    .RESET_B(_0050_),
    .Q(\hkspi.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6910_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0100_),
    .RESET_B(_0051_),
    .Q(\hkspi.count[2] ));
 sky130_fd_sc_hd__dfstp_2 _6911_ (.CLK(clknet_leaf_73_csclk),
    .D(net1944),
    .SET_B(net565),
    .Q(net293));
 sky130_fd_sc_hd__dfstp_2 _6912_ (.CLK(clknet_leaf_73_csclk),
    .D(net1285),
    .SET_B(net565),
    .Q(net294));
 sky130_fd_sc_hd__dfstp_4 _6913_ (.CLK(clknet_leaf_73_csclk),
    .D(net1149),
    .SET_B(net566),
    .Q(net270));
 sky130_fd_sc_hd__dfstp_2 _6914_ (.CLK(clknet_leaf_73_csclk),
    .D(net1584),
    .SET_B(net566),
    .Q(net271));
 sky130_fd_sc_hd__dfrtp_4 _6915_ (.CLK(clknet_leaf_73_csclk),
    .D(net1355),
    .RESET_B(net566),
    .Q(net272));
 sky130_fd_sc_hd__dfstp_4 _6916_ (.CLK(clknet_leaf_70_csclk),
    .D(net979),
    .SET_B(net566),
    .Q(net273));
 sky130_fd_sc_hd__dfstp_4 _6917_ (.CLK(clknet_leaf_70_csclk),
    .D(net2831),
    .SET_B(net566),
    .Q(net274));
 sky130_fd_sc_hd__dfstp_4 _6918_ (.CLK(clknet_leaf_70_csclk),
    .D(net2725),
    .SET_B(net566),
    .Q(net275));
 sky130_fd_sc_hd__dfstp_2 _6919_ (.CLK(clknet_leaf_74_csclk),
    .D(net1948),
    .SET_B(net565),
    .Q(net269));
 sky130_fd_sc_hd__dfstp_4 _6920_ (.CLK(clknet_leaf_73_csclk),
    .D(net1289),
    .SET_B(net565),
    .Q(net280));
 sky130_fd_sc_hd__dfstp_2 _6921_ (.CLK(clknet_leaf_74_csclk),
    .D(net1119),
    .SET_B(net565),
    .Q(net287));
 sky130_fd_sc_hd__dfstp_4 _6922_ (.CLK(clknet_leaf_74_csclk),
    .D(net1592),
    .SET_B(net565),
    .Q(net288));
 sky130_fd_sc_hd__dfstp_4 _6923_ (.CLK(clknet_leaf_73_csclk),
    .D(_0113_),
    .SET_B(net565),
    .Q(net289));
 sky130_fd_sc_hd__dfstp_4 _6924_ (.CLK(clknet_leaf_73_csclk),
    .D(net907),
    .SET_B(net565),
    .Q(net290));
 sky130_fd_sc_hd__dfstp_4 _6925_ (.CLK(clknet_leaf_73_csclk),
    .D(net2793),
    .SET_B(net565),
    .Q(net291));
 sky130_fd_sc_hd__dfstp_4 _6926_ (.CLK(clknet_leaf_73_csclk),
    .D(net2716),
    .SET_B(net565),
    .Q(net292));
 sky130_fd_sc_hd__dfstp_2 _6927_ (.CLK(clknet_leaf_69_csclk),
    .D(net1934),
    .SET_B(net575),
    .Q(net285));
 sky130_fd_sc_hd__dfstp_2 _6928_ (.CLK(clknet_leaf_69_csclk),
    .D(net1281),
    .SET_B(net575),
    .Q(net286));
 sky130_fd_sc_hd__dfstp_4 _6929_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(net3896),
    .SET_B(net563),
    .Q(\xfer_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6930_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0015_),
    .RESET_B(net565),
    .Q(\xfer_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6931_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0016_),
    .RESET_B(net567),
    .Q(\xfer_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6932_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0017_),
    .RESET_B(net567),
    .Q(\xfer_state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6933_ (.CLK(clknet_leaf_36_csclk),
    .D(net1504),
    .RESET_B(net603),
    .Q(\mgmt_gpio_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6934_ (.CLK(clknet_leaf_39_csclk),
    .D(net1850),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6935_ (.CLK(clknet_leaf_40_csclk),
    .D(net1424),
    .RESET_B(net594),
    .Q(\mgmt_gpio_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6936_ (.CLK(clknet_leaf_39_csclk),
    .D(net1493),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6937_ (.CLK(clknet_leaf_39_csclk),
    .D(net1614),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6938_ (.CLK(clknet_leaf_38_csclk),
    .D(net2023),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6939_ (.CLK(clknet_leaf_36_csclk),
    .D(net1035),
    .RESET_B(net603),
    .Q(\mgmt_gpio_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6940_ (.CLK(clknet_leaf_36_csclk),
    .D(net1518),
    .RESET_B(net604),
    .Q(\mgmt_gpio_data[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6941_ (.CLK(clknet_leaf_53_csclk),
    .D(net1846),
    .RESET_B(net582),
    .Q(\mgmt_gpio_data[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6942_ (.CLK(clknet_leaf_52_csclk),
    .D(net1506),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6943_ (.CLK(clknet_leaf_52_csclk),
    .D(net1307),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6944_ (.CLK(clknet_leaf_52_csclk),
    .D(net1442),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6945_ (.CLK(clknet_leaf_49_csclk),
    .D(net1219),
    .RESET_B(net583),
    .Q(\mgmt_gpio_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6946_ (.CLK(clknet_leaf_48_csclk),
    .D(net1842),
    .RESET_B(net583),
    .Q(\mgmt_gpio_data[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6947_ (.CLK(clknet_leaf_52_csclk),
    .D(net1670),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6948_ (.CLK(clknet_leaf_52_csclk),
    .D(net1499),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6949_ (.CLK(clknet_leaf_36_csclk),
    .D(net1163),
    .RESET_B(net604),
    .Q(\mgmt_gpio_data_buf[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6950_ (.CLK(clknet_leaf_38_csclk),
    .D(net1652),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data_buf[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6951_ (.CLK(clknet_leaf_39_csclk),
    .D(net874),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data_buf[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6952_ (.CLK(clknet_leaf_39_csclk),
    .D(net1029),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data_buf[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6953_ (.CLK(clknet_leaf_38_csclk),
    .D(net1272),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data_buf[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6954_ (.CLK(clknet_leaf_38_csclk),
    .D(net627),
    .RESET_B(net595),
    .Q(\mgmt_gpio_data_buf[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6955_ (.CLK(clknet_leaf_36_csclk),
    .D(net749),
    .RESET_B(net604),
    .Q(\mgmt_gpio_data_buf[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6956_ (.CLK(clknet_leaf_36_csclk),
    .D(net1237),
    .RESET_B(net604),
    .Q(\mgmt_gpio_data_buf[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6957_ (.CLK(clknet_leaf_71_csclk),
    .D(net1946),
    .RESET_B(net567),
    .Q(\gpio_configure[0][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6958_ (.CLK(clknet_leaf_71_csclk),
    .D(net1283),
    .RESET_B(net566),
    .Q(\gpio_configure[0][9] ));
 sky130_fd_sc_hd__dfrtp_4 _6959_ (.CLK(clknet_leaf_71_csclk),
    .D(net1113),
    .RESET_B(net567),
    .Q(\gpio_configure[0][10] ));
 sky130_fd_sc_hd__dfstp_2 _6960_ (.CLK(clknet_leaf_71_csclk),
    .D(net1596),
    .SET_B(net567),
    .Q(\gpio_configure[0][11] ));
 sky130_fd_sc_hd__dfstp_4 _6961_ (.CLK(clknet_leaf_71_csclk),
    .D(net1384),
    .SET_B(net566),
    .Q(\gpio_configure[0][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6962_ (.CLK(clknet_leaf_1_csclk),
    .D(net1901),
    .RESET_B(net572),
    .Q(\gpio_configure[1][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6963_ (.CLK(clknet_leaf_10_csclk),
    .D(net1762),
    .RESET_B(net590),
    .Q(\gpio_configure[1][9] ));
 sky130_fd_sc_hd__dfrtp_4 _6964_ (.CLK(clknet_leaf_0_csclk),
    .D(net2479),
    .RESET_B(net572),
    .Q(\gpio_configure[1][10] ));
 sky130_fd_sc_hd__dfstp_4 _6965_ (.CLK(clknet_leaf_1_csclk),
    .D(net1624),
    .SET_B(net570),
    .Q(\gpio_configure[1][11] ));
 sky130_fd_sc_hd__dfstp_2 _6966_ (.CLK(clknet_leaf_10_csclk),
    .D(net1473),
    .SET_B(net590),
    .Q(\gpio_configure[1][12] ));
 sky130_fd_sc_hd__dfrtp_4 _6967_ (.CLK(clknet_leaf_8_csclk),
    .D(net1650),
    .RESET_B(net589),
    .Q(\gpio_configure[2][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6968_ (.CLK(clknet_leaf_8_csclk),
    .D(net1709),
    .RESET_B(net588),
    .Q(\gpio_configure[2][9] ));
 sky130_fd_sc_hd__dfstp_4 _6969_ (.CLK(clknet_leaf_8_csclk),
    .D(net1520),
    .SET_B(net589),
    .Q(\gpio_configure[2][10] ));
 sky130_fd_sc_hd__dfrtp_4 _6970_ (.CLK(clknet_leaf_8_csclk),
    .D(net951),
    .RESET_B(net589),
    .Q(\gpio_configure[2][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6971_ (.CLK(clknet_leaf_8_csclk),
    .D(net1378),
    .RESET_B(net588),
    .Q(\gpio_configure[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0158_),
    .Q(net319));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0159_),
    .Q(net320));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0160_),
    .Q(net321));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0161_),
    .Q(net322));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0162_),
    .Q(net324));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0163_),
    .Q(net325));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0164_),
    .Q(net326));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0165_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0166_),
    .Q(net342));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0167_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0168_),
    .Q(net313));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0169_),
    .Q(net314));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0170_),
    .Q(net315));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0171_),
    .Q(net316));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0172_),
    .Q(net317));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0173_),
    .Q(net318));
 sky130_fd_sc_hd__dfrtp_4 _6988_ (.CLK(clknet_leaf_67_csclk),
    .D(net1950),
    .RESET_B(net568),
    .Q(\gpio_configure[3][8] ));
 sky130_fd_sc_hd__dfrtp_4 _6989_ (.CLK(clknet_leaf_67_csclk),
    .D(net1287),
    .RESET_B(net577),
    .Q(\gpio_configure[3][9] ));
 sky130_fd_sc_hd__dfrtp_4 _6990_ (.CLK(clknet_leaf_67_csclk),
    .D(net1137),
    .RESET_B(net577),
    .Q(\gpio_configure[3][10] ));
 sky130_fd_sc_hd__dfstp_4 _6991_ (.CLK(clknet_leaf_71_csclk),
    .D(net1598),
    .SET_B(net566),
    .Q(\gpio_configure[3][11] ));
 sky130_fd_sc_hd__dfrtp_4 _6992_ (.CLK(clknet_leaf_71_csclk),
    .D(net1370),
    .RESET_B(net568),
    .Q(\gpio_configure[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0179_),
    .Q(net312));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0180_),
    .Q(net323));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0181_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0182_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0183_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0184_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(clknet_4_2__leaf_wb_clk_i),
    .D(_0185_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0186_),
    .Q(net341));
 sky130_fd_sc_hd__dfrtp_4 _7001_ (.CLK(clknet_leaf_77_csclk),
    .D(net1921),
    .RESET_B(net572),
    .Q(\gpio_configure[4][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7002_ (.CLK(clknet_leaf_5_csclk),
    .D(net1293),
    .RESET_B(net574),
    .Q(\gpio_configure[4][9] ));
 sky130_fd_sc_hd__dfstp_2 _7003_ (.CLK(clknet_leaf_77_csclk),
    .D(net1221),
    .SET_B(net572),
    .Q(\gpio_configure[4][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7004_ (.CLK(clknet_leaf_5_csclk),
    .D(net1570),
    .RESET_B(net573),
    .Q(\gpio_configure[4][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7005_ (.CLK(clknet_leaf_5_csclk),
    .D(net1347),
    .RESET_B(net574),
    .Q(\gpio_configure[4][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7006_ (.CLK(clknet_leaf_4_csclk),
    .D(net1893),
    .RESET_B(net573),
    .Q(\gpio_configure[5][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7007_ (.CLK(clknet_leaf_2_csclk),
    .D(net1321),
    .RESET_B(net572),
    .Q(\gpio_configure[5][9] ));
 sky130_fd_sc_hd__dfstp_2 _7008_ (.CLK(clknet_leaf_0_csclk),
    .D(net2279),
    .SET_B(net572),
    .Q(\gpio_configure[5][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7009_ (.CLK(clknet_leaf_3_csclk),
    .D(net1556),
    .RESET_B(net573),
    .Q(\gpio_configure[5][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7010_ (.CLK(clknet_leaf_2_csclk),
    .D(net1410),
    .RESET_B(net573),
    .Q(\gpio_configure[5][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7011_ (.CLK(clknet_leaf_6_csclk),
    .D(net1917),
    .RESET_B(net572),
    .Q(\gpio_configure[6][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7012_ (.CLK(clknet_leaf_12_csclk),
    .D(net1760),
    .RESET_B(net589),
    .Q(\gpio_configure[6][9] ));
 sky130_fd_sc_hd__dfstp_2 _7013_ (.CLK(clknet_leaf_0_csclk),
    .D(net2456),
    .SET_B(net572),
    .Q(\gpio_configure[6][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7014_ (.CLK(clknet_leaf_10_csclk),
    .D(net1075),
    .RESET_B(net590),
    .Q(\gpio_configure[6][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7015_ (.CLK(clknet_leaf_10_csclk),
    .D(net1468),
    .RESET_B(net590),
    .Q(\gpio_configure[6][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7016_ (.CLK(clknet_leaf_6_csclk),
    .D(net1919),
    .RESET_B(net572),
    .Q(\gpio_configure[7][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7017_ (.CLK(clknet_leaf_4_csclk),
    .D(net690),
    .RESET_B(net573),
    .Q(\gpio_configure[7][9] ));
 sky130_fd_sc_hd__dfstp_2 _7018_ (.CLK(clknet_leaf_6_csclk),
    .D(net1197),
    .SET_B(net572),
    .Q(\gpio_configure[7][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7019_ (.CLK(clknet_leaf_4_csclk),
    .D(net1540),
    .RESET_B(net573),
    .Q(\gpio_configure[7][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7020_ (.CLK(clknet_leaf_4_csclk),
    .D(net1323),
    .RESET_B(net573),
    .Q(\gpio_configure[7][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7021_ (.CLK(clknet_leaf_67_csclk),
    .D(net1952),
    .RESET_B(net568),
    .Q(\gpio_configure[8][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7022_ (.CLK(clknet_leaf_67_csclk),
    .D(net1291),
    .RESET_B(net568),
    .Q(\gpio_configure[8][9] ));
 sky130_fd_sc_hd__dfstp_2 _7023_ (.CLK(clknet_leaf_71_csclk),
    .D(net1129),
    .SET_B(net568),
    .Q(\gpio_configure[8][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7024_ (.CLK(clknet_leaf_71_csclk),
    .D(net1576),
    .RESET_B(net568),
    .Q(\gpio_configure[8][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7025_ (.CLK(clknet_leaf_67_csclk),
    .D(net1374),
    .RESET_B(net568),
    .Q(\gpio_configure[8][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7026_ (.CLK(clknet_leaf_8_csclk),
    .D(net1644),
    .RESET_B(net590),
    .Q(\gpio_configure[9][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7027_ (.CLK(clknet_leaf_8_csclk),
    .D(net1717),
    .RESET_B(net589),
    .Q(\gpio_configure[9][9] ));
 sky130_fd_sc_hd__dfstp_4 _7028_ (.CLK(clknet_leaf_12_csclk),
    .D(net1586),
    .SET_B(net589),
    .Q(\gpio_configure[9][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7029_ (.CLK(clknet_leaf_8_csclk),
    .D(net939),
    .RESET_B(net590),
    .Q(\gpio_configure[9][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7030_ (.CLK(clknet_leaf_8_csclk),
    .D(net1390),
    .RESET_B(net590),
    .Q(\gpio_configure[9][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7031_ (.CLK(clknet_leaf_12_csclk),
    .D(net1689),
    .RESET_B(net589),
    .Q(\gpio_configure[10][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7032_ (.CLK(clknet_leaf_12_csclk),
    .D(net1756),
    .RESET_B(net589),
    .Q(\gpio_configure[10][9] ));
 sky130_fd_sc_hd__dfstp_4 _7033_ (.CLK(clknet_leaf_7_csclk),
    .D(net1532),
    .SET_B(net588),
    .Q(\gpio_configure[10][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7034_ (.CLK(clknet_leaf_12_csclk),
    .D(net2580),
    .RESET_B(net589),
    .Q(\gpio_configure[10][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7035_ (.CLK(clknet_leaf_8_csclk),
    .D(net1372),
    .RESET_B(net588),
    .Q(\gpio_configure[10][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7036_ (.CLK(clknet_leaf_77_csclk),
    .D(net1923),
    .RESET_B(net572),
    .Q(\gpio_configure[11][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7037_ (.CLK(clknet_leaf_0_csclk),
    .D(net1254),
    .RESET_B(net572),
    .Q(\gpio_configure[11][9] ));
 sky130_fd_sc_hd__dfstp_1 _7038_ (.CLK(clknet_leaf_0_csclk),
    .D(net2475),
    .SET_B(net572),
    .Q(\gpio_configure[11][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7039_ (.CLK(clknet_leaf_0_csclk),
    .D(net2595),
    .RESET_B(net572),
    .Q(\gpio_configure[11][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7040_ (.CLK(clknet_leaf_0_csclk),
    .D(net1345),
    .RESET_B(net572),
    .Q(\gpio_configure[11][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7041_ (.CLK(clknet_leaf_14_csclk),
    .D(net1695),
    .RESET_B(net592),
    .Q(\gpio_configure[12][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7042_ (.CLK(clknet_leaf_14_csclk),
    .D(net1241),
    .RESET_B(net591),
    .Q(\gpio_configure[12][9] ));
 sky130_fd_sc_hd__dfstp_4 _7043_ (.CLK(clknet_leaf_19_csclk),
    .D(net1606),
    .SET_B(net591),
    .Q(\gpio_configure[12][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7044_ (.CLK(clknet_leaf_14_csclk),
    .D(net1063),
    .RESET_B(net592),
    .Q(\gpio_configure[12][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7045_ (.CLK(clknet_leaf_13_csclk),
    .D(net785),
    .RESET_B(net591),
    .Q(\gpio_configure[12][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7046_ (.CLK(clknet_leaf_21_csclk),
    .D(net1719),
    .RESET_B(net588),
    .Q(\gpio_configure[29][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7047_ (.CLK(clknet_leaf_21_csclk),
    .D(net1766),
    .RESET_B(net588),
    .Q(\gpio_configure[29][9] ));
 sky130_fd_sc_hd__dfstp_4 _7048_ (.CLK(clknet_leaf_7_csclk),
    .D(net1530),
    .SET_B(net588),
    .Q(\gpio_configure[29][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7049_ (.CLK(clknet_leaf_7_csclk),
    .D(net995),
    .RESET_B(net588),
    .Q(\gpio_configure[29][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7050_ (.CLK(clknet_leaf_21_csclk),
    .D(net1481),
    .RESET_B(net593),
    .Q(\gpio_configure[29][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7051_ (.CLK(clknet_leaf_0_csclk),
    .D(net1889),
    .RESET_B(net572),
    .Q(\gpio_configure[23][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7052_ (.CLK(clknet_leaf_8_csclk),
    .D(net1703),
    .RESET_B(net590),
    .Q(\gpio_configure[23][9] ));
 sky130_fd_sc_hd__dfstp_2 _7053_ (.CLK(clknet_leaf_6_csclk),
    .D(net1033),
    .SET_B(net572),
    .Q(\gpio_configure[23][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7054_ (.CLK(clknet_leaf_4_csclk),
    .D(net997),
    .RESET_B(net573),
    .Q(\gpio_configure[23][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7055_ (.CLK(clknet_leaf_9_csclk),
    .D(net1436),
    .RESET_B(net590),
    .Q(\gpio_configure[23][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7056_ (.CLK(clknet_leaf_4_csclk),
    .D(net1764),
    .RESET_B(net573),
    .Q(\gpio_configure[27][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7057_ (.CLK(clknet_leaf_10_csclk),
    .D(net1750),
    .RESET_B(net590),
    .Q(\gpio_configure[27][9] ));
 sky130_fd_sc_hd__dfstp_1 _7058_ (.CLK(clknet_leaf_0_csclk),
    .D(net2212),
    .SET_B(net572),
    .Q(\gpio_configure[27][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7059_ (.CLK(clknet_leaf_3_csclk),
    .D(net1007),
    .RESET_B(net573),
    .Q(\gpio_configure[27][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7060_ (.CLK(clknet_leaf_4_csclk),
    .D(net1333),
    .RESET_B(net573),
    .Q(\gpio_configure[27][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7061_ (.CLK(clknet_leaf_1_csclk),
    .D(net1905),
    .RESET_B(net570),
    .Q(\gpio_configure[24][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7062_ (.CLK(clknet_leaf_3_csclk),
    .D(net668),
    .RESET_B(net573),
    .Q(\gpio_configure[24][9] ));
 sky130_fd_sc_hd__dfstp_2 _7063_ (.CLK(clknet_leaf_0_csclk),
    .D(net923),
    .SET_B(net572),
    .Q(\gpio_configure[24][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7064_ (.CLK(clknet_leaf_3_csclk),
    .D(net1538),
    .RESET_B(net573),
    .Q(\gpio_configure[24][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7065_ (.CLK(clknet_leaf_3_csclk),
    .D(net1325),
    .RESET_B(net573),
    .Q(\gpio_configure[24][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7066_ (.CLK(clknet_leaf_2_csclk),
    .D(net1885),
    .RESET_B(net571),
    .Q(\gpio_configure[26][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7067_ (.CLK(clknet_leaf_11_csclk),
    .D(net1796),
    .RESET_B(net606),
    .Q(\gpio_configure[26][9] ));
 sky130_fd_sc_hd__dfstp_2 _7068_ (.CLK(clknet_leaf_1_csclk),
    .D(net999),
    .SET_B(net570),
    .Q(\gpio_configure[26][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7069_ (.CLK(clknet_leaf_3_csclk),
    .D(net1009),
    .RESET_B(net571),
    .Q(\gpio_configure[26][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7070_ (.CLK(clknet_leaf_10_csclk),
    .D(net1460),
    .RESET_B(net590),
    .Q(\gpio_configure[26][12] ));
 sky130_fd_sc_hd__dfstp_4 _7071_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0004_),
    .SET_B(_0052_),
    .Q(\hkspi.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7072_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0005_),
    .RESET_B(_0053_),
    .Q(\hkspi.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7073_ (.CLK(clknet_2_0__leaf_mgmt_gpio_in[4]),
    .D(_0006_),
    .RESET_B(_0054_),
    .Q(\hkspi.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7074_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0007_),
    .RESET_B(_0055_),
    .Q(\hkspi.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7075_ (.CLK(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net3861),
    .RESET_B(_0056_),
    .Q(\hkspi.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7076_ (.CLK(clknet_leaf_35_csclk),
    .D(net1932),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7077_ (.CLK(clknet_leaf_35_csclk),
    .D(net1844),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7078_ (.CLK(clknet_leaf_35_csclk),
    .D(net1339),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7079_ (.CLK(clknet_leaf_35_csclk),
    .D(net1400),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7080_ (.CLK(clknet_leaf_15_csclk),
    .D(net1770),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7081_ (.CLK(clknet_leaf_16_csclk),
    .D(net1450),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7082_ (.CLK(clknet_leaf_16_csclk),
    .D(net1105),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7083_ (.CLK(clknet_leaf_29_csclk),
    .D(net1512),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[23] ));
 sky130_fd_sc_hd__dfrtp_4 _7084_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(_0265_),
    .RESET_B(net607),
    .Q(wbbd_busy));
 sky130_fd_sc_hd__dfrtp_1 _7085_ (.CLK(clknet_leaf_29_csclk),
    .D(net1852),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7086_ (.CLK(clknet_leaf_29_csclk),
    .D(net1633),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7087_ (.CLK(clknet_leaf_29_csclk),
    .D(net820),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7088_ (.CLK(clknet_leaf_29_csclk),
    .D(net878),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7089_ (.CLK(clknet_leaf_30_csclk),
    .D(net719),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7090_ (.CLK(clknet_leaf_30_csclk),
    .D(net810),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7091_ (.CLK(clknet_leaf_30_csclk),
    .D(net703),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[30] ));
 sky130_fd_sc_hd__dfrtp_1 _7092_ (.CLK(clknet_leaf_32_csclk),
    .D(net1172),
    .RESET_B(net603),
    .Q(\mgmt_gpio_data[31] ));
 sky130_fd_sc_hd__dfrtp_1 _7093_ (.CLK(clknet_leaf_35_csclk),
    .D(net1089),
    .RESET_B(net604),
    .Q(\mgmt_gpio_data_buf[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7094_ (.CLK(clknet_leaf_35_csclk),
    .D(net1648),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data_buf[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7095_ (.CLK(clknet_leaf_35_csclk),
    .D(net842),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data_buf[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7096_ (.CLK(clknet_leaf_35_csclk),
    .D(net884),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data_buf[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7097_ (.CLK(clknet_leaf_15_csclk),
    .D(net794),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data_buf[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7098_ (.CLK(clknet_leaf_15_csclk),
    .D(net1003),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data_buf[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7099_ (.CLK(clknet_leaf_16_csclk),
    .D(net760),
    .RESET_B(net601),
    .Q(\mgmt_gpio_data_buf[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7100_ (.CLK(clknet_leaf_28_csclk),
    .D(net1258),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data_buf[23] ));
 sky130_fd_sc_hd__dfstp_2 _7101_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(net3855),
    .SET_B(net607),
    .Q(\wbbd_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7102_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0000_),
    .RESET_B(net607),
    .Q(\wbbd_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7103_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0001_),
    .RESET_B(net608),
    .Q(\wbbd_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7104_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0002_),
    .RESET_B(net607),
    .Q(\wbbd_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7105_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(net3813),
    .RESET_B(net607),
    .Q(\wbbd_state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7106_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0003_),
    .RESET_B(net608),
    .Q(\wbbd_state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7107_ (.CLK(clknet_4_13__leaf_wb_clk_i),
    .D(_0011_),
    .RESET_B(net607),
    .Q(\wbbd_state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7108_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(net3810),
    .RESET_B(net607),
    .Q(\wbbd_state[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7109_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0012_),
    .RESET_B(net607),
    .Q(\wbbd_state[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7110_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(_0013_),
    .RESET_B(net607),
    .Q(\wbbd_state[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7111_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0010_),
    .RESET_B(net607),
    .Q(\wbbd_state[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7112_ (.CLK(clknet_leaf_12_csclk),
    .D(net1687),
    .RESET_B(net589),
    .Q(\gpio_configure[13][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7113_ (.CLK(clknet_leaf_8_csclk),
    .D(net1713),
    .RESET_B(net589),
    .Q(\gpio_configure[13][9] ));
 sky130_fd_sc_hd__dfstp_4 _7114_ (.CLK(clknet_leaf_13_csclk),
    .D(net1608),
    .SET_B(net589),
    .Q(\gpio_configure[13][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7115_ (.CLK(clknet_leaf_13_csclk),
    .D(net1107),
    .RESET_B(net589),
    .Q(\gpio_configure[13][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7116_ (.CLK(clknet_leaf_13_csclk),
    .D(net1477),
    .RESET_B(net588),
    .Q(\gpio_configure[13][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7117_ (.CLK(clknet_leaf_17_csclk),
    .D(net1701),
    .RESET_B(net598),
    .Q(\gpio_configure[37][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7118_ (.CLK(clknet_leaf_15_csclk),
    .D(net1774),
    .RESET_B(net601),
    .Q(\gpio_configure[37][9] ));
 sky130_fd_sc_hd__dfrtp_4 _7119_ (.CLK(clknet_leaf_17_csclk),
    .D(net1566),
    .RESET_B(net601),
    .Q(\gpio_configure[37][10] ));
 sky130_fd_sc_hd__dfstp_2 _7120_ (.CLK(clknet_leaf_17_csclk),
    .D(net1111),
    .SET_B(net601),
    .Q(\gpio_configure[37][11] ));
 sky130_fd_sc_hd__dfstp_2 _7121_ (.CLK(clknet_leaf_17_csclk),
    .D(net781),
    .SET_B(net598),
    .Q(\gpio_configure[37][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7122_ (.CLK(clknet_leaf_13_csclk),
    .D(net1705),
    .RESET_B(net591),
    .Q(\gpio_configure[14][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7123_ (.CLK(clknet_leaf_13_csclk),
    .D(net1768),
    .RESET_B(net591),
    .Q(\gpio_configure[14][9] ));
 sky130_fd_sc_hd__dfstp_4 _7124_ (.CLK(clknet_leaf_13_csclk),
    .D(net1600),
    .SET_B(net591),
    .Q(\gpio_configure[14][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7125_ (.CLK(clknet_leaf_13_csclk),
    .D(net2576),
    .RESET_B(net591),
    .Q(\gpio_configure[14][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7126_ (.CLK(clknet_leaf_13_csclk),
    .D(net2753),
    .RESET_B(net591),
    .Q(\gpio_configure[14][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7127_ (.CLK(clknet_leaf_18_csclk),
    .D(net1723),
    .RESET_B(net598),
    .Q(\gpio_configure[36][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7128_ (.CLK(clknet_leaf_18_csclk),
    .D(net1278),
    .RESET_B(net598),
    .Q(\gpio_configure[36][9] ));
 sky130_fd_sc_hd__dfrtp_4 _7129_ (.CLK(clknet_leaf_22_csclk),
    .D(net1578),
    .RESET_B(net593),
    .Q(\gpio_configure[36][10] ));
 sky130_fd_sc_hd__dfstp_2 _7130_ (.CLK(clknet_leaf_18_csclk),
    .D(net1135),
    .SET_B(net598),
    .Q(\gpio_configure[36][11] ));
 sky130_fd_sc_hd__dfstp_2 _7131_ (.CLK(clknet_leaf_18_csclk),
    .D(net792),
    .SET_B(net598),
    .Q(\gpio_configure[36][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7132_ (.CLK(clknet_leaf_7_csclk),
    .D(net1680),
    .RESET_B(net588),
    .Q(\gpio_configure[15][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7133_ (.CLK(clknet_leaf_20_csclk),
    .D(net1754),
    .RESET_B(net591),
    .Q(\gpio_configure[15][9] ));
 sky130_fd_sc_hd__dfstp_4 _7134_ (.CLK(clknet_leaf_13_csclk),
    .D(net1616),
    .SET_B(net588),
    .Q(\gpio_configure[15][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7135_ (.CLK(clknet_leaf_20_csclk),
    .D(net2606),
    .RESET_B(net588),
    .Q(\gpio_configure[15][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7136_ (.CLK(clknet_leaf_7_csclk),
    .D(net1422),
    .RESET_B(net588),
    .Q(\gpio_configure[15][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7137_ (.CLK(clknet_leaf_17_csclk),
    .D(net1699),
    .RESET_B(net601),
    .Q(\gpio_configure[35][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7138_ (.CLK(clknet_leaf_17_csclk),
    .D(net1260),
    .RESET_B(net598),
    .Q(\gpio_configure[35][9] ));
 sky130_fd_sc_hd__dfstp_4 _7139_ (.CLK(clknet_leaf_19_csclk),
    .D(net1618),
    .SET_B(net598),
    .Q(\gpio_configure[35][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7140_ (.CLK(clknet_leaf_19_csclk),
    .D(net1115),
    .RESET_B(net598),
    .Q(\gpio_configure[35][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7141_ (.CLK(clknet_leaf_15_csclk),
    .D(net1485),
    .RESET_B(net601),
    .Q(\gpio_configure[35][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7142_ (.CLK(clknet_leaf_77_csclk),
    .D(net1958),
    .RESET_B(net567),
    .Q(\gpio_configure[16][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7143_ (.CLK(clknet_leaf_76_csclk),
    .D(net1319),
    .RESET_B(net567),
    .Q(\gpio_configure[16][9] ));
 sky130_fd_sc_hd__dfstp_2 _7144_ (.CLK(clknet_leaf_77_csclk),
    .D(net2653),
    .SET_B(net567),
    .Q(\gpio_configure[16][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7145_ (.CLK(clknet_leaf_76_csclk),
    .D(net1626),
    .RESET_B(net567),
    .Q(\gpio_configure[16][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7146_ (.CLK(clknet_leaf_76_csclk),
    .D(net1396),
    .RESET_B(net567),
    .Q(\gpio_configure[16][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7147_ (.CLK(clknet_leaf_17_csclk),
    .D(net1697),
    .RESET_B(net598),
    .Q(\gpio_configure[34][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7148_ (.CLK(clknet_leaf_18_csclk),
    .D(net1295),
    .RESET_B(net598),
    .Q(\gpio_configure[34][9] ));
 sky130_fd_sc_hd__dfstp_2 _7149_ (.CLK(clknet_leaf_17_csclk),
    .D(net1582),
    .SET_B(net598),
    .Q(\gpio_configure[34][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7150_ (.CLK(clknet_leaf_18_csclk),
    .D(net1133),
    .RESET_B(net598),
    .Q(\gpio_configure[34][11] ));
 sky130_fd_sc_hd__dfrtp_2 _7151_ (.CLK(clknet_leaf_21_csclk),
    .D(net1483),
    .RESET_B(net593),
    .Q(\gpio_configure[34][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7152_ (.CLK(clknet_leaf_19_csclk),
    .D(net1711),
    .RESET_B(net591),
    .Q(\gpio_configure[17][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7153_ (.CLK(clknet_leaf_19_csclk),
    .D(net1266),
    .RESET_B(net591),
    .Q(\gpio_configure[17][9] ));
 sky130_fd_sc_hd__dfstp_4 _7154_ (.CLK(clknet_leaf_19_csclk),
    .D(net1612),
    .SET_B(net591),
    .Q(\gpio_configure[17][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7155_ (.CLK(clknet_leaf_19_csclk),
    .D(net2620),
    .RESET_B(net591),
    .Q(\gpio_configure[17][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7156_ (.CLK(clknet_leaf_19_csclk),
    .D(net2732),
    .RESET_B(net598),
    .Q(\gpio_configure[17][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7157_ (.CLK(clknet_leaf_1_csclk),
    .D(net1903),
    .RESET_B(net571),
    .Q(\gpio_configure[33][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7158_ (.CLK(clknet_leaf_2_csclk),
    .D(net1315),
    .RESET_B(net571),
    .Q(\gpio_configure[33][9] ));
 sky130_fd_sc_hd__dfstp_2 _7159_ (.CLK(clknet_leaf_1_csclk),
    .D(net965),
    .SET_B(net571),
    .Q(\gpio_configure[33][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7160_ (.CLK(clknet_leaf_3_csclk),
    .D(net1552),
    .RESET_B(net571),
    .Q(\gpio_configure[33][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7161_ (.CLK(clknet_leaf_2_csclk),
    .D(net1404),
    .RESET_B(net571),
    .Q(\gpio_configure[33][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7162_ (.CLK(clknet_leaf_5_csclk),
    .D(net1879),
    .RESET_B(net573),
    .Q(\gpio_configure[18][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7163_ (.CLK(clknet_leaf_9_csclk),
    .D(net1748),
    .RESET_B(net590),
    .Q(\gpio_configure[18][9] ));
 sky130_fd_sc_hd__dfstp_1 _7164_ (.CLK(clknet_leaf_0_csclk),
    .D(net957),
    .SET_B(net572),
    .Q(\gpio_configure[18][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7165_ (.CLK(clknet_leaf_4_csclk),
    .D(net1049),
    .RESET_B(net573),
    .Q(\gpio_configure[18][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7166_ (.CLK(clknet_leaf_9_csclk),
    .D(net1458),
    .RESET_B(net590),
    .Q(\gpio_configure[18][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7167_ (.CLK(clknet_leaf_4_csclk),
    .D(net1897),
    .RESET_B(net573),
    .Q(\gpio_configure[32][8] ));
 sky130_fd_sc_hd__dfrtp_2 _7168_ (.CLK(clknet_leaf_9_csclk),
    .D(net1742),
    .RESET_B(net590),
    .Q(\gpio_configure[32][9] ));
 sky130_fd_sc_hd__dfstp_2 _7169_ (.CLK(clknet_leaf_4_csclk),
    .D(net2300),
    .SET_B(net573),
    .Q(\gpio_configure[32][10] ));
 sky130_fd_sc_hd__dfrtp_2 _7170_ (.CLK(clknet_leaf_4_csclk),
    .D(net1542),
    .RESET_B(net574),
    .Q(\gpio_configure[32][11] ));
 sky130_fd_sc_hd__dfrtp_2 _7171_ (.CLK(clknet_leaf_9_csclk),
    .D(net1454),
    .RESET_B(net590),
    .Q(\gpio_configure[32][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7172_ (.CLK(clknet_leaf_7_csclk),
    .D(net1678),
    .RESET_B(net588),
    .Q(\gpio_configure[19][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7173_ (.CLK(clknet_leaf_7_csclk),
    .D(net1732),
    .RESET_B(net588),
    .Q(\gpio_configure[19][9] ));
 sky130_fd_sc_hd__dfstp_4 _7174_ (.CLK(clknet_leaf_7_csclk),
    .D(net1536),
    .SET_B(net588),
    .Q(\gpio_configure[19][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7175_ (.CLK(clknet_leaf_7_csclk),
    .D(net1001),
    .RESET_B(net588),
    .Q(\gpio_configure[19][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7176_ (.CLK(clknet_leaf_7_csclk),
    .D(net1440),
    .RESET_B(net590),
    .Q(\gpio_configure[19][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7177_ (.CLK(clknet_leaf_1_csclk),
    .D(net1899),
    .RESET_B(net571),
    .Q(\gpio_configure[31][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7178_ (.CLK(clknet_leaf_11_csclk),
    .D(net1329),
    .RESET_B(net606),
    .Q(\gpio_configure[31][9] ));
 sky130_fd_sc_hd__dfstp_2 _7179_ (.CLK(clknet_leaf_1_csclk),
    .D(net977),
    .SET_B(net571),
    .Q(\gpio_configure[31][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7180_ (.CLK(clknet_leaf_3_csclk),
    .D(net1550),
    .RESET_B(net571),
    .Q(\gpio_configure[31][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7181_ (.CLK(clknet_leaf_3_csclk),
    .D(net751),
    .RESET_B(net571),
    .Q(\gpio_configure[31][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7182_ (.CLK(clknet_leaf_20_csclk),
    .D(net1685),
    .RESET_B(net588),
    .Q(\gpio_configure[20][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7183_ (.CLK(clknet_leaf_20_csclk),
    .D(net1752),
    .RESET_B(net588),
    .Q(\gpio_configure[20][9] ));
 sky130_fd_sc_hd__dfstp_4 _7184_ (.CLK(clknet_leaf_20_csclk),
    .D(net1562),
    .SET_B(net588),
    .Q(\gpio_configure[20][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7185_ (.CLK(clknet_leaf_20_csclk),
    .D(net1059),
    .RESET_B(net591),
    .Q(\gpio_configure[20][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7186_ (.CLK(clknet_leaf_20_csclk),
    .D(net1462),
    .RESET_B(net589),
    .Q(\gpio_configure[20][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7187_ (.CLK(clknet_leaf_1_csclk),
    .D(net1909),
    .RESET_B(net571),
    .Q(\gpio_configure[30][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7188_ (.CLK(clknet_leaf_3_csclk),
    .D(net2351),
    .RESET_B(net574),
    .Q(\gpio_configure[30][9] ));
 sky130_fd_sc_hd__dfstp_2 _7189_ (.CLK(clknet_leaf_0_csclk),
    .D(net949),
    .SET_B(net574),
    .Q(\gpio_configure[30][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7190_ (.CLK(clknet_leaf_3_csclk),
    .D(net1544),
    .RESET_B(net587),
    .Q(\gpio_configure[30][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7191_ (.CLK(clknet_leaf_2_csclk),
    .D(net1398),
    .RESET_B(net573),
    .Q(\gpio_configure[30][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7192_ (.CLK(clknet_leaf_5_csclk),
    .D(net1911),
    .RESET_B(net574),
    .Q(\gpio_configure[21][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7193_ (.CLK(clknet_leaf_9_csclk),
    .D(net1746),
    .RESET_B(net590),
    .Q(\gpio_configure[21][9] ));
 sky130_fd_sc_hd__dfstp_1 _7194_ (.CLK(clknet_leaf_6_csclk),
    .D(net1073),
    .SET_B(net574),
    .Q(\gpio_configure[21][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7195_ (.CLK(clknet_leaf_5_csclk),
    .D(net1031),
    .RESET_B(net574),
    .Q(\gpio_configure[21][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7196_ (.CLK(clknet_leaf_8_csclk),
    .D(net1388),
    .RESET_B(net590),
    .Q(\gpio_configure[21][12] ));
 sky130_fd_sc_hd__dfrtp_4 _7197_ (.CLK(clknet_leaf_15_csclk),
    .D(net1721),
    .RESET_B(net592),
    .Q(\gpio_configure[22][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7198_ (.CLK(clknet_leaf_14_csclk),
    .D(net1249),
    .RESET_B(net592),
    .Q(\gpio_configure[22][9] ));
 sky130_fd_sc_hd__dfstp_4 _7199_ (.CLK(clknet_leaf_14_csclk),
    .D(net1572),
    .SET_B(net592),
    .Q(\gpio_configure[22][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7200_ (.CLK(clknet_leaf_14_csclk),
    .D(net1067),
    .RESET_B(net592),
    .Q(\gpio_configure[22][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7201_ (.CLK(clknet_leaf_14_csclk),
    .D(net1448),
    .RESET_B(net592),
    .Q(\gpio_configure[22][12] ));
 sky130_fd_sc_hd__dfrtp_1 _7202_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0372_),
    .RESET_B(net608),
    .Q(\wbbd_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7203_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0373_),
    .RESET_B(net608),
    .Q(\wbbd_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7204_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0374_),
    .RESET_B(net608),
    .Q(\wbbd_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7205_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0375_),
    .RESET_B(net608),
    .Q(\wbbd_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7206_ (.CLK(clknet_4_9__leaf_wb_clk_i),
    .D(_0376_),
    .RESET_B(net608),
    .Q(\wbbd_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7207_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_0377_),
    .RESET_B(net608),
    .Q(\wbbd_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7208_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0378_),
    .RESET_B(net608),
    .Q(\wbbd_addr[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7209_ (.CLK(clknet_leaf_5_csclk),
    .D(net1907),
    .RESET_B(net573),
    .Q(\gpio_configure[28][8] ));
 sky130_fd_sc_hd__dfrtp_4 _7210_ (.CLK(clknet_leaf_9_csclk),
    .D(net1738),
    .RESET_B(net590),
    .Q(\gpio_configure[28][9] ));
 sky130_fd_sc_hd__dfstp_1 _7211_ (.CLK(clknet_leaf_6_csclk),
    .D(net1043),
    .SET_B(net574),
    .Q(\gpio_configure[28][10] ));
 sky130_fd_sc_hd__dfrtp_4 _7212_ (.CLK(clknet_leaf_5_csclk),
    .D(net1041),
    .RESET_B(net574),
    .Q(\gpio_configure[28][11] ));
 sky130_fd_sc_hd__dfrtp_4 _7213_ (.CLK(clknet_leaf_9_csclk),
    .D(net1444),
    .RESET_B(net590),
    .Q(\gpio_configure[28][12] ));
 sky130_fd_sc_hd__dfrtn_1 _7214_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0384_),
    .RESET_B(_0057_),
    .Q(\hkspi.ldata[0] ));
 sky130_fd_sc_hd__dfrtn_1 _7215_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(net3801),
    .RESET_B(_0058_),
    .Q(\hkspi.ldata[1] ));
 sky130_fd_sc_hd__dfrtn_1 _7216_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0386_),
    .RESET_B(_0059_),
    .Q(\hkspi.ldata[2] ));
 sky130_fd_sc_hd__dfrtn_1 _7217_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(net3804),
    .RESET_B(_0060_),
    .Q(\hkspi.ldata[3] ));
 sky130_fd_sc_hd__dfrtn_1 _7218_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(_0388_),
    .RESET_B(_0061_),
    .Q(\hkspi.ldata[4] ));
 sky130_fd_sc_hd__dfrtn_1 _7219_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(net3807),
    .RESET_B(_0062_),
    .Q(\hkspi.ldata[5] ));
 sky130_fd_sc_hd__dfrtn_1 _7220_ (.CLK_N(clknet_2_2__leaf_mgmt_gpio_in[4]),
    .D(net3799),
    .RESET_B(_0063_),
    .Q(\hkspi.ldata[6] ));
 sky130_fd_sc_hd__dfrtn_1 _7221_ (.CLK_N(clknet_2_1__leaf_mgmt_gpio_in[4]),
    .D(_0391_),
    .RESET_B(_0064_),
    .Q(\hkspi.SDO ));
 sky130_fd_sc_hd__dfrtp_4 _7222_ (.CLK(clknet_leaf_75_csclk),
    .D(net1927),
    .RESET_B(net564),
    .Q(net265));
 sky130_fd_sc_hd__dfstp_2 _7223_ (.CLK(clknet_leaf_75_csclk),
    .D(net1301),
    .SET_B(net564),
    .Q(net259));
 sky130_fd_sc_hd__dfrtp_4 _7224_ (.CLK(clknet_leaf_75_csclk),
    .D(net1925),
    .RESET_B(net564),
    .Q(net260));
 sky130_fd_sc_hd__dfrtp_4 _7225_ (.CLK(clknet_leaf_75_csclk),
    .D(net1303),
    .RESET_B(net564),
    .Q(net261));
 sky130_fd_sc_hd__dfstp_4 _7226_ (.CLK(clknet_leaf_75_csclk),
    .D(net1170),
    .SET_B(net564),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_4 _7227_ (.CLK(clknet_leaf_75_csclk),
    .D(net1580),
    .RESET_B(net565),
    .Q(net263));
 sky130_fd_sc_hd__dfrtp_4 _7228_ (.CLK(clknet_leaf_75_csclk),
    .D(net1363),
    .RESET_B(net564),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_4 _7229_ (.CLK(clknet_leaf_74_csclk),
    .D(net1854),
    .RESET_B(net564),
    .Q(net266));
 sky130_fd_sc_hd__dfstp_4 _7230_ (.CLK(clknet_leaf_74_csclk),
    .D(net1299),
    .SET_B(net564),
    .Q(net267));
 sky130_fd_sc_hd__dfrtp_4 _7231_ (.CLK(clknet_leaf_75_csclk),
    .D(net1145),
    .RESET_B(net564),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_4 _7232_ (.CLK(clknet_leaf_74_csclk),
    .D(net1564),
    .RESET_B(net565),
    .Q(net255));
 sky130_fd_sc_hd__dfstp_4 _7233_ (.CLK(clknet_leaf_74_csclk),
    .D(net1376),
    .SET_B(net565),
    .Q(net256));
 sky130_fd_sc_hd__dfrtp_4 _7234_ (.CLK(clknet_leaf_74_csclk),
    .D(net894),
    .RESET_B(net565),
    .Q(net257));
 sky130_fd_sc_hd__dfstp_2 _7235_ (.CLK(clknet_leaf_70_csclk),
    .D(net1956),
    .SET_B(net566),
    .Q(net276));
 sky130_fd_sc_hd__dfstp_2 _7236_ (.CLK(clknet_leaf_69_csclk),
    .D(net1270),
    .SET_B(net575),
    .Q(net277));
 sky130_fd_sc_hd__dfstp_2 _7237_ (.CLK(clknet_leaf_70_csclk),
    .D(net1199),
    .SET_B(net566),
    .Q(net278));
 sky130_fd_sc_hd__dfstp_2 _7238_ (.CLK(clknet_leaf_70_csclk),
    .D(net1630),
    .SET_B(net566),
    .Q(net279));
 sky130_fd_sc_hd__dfstp_1 _7239_ (.CLK(clknet_leaf_70_csclk),
    .D(net1412),
    .SET_B(net566),
    .Q(net281));
 sky130_fd_sc_hd__dfstp_4 _7240_ (.CLK(clknet_leaf_69_csclk),
    .D(net898),
    .SET_B(net575),
    .Q(net282));
 sky130_fd_sc_hd__dfstp_2 _7241_ (.CLK(clknet_leaf_69_csclk),
    .D(net1470),
    .SET_B(net575),
    .Q(net283));
 sky130_fd_sc_hd__dfstp_4 _7242_ (.CLK(clknet_leaf_69_csclk),
    .D(net2713),
    .SET_B(net575),
    .Q(net284));
 sky130_fd_sc_hd__dfstp_4 _7243_ (.CLK(clknet_leaf_69_csclk),
    .D(net3783),
    .SET_B(net575),
    .Q(net258));
 sky130_fd_sc_hd__dfrtp_4 _7244_ (.CLK(clknet_leaf_54_csclk),
    .D(net1594),
    .RESET_B(net579),
    .Q(net295));
 sky130_fd_sc_hd__dfrtp_4 _7245_ (.CLK(clknet_leaf_54_csclk),
    .D(net1097),
    .RESET_B(net582),
    .Q(net296));
 sky130_fd_sc_hd__dfrtp_4 _7246_ (.CLK(clknet_leaf_54_csclk),
    .D(net2045),
    .RESET_B(net579),
    .Q(net297));
 sky130_fd_sc_hd__dfrtp_4 _7247_ (.CLK(clknet_leaf_53_csclk),
    .D(net1015),
    .RESET_B(net582),
    .Q(net298));
 sky130_fd_sc_hd__dfrtp_2 _7248_ (.CLK(clknet_leaf_76_csclk),
    .D(net1942),
    .RESET_B(net563),
    .Q(reset_reg));
 sky130_fd_sc_hd__dfrtp_4 _7249_ (.CLK(clknet_leaf_76_csclk),
    .D(net1868),
    .RESET_B(net567),
    .Q(irq_spi));
 sky130_fd_sc_hd__dfrtp_2 _7250_ (.CLK(clknet_leaf_74_csclk),
    .D(net1361),
    .RESET_B(net565),
    .Q(serial_bb_clock));
 sky130_fd_sc_hd__dfrtp_4 _7251_ (.CLK(clknet_leaf_72_csclk),
    .D(net1640),
    .RESET_B(net565),
    .Q(serial_bb_load));
 sky130_fd_sc_hd__dfrtp_4 _7252_ (.CLK(clknet_leaf_72_csclk),
    .D(net1203),
    .RESET_B(net565),
    .Q(serial_bb_resetn));
 sky130_fd_sc_hd__dfrtp_1 _7253_ (.CLK(clknet_leaf_72_csclk),
    .D(net2338),
    .RESET_B(net565),
    .Q(serial_bb_data_1));
 sky130_fd_sc_hd__dfrtp_1 _7254_ (.CLK(clknet_leaf_72_csclk),
    .D(net1491),
    .RESET_B(net565),
    .Q(serial_bb_data_2));
 sky130_fd_sc_hd__dfrtp_4 _7255_ (.CLK(clknet_leaf_74_csclk),
    .D(net1274),
    .RESET_B(net569),
    .Q(serial_bb_enable));
 sky130_fd_sc_hd__dfrtp_4 _7256_ (.CLK(clknet_leaf_76_csclk),
    .D(_0426_),
    .RESET_B(net567),
    .Q(serial_xfer));
 sky130_fd_sc_hd__dfrtp_4 _7257_ (.CLK(clknet_leaf_37_csclk),
    .D(net3624),
    .RESET_B(net595),
    .Q(hkspi_disable));
 sky130_fd_sc_hd__dfrtp_4 _7258_ (.CLK(clknet_leaf_37_csclk),
    .D(net2186),
    .RESET_B(net604),
    .Q(\clk1_output_dest[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7259_ (.CLK(clknet_leaf_32_csclk),
    .D(net733),
    .RESET_B(net603),
    .Q(\clk1_output_dest[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7260_ (.CLK(clknet_leaf_37_csclk),
    .D(net1664),
    .RESET_B(net604),
    .Q(\clk2_output_dest[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7261_ (.CLK(clknet_leaf_33_csclk),
    .D(net973),
    .RESET_B(net603),
    .Q(\clk2_output_dest[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7262_ (.CLK(clknet_leaf_37_csclk),
    .D(net1093),
    .RESET_B(net604),
    .Q(trap_output_dest));
 sky130_fd_sc_hd__dfrtp_1 _7263_ (.CLK(clknet_leaf_72_csclk),
    .D(net1915),
    .RESET_B(net569),
    .Q(irq_1_inputsrc));
 sky130_fd_sc_hd__dfrtp_1 _7264_ (.CLK(clknet_leaf_72_csclk),
    .D(net1327),
    .RESET_B(net567),
    .Q(irq_2_inputsrc));
 sky130_fd_sc_hd__dfrtp_1 _7265_ (.CLK(clknet_leaf_76_csclk),
    .D(net1938),
    .RESET_B(net563),
    .Q(\mgmt_gpio_data[32] ));
 sky130_fd_sc_hd__dfrtp_1 _7266_ (.CLK(clknet_leaf_76_csclk),
    .D(net1309),
    .RESET_B(net563),
    .Q(\mgmt_gpio_data[33] ));
 sky130_fd_sc_hd__dfrtp_1 _7267_ (.CLK(clknet_3_7_0_csclk),
    .D(net1510),
    .RESET_B(net605),
    .Q(\mgmt_gpio_data[34] ));
 sky130_fd_sc_hd__dfrtp_1 _7268_ (.CLK(clknet_leaf_1_csclk),
    .D(net1574),
    .RESET_B(net571),
    .Q(\mgmt_gpio_data[35] ));
 sky130_fd_sc_hd__dfrtp_1 _7269_ (.CLK(clknet_leaf_30_csclk),
    .D(net1251),
    .RESET_B(net600),
    .Q(\mgmt_gpio_data[36] ));
 sky130_fd_sc_hd__dfrtp_1 _7270_ (.CLK(clknet_leaf_30_csclk),
    .D(net2082),
    .RESET_B(net602),
    .Q(\mgmt_gpio_data[37] ));
 sky130_fd_sc_hd__dfrtp_1 _7271_ (.CLK(clknet_leaf_53_csclk),
    .D(net1676),
    .RESET_B(net582),
    .Q(\mgmt_gpio_data_buf[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7272_ (.CLK(clknet_leaf_52_csclk),
    .D(net1125),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data_buf[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7273_ (.CLK(clknet_leaf_52_csclk),
    .D(net2057),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data_buf[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7274_ (.CLK(clknet_leaf_52_csclk),
    .D(net911),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data_buf[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7275_ (.CLK(clknet_leaf_49_csclk),
    .D(net776),
    .RESET_B(net583),
    .Q(\mgmt_gpio_data_buf[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7276_ (.CLK(clknet_leaf_48_csclk),
    .D(net941),
    .RESET_B(net583),
    .Q(\mgmt_gpio_data_buf[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7277_ (.CLK(clknet_leaf_52_csclk),
    .D(net1380),
    .RESET_B(net580),
    .Q(\mgmt_gpio_data_buf[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7278_ (.CLK(clknet_leaf_52_csclk),
    .D(net1061),
    .RESET_B(net582),
    .Q(\mgmt_gpio_data_buf[7] ));
 sky130_fd_sc_hd__dfstp_2 _7279_ (.CLK(clknet_leaf_58_csclk),
    .D(net1662),
    .SET_B(net576),
    .Q(\gpio_configure[0][0] ));
 sky130_fd_sc_hd__dfstp_2 _7280_ (.CLK(clknet_leaf_58_csclk),
    .D(net1217),
    .SET_B(net576),
    .Q(\gpio_configure[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7281_ (.CLK(clknet_leaf_59_csclk),
    .D(net2149),
    .RESET_B(net576),
    .Q(\gpio_configure[0][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7282_ (.CLK(clknet_leaf_58_csclk),
    .D(net2487),
    .RESET_B(net576),
    .Q(\gpio_configure[0][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7283_ (.CLK(clknet_leaf_58_csclk),
    .D(net725),
    .RESET_B(net576),
    .Q(\gpio_configure[0][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7284_ (.CLK(clknet_leaf_58_csclk),
    .D(net1548),
    .RESET_B(net579),
    .Q(\gpio_configure[0][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7285_ (.CLK(clknet_leaf_57_csclk),
    .D(net1464),
    .RESET_B(net579),
    .Q(\gpio_configure[0][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7286_ (.CLK(clknet_leaf_58_csclk),
    .D(net2845),
    .RESET_B(net579),
    .Q(\gpio_configure[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _7287_ (.CLK(clknet_leaf_69_csclk),
    .D(net1691),
    .SET_B(net575),
    .Q(\gpio_configure[1][0] ));
 sky130_fd_sc_hd__dfstp_4 _7288_ (.CLK(clknet_leaf_69_csclk),
    .D(net1256),
    .SET_B(net575),
    .Q(\gpio_configure[1][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7289_ (.CLK(clknet_leaf_59_csclk),
    .D(net2096),
    .RESET_B(net575),
    .Q(\gpio_configure[1][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7290_ (.CLK(clknet_leaf_55_csclk),
    .D(net919),
    .RESET_B(net581),
    .Q(\gpio_configure[1][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7291_ (.CLK(clknet_leaf_60_csclk),
    .D(net709),
    .RESET_B(net577),
    .Q(\gpio_configure[1][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7292_ (.CLK(clknet_leaf_54_csclk),
    .D(net1514),
    .RESET_B(net579),
    .Q(\gpio_configure[1][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7293_ (.CLK(clknet_leaf_54_csclk),
    .D(net1343),
    .RESET_B(net579),
    .Q(\gpio_configure[1][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7294_ (.CLK(clknet_leaf_54_csclk),
    .D(net1017),
    .RESET_B(net579),
    .Q(\gpio_configure[1][7] ));
 sky130_fd_sc_hd__dfstp_2 _7295_ (.CLK(clknet_leaf_60_csclk),
    .D(net1635),
    .SET_B(net577),
    .Q(\gpio_configure[2][0] ));
 sky130_fd_sc_hd__dfstp_2 _7296_ (.CLK(clknet_leaf_60_csclk),
    .D(net1161),
    .SET_B(net577),
    .Q(\gpio_configure[2][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7297_ (.CLK(clknet_leaf_60_csclk),
    .D(net2065),
    .RESET_B(net577),
    .Q(\gpio_configure[2][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7298_ (.CLK(clknet_leaf_55_csclk),
    .D(net931),
    .RESET_B(net580),
    .Q(\gpio_configure[2][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7299_ (.CLK(clknet_leaf_57_csclk),
    .D(net753),
    .RESET_B(net576),
    .Q(\gpio_configure[2][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7300_ (.CLK(clknet_leaf_55_csclk),
    .D(net1524),
    .RESET_B(net582),
    .Q(\gpio_configure[2][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7301_ (.CLK(clknet_leaf_51_csclk),
    .D(net1432),
    .RESET_B(net580),
    .Q(\gpio_configure[2][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7302_ (.CLK(clknet_leaf_55_csclk),
    .D(net1083),
    .RESET_B(net579),
    .Q(\gpio_configure[2][7] ));
 sky130_fd_sc_hd__dfstp_4 _7303_ (.CLK(clknet_leaf_58_csclk),
    .D(net1654),
    .SET_B(net576),
    .Q(\gpio_configure[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _7304_ (.CLK(clknet_leaf_56_csclk),
    .D(net1213),
    .RESET_B(net577),
    .Q(\gpio_configure[3][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7305_ (.CLK(clknet_leaf_59_csclk),
    .D(net2078),
    .RESET_B(net576),
    .Q(\gpio_configure[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7306_ (.CLK(clknet_leaf_55_csclk),
    .D(net2391),
    .RESET_B(net580),
    .Q(\gpio_configure[3][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7307_ (.CLK(clknet_leaf_59_csclk),
    .D(net713),
    .RESET_B(net576),
    .Q(\gpio_configure[3][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7308_ (.CLK(clknet_leaf_56_csclk),
    .D(net1546),
    .RESET_B(net581),
    .Q(\gpio_configure[3][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7309_ (.CLK(clknet_leaf_58_csclk),
    .D(net1416),
    .RESET_B(net579),
    .Q(\gpio_configure[3][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7310_ (.CLK(clknet_leaf_56_csclk),
    .D(net1139),
    .RESET_B(net581),
    .Q(\gpio_configure[3][7] ));
 sky130_fd_sc_hd__dfstp_4 _7311_ (.CLK(clknet_leaf_48_csclk),
    .D(_0481_),
    .SET_B(net584),
    .Q(\gpio_configure[4][0] ));
 sky130_fd_sc_hd__dfstp_2 _7312_ (.CLK(clknet_leaf_47_csclk),
    .D(net1229),
    .SET_B(net584),
    .Q(\gpio_configure[4][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7313_ (.CLK(clknet_leaf_48_csclk),
    .D(net890),
    .RESET_B(net583),
    .Q(\gpio_configure[4][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7314_ (.CLK(clknet_leaf_51_csclk),
    .D(net969),
    .RESET_B(net580),
    .Q(\gpio_configure[4][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7315_ (.CLK(clknet_leaf_50_csclk),
    .D(net762),
    .RESET_B(net583),
    .Q(\gpio_configure[4][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7316_ (.CLK(clknet_leaf_50_csclk),
    .D(net1622),
    .RESET_B(net580),
    .Q(\gpio_configure[4][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7317_ (.CLK(clknet_leaf_50_csclk),
    .D(net1489),
    .RESET_B(net580),
    .Q(\gpio_configure[4][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7318_ (.CLK(clknet_leaf_47_csclk),
    .D(net1109),
    .RESET_B(net584),
    .Q(\gpio_configure[4][7] ));
 sky130_fd_sc_hd__dfstp_4 _7319_ (.CLK(clknet_leaf_61_csclk),
    .D(net1660),
    .SET_B(net578),
    .Q(\gpio_configure[5][0] ));
 sky130_fd_sc_hd__dfstp_4 _7320_ (.CLK(clknet_leaf_61_csclk),
    .D(net1201),
    .SET_B(net578),
    .Q(\gpio_configure[5][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7321_ (.CLK(clknet_leaf_63_csclk),
    .D(net1057),
    .RESET_B(net586),
    .Q(\gpio_configure[5][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7322_ (.CLK(clknet_leaf_49_csclk),
    .D(net1190),
    .RESET_B(net583),
    .Q(\gpio_configure[5][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7323_ (.CLK(clknet_leaf_61_csclk),
    .D(net723),
    .RESET_B(net578),
    .Q(\gpio_configure[5][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7324_ (.CLK(clknet_leaf_51_csclk),
    .D(net1526),
    .RESET_B(net580),
    .Q(\gpio_configure[5][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7325_ (.CLK(clknet_leaf_49_csclk),
    .D(net1466),
    .RESET_B(net583),
    .Q(\gpio_configure[5][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7326_ (.CLK(clknet_leaf_50_csclk),
    .D(net1195),
    .RESET_B(net583),
    .Q(\gpio_configure[5][7] ));
 sky130_fd_sc_hd__dfstp_2 _7327_ (.CLK(clknet_leaf_59_csclk),
    .D(net1848),
    .SET_B(net575),
    .Q(\gpio_configure[6][0] ));
 sky130_fd_sc_hd__dfstp_4 _7328_ (.CLK(clknet_leaf_59_csclk),
    .D(net1157),
    .SET_B(net576),
    .Q(\gpio_configure[6][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7329_ (.CLK(clknet_leaf_59_csclk),
    .D(net2049),
    .RESET_B(net576),
    .Q(\gpio_configure[6][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7330_ (.CLK(clknet_leaf_54_csclk),
    .D(net868),
    .RESET_B(net582),
    .Q(\gpio_configure[6][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7331_ (.CLK(clknet_leaf_69_csclk),
    .D(net1341),
    .RESET_B(net575),
    .Q(\gpio_configure[6][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7332_ (.CLK(clknet_leaf_54_csclk),
    .D(net1516),
    .RESET_B(net579),
    .Q(\gpio_configure[6][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7333_ (.CLK(clknet_leaf_53_csclk),
    .D(net1446),
    .RESET_B(net579),
    .Q(\gpio_configure[6][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7334_ (.CLK(clknet_leaf_54_csclk),
    .D(net1013),
    .RESET_B(net579),
    .Q(\gpio_configure[6][7] ));
 sky130_fd_sc_hd__dfstp_2 _7335_ (.CLK(clknet_leaf_60_csclk),
    .D(net1642),
    .SET_B(net577),
    .Q(\gpio_configure[7][0] ));
 sky130_fd_sc_hd__dfstp_4 _7336_ (.CLK(clknet_leaf_51_csclk),
    .D(net2939),
    .SET_B(net580),
    .Q(\gpio_configure[7][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7337_ (.CLK(clknet_leaf_60_csclk),
    .D(net2061),
    .RESET_B(net578),
    .Q(\gpio_configure[7][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7338_ (.CLK(clknet_leaf_41_csclk),
    .D(net2429),
    .RESET_B(net594),
    .Q(\gpio_configure[7][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7339_ (.CLK(clknet_leaf_61_csclk),
    .D(net731),
    .RESET_B(net578),
    .Q(\gpio_configure[7][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7340_ (.CLK(clknet_leaf_46_csclk),
    .D(net2319),
    .RESET_B(net584),
    .Q(\gpio_configure[7][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7341_ (.CLK(clknet_leaf_50_csclk),
    .D(net1501),
    .RESET_B(net580),
    .Q(\gpio_configure[7][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7342_ (.CLK(clknet_leaf_41_csclk),
    .D(net2889),
    .RESET_B(net594),
    .Q(\gpio_configure[7][7] ));
 sky130_fd_sc_hd__dfstp_2 _7343_ (.CLK(clknet_leaf_68_csclk),
    .D(net1940),
    .SET_B(net577),
    .Q(\gpio_configure[8][0] ));
 sky130_fd_sc_hd__dfstp_2 _7344_ (.CLK(clknet_leaf_60_csclk),
    .D(net1186),
    .SET_B(net578),
    .Q(\gpio_configure[8][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7345_ (.CLK(clknet_leaf_68_csclk),
    .D(net1184),
    .RESET_B(net577),
    .Q(\gpio_configure[8][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7346_ (.CLK(clknet_leaf_51_csclk),
    .D(net630),
    .RESET_B(net580),
    .Q(\gpio_configure[8][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7347_ (.CLK(clknet_leaf_60_csclk),
    .D(net711),
    .RESET_B(net577),
    .Q(\gpio_configure[8][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7348_ (.CLK(clknet_leaf_50_csclk),
    .D(net1628),
    .RESET_B(net580),
    .Q(\gpio_configure[8][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7349_ (.CLK(clknet_leaf_55_csclk),
    .D(net1408),
    .RESET_B(net581),
    .Q(\gpio_configure[8][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7350_ (.CLK(clknet_leaf_51_csclk),
    .D(net1085),
    .RESET_B(net581),
    .Q(\gpio_configure[8][7] ));
 sky130_fd_sc_hd__dfstp_2 _7351_ (.CLK(clknet_leaf_18_csclk),
    .D(net1913),
    .SET_B(net598),
    .Q(\gpio_configure[9][0] ));
 sky130_fd_sc_hd__dfstp_2 _7352_ (.CLK(clknet_leaf_27_csclk),
    .D(net1736),
    .SET_B(net598),
    .Q(\gpio_configure[9][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7353_ (.CLK(clknet_leaf_50_csclk),
    .D(net2200),
    .RESET_B(net583),
    .Q(\gpio_configure[9][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7354_ (.CLK(clknet_leaf_38_csclk),
    .D(net2528),
    .RESET_B(net595),
    .Q(\gpio_configure[9][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7355_ (.CLK(clknet_leaf_27_csclk),
    .D(net2736),
    .RESET_B(net599),
    .Q(\gpio_configure[9][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7356_ (.CLK(clknet_leaf_49_csclk),
    .D(net1672),
    .RESET_B(net583),
    .Q(\gpio_configure[9][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7357_ (.CLK(clknet_leaf_49_csclk),
    .D(net1479),
    .RESET_B(net583),
    .Q(\gpio_configure[9][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7358_ (.CLK(clknet_leaf_41_csclk),
    .D(net1215),
    .RESET_B(net594),
    .Q(\gpio_configure[9][7] ));
 sky130_fd_sc_hd__dfstp_2 _7359_ (.CLK(clknet_leaf_59_csclk),
    .D(net1638),
    .SET_B(net575),
    .Q(\gpio_configure[10][0] ));
 sky130_fd_sc_hd__dfstp_2 _7360_ (.CLK(clknet_leaf_68_csclk),
    .D(net1311),
    .SET_B(net577),
    .Q(\gpio_configure[10][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7361_ (.CLK(clknet_leaf_68_csclk),
    .D(net2587),
    .RESET_B(net575),
    .Q(\gpio_configure[10][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7362_ (.CLK(clknet_leaf_54_csclk),
    .D(net2270),
    .RESET_B(net579),
    .Q(\gpio_configure[10][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7363_ (.CLK(clknet_leaf_69_csclk),
    .D(net1351),
    .RESET_B(net575),
    .Q(\gpio_configure[10][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7364_ (.CLK(clknet_leaf_55_csclk),
    .D(net1522),
    .RESET_B(net581),
    .Q(\gpio_configure[10][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7365_ (.CLK(clknet_leaf_54_csclk),
    .D(net1357),
    .RESET_B(net579),
    .Q(\gpio_configure[10][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7366_ (.CLK(clknet_leaf_54_csclk),
    .D(net2797),
    .RESET_B(net579),
    .Q(\gpio_configure[10][7] ));
 sky130_fd_sc_hd__dfstp_4 _7367_ (.CLK(clknet_leaf_38_csclk),
    .D(net3590),
    .SET_B(net595),
    .Q(\gpio_configure[11][0] ));
 sky130_fd_sc_hd__dfstp_1 _7368_ (.CLK(clknet_leaf_45_csclk),
    .D(net699),
    .SET_B(net586),
    .Q(\gpio_configure[11][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7369_ (.CLK(clknet_leaf_62_csclk),
    .D(net1039),
    .RESET_B(net586),
    .Q(\gpio_configure[11][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7370_ (.CLK(clknet_leaf_38_csclk),
    .D(net913),
    .RESET_B(net595),
    .Q(\gpio_configure[11][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7371_ (.CLK(clknet_leaf_24_csclk),
    .D(net1331),
    .RESET_B(net593),
    .Q(\gpio_configure[11][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7372_ (.CLK(clknet_leaf_50_csclk),
    .D(net1602),
    .RESET_B(net583),
    .Q(\gpio_configure[11][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7373_ (.CLK(clknet_leaf_49_csclk),
    .D(net1508),
    .RESET_B(net583),
    .Q(\gpio_configure[11][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7374_ (.CLK(clknet_leaf_47_csclk),
    .D(net1121),
    .RESET_B(net584),
    .Q(\gpio_configure[11][7] ));
 sky130_fd_sc_hd__dfstp_2 _7375_ (.CLK(clknet_leaf_23_csclk),
    .D(net1887),
    .SET_B(net593),
    .Q(\gpio_configure[12][0] ));
 sky130_fd_sc_hd__dfstp_4 _7376_ (.CLK(clknet_leaf_27_csclk),
    .D(net1725),
    .SET_B(net599),
    .Q(\gpio_configure[12][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7377_ (.CLK(clknet_leaf_24_csclk),
    .D(net2216),
    .RESET_B(net593),
    .Q(\gpio_configure[12][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7378_ (.CLK(clknet_leaf_38_csclk),
    .D(net2521),
    .RESET_B(net595),
    .Q(\gpio_configure[12][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7379_ (.CLK(clknet_leaf_24_csclk),
    .D(net1335),
    .RESET_B(net593),
    .Q(\gpio_configure[12][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7380_ (.CLK(clknet_leaf_48_csclk),
    .D(net1620),
    .RESET_B(net583),
    .Q(\gpio_configure[12][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7381_ (.CLK(clknet_leaf_49_csclk),
    .D(net1487),
    .RESET_B(net583),
    .Q(\gpio_configure[12][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7382_ (.CLK(clknet_leaf_46_csclk),
    .D(net2236),
    .RESET_B(net584),
    .Q(\gpio_configure[12][7] ));
 sky130_fd_sc_hd__dfstp_4 _7383_ (.CLK(clknet_leaf_38_csclk),
    .D(net1856),
    .SET_B(net595),
    .Q(\gpio_configure[13][0] ));
 sky130_fd_sc_hd__dfstp_2 _7384_ (.CLK(clknet_leaf_48_csclk),
    .D(net674),
    .SET_B(net584),
    .Q(\gpio_configure[13][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7385_ (.CLK(clknet_leaf_48_csclk),
    .D(net888),
    .RESET_B(net583),
    .Q(\gpio_configure[13][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7386_ (.CLK(clknet_leaf_38_csclk),
    .D(net915),
    .RESET_B(net596),
    .Q(\gpio_configure[13][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7387_ (.CLK(clknet_leaf_38_csclk),
    .D(net1262),
    .RESET_B(net595),
    .Q(\gpio_configure[13][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7388_ (.CLK(clknet_leaf_48_csclk),
    .D(net1590),
    .RESET_B(net583),
    .Q(\gpio_configure[13][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7389_ (.CLK(clknet_leaf_48_csclk),
    .D(net1418),
    .RESET_B(net584),
    .Q(\gpio_configure[13][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7390_ (.CLK(clknet_leaf_47_csclk),
    .D(net1207),
    .RESET_B(net584),
    .Q(\gpio_configure[13][7] ));
 sky130_fd_sc_hd__dfstp_4 _7391_ (.CLK(clknet_leaf_24_csclk),
    .D(net2665),
    .SET_B(net593),
    .Q(\gpio_configure[14][0] ));
 sky130_fd_sc_hd__dfstp_4 _7392_ (.CLK(clknet_leaf_25_csclk),
    .D(net2851),
    .SET_B(net599),
    .Q(\gpio_configure[14][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7393_ (.CLK(clknet_leaf_23_csclk),
    .D(net1558),
    .RESET_B(net593),
    .Q(\gpio_configure[14][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7394_ (.CLK(clknet_leaf_37_csclk),
    .D(net2400),
    .RESET_B(net604),
    .Q(\gpio_configure[14][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7395_ (.CLK(clknet_leaf_18_csclk),
    .D(net2769),
    .RESET_B(net598),
    .Q(\gpio_configure[14][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7396_ (.CLK(clknet_leaf_46_csclk),
    .D(net1610),
    .RESET_B(net584),
    .Q(\gpio_configure[14][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7397_ (.CLK(clknet_leaf_46_csclk),
    .D(net1438),
    .RESET_B(net584),
    .Q(\gpio_configure[14][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7398_ (.CLK(clknet_leaf_47_csclk),
    .D(net1235),
    .RESET_B(net585),
    .Q(\gpio_configure[14][7] ));
 sky130_fd_sc_hd__dfstp_4 _7399_ (.CLK(clknet_leaf_63_csclk),
    .D(net1758),
    .SET_B(net586),
    .Q(\gpio_configure[15][0] ));
 sky130_fd_sc_hd__dfstp_4 _7400_ (.CLK(clknet_leaf_62_csclk),
    .D(net1349),
    .SET_B(net578),
    .Q(\gpio_configure[15][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7401_ (.CLK(clknet_leaf_62_csclk),
    .D(net1027),
    .RESET_B(net586),
    .Q(\gpio_configure[15][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7402_ (.CLK(clknet_leaf_41_csclk),
    .D(net985),
    .RESET_B(net594),
    .Q(\gpio_configure[15][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7403_ (.CLK(clknet_leaf_45_csclk),
    .D(net1353),
    .RESET_B(net593),
    .Q(\gpio_configure[15][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7404_ (.CLK(clknet_leaf_55_csclk),
    .D(net1528),
    .RESET_B(net581),
    .Q(\gpio_configure[15][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7405_ (.CLK(clknet_leaf_48_csclk),
    .D(net1420),
    .RESET_B(net584),
    .Q(\gpio_configure[15][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7406_ (.CLK(clknet_leaf_55_csclk),
    .D(net1079),
    .RESET_B(net581),
    .Q(\gpio_configure[15][7] ));
 sky130_fd_sc_hd__dfstp_4 _7407_ (.CLK(clknet_leaf_67_csclk),
    .D(net1954),
    .SET_B(net577),
    .Q(\gpio_configure[16][0] ));
 sky130_fd_sc_hd__dfstp_2 _7408_ (.CLK(clknet_leaf_67_csclk),
    .D(net1297),
    .SET_B(net577),
    .Q(\gpio_configure[16][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7409_ (.CLK(clknet_leaf_67_csclk),
    .D(net2591),
    .RESET_B(net577),
    .Q(\gpio_configure[16][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7410_ (.CLK(clknet_leaf_51_csclk),
    .D(net2483),
    .RESET_B(net581),
    .Q(\gpio_configure[16][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7411_ (.CLK(clknet_leaf_61_csclk),
    .D(net729),
    .RESET_B(net578),
    .Q(\gpio_configure[16][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7412_ (.CLK(clknet_leaf_51_csclk),
    .D(net1534),
    .RESET_B(net581),
    .Q(\gpio_configure[16][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7413_ (.CLK(clknet_leaf_50_csclk),
    .D(net1497),
    .RESET_B(net581),
    .Q(\gpio_configure[16][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7414_ (.CLK(clknet_leaf_50_csclk),
    .D(net1227),
    .RESET_B(net581),
    .Q(\gpio_configure[16][7] ));
 sky130_fd_sc_hd__dfstp_2 _7415_ (.CLK(clknet_leaf_22_csclk),
    .D(net1727),
    .SET_B(net593),
    .Q(\gpio_configure[17][0] ));
 sky130_fd_sc_hd__dfstp_2 _7416_ (.CLK(clknet_leaf_66_csclk),
    .D(net1394),
    .SET_B(net586),
    .Q(\gpio_configure[17][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7417_ (.CLK(clknet_leaf_66_csclk),
    .D(net1174),
    .RESET_B(net586),
    .Q(\gpio_configure[17][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7418_ (.CLK(clknet_leaf_41_csclk),
    .D(net991),
    .RESET_B(net594),
    .Q(\gpio_configure[17][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7419_ (.CLK(clknet_leaf_23_csclk),
    .D(net1392),
    .RESET_B(net593),
    .Q(\gpio_configure[17][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7420_ (.CLK(clknet_leaf_46_csclk),
    .D(net1604),
    .RESET_B(net584),
    .Q(\gpio_configure[17][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7421_ (.CLK(clknet_leaf_46_csclk),
    .D(net1434),
    .RESET_B(net585),
    .Q(\gpio_configure[17][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7422_ (.CLK(clknet_leaf_50_csclk),
    .D(net1225),
    .RESET_B(net583),
    .Q(\gpio_configure[17][7] ));
 sky130_fd_sc_hd__dfstp_1 _7423_ (.CLK(clknet_leaf_23_csclk),
    .D(net1891),
    .SET_B(net593),
    .Q(\gpio_configure[18][0] ));
 sky130_fd_sc_hd__dfstp_2 _7424_ (.CLK(clknet_leaf_62_csclk),
    .D(net1337),
    .SET_B(net586),
    .Q(\gpio_configure[18][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7425_ (.CLK(clknet_leaf_64_csclk),
    .D(net1123),
    .RESET_B(net586),
    .Q(\gpio_configure[18][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7426_ (.CLK(clknet_leaf_40_csclk),
    .D(net1055),
    .RESET_B(net594),
    .Q(\gpio_configure[18][3] ));
 sky130_fd_sc_hd__dfrtp_2 _7427_ (.CLK(clknet_leaf_23_csclk),
    .D(net1386),
    .RESET_B(net593),
    .Q(\gpio_configure[18][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7428_ (.CLK(clknet_leaf_47_csclk),
    .D(net2175),
    .RESET_B(net584),
    .Q(\gpio_configure[18][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7429_ (.CLK(clknet_leaf_49_csclk),
    .D(net1475),
    .RESET_B(net583),
    .Q(\gpio_configure[18][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7430_ (.CLK(clknet_leaf_41_csclk),
    .D(net1205),
    .RESET_B(net594),
    .Q(\gpio_configure[18][7] ));
 sky130_fd_sc_hd__dfstp_2 _7431_ (.CLK(clknet_leaf_44_csclk),
    .D(net1883),
    .SET_B(net593),
    .Q(\gpio_configure[19][0] ));
 sky130_fd_sc_hd__dfstp_2 _7432_ (.CLK(clknet_leaf_45_csclk),
    .D(net1715),
    .SET_B(net593),
    .Q(\gpio_configure[19][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7433_ (.CLK(clknet_leaf_63_csclk),
    .D(net1045),
    .RESET_B(net586),
    .Q(\gpio_configure[19][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7434_ (.CLK(clknet_leaf_40_csclk),
    .D(net1065),
    .RESET_B(net594),
    .Q(\gpio_configure[19][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7435_ (.CLK(clknet_leaf_44_csclk),
    .D(net1382),
    .RESET_B(net593),
    .Q(\gpio_configure[19][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7436_ (.CLK(clknet_leaf_40_csclk),
    .D(net876),
    .RESET_B(net594),
    .Q(\gpio_configure[19][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7437_ (.CLK(clknet_leaf_48_csclk),
    .D(net1430),
    .RESET_B(net584),
    .Q(\gpio_configure[19][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7438_ (.CLK(clknet_leaf_47_csclk),
    .D(net2160),
    .RESET_B(net585),
    .Q(\gpio_configure[19][7] ));
 sky130_fd_sc_hd__dfstp_4 _7439_ (.CLK(clknet_leaf_16_csclk),
    .D(net1707),
    .SET_B(net601),
    .Q(\gpio_configure[20][0] ));
 sky130_fd_sc_hd__dfstp_4 _7440_ (.CLK(clknet_leaf_28_csclk),
    .D(net1740),
    .SET_B(net600),
    .Q(\gpio_configure[20][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7441_ (.CLK(clknet_leaf_17_csclk),
    .D(net1568),
    .RESET_B(net598),
    .Q(\gpio_configure[20][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7442_ (.CLK(clknet_leaf_29_csclk),
    .D(net870),
    .RESET_B(net600),
    .Q(\gpio_configure[20][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7443_ (.CLK(clknet_leaf_16_csclk),
    .D(net772),
    .RESET_B(net601),
    .Q(\gpio_configure[20][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7444_ (.CLK(clknet_leaf_31_csclk),
    .D(net2126),
    .RESET_B(net599),
    .Q(\gpio_configure[20][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7445_ (.CLK(clknet_leaf_33_csclk),
    .D(net747),
    .RESET_B(net605),
    .Q(\gpio_configure[20][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7446_ (.CLK(clknet_leaf_32_csclk),
    .D(net2103),
    .RESET_B(net603),
    .Q(\gpio_configure[20][7] ));
 sky130_fd_sc_hd__dfstp_4 _7447_ (.CLK(clknet_leaf_17_csclk),
    .D(net2685),
    .SET_B(net598),
    .Q(\gpio_configure[21][0] ));
 sky130_fd_sc_hd__dfstp_4 _7448_ (.CLK(clknet_leaf_28_csclk),
    .D(net3284),
    .SET_B(net600),
    .Q(\gpio_configure[21][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7449_ (.CLK(clknet_leaf_16_csclk),
    .D(net935),
    .RESET_B(net601),
    .Q(\gpio_configure[21][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7450_ (.CLK(clknet_leaf_16_csclk),
    .D(net1053),
    .RESET_B(net601),
    .Q(\gpio_configure[21][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7451_ (.CLK(clknet_leaf_16_csclk),
    .D(net766),
    .RESET_B(net601),
    .Q(\gpio_configure[21][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7452_ (.CLK(clknet_leaf_43_csclk),
    .D(net2193),
    .RESET_B(net596),
    .Q(\gpio_configure[21][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7453_ (.CLK(clknet_leaf_43_csclk),
    .D(net745),
    .RESET_B(net596),
    .Q(\gpio_configure[21][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7454_ (.CLK(clknet_leaf_43_csclk),
    .D(net1182),
    .RESET_B(net596),
    .Q(\gpio_configure[21][7] ));
 sky130_fd_sc_hd__dfstp_2 _7455_ (.CLK(clknet_leaf_24_csclk),
    .D(net1861),
    .SET_B(net593),
    .Q(\gpio_configure[22][0] ));
 sky130_fd_sc_hd__dfstp_2 _7456_ (.CLK(clknet_leaf_46_csclk),
    .D(net688),
    .SET_B(net585),
    .Q(\gpio_configure[22][1] ));
 sky130_fd_sc_hd__dfrtp_2 _7457_ (.CLK(clknet_leaf_63_csclk),
    .D(net1037),
    .RESET_B(net586),
    .Q(\gpio_configure[22][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7458_ (.CLK(clknet_leaf_25_csclk),
    .D(net925),
    .RESET_B(net593),
    .Q(\gpio_configure[22][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7459_ (.CLK(clknet_leaf_24_csclk),
    .D(net1317),
    .RESET_B(net593),
    .Q(\gpio_configure[22][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7460_ (.CLK(clknet_leaf_46_csclk),
    .D(net963),
    .RESET_B(net584),
    .Q(\gpio_configure[22][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7461_ (.CLK(clknet_leaf_50_csclk),
    .D(net1414),
    .RESET_B(net585),
    .Q(\gpio_configure[22][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7462_ (.CLK(clknet_leaf_42_csclk),
    .D(net1127),
    .RESET_B(net594),
    .Q(\gpio_configure[22][7] ));
 sky130_fd_sc_hd__dfstp_4 _7463_ (.CLK(clknet_leaf_31_csclk),
    .D(net3575),
    .SET_B(net599),
    .Q(\gpio_configure[23][0] ));
 sky130_fd_sc_hd__dfstp_4 _7464_ (.CLK(clknet_leaf_30_csclk),
    .D(net1646),
    .SET_B(net600),
    .Q(\gpio_configure[23][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7465_ (.CLK(clknet_leaf_27_csclk),
    .D(net947),
    .RESET_B(net602),
    .Q(\gpio_configure[23][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7466_ (.CLK(clknet_leaf_30_csclk),
    .D(net862),
    .RESET_B(net600),
    .Q(\gpio_configure[23][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7467_ (.CLK(clknet_leaf_16_csclk),
    .D(net1365),
    .RESET_B(net601),
    .Q(\gpio_configure[23][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7468_ (.CLK(clknet_leaf_31_csclk),
    .D(net2107),
    .RESET_B(net599),
    .Q(\gpio_configure[23][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7469_ (.CLK(clknet_leaf_32_csclk),
    .D(net737),
    .RESET_B(net603),
    .Q(\gpio_configure[23][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7470_ (.CLK(clknet_leaf_32_csclk),
    .D(net1168),
    .RESET_B(net603),
    .Q(\gpio_configure[23][7] ));
 sky130_fd_sc_hd__dfstp_2 _7471_ (.CLK(clknet_leaf_23_csclk),
    .D(net1895),
    .SET_B(net597),
    .Q(\gpio_configure[24][0] ));
 sky130_fd_sc_hd__dfstp_2 _7472_ (.CLK(clknet_leaf_61_csclk),
    .D(net1193),
    .SET_B(net578),
    .Q(\gpio_configure[24][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7473_ (.CLK(clknet_leaf_61_csclk),
    .D(net2053),
    .RESET_B(net577),
    .Q(\gpio_configure[24][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7474_ (.CLK(clknet_leaf_33_csclk),
    .D(net1025),
    .RESET_B(net603),
    .Q(\gpio_configure[24][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7475_ (.CLK(clknet_leaf_27_csclk),
    .D(net1367),
    .RESET_B(net599),
    .Q(\gpio_configure[24][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7476_ (.CLK(clknet_leaf_62_csclk),
    .D(net1682),
    .RESET_B(net581),
    .Q(\gpio_configure[24][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7477_ (.CLK(clknet_leaf_50_csclk),
    .D(net1495),
    .RESET_B(net585),
    .Q(\gpio_configure[24][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7478_ (.CLK(clknet_leaf_50_csclk),
    .D(net1231),
    .RESET_B(net581),
    .Q(\gpio_configure[24][7] ));
 sky130_fd_sc_hd__dfstp_2 _7479_ (.CLK(clknet_leaf_25_csclk),
    .D(net1099),
    .SET_B(net599),
    .Q(\gpio_configure[25][0] ));
 sky130_fd_sc_hd__dfstp_4 _7480_ (.CLK(clknet_leaf_31_csclk),
    .D(_0650_),
    .SET_B(net600),
    .Q(\gpio_configure[25][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7481_ (.CLK(clknet_leaf_26_csclk),
    .D(net2118),
    .RESET_B(net599),
    .Q(\gpio_configure[25][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7482_ (.CLK(clknet_leaf_31_csclk),
    .D(net856),
    .RESET_B(net605),
    .Q(\gpio_configure[25][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7483_ (.CLK(clknet_leaf_28_csclk),
    .D(net1406),
    .RESET_B(net600),
    .Q(\gpio_configure[25][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7484_ (.CLK(clknet_leaf_32_csclk),
    .D(net852),
    .RESET_B(net603),
    .Q(\gpio_configure[25][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7485_ (.CLK(clknet_leaf_31_csclk),
    .D(net705),
    .RESET_B(net603),
    .Q(\gpio_configure[25][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7486_ (.CLK(clknet_leaf_37_csclk),
    .D(net1180),
    .RESET_B(net603),
    .Q(\gpio_configure[25][7] ));
 sky130_fd_sc_hd__dfstp_2 _7487_ (.CLK(clknet_leaf_24_csclk),
    .D(net1873),
    .SET_B(net597),
    .Q(\gpio_configure[26][0] ));
 sky130_fd_sc_hd__dfstp_4 _7488_ (.CLK(clknet_leaf_26_csclk),
    .D(net1668),
    .SET_B(net599),
    .Q(\gpio_configure[26][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7489_ (.CLK(clknet_leaf_64_csclk),
    .D(net1051),
    .RESET_B(net586),
    .Q(\gpio_configure[26][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7490_ (.CLK(clknet_leaf_32_csclk),
    .D(net955),
    .RESET_B(net603),
    .Q(\gpio_configure[26][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7491_ (.CLK(clknet_leaf_26_csclk),
    .D(net2698),
    .RESET_B(net599),
    .Q(\gpio_configure[26][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7492_ (.CLK(clknet_leaf_42_csclk),
    .D(net2074),
    .RESET_B(net594),
    .Q(\gpio_configure[26][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7493_ (.CLK(clknet_leaf_46_csclk),
    .D(net1426),
    .RESET_B(net585),
    .Q(\gpio_configure[26][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7494_ (.CLK(clknet_leaf_42_csclk),
    .D(net1117),
    .RESET_B(net594),
    .Q(\gpio_configure[26][7] ));
 sky130_fd_sc_hd__dfstp_2 _7495_ (.CLK(clknet_leaf_68_csclk),
    .D(net1729),
    .SET_B(net577),
    .Q(\gpio_configure[27][0] ));
 sky130_fd_sc_hd__dfstp_1 _7496_ (.CLK(clknet_3_3_0_csclk),
    .D(net1734),
    .SET_B(net586),
    .Q(\gpio_configure[27][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7497_ (.CLK(clknet_leaf_60_csclk),
    .D(net900),
    .RESET_B(net577),
    .Q(\gpio_configure[27][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7498_ (.CLK(clknet_leaf_29_csclk),
    .D(net866),
    .RESET_B(net602),
    .Q(\gpio_configure[27][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7499_ (.CLK(clknet_leaf_61_csclk),
    .D(net727),
    .RESET_B(net578),
    .Q(\gpio_configure[27][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7500_ (.CLK(clknet_leaf_43_csclk),
    .D(net850),
    .RESET_B(net596),
    .Q(\gpio_configure[27][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7501_ (.CLK(clknet_leaf_55_csclk),
    .D(net1402),
    .RESET_B(net581),
    .Q(\gpio_configure[27][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7502_ (.CLK(clknet_leaf_42_csclk),
    .D(net1151),
    .RESET_B(net594),
    .Q(\gpio_configure[27][7] ));
 sky130_fd_sc_hd__dfstp_4 _7503_ (.CLK(clknet_leaf_28_csclk),
    .D(net1268),
    .SET_B(net601),
    .Q(\gpio_configure[28][0] ));
 sky130_fd_sc_hd__dfstp_4 _7504_ (.CLK(clknet_leaf_28_csclk),
    .D(net1744),
    .SET_B(net600),
    .Q(\gpio_configure[28][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7505_ (.CLK(clknet_leaf_16_csclk),
    .D(net1560),
    .RESET_B(net601),
    .Q(\gpio_configure[28][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7506_ (.CLK(clknet_leaf_29_csclk),
    .D(net872),
    .RESET_B(net602),
    .Q(\gpio_configure[28][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7507_ (.CLK(clknet_leaf_28_csclk),
    .D(net787),
    .RESET_B(net600),
    .Q(\gpio_configure[28][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7508_ (.CLK(clknet_leaf_25_csclk),
    .D(net2179),
    .RESET_B(net603),
    .Q(\gpio_configure[28][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7509_ (.CLK(clknet_leaf_31_csclk),
    .D(net2289),
    .RESET_B(net605),
    .Q(\gpio_configure[28][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7510_ (.CLK(clknet_leaf_32_csclk),
    .D(net1188),
    .RESET_B(net603),
    .Q(\gpio_configure[28][7] ));
 sky130_fd_sc_hd__dfstp_4 _7511_ (.CLK(clknet_leaf_26_csclk),
    .D(net3583),
    .SET_B(net599),
    .Q(\gpio_configure[29][0] ));
 sky130_fd_sc_hd__dfstp_4 _7512_ (.CLK(clknet_leaf_29_csclk),
    .D(net3224),
    .SET_B(net602),
    .Q(\gpio_configure[29][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7513_ (.CLK(clknet_leaf_29_csclk),
    .D(net2142),
    .RESET_B(net602),
    .Q(\gpio_configure[29][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7514_ (.CLK(clknet_leaf_31_csclk),
    .D(net2168),
    .RESET_B(net602),
    .Q(\gpio_configure[29][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7515_ (.CLK(clknet_leaf_30_csclk),
    .D(net1245),
    .RESET_B(net600),
    .Q(\gpio_configure[29][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7516_ (.CLK(clknet_leaf_31_csclk),
    .D(net2086),
    .RESET_B(net603),
    .Q(\gpio_configure[29][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7517_ (.CLK(clknet_leaf_31_csclk),
    .D(net686),
    .RESET_B(net605),
    .Q(\gpio_configure[29][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7518_ (.CLK(clknet_leaf_31_csclk),
    .D(net1069),
    .RESET_B(net603),
    .Q(\gpio_configure[29][7] ));
 sky130_fd_sc_hd__dfstp_4 _7519_ (.CLK(clknet_leaf_27_csclk),
    .D(net1239),
    .SET_B(net602),
    .Q(\gpio_configure[30][0] ));
 sky130_fd_sc_hd__dfstp_4 _7520_ (.CLK(clknet_leaf_26_csclk),
    .D(net1666),
    .SET_B(net599),
    .Q(\gpio_configure[30][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7521_ (.CLK(clknet_leaf_28_csclk),
    .D(net987),
    .RESET_B(net600),
    .Q(\gpio_configure[30][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7522_ (.CLK(clknet_leaf_33_csclk),
    .D(net975),
    .RESET_B(net605),
    .Q(\gpio_configure[30][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7523_ (.CLK(clknet_leaf_27_csclk),
    .D(net1359),
    .RESET_B(net599),
    .Q(\gpio_configure[30][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7524_ (.CLK(clknet_leaf_43_csclk),
    .D(net840),
    .RESET_B(net596),
    .Q(\gpio_configure[30][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7525_ (.CLK(clknet_leaf_43_csclk),
    .D(net741),
    .RESET_B(net596),
    .Q(\gpio_configure[30][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7526_ (.CLK(clknet_leaf_43_csclk),
    .D(net650),
    .RESET_B(net596),
    .Q(\gpio_configure[30][7] ));
 sky130_fd_sc_hd__dfstp_4 _7527_ (.CLK(clknet_leaf_26_csclk),
    .D(net1865),
    .SET_B(net599),
    .Q(\gpio_configure[31][0] ));
 sky130_fd_sc_hd__dfstp_4 _7528_ (.CLK(clknet_leaf_26_csclk),
    .D(net2691),
    .SET_B(net599),
    .Q(\gpio_configure[31][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7529_ (.CLK(clknet_leaf_27_csclk),
    .D(net937),
    .RESET_B(net599),
    .Q(\gpio_configure[31][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7530_ (.CLK(clknet_leaf_30_csclk),
    .D(net2229),
    .RESET_B(net600),
    .Q(\gpio_configure[31][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7531_ (.CLK(clknet_leaf_26_csclk),
    .D(net735),
    .RESET_B(net599),
    .Q(\gpio_configure[31][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7532_ (.CLK(clknet_leaf_25_csclk),
    .D(net2156),
    .RESET_B(net596),
    .Q(\gpio_configure[31][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7533_ (.CLK(clknet_leaf_37_csclk),
    .D(net743),
    .RESET_B(net596),
    .Q(\gpio_configure[31][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7534_ (.CLK(clknet_leaf_25_csclk),
    .D(net2122),
    .RESET_B(net596),
    .Q(\gpio_configure[31][7] ));
 sky130_fd_sc_hd__dfstp_2 _7535_ (.CLK(clknet_leaf_68_csclk),
    .D(net1936),
    .SET_B(net577),
    .Q(\gpio_configure[32][0] ));
 sky130_fd_sc_hd__dfstp_2 _7536_ (.CLK(clknet_leaf_60_csclk),
    .D(net1165),
    .SET_B(net578),
    .Q(\gpio_configure[32][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7537_ (.CLK(clknet_leaf_68_csclk),
    .D(net1176),
    .RESET_B(net577),
    .Q(\gpio_configure[32][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7538_ (.CLK(clknet_leaf_56_csclk),
    .D(net1005),
    .RESET_B(net581),
    .Q(\gpio_configure[32][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7539_ (.CLK(clknet_leaf_60_csclk),
    .D(net717),
    .RESET_B(net578),
    .Q(\gpio_configure[32][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7540_ (.CLK(clknet_leaf_56_csclk),
    .D(net1554),
    .RESET_B(net581),
    .Q(\gpio_configure[32][5] ));
 sky130_fd_sc_hd__dfrtp_2 _7541_ (.CLK(clknet_leaf_56_csclk),
    .D(net1456),
    .RESET_B(net581),
    .Q(\gpio_configure[32][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7542_ (.CLK(clknet_leaf_56_csclk),
    .D(net1159),
    .RESET_B(net581),
    .Q(\gpio_configure[32][7] ));
 sky130_fd_sc_hd__dfstp_2 _7543_ (.CLK(clknet_leaf_39_csclk),
    .D(net1875),
    .SET_B(net595),
    .Q(\gpio_configure[33][0] ));
 sky130_fd_sc_hd__dfstp_2 _7544_ (.CLK(clknet_leaf_42_csclk),
    .D(net1658),
    .SET_B(net594),
    .Q(\gpio_configure[33][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7545_ (.CLK(clknet_leaf_42_csclk),
    .D(net2164),
    .RESET_B(net594),
    .Q(\gpio_configure[33][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7546_ (.CLK(clknet_leaf_42_csclk),
    .D(net927),
    .RESET_B(net594),
    .Q(\gpio_configure[33][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7547_ (.CLK(clknet_leaf_41_csclk),
    .D(net1305),
    .RESET_B(net597),
    .Q(\gpio_configure[33][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7548_ (.CLK(clknet_leaf_40_csclk),
    .D(net2260),
    .RESET_B(net597),
    .Q(\gpio_configure[33][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7549_ (.CLK(clknet_leaf_41_csclk),
    .D(net758),
    .RESET_B(net594),
    .Q(\gpio_configure[33][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7550_ (.CLK(clknet_leaf_41_csclk),
    .D(net1209),
    .RESET_B(net594),
    .Q(\gpio_configure[33][7] ));
 sky130_fd_sc_hd__dfstp_1 _7551_ (.CLK(clknet_leaf_39_csclk),
    .D(net1877),
    .SET_B(net595),
    .Q(\gpio_configure[34][0] ));
 sky130_fd_sc_hd__dfstp_1 _7552_ (.CLK(clknet_leaf_46_csclk),
    .D(net1243),
    .SET_B(net584),
    .Q(\gpio_configure[34][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7553_ (.CLK(clknet_leaf_48_csclk),
    .D(net638),
    .RESET_B(net585),
    .Q(\gpio_configure[34][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7554_ (.CLK(clknet_leaf_38_csclk),
    .D(net989),
    .RESET_B(net595),
    .Q(\gpio_configure[34][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7555_ (.CLK(clknet_leaf_41_csclk),
    .D(net1313),
    .RESET_B(net594),
    .Q(\gpio_configure[34][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7556_ (.CLK(clknet_leaf_40_csclk),
    .D(net880),
    .RESET_B(net597),
    .Q(\gpio_configure[34][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7557_ (.CLK(clknet_leaf_48_csclk),
    .D(net1428),
    .RESET_B(net584),
    .Q(\gpio_configure[34][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7558_ (.CLK(clknet_leaf_47_csclk),
    .D(net656),
    .RESET_B(net585),
    .Q(\gpio_configure[34][7] ));
 sky130_fd_sc_hd__dfstp_4 _7559_ (.CLK(clknet_leaf_27_csclk),
    .D(net1881),
    .SET_B(net602),
    .Q(\gpio_configure[35][0] ));
 sky130_fd_sc_hd__dfstp_2 _7560_ (.CLK(clknet_leaf_26_csclk),
    .D(net1656),
    .SET_B(net599),
    .Q(\gpio_configure[35][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7561_ (.CLK(clknet_leaf_27_csclk),
    .D(net933),
    .RESET_B(net598),
    .Q(\gpio_configure[35][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7562_ (.CLK(clknet_leaf_25_csclk),
    .D(net921),
    .RESET_B(net599),
    .Q(\gpio_configure[35][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7563_ (.CLK(clknet_leaf_27_csclk),
    .D(net770),
    .RESET_B(net602),
    .Q(\gpio_configure[35][4] ));
 sky130_fd_sc_hd__dfrtp_4 _7564_ (.CLK(clknet_leaf_25_csclk),
    .D(net834),
    .RESET_B(net603),
    .Q(\gpio_configure[35][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7565_ (.CLK(clknet_leaf_31_csclk),
    .D(net697),
    .RESET_B(net603),
    .Q(\gpio_configure[35][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7566_ (.CLK(clknet_leaf_25_csclk),
    .D(net642),
    .RESET_B(net603),
    .Q(\gpio_configure[35][7] ));
 sky130_fd_sc_hd__dfstp_1 _7567_ (.CLK(clknet_leaf_43_csclk),
    .D(net1871),
    .SET_B(net596),
    .Q(\gpio_configure[36][0] ));
 sky130_fd_sc_hd__dfstp_2 _7568_ (.CLK(clknet_leaf_42_csclk),
    .D(net1674),
    .SET_B(net596),
    .Q(\gpio_configure[36][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7569_ (.CLK(clknet_leaf_44_csclk),
    .D(net929),
    .RESET_B(net597),
    .Q(\gpio_configure[36][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7570_ (.CLK(clknet_leaf_43_csclk),
    .D(net1011),
    .RESET_B(net596),
    .Q(\gpio_configure[36][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7571_ (.CLK(clknet_leaf_38_csclk),
    .D(net1264),
    .RESET_B(net596),
    .Q(\gpio_configure[36][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7572_ (.CLK(clknet_leaf_43_csclk),
    .D(net858),
    .RESET_B(net596),
    .Q(\gpio_configure[36][5] ));
 sky130_fd_sc_hd__dfrtp_4 _7573_ (.CLK(clknet_leaf_42_csclk),
    .D(net739),
    .RESET_B(net597),
    .Q(\gpio_configure[36][6] ));
 sky130_fd_sc_hd__dfrtp_2 _7574_ (.CLK(clknet_leaf_42_csclk),
    .D(net1141),
    .RESET_B(net597),
    .Q(\gpio_configure[36][7] ));
 sky130_fd_sc_hd__dfstp_2 _7575_ (.CLK(clknet_leaf_38_csclk),
    .D(net1859),
    .SET_B(net595),
    .Q(\gpio_configure[37][0] ));
 sky130_fd_sc_hd__dfstp_1 _7576_ (.CLK(clknet_leaf_46_csclk),
    .D(net692),
    .SET_B(net585),
    .Q(\gpio_configure[37][1] ));
 sky130_fd_sc_hd__dfrtp_4 _7577_ (.CLK(clknet_leaf_48_csclk),
    .D(net633),
    .RESET_B(net584),
    .Q(\gpio_configure[37][2] ));
 sky130_fd_sc_hd__dfrtp_4 _7578_ (.CLK(clknet_leaf_37_csclk),
    .D(net902),
    .RESET_B(net604),
    .Q(\gpio_configure[37][3] ));
 sky130_fd_sc_hd__dfrtp_4 _7579_ (.CLK(clknet_leaf_42_csclk),
    .D(net1276),
    .RESET_B(net597),
    .Q(\gpio_configure[37][4] ));
 sky130_fd_sc_hd__dfrtp_2 _7580_ (.CLK(clknet_leaf_42_csclk),
    .D(net832),
    .RESET_B(net596),
    .Q(\gpio_configure[37][5] ));
 sky130_fd_sc_hd__dfrtp_1 _7581_ (.CLK(clknet_leaf_46_csclk),
    .D(net1452),
    .RESET_B(net584),
    .Q(\gpio_configure[37][6] ));
 sky130_fd_sc_hd__dfrtp_4 _7582_ (.CLK(clknet_leaf_47_csclk),
    .D(net662),
    .RESET_B(net585),
    .Q(\gpio_configure[37][7] ));
 sky130_fd_sc_hd__dfrtp_4 _7583_ (.CLK(clknet_4_3__leaf_wb_clk_i),
    .D(_0753_),
    .RESET_B(net563),
    .Q(serial_busy));
 sky130_fd_sc_hd__dfrtp_4 _7584_ (.CLK(clknet_4_3__leaf_wb_clk_i),
    .D(_0754_),
    .RESET_B(net564),
    .Q(\xfer_count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7585_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0755_),
    .RESET_B(net564),
    .Q(\xfer_count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7586_ (.CLK(clknet_4_3__leaf_wb_clk_i),
    .D(_0756_),
    .RESET_B(net564),
    .Q(\xfer_count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7587_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0757_),
    .RESET_B(net564),
    .Q(\xfer_count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7588_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0758_),
    .RESET_B(net567),
    .Q(\pad_count_1[0] ));
 sky130_fd_sc_hd__dfstp_4 _7589_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_0759_),
    .SET_B(net567),
    .Q(\pad_count_1[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7590_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_0760_),
    .RESET_B(net567),
    .Q(\pad_count_1[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7591_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_0761_),
    .RESET_B(net568),
    .Q(\pad_count_1[3] ));
 sky130_fd_sc_hd__dfstp_4 _7592_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_0762_),
    .SET_B(net568),
    .Q(\pad_count_1[4] ));
 sky130_fd_sc_hd__dfstp_4 _7593_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_0763_),
    .SET_B(net567),
    .Q(\pad_count_2[0] ));
 sky130_fd_sc_hd__dfstp_4 _7594_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0764_),
    .SET_B(net568),
    .Q(\pad_count_2[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7595_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0765_),
    .RESET_B(net567),
    .Q(\pad_count_2[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7596_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0766_),
    .RESET_B(net567),
    .Q(\pad_count_2[3] ));
 sky130_fd_sc_hd__dfstp_4 _7597_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0767_),
    .SET_B(net568),
    .Q(\pad_count_2[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7598_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(_0768_),
    .RESET_B(net568),
    .Q(\pad_count_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7599_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(net622),
    .RESET_B(net566),
    .Q(serial_resetn_pre));
 sky130_fd_sc_hd__conb_1 _7599__622 (.HI(net622));
 sky130_fd_sc_hd__dfrtp_1 _7600_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(_0769_),
    .RESET_B(net567),
    .Q(serial_clock_pre));
 sky130_fd_sc_hd__dfrtp_1 _7601_ (.CLK(clknet_4_0__leaf_wb_clk_i),
    .D(net3870),
    .RESET_B(net569),
    .Q(serial_load_pre));
 sky130_fd_sc_hd__dfrtp_1 _7602_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(_0771_),
    .RESET_B(net575),
    .Q(\serial_data_staging_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7603_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(_0772_),
    .RESET_B(net575),
    .Q(\serial_data_staging_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7604_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(_0773_),
    .RESET_B(net576),
    .Q(\serial_data_staging_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7605_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(net3832),
    .RESET_B(net576),
    .Q(\serial_data_staging_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7606_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(net3824),
    .RESET_B(net576),
    .Q(\serial_data_staging_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7607_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0776_),
    .RESET_B(net579),
    .Q(\serial_data_staging_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7608_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0777_),
    .RESET_B(net579),
    .Q(\serial_data_staging_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7609_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0778_),
    .RESET_B(net575),
    .Q(\serial_data_staging_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7610_ (.CLK(clknet_4_6__leaf_wb_clk_i),
    .D(net3820),
    .RESET_B(net568),
    .Q(\serial_data_staging_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7611_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(_0780_),
    .RESET_B(net566),
    .Q(\serial_data_staging_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7612_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(net3840),
    .RESET_B(net566),
    .Q(\serial_data_staging_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7613_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(_0782_),
    .RESET_B(net566),
    .Q(\serial_data_staging_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7614_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(net3859),
    .RESET_B(net566),
    .Q(\serial_data_staging_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7615_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(net3838),
    .RESET_B(net576),
    .Q(\serial_data_staging_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7616_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(net3818),
    .RESET_B(net576),
    .Q(\serial_data_staging_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7617_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0786_),
    .RESET_B(net576),
    .Q(\serial_data_staging_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7618_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(net3827),
    .RESET_B(net576),
    .Q(\serial_data_staging_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7619_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0788_),
    .RESET_B(net579),
    .Q(\serial_data_staging_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7620_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(_0789_),
    .RESET_B(net582),
    .Q(\serial_data_staging_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7621_ (.CLK(clknet_4_5__leaf_wb_clk_i),
    .D(net3836),
    .RESET_B(net579),
    .Q(\serial_data_staging_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7622_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(_0791_),
    .RESET_B(net575),
    .Q(\serial_data_staging_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7623_ (.CLK(clknet_4_4__leaf_wb_clk_i),
    .D(_0792_),
    .RESET_B(net575),
    .Q(\serial_data_staging_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7624_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(net3815),
    .RESET_B(net569),
    .Q(\serial_data_staging_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7625_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(_0794_),
    .RESET_B(net566),
    .Q(\serial_data_staging_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7626_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(_0795_),
    .RESET_B(net569),
    .Q(\serial_data_staging_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7627_ (.CLK(clknet_4_7__leaf_wb_clk_i),
    .D(_0796_),
    .RESET_B(net566),
    .Q(\serial_data_staging_2[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7628_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(net3884),
    .RESET_B(net607),
    .Q(net311));
 sky130_fd_sc_hd__dfxtp_1 _7629_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0798_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_4_11__leaf_wb_clk_i),
    .D(_0799_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0800_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0801_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_4_8__leaf_wb_clk_i),
    .D(_0802_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0803_),
    .Q(net333));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0804_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_4_10__leaf_wb_clk_i),
    .D(_0805_),
    .Q(net336));
 sky130_fd_sc_hd__dfrtp_1 _7637_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0806_),
    .RESET_B(net607),
    .Q(\wbbd_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7638_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0807_),
    .RESET_B(net607),
    .Q(\wbbd_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7639_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0808_),
    .RESET_B(net607),
    .Q(\wbbd_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7640_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0809_),
    .RESET_B(net607),
    .Q(\wbbd_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7641_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0810_),
    .RESET_B(net607),
    .Q(\wbbd_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7642_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0811_),
    .RESET_B(net607),
    .Q(\wbbd_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7643_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(_0812_),
    .RESET_B(net607),
    .Q(\wbbd_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7644_ (.CLK(clknet_4_15__leaf_wb_clk_i),
    .D(_0813_),
    .RESET_B(net608),
    .Q(\wbbd_data[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7645_ (.CLK(clknet_4_13__leaf_wb_clk_i),
    .D(_0814_),
    .RESET_B(net607),
    .Q(wbbd_sck));
 sky130_fd_sc_hd__dfrtp_1 _7646_ (.CLK(clknet_4_14__leaf_wb_clk_i),
    .D(_0815_),
    .RESET_B(net608),
    .Q(wbbd_write));
 sky130_fd_sc_hd__clkbuf_2 _7648_ (.A(irq_spi),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 _7649_ (.A(\mgmt_gpio_data[2] ),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 _7650_ (.A(\mgmt_gpio_data[3] ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 _7651_ (.A(\mgmt_gpio_data[4] ),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 _7652_ (.A(\mgmt_gpio_data[5] ),
    .X(net242));
 sky130_fd_sc_hd__buf_2 _7653_ (.A(\mgmt_gpio_data[7] ),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 _7654_ (.A(\mgmt_gpio_data[11] ),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 _7655_ (.A(\mgmt_gpio_data[12] ),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 _7656_ (.A(\mgmt_gpio_data[16] ),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 _7657_ (.A(\mgmt_gpio_data[17] ),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 _7658_ (.A(\mgmt_gpio_data[18] ),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 _7659_ (.A(\mgmt_gpio_data[19] ),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 _7660_ (.A(\mgmt_gpio_data[20] ),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 _7661_ (.A(\mgmt_gpio_data[21] ),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 _7662_ (.A(\mgmt_gpio_data[22] ),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 _7663_ (.A(\mgmt_gpio_data[23] ),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 _7664_ (.A(\mgmt_gpio_data[24] ),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 _7665_ (.A(\mgmt_gpio_data[25] ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 _7666_ (.A(\mgmt_gpio_data[26] ),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 _7667_ (.A(\mgmt_gpio_data[27] ),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 _7668_ (.A(\mgmt_gpio_data[28] ),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 _7669_ (.A(\mgmt_gpio_data[29] ),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 _7670_ (.A(\mgmt_gpio_data[34] ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _7671_ (.A(net87),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 _7672_ (.A(net65),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 _7673_ (.A(net66),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1111_ (.A(_1111_),
    .X(clknet_0__1111_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_csclk (.A(csclk),
    .X(clknet_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_mgmt_gpio_in[4]  (.A(mgmt_gpio_in[4]),
    .X(clknet_0_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock (.A(user_clock),
    .X(clknet_0_user_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wbbd_sck (.A(wbbd_sck),
    .X(clknet_0_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1111_ (.A(clknet_0__1111_),
    .X(clknet_1_0__leaf__1111_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_user_clock (.A(clknet_0_user_clock),
    .X(clknet_1_0__leaf_user_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_0__leaf_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1111_ (.A(clknet_0__1111_),
    .X(clknet_1_1__leaf__1111_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_user_clock (.A(clknet_0_user_clock),
    .X(clknet_1_1__leaf_user_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wbbd_sck (.A(clknet_0_wbbd_sck),
    .X(clknet_1_1__leaf_wbbd_sck));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_0__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_1__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_2__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_mgmt_gpio_in[4]  (.A(clknet_0_mgmt_gpio_in[4]),
    .X(clknet_2_3__leaf_mgmt_gpio_in[4]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_0_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_1_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_2_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_3_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_4_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_5_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_6_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_csclk (.A(clknet_0_csclk),
    .X(clknet_3_7_0_csclk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_10__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_11__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_12__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_14__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_15__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_8__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_9__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_0_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_10_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_11_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_12_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_13_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_14_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_15_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_16_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_17_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_18_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_19_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_1_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_20_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_21_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_22_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_23_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_24_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_25_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_26_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_27_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_csclk (.A(clknet_3_5_0_csclk),
    .X(clknet_leaf_28_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_29_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_2_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_30_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_31_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_32_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_33_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_35_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_36_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_csclk (.A(clknet_3_7_0_csclk),
    .X(clknet_leaf_37_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_38_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_39_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_3_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_40_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_41_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_42_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_43_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_44_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_45_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_46_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_csclk (.A(clknet_3_6_0_csclk),
    .X(clknet_leaf_47_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_48_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_49_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_4_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_50_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_51_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_52_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_53_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_54_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_55_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_56_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_57_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_58_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_59_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_5_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_60_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_csclk (.A(clknet_3_2_0_csclk),
    .X(clknet_leaf_61_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_62_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_63_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_64_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_csclk (.A(clknet_3_3_0_csclk),
    .X(clknet_leaf_66_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_67_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_68_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_69_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_6_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_70_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_71_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_72_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_73_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_74_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_csclk (.A(clknet_3_0_0_csclk),
    .X(clknet_leaf_75_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_76_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_csclk (.A(clknet_3_1_0_csclk),
    .X(clknet_leaf_77_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_7_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_8_csclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_csclk (.A(clknet_3_4_0_csclk),
    .X(clknet_leaf_9_csclk));
 sky130_fd_sc_hd__buf_12 fanout353 (.A(_2681_),
    .X(net353));
 sky130_fd_sc_hd__buf_12 fanout354 (.A(net679),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_16 fanout355 (.A(net679),
    .X(net355));
 sky130_fd_sc_hd__buf_12 fanout356 (.A(net2115),
    .X(net356));
 sky130_fd_sc_hd__buf_12 fanout357 (.A(net359),
    .X(net357));
 sky130_fd_sc_hd__buf_12 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_12 fanout359 (.A(net1024),
    .X(net359));
 sky130_fd_sc_hd__buf_12 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_6 fanout361 (.A(_1729_),
    .X(net361));
 sky130_fd_sc_hd__buf_6 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_4 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_12 fanout369 (.A(_1421_),
    .X(net369));
 sky130_fd_sc_hd__buf_12 fanout370 (.A(_0958_),
    .X(net370));
 sky130_fd_sc_hd__buf_8 fanout371 (.A(_0958_),
    .X(net371));
 sky130_fd_sc_hd__buf_12 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__buf_12 fanout373 (.A(_0940_),
    .X(net373));
 sky130_fd_sc_hd__buf_12 fanout374 (.A(_0931_),
    .X(net374));
 sky130_fd_sc_hd__buf_12 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_12 fanout376 (.A(_0897_),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_16 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_16 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_12 fanout379 (.A(net2453),
    .X(net379));
 sky130_fd_sc_hd__buf_8 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_8 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_8 fanout382 (.A(net756),
    .X(net382));
 sky130_fd_sc_hd__buf_12 fanout383 (.A(_0875_),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_16 fanout384 (.A(_0875_),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_16 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_8 fanout386 (.A(net905),
    .X(net386));
 sky130_fd_sc_hd__buf_12 fanout387 (.A(_0867_),
    .X(net387));
 sky130_fd_sc_hd__buf_12 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_12 fanout389 (.A(_0855_),
    .X(net389));
 sky130_fd_sc_hd__buf_12 fanout390 (.A(net2849),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_16 fanout391 (.A(net2849),
    .X(net391));
 sky130_fd_sc_hd__buf_6 fanout392 (.A(net2849),
    .X(net392));
 sky130_fd_sc_hd__buf_12 fanout394 (.A(_1864_),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_16 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_8 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_12 fanout403 (.A(net406),
    .X(net403));
 sky130_fd_sc_hd__buf_12 fanout407 (.A(net2091),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_16 fanout408 (.A(net2091),
    .X(net408));
 sky130_fd_sc_hd__buf_12 fanout409 (.A(net2210),
    .X(net409));
 sky130_fd_sc_hd__buf_12 fanout410 (.A(net412),
    .X(net410));
 sky130_fd_sc_hd__buf_12 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_12 fanout412 (.A(_0872_),
    .X(net412));
 sky130_fd_sc_hd__buf_12 fanout413 (.A(net695),
    .X(net413));
 sky130_fd_sc_hd__buf_8 fanout414 (.A(net695),
    .X(net414));
 sky130_fd_sc_hd__buf_12 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_12 fanout416 (.A(_0863_),
    .X(net416));
 sky130_fd_sc_hd__buf_12 fanout417 (.A(net645),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(net645),
    .X(net418));
 sky130_fd_sc_hd__buf_12 fanout419 (.A(net2070),
    .X(net419));
 sky130_fd_sc_hd__buf_12 fanout420 (.A(net660),
    .X(net420));
 sky130_fd_sc_hd__buf_12 fanout421 (.A(net659),
    .X(net421));
 sky130_fd_sc_hd__buf_12 fanout422 (.A(_2719_),
    .X(net422));
 sky130_fd_sc_hd__buf_12 fanout423 (.A(_2686_),
    .X(net423));
 sky130_fd_sc_hd__buf_6 fanout425 (.A(_1865_),
    .X(net425));
 sky130_fd_sc_hd__buf_12 fanout430 (.A(_3033_),
    .X(net430));
 sky130_fd_sc_hd__buf_12 fanout431 (.A(_3029_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_16 fanout432 (.A(_3004_),
    .X(net432));
 sky130_fd_sc_hd__buf_4 fanout433 (.A(_3004_),
    .X(net433));
 sky130_fd_sc_hd__buf_12 fanout434 (.A(_3004_),
    .X(net434));
 sky130_fd_sc_hd__buf_12 fanout435 (.A(_3002_),
    .X(net435));
 sky130_fd_sc_hd__buf_12 fanout436 (.A(_2706_),
    .X(net436));
 sky130_fd_sc_hd__buf_12 fanout437 (.A(_2691_),
    .X(net437));
 sky130_fd_sc_hd__buf_8 fanout438 (.A(_2691_),
    .X(net438));
 sky130_fd_sc_hd__buf_12 fanout439 (.A(_2672_),
    .X(net439));
 sky130_fd_sc_hd__buf_8 fanout440 (.A(_2672_),
    .X(net440));
 sky130_fd_sc_hd__buf_12 fanout441 (.A(_2663_),
    .X(net441));
 sky130_fd_sc_hd__buf_12 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_12 fanout443 (.A(_2657_),
    .X(net443));
 sky130_fd_sc_hd__buf_12 fanout444 (.A(_2648_),
    .X(net444));
 sky130_fd_sc_hd__buf_6 fanout445 (.A(_2648_),
    .X(net445));
 sky130_fd_sc_hd__buf_12 fanout446 (.A(_2647_),
    .X(net446));
 sky130_fd_sc_hd__buf_12 fanout447 (.A(_2646_),
    .X(net447));
 sky130_fd_sc_hd__buf_12 fanout448 (.A(_1861_),
    .X(net448));
 sky130_fd_sc_hd__buf_8 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_8 fanout458 (.A(_1709_),
    .X(net458));
 sky130_fd_sc_hd__buf_12 fanout465 (.A(net641),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_16 fanout466 (.A(net641),
    .X(net466));
 sky130_fd_sc_hd__buf_6 fanout467 (.A(net2100),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_16 fanout468 (.A(net685),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net685),
    .X(net469));
 sky130_fd_sc_hd__buf_6 fanout470 (.A(net2286),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_16 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_16 fanout472 (.A(net2017),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_16 fanout473 (.A(net2017),
    .X(net473));
 sky130_fd_sc_hd__buf_12 fanout474 (.A(net708),
    .X(net474));
 sky130_fd_sc_hd__buf_6 fanout475 (.A(net2696),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_16 fanout476 (.A(net478),
    .X(net476));
 sky130_fd_sc_hd__buf_12 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__buf_12 fanout478 (.A(net2696),
    .X(net478));
 sky130_fd_sc_hd__buf_12 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_12 fanout480 (.A(net2027),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_16 fanout481 (.A(net2027),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_8 fanout482 (.A(net2027),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_16 fanout483 (.A(net2027),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_16 fanout484 (.A(net2033),
    .X(net484));
 sky130_fd_sc_hd__buf_6 fanout485 (.A(net2033),
    .X(net485));
 sky130_fd_sc_hd__buf_12 fanout486 (.A(net2033),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_16 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_12 fanout488 (.A(net2033),
    .X(net488));
 sky130_fd_sc_hd__buf_12 fanout489 (.A(net667),
    .X(net489));
 sky130_fd_sc_hd__buf_12 fanout490 (.A(net667),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_16 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_12 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_6 fanout493 (.A(net667),
    .X(net493));
 sky130_fd_sc_hd__buf_6 fanout494 (.A(net2348),
    .X(net494));
 sky130_fd_sc_hd__buf_12 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_16 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_12 fanout497 (.A(net1088),
    .X(net497));
 sky130_fd_sc_hd__buf_12 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_12 fanout499 (.A(net1088),
    .X(net499));
 sky130_fd_sc_hd__buf_6 fanout500 (.A(net2663),
    .X(net500));
 sky130_fd_sc_hd__buf_12 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_12 fanout502 (.A(net671),
    .X(net502));
 sky130_fd_sc_hd__buf_12 fanout503 (.A(net671),
    .X(net503));
 sky130_fd_sc_hd__buf_12 fanout504 (.A(net672),
    .X(net504));
 sky130_fd_sc_hd__buf_6 fanout505 (.A(net671),
    .X(net505));
 sky130_fd_sc_hd__buf_6 fanout506 (.A(net2042),
    .X(net506));
 sky130_fd_sc_hd__buf_12 fanout510 (.A(net512),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_16 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__buf_12 fanout512 (.A(_0827_),
    .X(net512));
 sky130_fd_sc_hd__buf_12 fanout513 (.A(_0824_),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_16 fanout514 (.A(\pad_count_2[3] ),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_16 fanout515 (.A(\pad_count_2[2] ),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_16 fanout516 (.A(\pad_count_1[4] ),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(\pad_count_1[4] ),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_16 fanout518 (.A(\pad_count_1[4] ),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_16 fanout519 (.A(\pad_count_1[4] ),
    .X(net519));
 sky130_fd_sc_hd__buf_12 fanout520 (.A(\pad_count_1[3] ),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_8 fanout521 (.A(\pad_count_1[3] ),
    .X(net521));
 sky130_fd_sc_hd__buf_12 fanout522 (.A(\pad_count_1[2] ),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_8 fanout523 (.A(\pad_count_1[2] ),
    .X(net523));
 sky130_fd_sc_hd__buf_12 fanout524 (.A(net2935),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_16 fanout525 (.A(net3907),
    .X(net525));
 sky130_fd_sc_hd__buf_12 fanout526 (.A(\xfer_state[2] ),
    .X(net526));
 sky130_fd_sc_hd__buf_12 fanout527 (.A(\xfer_state[1] ),
    .X(net527));
 sky130_fd_sc_hd__buf_8 fanout528 (.A(\xfer_state[1] ),
    .X(net528));
 sky130_fd_sc_hd__buf_12 fanout531 (.A(_1891_),
    .X(net531));
 sky130_fd_sc_hd__buf_12 fanout532 (.A(_1875_),
    .X(net532));
 sky130_fd_sc_hd__buf_12 fanout535 (.A(_1844_),
    .X(net535));
 sky130_fd_sc_hd__buf_12 fanout542 (.A(net544),
    .X(net542));
 sky130_fd_sc_hd__buf_12 fanout543 (.A(_1708_),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_16 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_12 fanout558 (.A(_1585_),
    .X(net558));
 sky130_fd_sc_hd__buf_12 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__buf_12 fanout562 (.A(net99),
    .X(net562));
 sky130_fd_sc_hd__buf_8 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_16 fanout564 (.A(net569),
    .X(net564));
 sky130_fd_sc_hd__buf_12 fanout565 (.A(net569),
    .X(net565));
 sky130_fd_sc_hd__buf_12 fanout566 (.A(net569),
    .X(net566));
 sky130_fd_sc_hd__buf_12 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__buf_6 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_12 fanout569 (.A(net587),
    .X(net569));
 sky130_fd_sc_hd__buf_6 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_12 fanout571 (.A(net587),
    .X(net571));
 sky130_fd_sc_hd__buf_12 fanout572 (.A(net574),
    .X(net572));
 sky130_fd_sc_hd__buf_12 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__buf_8 fanout574 (.A(net587),
    .X(net574));
 sky130_fd_sc_hd__buf_12 fanout575 (.A(net587),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_16 fanout576 (.A(net587),
    .X(net576));
 sky130_fd_sc_hd__buf_12 fanout577 (.A(net587),
    .X(net577));
 sky130_fd_sc_hd__buf_6 fanout578 (.A(net587),
    .X(net578));
 sky130_fd_sc_hd__buf_12 fanout579 (.A(net582),
    .X(net579));
 sky130_fd_sc_hd__buf_12 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__buf_12 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_8 fanout582 (.A(net587),
    .X(net582));
 sky130_fd_sc_hd__buf_12 fanout583 (.A(net585),
    .X(net583));
 sky130_fd_sc_hd__buf_12 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_16 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_16 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__buf_12 fanout587 (.A(net606),
    .X(net587));
 sky130_fd_sc_hd__buf_12 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_16 fanout589 (.A(net606),
    .X(net589));
 sky130_fd_sc_hd__buf_12 fanout590 (.A(net606),
    .X(net590));
 sky130_fd_sc_hd__buf_12 fanout591 (.A(net606),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_8 fanout592 (.A(net606),
    .X(net592));
 sky130_fd_sc_hd__buf_12 fanout593 (.A(net597),
    .X(net593));
 sky130_fd_sc_hd__buf_12 fanout594 (.A(net597),
    .X(net594));
 sky130_fd_sc_hd__buf_12 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_12 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_12 fanout597 (.A(net606),
    .X(net597));
 sky130_fd_sc_hd__buf_12 fanout598 (.A(net602),
    .X(net598));
 sky130_fd_sc_hd__buf_12 fanout599 (.A(net602),
    .X(net599));
 sky130_fd_sc_hd__buf_12 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_12 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_12 fanout602 (.A(net606),
    .X(net602));
 sky130_fd_sc_hd__buf_12 fanout603 (.A(net605),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_8 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__buf_12 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_12 fanout606 (.A(net75),
    .X(net606));
 sky130_fd_sc_hd__buf_12 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_12 fanout608 (.A(net164),
    .X(net608));
 sky130_fd_sc_hd__buf_12 fanout609 (.A(net128),
    .X(net609));
 sky130_fd_sc_hd__buf_12 fanout610 (.A(net127),
    .X(net610));
 sky130_fd_sc_hd__buf_12 fanout611 (.A(net613),
    .X(net611));
 sky130_fd_sc_hd__buf_12 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__buf_8 fanout613 (.A(net126),
    .X(net613));
 sky130_fd_sc_hd__buf_12 fanout614 (.A(net125),
    .X(net614));
 sky130_fd_sc_hd__buf_12 fanout615 (.A(net124),
    .X(net615));
 sky130_fd_sc_hd__buf_12 fanout616 (.A(net124),
    .X(net616));
 sky130_fd_sc_hd__buf_12 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__buf_12 fanout618 (.A(net121),
    .X(net618));
 sky130_fd_sc_hd__buf_12 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__buf_8 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_12 fanout621 (.A(net110),
    .X(net621));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1 (.A(net2014),
    .X(net625));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold10 (.A(net2066),
    .X(net634));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold100 (.A(net2974),
    .X(net724));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1000 (.A(net3029),
    .X(net1624));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1001 (.A(net3042),
    .X(net1625));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1002 (.A(_0315_),
    .X(net1626));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1003 (.A(net3046),
    .X(net1627));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1004 (.A(_0518_),
    .X(net1628));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1005 (.A(net3101),
    .X(net1629));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1006 (.A(_0408_),
    .X(net1630));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1007 (.A(net3222),
    .X(net1631));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1008 (.A(net3449),
    .X(net1632));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1009 (.A(_0267_),
    .X(net1633));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold101 (.A(net2976),
    .X(net725));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1010 (.A(net3380),
    .X(net1634));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1011 (.A(_0465_),
    .X(net1635));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1012 (.A(net3227),
    .X(net1636));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1013 (.A(net3367),
    .X(net1637));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1014 (.A(_0529_),
    .X(net1638));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1015 (.A(net3088),
    .X(net1639));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1016 (.A(net3090),
    .X(net1640));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1017 (.A(net3341),
    .X(net1641));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1018 (.A(net3343),
    .X(net1642));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1019 (.A(net3403),
    .X(net1643));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold102 (.A(net2940),
    .X(net726));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1020 (.A(_0212_),
    .X(net1644));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1021 (.A(net3508),
    .X(net1645));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1022 (.A(net3510),
    .X(net1646));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1023 (.A(net3458),
    .X(net1647));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1024 (.A(net3460),
    .X(net1648));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1025 (.A(net3394),
    .X(net1649));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1026 (.A(_0153_),
    .X(net1650));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1027 (.A(net3521),
    .X(net1651));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1028 (.A(net3523),
    .X(net1652));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1029 (.A(net3365),
    .X(net1653));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold103 (.A(_0669_),
    .X(net727));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1030 (.A(_0473_),
    .X(net1654));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1031 (.A(net3531),
    .X(net1655));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1032 (.A(_0730_),
    .X(net1656));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1033 (.A(net3528),
    .X(net1657));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1034 (.A(net3530),
    .X(net1658));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1035 (.A(net3361),
    .X(net1659));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1036 (.A(_0489_),
    .X(net1660));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1037 (.A(net3358),
    .X(net1661));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1038 (.A(net3360),
    .X(net1662));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1039 (.A(net3513),
    .X(net1663));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold104 (.A(net3025),
    .X(net728));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1040 (.A(net3515),
    .X(net1664));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1041 (.A(net3502),
    .X(net1665));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1042 (.A(_0690_),
    .X(net1666));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1043 (.A(net3511),
    .X(net1667));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1044 (.A(_0658_),
    .X(net1668));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1045 (.A(net3478),
    .X(net1669));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1046 (.A(net3480),
    .X(net1670));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1047 (.A(net3183),
    .X(net1671));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1048 (.A(_0526_),
    .X(net1672));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1049 (.A(net3543),
    .X(net1673));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold105 (.A(_0581_),
    .X(net729));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1050 (.A(_0738_),
    .X(net1674));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1051 (.A(net3372),
    .X(net1675));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1052 (.A(net3374),
    .X(net1676));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1053 (.A(net3398),
    .X(net1677));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1054 (.A(net3400),
    .X(net1678));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1055 (.A(net3396),
    .X(net1679));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1056 (.A(_0302_),
    .X(net1680));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1057 (.A(net3194),
    .X(net1681));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1058 (.A(net3196),
    .X(net1682));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1059 (.A(net3215),
    .X(net1683));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold106 (.A(net2983),
    .X(net730));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1060 (.A(net3416),
    .X(net1684));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1061 (.A(net3418),
    .X(net1685));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1062 (.A(net3422),
    .X(net1686));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1063 (.A(_0282_),
    .X(net1687));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1064 (.A(net3445),
    .X(net1688));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1065 (.A(_0217_),
    .X(net1689));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1066 (.A(net3435),
    .X(net1690));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1067 (.A(_0457_),
    .X(net1691));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1068 (.A(net3465),
    .X(net1692));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1069 (.A(net3467),
    .X(net1693));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold107 (.A(net2985),
    .X(net731));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1070 (.A(net3456),
    .X(net1694));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1071 (.A(_0227_),
    .X(net1695));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1072 (.A(net3488),
    .X(net1696));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1073 (.A(_0317_),
    .X(net1697));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1074 (.A(net3427),
    .X(net1698));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1075 (.A(_0307_),
    .X(net1699));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1076 (.A(net3437),
    .X(net1700));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1077 (.A(_0287_),
    .X(net1701));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1078 (.A(net3550),
    .X(net1702));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1079 (.A(net3552),
    .X(net1703));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold108 (.A(net2702),
    .X(net732));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1080 (.A(net3526),
    .X(net1704));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1081 (.A(_0292_),
    .X(net1705));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1082 (.A(net3453),
    .X(net1706));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1083 (.A(net3455),
    .X(net1707));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1084 (.A(net3541),
    .X(net1708));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1085 (.A(_0154_),
    .X(net1709));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1086 (.A(net3490),
    .X(net1710));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1087 (.A(_0322_),
    .X(net1711));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1088 (.A(net3553),
    .X(net1712));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1089 (.A(_0283_),
    .X(net1713));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold109 (.A(net2704),
    .X(net733));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1090 (.A(net3545),
    .X(net1714));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1091 (.A(net3547),
    .X(net1715));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1092 (.A(net3557),
    .X(net1716));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1093 (.A(_0213_),
    .X(net1717));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1094 (.A(net3496),
    .X(net1718));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1095 (.A(_0232_),
    .X(net1719));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1096 (.A(net3516),
    .X(net1720));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1097 (.A(net3518),
    .X(net1721));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1098 (.A(net3498),
    .X(net1722));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1099 (.A(_0297_),
    .X(net1723));
 sky130_fd_sc_hd__clkbuf_2 hold11 (.A(net2068),
    .X(net635));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold110 (.A(net2699),
    .X(net734));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1100 (.A(net3555),
    .X(net1724));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1101 (.A(_0546_),
    .X(net1725));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1102 (.A(net3481),
    .X(net1726));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1103 (.A(net3483),
    .X(net1727));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1104 (.A(net3504),
    .X(net1728));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1105 (.A(_0665_),
    .X(net1729));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1106 (.A(net3282),
    .X(net1730));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1107 (.A(net3617),
    .X(net1731));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1108 (.A(net3619),
    .X(net1732));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1109 (.A(net3571),
    .X(net1733));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold111 (.A(net2701),
    .X(net735));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1110 (.A(_0666_),
    .X(net1734));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1111 (.A(net3615),
    .X(net1735));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1112 (.A(_0522_),
    .X(net1736));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1113 (.A(net3559),
    .X(net1737));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1114 (.A(_0380_),
    .X(net1738));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1115 (.A(net3627),
    .X(net1739));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1116 (.A(net3629),
    .X(net1740));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1117 (.A(net3586),
    .X(net1741));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1118 (.A(_0338_),
    .X(net1742));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1119 (.A(net3584),
    .X(net1743));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold112 (.A(net2379),
    .X(net736));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1120 (.A(_0674_),
    .X(net1744));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1121 (.A(net3599),
    .X(net1745));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1122 (.A(net3601),
    .X(net1746));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1123 (.A(net3605),
    .X(net1747));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1124 (.A(net3607),
    .X(net1748));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1125 (.A(net3339),
    .X(net1749));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1126 (.A(_0243_),
    .X(net1750));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1127 (.A(net3602),
    .X(net1751));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1128 (.A(net3604),
    .X(net1752));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1129 (.A(net3597),
    .X(net1753));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold113 (.A(net2381),
    .X(net737));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1130 (.A(_0303_),
    .X(net1754));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1131 (.A(net3643),
    .X(net1755));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1132 (.A(_0218_),
    .X(net1756));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1133 (.A(net3533),
    .X(net1757));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1134 (.A(_0569_),
    .X(net1758));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1135 (.A(net3630),
    .X(net1759));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1136 (.A(_0198_),
    .X(net1760));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1137 (.A(net3594),
    .X(net1761));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1138 (.A(net3596),
    .X(net1762));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1139 (.A(net3327),
    .X(net1763));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold114 (.A(net2538),
    .X(net738));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1140 (.A(_0242_),
    .X(net1764));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1141 (.A(net3645),
    .X(net1765));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1142 (.A(_0233_),
    .X(net1766));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1143 (.A(net3611),
    .X(net1767));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1144 (.A(_0293_),
    .X(net1768));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1145 (.A(net3576),
    .X(net1769));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1146 (.A(net3578),
    .X(net1770));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1147 (.A(net3608),
    .X(net1771));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1148 (.A(net3610),
    .X(net1772));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1149 (.A(net3659),
    .X(net1773));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold115 (.A(net2540),
    .X(net739));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1150 (.A(_0288_),
    .X(net1774));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1151 (.A(net3433),
    .X(net1775));
 sky130_fd_sc_hd__buf_12 hold1152 (.A(net1776),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1153 (.A(net3387),
    .X(net1777));
 sky130_fd_sc_hd__buf_12 hold1154 (.A(net1778),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1155 (.A(net3409),
    .X(net1779));
 sky130_fd_sc_hd__buf_12 hold1156 (.A(net1780),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1157 (.A(net3474),
    .X(net1781));
 sky130_fd_sc_hd__buf_12 hold1158 (.A(net1782),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1159 (.A(net3420),
    .X(net1783));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold116 (.A(net2433),
    .X(net740));
 sky130_fd_sc_hd__buf_12 hold1160 (.A(net1784),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1161 (.A(net3392),
    .X(net1785));
 sky130_fd_sc_hd__buf_12 hold1162 (.A(net1786),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1163 (.A(net3430),
    .X(net1787));
 sky130_fd_sc_hd__buf_12 hold1164 (.A(net1788),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1165 (.A(net3411),
    .X(net1789));
 sky130_fd_sc_hd__buf_12 hold1166 (.A(net1790),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1167 (.A(net3443),
    .X(net1791));
 sky130_fd_sc_hd__buf_12 hold1168 (.A(net1792),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1169 (.A(net3406),
    .X(net1793));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold117 (.A(_0695_),
    .X(net741));
 sky130_fd_sc_hd__buf_12 hold1170 (.A(net1794),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1171 (.A(net3681),
    .X(net1795));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1172 (.A(_0253_),
    .X(net1796));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1173 (.A(net3425),
    .X(net1797));
 sky130_fd_sc_hd__buf_12 hold1174 (.A(net1798),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1175 (.A(net3414),
    .X(net1799));
 sky130_fd_sc_hd__buf_12 hold1176 (.A(net1800),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1177 (.A(net3452),
    .X(net1801));
 sky130_fd_sc_hd__buf_12 hold1178 (.A(net1802),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1179 (.A(net3487),
    .X(net1803));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold118 (.A(net2357),
    .X(net742));
 sky130_fd_sc_hd__buf_12 hold1180 (.A(net1804),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1181 (.A(net3538),
    .X(net1805));
 sky130_fd_sc_hd__buf_12 hold1182 (.A(net1806),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1183 (.A(net3462),
    .X(net1807));
 sky130_fd_sc_hd__buf_12 hold1184 (.A(net1808),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1185 (.A(net3507),
    .X(net1809));
 sky130_fd_sc_hd__buf_12 hold1186 (.A(net1810),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1187 (.A(net3472),
    .X(net1811));
 sky130_fd_sc_hd__buf_12 hold1188 (.A(net1812),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1189 (.A(net3440),
    .X(net1813));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold119 (.A(net2359),
    .X(net743));
 sky130_fd_sc_hd__buf_12 hold1190 (.A(net1814),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1191 (.A(net3448),
    .X(net1815));
 sky130_fd_sc_hd__buf_12 hold1192 (.A(net1816),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1193 (.A(net3525),
    .X(net1817));
 sky130_fd_sc_hd__buf_12 hold1194 (.A(net1818),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1195 (.A(net3536),
    .X(net1819));
 sky130_fd_sc_hd__buf_12 hold1196 (.A(net1820),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1197 (.A(net3540),
    .X(net1821));
 sky130_fd_sc_hd__buf_12 hold1198 (.A(net1822),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1199 (.A(net3501),
    .X(net1823));
 sky130_fd_sc_hd__clkbuf_4 hold12 (.A(_0890_),
    .X(net636));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold120 (.A(net2492),
    .X(net744));
 sky130_fd_sc_hd__buf_12 hold1200 (.A(net1824),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1201 (.A(net3485),
    .X(net1825));
 sky130_fd_sc_hd__buf_12 hold1202 (.A(net1826),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1203 (.A(net3477),
    .X(net1827));
 sky130_fd_sc_hd__buf_12 hold1204 (.A(net1828),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1205 (.A(net3495),
    .X(net1829));
 sky130_fd_sc_hd__buf_12 hold1206 (.A(net1830),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1207 (.A(net3493),
    .X(net1831));
 sky130_fd_sc_hd__buf_12 hold1208 (.A(net1832),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1209 (.A(net3549),
    .X(net1833));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold121 (.A(net2494),
    .X(net745));
 sky130_fd_sc_hd__buf_12 hold1210 (.A(net1834),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1211 (.A(net3464),
    .X(net1835));
 sky130_fd_sc_hd__buf_12 hold1212 (.A(net1836),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1213 (.A(net3520),
    .X(net1837));
 sky130_fd_sc_hd__buf_12 hold1214 (.A(net1838),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__dlygate4sd1_1 hold1215 (.A(net3705),
    .X(net1839));
 sky130_fd_sc_hd__buf_12 hold1216 (.A(net1840),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1217 (.A(net3377),
    .X(net1841));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1218 (.A(net3379),
    .X(net1842));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1219 (.A(net3638),
    .X(net1843));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold122 (.A(net2495),
    .X(net746));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1220 (.A(_0258_),
    .X(net1844));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1221 (.A(net3683),
    .X(net1845));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1222 (.A(net3685),
    .X(net1846));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1223 (.A(net3657),
    .X(net1847));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1224 (.A(_0497_),
    .X(net1848));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1225 (.A(net3691),
    .X(net1849));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1226 (.A(_0120_),
    .X(net1850));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1227 (.A(net3625),
    .X(net1851));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1228 (.A(_0266_),
    .X(net1852));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1229 (.A(net3674),
    .X(net1853));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold123 (.A(net2497),
    .X(net747));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1230 (.A(net3676),
    .X(net1854));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1231 (.A(net3702),
    .X(net1855));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1232 (.A(_0553_),
    .X(net1856));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1233 (.A(net3588),
    .X(net1857));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1234 (.A(net3712),
    .X(net1858));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1235 (.A(_0745_),
    .X(net1859));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1236 (.A(net3698),
    .X(net1860));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1237 (.A(_0625_),
    .X(net1861));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1238 (.A(net3581),
    .X(net1862));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1239 (.A(net3573),
    .X(net1863));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold124 (.A(net2541),
    .X(net748));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1240 (.A(net3706),
    .X(net1864));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1241 (.A(_0697_),
    .X(net1865));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1242 (.A(net3563),
    .X(net1866));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1243 (.A(_2586_),
    .X(net1867));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1244 (.A(_0419_),
    .X(net1868));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1245 (.A(net3622),
    .X(net1869));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1246 (.A(net3708),
    .X(net1870));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1247 (.A(_0737_),
    .X(net1871));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1248 (.A(net3717),
    .X(net1872));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1249 (.A(_0657_),
    .X(net1873));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold125 (.A(net2543),
    .X(net749));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1250 (.A(net3719),
    .X(net1874));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1251 (.A(net3721),
    .X(net1875));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1252 (.A(net3732),
    .X(net1876));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1253 (.A(net3734),
    .X(net1877));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1254 (.A(net3688),
    .X(net1878));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1255 (.A(net3690),
    .X(net1879));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1256 (.A(net3772),
    .X(net1880));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1257 (.A(_0729_),
    .X(net1881));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1258 (.A(net3740),
    .X(net1882));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1259 (.A(net3742),
    .X(net1883));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold126 (.A(net3152),
    .X(net750));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1260 (.A(net3693),
    .X(net1884));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1261 (.A(_0252_),
    .X(net1885));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1262 (.A(net3700),
    .X(net1886));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1263 (.A(_0545_),
    .X(net1887));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1264 (.A(net3765),
    .X(net1888));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1265 (.A(net3767),
    .X(net1889));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1266 (.A(net3743),
    .X(net1890));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1267 (.A(net3745),
    .X(net1891));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1268 (.A(net3722),
    .X(net1892));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1269 (.A(_0192_),
    .X(net1893));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold127 (.A(_0351_),
    .X(net751));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1270 (.A(net3776),
    .X(net1894));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1271 (.A(net3778),
    .X(net1895));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1272 (.A(net3735),
    .X(net1896));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1273 (.A(_0337_),
    .X(net1897));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1274 (.A(net3763),
    .X(net1898));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1275 (.A(_0347_),
    .X(net1899));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1276 (.A(net3737),
    .X(net1900));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1277 (.A(net3739),
    .X(net1901));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1278 (.A(net3724),
    .X(net1902));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1279 (.A(_0327_),
    .X(net1903));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold128 (.A(net3141),
    .X(net752));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1280 (.A(net3760),
    .X(net1904));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1281 (.A(net3762),
    .X(net1905));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1282 (.A(net3728),
    .X(net1906));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1283 (.A(_0379_),
    .X(net1907));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1284 (.A(net3774),
    .X(net1908));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1285 (.A(_0357_),
    .X(net1909));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1286 (.A(net3714),
    .X(net1910));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1287 (.A(net3716),
    .X(net1911));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1288 (.A(net3768),
    .X(net1912));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1289 (.A(_0521_),
    .X(net1913));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold129 (.A(_0469_),
    .X(net753));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1290 (.A(net3669),
    .X(net1914));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1291 (.A(net3671),
    .X(net1915));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1292 (.A(net3770),
    .X(net1916));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1293 (.A(_0197_),
    .X(net1917));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1294 (.A(net3710),
    .X(net1918));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1295 (.A(_0202_),
    .X(net1919));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1296 (.A(net3784),
    .X(net1920));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1297 (.A(_0187_),
    .X(net1921));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1298 (.A(net3726),
    .X(net1922));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1299 (.A(_0222_),
    .X(net1923));
 sky130_fd_sc_hd__clkbuf_8 hold13 (.A(_2628_),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_2 hold130 (.A(net2111),
    .X(net754));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1300 (.A(net3652),
    .X(net1924));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1301 (.A(net3654),
    .X(net1925));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1302 (.A(net3749),
    .X(net1926));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1303 (.A(net3751),
    .X(net1927));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1304 (.A(net3781),
    .X(net1928));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1305 (.A(net3754),
    .X(net1929));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1306 (.A(net3756),
    .X(net1930));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1307 (.A(net3568),
    .X(net1931));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1308 (.A(net3570),
    .X(net1932));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1309 (.A(net3757),
    .X(net1933));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold131 (.A(net2113),
    .X(net755));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1310 (.A(net3759),
    .X(net1934));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1311 (.A(net3786),
    .X(net1935));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1312 (.A(_0705_),
    .X(net1936));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1313 (.A(net3686),
    .X(net1937));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1314 (.A(_0435_),
    .X(net1938));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1315 (.A(net3788),
    .X(net1939));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1316 (.A(_0513_),
    .X(net1940));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1317 (.A(net3695),
    .X(net1941));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1318 (.A(net3697),
    .X(net1942));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1319 (.A(net3790),
    .X(net1943));
 sky130_fd_sc_hd__buf_4 hold132 (.A(_0883_),
    .X(net756));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1320 (.A(_0101_),
    .X(net1944));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1321 (.A(net3746),
    .X(net1945));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1322 (.A(net3748),
    .X(net1946));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1323 (.A(net3794),
    .X(net1947));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1324 (.A(_0109_),
    .X(net1948));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1325 (.A(net3779),
    .X(net1949));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1326 (.A(_0174_),
    .X(net1950));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1327 (.A(net3730),
    .X(net1951));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1328 (.A(_0207_),
    .X(net1952));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1329 (.A(net3796),
    .X(net1953));
 sky130_fd_sc_hd__buf_4 hold133 (.A(_2627_),
    .X(net757));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1330 (.A(_0577_),
    .X(net1954));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1331 (.A(net3792),
    .X(net1955));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1332 (.A(_0405_),
    .X(net1956));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1333 (.A(net3752),
    .X(net1957));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1334 (.A(_0312_),
    .X(net1958));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1335 (.A(net3432),
    .X(net1959));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1336 (.A(net3386),
    .X(net1960));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1337 (.A(net3408),
    .X(net1961));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1338 (.A(net3419),
    .X(net1962));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1339 (.A(net3391),
    .X(net1963));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold134 (.A(net2531),
    .X(net758));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1340 (.A(net3429),
    .X(net1964));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1341 (.A(net3473),
    .X(net1965));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1342 (.A(net3442),
    .X(net1966));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1343 (.A(net3405),
    .X(net1967));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1344 (.A(net3410),
    .X(net1968));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1345 (.A(net3506),
    .X(net1969));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1346 (.A(net3413),
    .X(net1970));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1347 (.A(net3424),
    .X(net1971));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1348 (.A(net3451),
    .X(net1972));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1349 (.A(net3461),
    .X(net1973));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold135 (.A(net2626),
    .X(net759));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1350 (.A(net3486),
    .X(net1974));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1351 (.A(net3471),
    .X(net1975));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1352 (.A(net3439),
    .X(net1976));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1353 (.A(net3447),
    .X(net1977));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1354 (.A(net3524),
    .X(net1978));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1355 (.A(net3500),
    .X(net1979));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1356 (.A(net3484),
    .X(net1980));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1357 (.A(net3476),
    .X(net1981));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1358 (.A(net3494),
    .X(net1982));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1359 (.A(net3492),
    .X(net1983));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold136 (.A(net2628),
    .X(net760));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1360 (.A(net3463),
    .X(net1984));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1361 (.A(net3519),
    .X(net1985));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1362 (.A(net3537),
    .X(net1986));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1363 (.A(net3535),
    .X(net1987));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1364 (.A(net3539),
    .X(net1988));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1365 (.A(net3548),
    .X(net1989));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1366 (.A(net3704),
    .X(net1990));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1367 (.A(\mgmt_gpio_data_buf[13] ),
    .X(net1991));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1368 (.A(net2018),
    .X(net1992));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1369 (.A(net2742),
    .X(net1993));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold137 (.A(net3074),
    .X(net761));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1370 (.A(\gpio_configure[37][2] ),
    .X(net1994));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1371 (.A(net2034),
    .X(net1995));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1372 (.A(net2201),
    .X(net1996));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1373 (.A(net2529),
    .X(net1997));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1374 (.A(net2036),
    .X(net1998));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1375 (.A(net2038),
    .X(net1999));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1376 (.A(net2119),
    .X(net2000));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1377 (.A(\gpio_configure[30][9] ),
    .X(net2001));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1378 (.A(net2392),
    .X(net2002));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1379 (.A(net2130),
    .X(net2003));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold138 (.A(_0485_),
    .X(net762));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1380 (.A(net2415),
    .X(net2004));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1381 (.A(net2905),
    .X(net2005));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1382 (.A(\gpio_configure[8][3] ),
    .X(net2006));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1383 (.A(net2028),
    .X(net2007));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1384 (.A(net2323),
    .X(net2008));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1385 (.A(net2760),
    .X(net2009));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1386 (.A(net2550),
    .X(net2010));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1387 (.A(net2368),
    .X(net2011));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1388 (.A(net2770),
    .X(net2012));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1389 (.A(\gpio_configure[14][1] ),
    .X(net2013));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold139 (.A(net2733),
    .X(net763));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1390 (.A(\hkspi.odata[5] ),
    .X(net2014));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1391 (.A(net625),
    .X(net2015));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1392 (.A(_1467_),
    .X(net2016));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1393 (.A(net626),
    .X(net2017));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1394 (.A(_0140_),
    .X(net2018));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1395 (.A(net1992),
    .X(net2019));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1396 (.A(\mgmt_gpio_data[13] ),
    .X(net2020));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1397 (.A(net714),
    .X(net2021));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1398 (.A(_0124_),
    .X(net2022));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1399 (.A(net715),
    .X(net2023));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold14 (.A(net1999),
    .X(net638));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold140 (.A(net2735),
    .X(net764));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1400 (.A(\hkspi.odata[3] ),
    .X(net2024));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1401 (.A(net628),
    .X(net2025));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1402 (.A(_1464_),
    .X(net2026));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1403 (.A(net629),
    .X(net2027));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1404 (.A(_0516_),
    .X(net2028));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1405 (.A(net2007),
    .X(net2029));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1406 (.A(\hkspi.odata[2] ),
    .X(net2030));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1407 (.A(net631),
    .X(net2031));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1408 (.A(_1463_),
    .X(net2032));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1409 (.A(net632),
    .X(net2033));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold141 (.A(net2773),
    .X(net765));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1410 (.A(_0747_),
    .X(net2034));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1411 (.A(net1995),
    .X(net2035));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1412 (.A(\gpio_configure[34][2] ),
    .X(net2036));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1413 (.A(net1998),
    .X(net2037));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1414 (.A(_0723_),
    .X(net2038));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1415 (.A(wbbd_write),
    .X(net2039));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1416 (.A(net669),
    .X(net2040));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1417 (.A(_1459_),
    .X(net2041));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1418 (.A(net670),
    .X(net2042));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1419 (.A(_2584_),
    .X(net2043));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold142 (.A(net2775),
    .X(net766));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1420 (.A(_0416_),
    .X(net2044));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1421 (.A(net800),
    .X(net2045));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1422 (.A(\gpio_configure[6][2] ),
    .X(net2046));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1423 (.A(net817),
    .X(net2047));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1424 (.A(_0499_),
    .X(net2048));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1425 (.A(net818),
    .X(net2049));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1426 (.A(\gpio_configure[24][2] ),
    .X(net2050));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1427 (.A(net845),
    .X(net2051));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1428 (.A(_0643_),
    .X(net2052));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1429 (.A(net846),
    .X(net2053));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold143 (.A(net2720),
    .X(net767));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1430 (.A(\mgmt_gpio_data_buf[2] ),
    .X(net2054));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1431 (.A(net805),
    .X(net2055));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1432 (.A(_0443_),
    .X(net2056));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1433 (.A(net806),
    .X(net2057));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1434 (.A(\gpio_configure[7][2] ),
    .X(net2058));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1435 (.A(net825),
    .X(net2059));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1436 (.A(_0507_),
    .X(net2060));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1437 (.A(net826),
    .X(net2061));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1438 (.A(\gpio_configure[2][2] ),
    .X(net2062));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1439 (.A(net815),
    .X(net2063));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold144 (.A(net2722),
    .X(net768));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1440 (.A(_0467_),
    .X(net2064));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1441 (.A(net816),
    .X(net2065));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1442 (.A(\wbbd_addr[0] ),
    .X(net2066));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1443 (.A(net634),
    .X(net2067));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1444 (.A(_0850_),
    .X(net2068));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1445 (.A(net635),
    .X(net2069));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1446 (.A(_0854_),
    .X(net2070));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1447 (.A(_0952_),
    .X(net2071));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1448 (.A(_2620_),
    .X(net2072));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1449 (.A(_0662_),
    .X(net2073));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold145 (.A(net2763),
    .X(net769));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1450 (.A(net812),
    .X(net2074));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1451 (.A(\gpio_configure[3][2] ),
    .X(net2075));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1452 (.A(net813),
    .X(net2076));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1453 (.A(_0475_),
    .X(net2077));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1454 (.A(net814),
    .X(net2078));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1455 (.A(\mgmt_gpio_data[37] ),
    .X(net2079));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1456 (.A(net801),
    .X(net2080));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1457 (.A(_0440_),
    .X(net2081));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1458 (.A(net802),
    .X(net2082));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1459 (.A(\gpio_configure[29][5] ),
    .X(net2083));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold146 (.A(net2765),
    .X(net770));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1460 (.A(net795),
    .X(net2084));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1461 (.A(_0686_),
    .X(net2085));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1462 (.A(net796),
    .X(net2086));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1463 (.A(\wbbd_addr[3] ),
    .X(net2087));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1464 (.A(net693),
    .X(net2088));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1465 (.A(_0844_),
    .X(net2089));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1466 (.A(net694),
    .X(net2090));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1467 (.A(_0887_),
    .X(net2091));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1468 (.A(net407),
    .X(net2092));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1469 (.A(_0926_),
    .X(net2093));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold147 (.A(net2726),
    .X(net771));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1470 (.A(_2595_),
    .X(net2094));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1471 (.A(_0459_),
    .X(net2095));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1472 (.A(net822),
    .X(net2096));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1473 (.A(\hkspi.odata[7] ),
    .X(net2097));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1474 (.A(net639),
    .X(net2098));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1475 (.A(_1469_),
    .X(net2099));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1476 (.A(net640),
    .X(net2100));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1477 (.A(net467),
    .X(net2101));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1478 (.A(_0616_),
    .X(net2102));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1479 (.A(net652),
    .X(net2103));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold148 (.A(net2728),
    .X(net772));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1480 (.A(\gpio_configure[23][5] ),
    .X(net2104));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1481 (.A(net803),
    .X(net2105));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1482 (.A(_0638_),
    .X(net2106));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1483 (.A(net804),
    .X(net2107));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1484 (.A(\mgmt_gpio_data[29] ),
    .X(net2108));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1485 (.A(net809),
    .X(net2109));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1486 (.A(_0271_),
    .X(net2110));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1487 (.A(\wbbd_addr[4] ),
    .X(net2111));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1488 (.A(net754),
    .X(net2112));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1489 (.A(_0841_),
    .X(net2113));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold149 (.A(net2750),
    .X(net773));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1490 (.A(_0879_),
    .X(net2114));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1491 (.A(net679),
    .X(net2115));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1492 (.A(_2619_),
    .X(net2116));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1493 (.A(_0651_),
    .X(net2117));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1494 (.A(net838),
    .X(net2118));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1495 (.A(\gpio_configure[31][7] ),
    .X(net2119));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1496 (.A(net2000),
    .X(net2120));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1497 (.A(_0704_),
    .X(net2121));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1498 (.A(net648),
    .X(net2122));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1499 (.A(\gpio_configure[20][5] ),
    .X(net2123));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold15 (.A(net2097),
    .X(net639));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold150 (.A(net2752),
    .X(net774));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1500 (.A(net797),
    .X(net2124));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1501 (.A(_0614_),
    .X(net2125));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1502 (.A(net798),
    .X(net2126));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1503 (.A(\gpio_configure[27][5] ),
    .X(net2127));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1504 (.A(net849),
    .X(net2128));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1505 (.A(_0670_),
    .X(net2129));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1506 (.A(\gpio_configure[35][7] ),
    .X(net2130));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1507 (.A(net2003),
    .X(net2131));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1508 (.A(_0736_),
    .X(net2132));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1509 (.A(\gpio_configure[30][7] ),
    .X(net2133));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold151 (.A(net3172),
    .X(net775));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1510 (.A(net649),
    .X(net2134));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1511 (.A(_0696_),
    .X(net2135));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1512 (.A(\gpio_configure[35][5] ),
    .X(net2136));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1513 (.A(net833),
    .X(net2137));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1514 (.A(_0734_),
    .X(net2138));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1515 (.A(\gpio_configure[29][2] ),
    .X(net2139));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1516 (.A(net807),
    .X(net2140));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1517 (.A(_0683_),
    .X(net2141));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1518 (.A(net808),
    .X(net2142));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1519 (.A(\mgmt_gpio_data_buf[18] ),
    .X(net2143));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold152 (.A(net3174),
    .X(net776));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1520 (.A(net841),
    .X(net2144));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1521 (.A(_0276_),
    .X(net2145));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1522 (.A(\gpio_configure[0][2] ),
    .X(net2146));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1523 (.A(net827),
    .X(net2147));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1524 (.A(_0451_),
    .X(net2148));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1525 (.A(net828),
    .X(net2149));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1526 (.A(\gpio_configure[34][7] ),
    .X(net2150));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1527 (.A(net655),
    .X(net2151));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1528 (.A(_0728_),
    .X(net2152));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1529 (.A(\gpio_configure[31][5] ),
    .X(net2153));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold153 (.A(\hkspi.addr[0] ),
    .X(net777));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1530 (.A(net835),
    .X(net2154));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1531 (.A(_0702_),
    .X(net2155));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1532 (.A(net836),
    .X(net2156));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1533 (.A(\gpio_configure[19][7] ),
    .X(net2157));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1534 (.A(net653),
    .X(net2158));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1535 (.A(_0608_),
    .X(net2159));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1536 (.A(net654),
    .X(net2160));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1537 (.A(\gpio_configure[33][2] ),
    .X(net2161));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1538 (.A(net823),
    .X(net2162));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1539 (.A(_0715_),
    .X(net2163));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold154 (.A(_0849_),
    .X(net778));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1540 (.A(net824),
    .X(net2164));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1541 (.A(\gpio_configure[29][3] ),
    .X(net2165));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1542 (.A(net853),
    .X(net2166));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1543 (.A(_0684_),
    .X(net2167));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1544 (.A(net854),
    .X(net2168));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1545 (.A(\gpio_configure[37][5] ),
    .X(net2169));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1546 (.A(net831),
    .X(net2170));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1547 (.A(_0750_),
    .X(net2171));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1548 (.A(\gpio_configure[18][5] ),
    .X(net2172));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1549 (.A(net895),
    .X(net2173));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold155 (.A(_0851_),
    .X(net779));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1550 (.A(_0598_),
    .X(net2174));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1551 (.A(net896),
    .X(net2175));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1552 (.A(\gpio_configure[28][5] ),
    .X(net2176));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1553 (.A(net829),
    .X(net2177));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1554 (.A(_0678_),
    .X(net2178));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1555 (.A(net830),
    .X(net2179));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1556 (.A(\mgmt_gpio_data[26] ),
    .X(net2180));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1557 (.A(net819),
    .X(net2181));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1558 (.A(_0268_),
    .X(net2182));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1559 (.A(\clk1_output_dest[0] ),
    .X(net2183));
 sky130_fd_sc_hd__buf_2 hold156 (.A(_1544_),
    .X(net780));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1560 (.A(net847),
    .X(net2184));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1561 (.A(_0428_),
    .X(net2185));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1562 (.A(net848),
    .X(net2186));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1563 (.A(\gpio_configure[30][5] ),
    .X(net2187));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1564 (.A(net839),
    .X(net2188));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1565 (.A(_0694_),
    .X(net2189));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1566 (.A(\gpio_configure[21][5] ),
    .X(net2190));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1567 (.A(net843),
    .X(net2191));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1568 (.A(_0622_),
    .X(net2192));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1569 (.A(net844),
    .X(net2193));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold157 (.A(net2762),
    .X(net781));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1570 (.A(\gpio_configure[27][3] ),
    .X(net2194));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1571 (.A(net865),
    .X(net2195));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1572 (.A(_0668_),
    .X(net2196));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1573 (.A(\gpio_configure[9][2] ),
    .X(net2197));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1574 (.A(net891),
    .X(net2198));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1575 (.A(_0523_),
    .X(net2199));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1576 (.A(net892),
    .X(net2200));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1577 (.A(\gpio_configure[37][7] ),
    .X(net2201));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1578 (.A(net1996),
    .X(net2202));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1579 (.A(_0752_),
    .X(net2203));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold158 (.A(net2729),
    .X(net782));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1580 (.A(\gpio_configure[25][5] ),
    .X(net2204));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1581 (.A(net851),
    .X(net2205));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1582 (.A(\wbbd_addr[1] ),
    .X(net2206));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1583 (.A(net643),
    .X(net2207));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1584 (.A(_0853_),
    .X(net2208));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1585 (.A(net644),
    .X(net2209));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1586 (.A(_0885_),
    .X(net2210));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1587 (.A(_0244_),
    .X(net2211));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1588 (.A(net981),
    .X(net2212));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1589 (.A(\gpio_configure[12][2] ),
    .X(net2213));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold159 (.A(net2731),
    .X(net783));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1590 (.A(net863),
    .X(net2214));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1591 (.A(_0547_),
    .X(net2215));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1592 (.A(net864),
    .X(net2216));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1593 (.A(\gpio_configure[24][10] ),
    .X(net2217));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1594 (.A(net922),
    .X(net2218));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1595 (.A(_0249_),
    .X(net2219));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1596 (.A(\gpio_configure[4][2] ),
    .X(net2220));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1597 (.A(net889),
    .X(net2221));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1598 (.A(_0483_),
    .X(net2222));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1599 (.A(\gpio_configure[13][2] ),
    .X(net2223));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold16 (.A(net2099),
    .X(net640));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold160 (.A(net2779),
    .X(net784));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1600 (.A(net887),
    .X(net2224));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1601 (.A(_0555_),
    .X(net2225));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1602 (.A(\gpio_configure[31][3] ),
    .X(net2226));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1603 (.A(net859),
    .X(net2227));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1604 (.A(_0700_),
    .X(net2228));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1605 (.A(net860),
    .X(net2229));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1606 (.A(\gpio_configure[27][2] ),
    .X(net2230));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1607 (.A(net899),
    .X(net2231));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1608 (.A(_0667_),
    .X(net2232));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1609 (.A(\gpio_configure[12][7] ),
    .X(net2233));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold161 (.A(net2781),
    .X(net785));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1610 (.A(net663),
    .X(net2234));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1611 (.A(_0552_),
    .X(net2235));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1612 (.A(net664),
    .X(net2236));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1613 (.A(\gpio_configure[34][5] ),
    .X(net2237));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1614 (.A(net879),
    .X(net2238));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1615 (.A(_0726_),
    .X(net2239));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1616 (.A(\mgmt_gpio_data_buf[19] ),
    .X(net2240));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1617 (.A(net883),
    .X(net2241));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1618 (.A(_0277_),
    .X(net2242));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1619 (.A(\gpio_configure[25][3] ),
    .X(net2243));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold162 (.A(net2748),
    .X(net786));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1620 (.A(net855),
    .X(net2244));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1621 (.A(\gpio_configure[6][3] ),
    .X(net2245));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1622 (.A(net867),
    .X(net2246));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1623 (.A(_0500_),
    .X(net2247));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1624 (.A(\mgmt_gpio_data_buf[10] ),
    .X(net2248));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1625 (.A(net873),
    .X(net2249));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1626 (.A(_0137_),
    .X(net2250));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1627 (.A(\gpio_configure[28][3] ),
    .X(net2251));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1628 (.A(net871),
    .X(net2252));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1629 (.A(_0676_),
    .X(net2253));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold163 (.A(_0677_),
    .X(net787));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1630 (.A(\gpio_configure[30][10] ),
    .X(net2254));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1631 (.A(net948),
    .X(net2255));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1632 (.A(_0359_),
    .X(net2256));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1633 (.A(\gpio_configure[33][5] ),
    .X(net2257));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1634 (.A(net885),
    .X(net2258));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1635 (.A(_0718_),
    .X(net2259));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1636 (.A(net886),
    .X(net2260));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1637 (.A(\mgmt_gpio_data[27] ),
    .X(net2261));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1638 (.A(net877),
    .X(net2262));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1639 (.A(_0269_),
    .X(net2263));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold164 (.A(net2766),
    .X(net788));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1640 (.A(\gpio_configure[33][10] ),
    .X(net2264));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1641 (.A(net964),
    .X(net2265));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1642 (.A(_0329_),
    .X(net2266));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1643 (.A(\gpio_configure[10][3] ),
    .X(net2267));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1644 (.A(net881),
    .X(net2268));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1645 (.A(_0532_),
    .X(net2269));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1646 (.A(net882),
    .X(net2270));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1647 (.A(net282),
    .X(net2271));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1648 (.A(net897),
    .X(net2272));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1649 (.A(_0410_),
    .X(net2273));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold165 (.A(net2768),
    .X(net789));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1650 (.A(\gpio_configure[26][10] ),
    .X(net2274));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1651 (.A(net998),
    .X(net2275));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1652 (.A(\gpio_configure[5][10] ),
    .X(net2276));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1653 (.A(net944),
    .X(net2277));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1654 (.A(_0194_),
    .X(net2278));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1655 (.A(net945),
    .X(net2279));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1656 (.A(\gpio_configure[13][3] ),
    .X(net2280));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1657 (.A(net914),
    .X(net2281));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1658 (.A(_0556_),
    .X(net2282));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1659 (.A(\hkspi.odata[6] ),
    .X(net2283));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold166 (.A(\wbbd_data[4] ),
    .X(net790));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1660 (.A(net683),
    .X(net2284));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1661 (.A(_1468_),
    .X(net2285));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1662 (.A(net684),
    .X(net2286));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1663 (.A(net470),
    .X(net2287));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1664 (.A(_0679_),
    .X(net2288));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1665 (.A(net701),
    .X(net2289));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1666 (.A(\gpio_configure[20][3] ),
    .X(net2290));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1667 (.A(net869),
    .X(net2291));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1668 (.A(_0612_),
    .X(net2292));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1669 (.A(net290),
    .X(net2293));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold167 (.A(net2694),
    .X(net791));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1670 (.A(_0114_),
    .X(net2294));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1671 (.A(\wbbd_addr[2] ),
    .X(net2295));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1672 (.A(net657),
    .X(net2296));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1673 (.A(_0846_),
    .X(net2297));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1674 (.A(net658),
    .X(net2298));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1675 (.A(_0339_),
    .X(net2299));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1676 (.A(net943),
    .X(net2300));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1677 (.A(\gpio_configure[36][5] ),
    .X(net2301));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1678 (.A(net857),
    .X(net2302));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1679 (.A(_0742_),
    .X(net2303));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold168 (.A(net2772),
    .X(net792));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1680 (.A(\gpio_configure[19][5] ),
    .X(net2304));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1681 (.A(net875),
    .X(net2305));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1682 (.A(_0606_),
    .X(net2306));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1683 (.A(\gpio_configure[22][5] ),
    .X(net2307));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1684 (.A(net962),
    .X(net2308));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1685 (.A(_0630_),
    .X(net2309));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1686 (.A(net257),
    .X(net2310));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1687 (.A(net893),
    .X(net2311));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1688 (.A(_0404_),
    .X(net2312));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1689 (.A(\mgmt_gpio_data[30] ),
    .X(net2313));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold169 (.A(net2782),
    .X(net793));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1690 (.A(net702),
    .X(net2314));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1691 (.A(_0272_),
    .X(net2315));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1692 (.A(\gpio_configure[7][5] ),
    .X(net2316));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1693 (.A(net982),
    .X(net2317));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1694 (.A(_0510_),
    .X(net2318));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1695 (.A(net983),
    .X(net2319));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1696 (.A(\gpio_configure[11][2] ),
    .X(net2320));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1697 (.A(net1038),
    .X(net2321));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1698 (.A(_0539_),
    .X(net2322));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1699 (.A(\gpio_configure[29][6] ),
    .X(net2323));
 sky130_fd_sc_hd__buf_8 hold17 (.A(net2101),
    .X(net641));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold170 (.A(net2784),
    .X(net794));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1700 (.A(net2008),
    .X(net2324));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1701 (.A(_0687_),
    .X(net2325));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1702 (.A(\gpio_configure[31][2] ),
    .X(net2326));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1703 (.A(net936),
    .X(net2327));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1704 (.A(_0699_),
    .X(net2328));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1705 (.A(\gpio_configure[11][3] ),
    .X(net2329));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1706 (.A(net912),
    .X(net2330));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1707 (.A(_0540_),
    .X(net2331));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1708 (.A(\gpio_configure[18][10] ),
    .X(net2332));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1709 (.A(net956),
    .X(net2333));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold171 (.A(net2083),
    .X(net795));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1710 (.A(_0334_),
    .X(net2334));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1711 (.A(serial_bb_data_1),
    .X(net2335));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1712 (.A(net960),
    .X(net2336));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1713 (.A(_0423_),
    .X(net2337));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1714 (.A(net961),
    .X(net2338));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1715 (.A(\gpio_configure[2][3] ),
    .X(net2339));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1716 (.A(net930),
    .X(net2340));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1717 (.A(_0468_),
    .X(net2341));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1718 (.A(\gpio_configure[37][3] ),
    .X(net2342));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1719 (.A(net901),
    .X(net2343));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold172 (.A(net2085),
    .X(net796));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1720 (.A(_0748_),
    .X(net2344));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1721 (.A(\hkspi.odata[1] ),
    .X(net2345));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1722 (.A(net665),
    .X(net2346));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1723 (.A(_1462_),
    .X(net2347));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1724 (.A(net666),
    .X(net2348));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1725 (.A(net494),
    .X(net2349));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1726 (.A(_0358_),
    .X(net2350));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1727 (.A(net682),
    .X(net2351));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1728 (.A(\gpio_configure[31][10] ),
    .X(net2352));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1729 (.A(net976),
    .X(net2353));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold173 (.A(net2123),
    .X(net797));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1730 (.A(\mgmt_gpio_data_buf[5] ),
    .X(net2354));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1731 (.A(net940),
    .X(net2355));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1732 (.A(_0446_),
    .X(net2356));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1733 (.A(\gpio_configure[31][6] ),
    .X(net2357));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1734 (.A(net742),
    .X(net2358));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1735 (.A(_0703_),
    .X(net2359));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1736 (.A(\gpio_configure[23][10] ),
    .X(net2360));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1737 (.A(net1032),
    .X(net2361));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1738 (.A(_0239_),
    .X(net2362));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1739 (.A(\gpio_configure[23][3] ),
    .X(net2363));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold174 (.A(net2125),
    .X(net798));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1740 (.A(net861),
    .X(net2364));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1741 (.A(_0636_),
    .X(net2365));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1742 (.A(\gpio_configure[27][11] ),
    .X(net2366));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1743 (.A(net1006),
    .X(net2367));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1744 (.A(\gpio_configure[13][1] ),
    .X(net2368));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1745 (.A(net2011),
    .X(net2369));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1746 (.A(_0554_),
    .X(net2370));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1747 (.A(\gpio_configure[35][3] ),
    .X(net2371));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1748 (.A(net920),
    .X(net2372));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1749 (.A(_0732_),
    .X(net2373));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold175 (.A(net297),
    .X(net799));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1750 (.A(\gpio_configure[25][6] ),
    .X(net2374));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1751 (.A(net704),
    .X(net2375));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1752 (.A(\gpio_configure[11][1] ),
    .X(net2376));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1753 (.A(net698),
    .X(net2377));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1754 (.A(_0538_),
    .X(net2378));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1755 (.A(\gpio_configure[23][6] ),
    .X(net2379));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1756 (.A(net736),
    .X(net2380));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1757 (.A(_0639_),
    .X(net2381));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1758 (.A(\gpio_configure[37][1] ),
    .X(net2382));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1759 (.A(net691),
    .X(net2383));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold176 (.A(net2044),
    .X(net800));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1760 (.A(_0746_),
    .X(net2384));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1761 (.A(\gpio_configure[33][3] ),
    .X(net2385));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1762 (.A(net926),
    .X(net2386));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1763 (.A(_0716_),
    .X(net2387));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1764 (.A(\gpio_configure[3][3] ),
    .X(net2388));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1765 (.A(net908),
    .X(net2389));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1766 (.A(_0476_),
    .X(net2390));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1767 (.A(net909),
    .X(net2391));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1768 (.A(\gpio_configure[24][9] ),
    .X(net2392));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1769 (.A(net2002),
    .X(net2393));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold177 (.A(net2079),
    .X(net801));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1770 (.A(_0248_),
    .X(net2394));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1771 (.A(\gpio_configure[1][3] ),
    .X(net2395));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1772 (.A(net918),
    .X(net2396));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1773 (.A(\gpio_configure[14][3] ),
    .X(net2397));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1774 (.A(net958),
    .X(net2398));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1775 (.A(_0564_),
    .X(net2399));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1776 (.A(net959),
    .X(net2400));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1777 (.A(\gpio_configure[36][3] ),
    .X(net2401));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1778 (.A(net1010),
    .X(net2402));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1779 (.A(_0740_),
    .X(net2403));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold178 (.A(net2081),
    .X(net802));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1780 (.A(\mgmt_gpio_data_buf[21] ),
    .X(net2404));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1781 (.A(net1002),
    .X(net2405));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1782 (.A(_0279_),
    .X(net2406));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1783 (.A(\gpio_configure[28][10] ),
    .X(net2407));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1784 (.A(net1042),
    .X(net2408));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1785 (.A(\gpio_configure[35][2] ),
    .X(net2409));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1786 (.A(net932),
    .X(net2410));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1787 (.A(_0731_),
    .X(net2411));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1788 (.A(\gpio_configure[15][2] ),
    .X(net2412));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1789 (.A(net1026),
    .X(net2413));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold179 (.A(net2104),
    .X(net803));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1790 (.A(_0571_),
    .X(net2414));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1791 (.A(\gpio_configure[35][6] ),
    .X(net2415));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1792 (.A(net2004),
    .X(net2416));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1793 (.A(_0735_),
    .X(net2417));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1794 (.A(\gpio_configure[34][3] ),
    .X(net2418));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1795 (.A(net988),
    .X(net2419));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1796 (.A(_0724_),
    .X(net2420));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1797 (.A(\gpio_configure[26][3] ),
    .X(net2421));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1798 (.A(net954),
    .X(net2422));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1799 (.A(\gpio_configure[4][3] ),
    .X(net2423));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold18 (.A(net2132),
    .X(net642));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold180 (.A(net2106),
    .X(net804));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1800 (.A(net968),
    .X(net2424));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1801 (.A(_0484_),
    .X(net2425));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1802 (.A(\gpio_configure[7][3] ),
    .X(net2426));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1803 (.A(net992),
    .X(net2427));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1804 (.A(_0508_),
    .X(net2428));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1805 (.A(net993),
    .X(net2429));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1806 (.A(\gpio_configure[22][2] ),
    .X(net2430));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1807 (.A(net1036),
    .X(net2431));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1808 (.A(_0627_),
    .X(net2432));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1809 (.A(\gpio_configure[30][6] ),
    .X(net2433));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold181 (.A(net2054),
    .X(net805));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1810 (.A(net740),
    .X(net2434));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1811 (.A(\gpio_configure[23][11] ),
    .X(net2435));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1812 (.A(net996),
    .X(net2436));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1813 (.A(_0240_),
    .X(net2437));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1814 (.A(\gpio_configure[19][2] ),
    .X(net2438));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1815 (.A(net1044),
    .X(net2439));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1816 (.A(_0603_),
    .X(net2440));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1817 (.A(\gpio_configure[19][11] ),
    .X(net2441));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1818 (.A(net1000),
    .X(net2442));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1819 (.A(_0345_),
    .X(net2443));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold182 (.A(net2056),
    .X(net806));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1820 (.A(\gpio_configure[36][2] ),
    .X(net2444));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1821 (.A(net928),
    .X(net2445));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1822 (.A(_0739_),
    .X(net2446));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1823 (.A(\gpio_configure[32][3] ),
    .X(net2447));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1824 (.A(net1004),
    .X(net2448));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1825 (.A(\hkspi.addr[5] ),
    .X(net2449));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1826 (.A(_0831_),
    .X(net2450));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1827 (.A(_0832_),
    .X(net2451));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1828 (.A(net904),
    .X(net2452));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1829 (.A(_0894_),
    .X(net2453));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold183 (.A(net2139),
    .X(net807));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1830 (.A(net379),
    .X(net2454));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1831 (.A(_0199_),
    .X(net2455));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1832 (.A(net1095),
    .X(net2456));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1833 (.A(\gpio_configure[2][11] ),
    .X(net2457));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1834 (.A(net950),
    .X(net2458));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1835 (.A(\mgmt_gpio_data_buf[3] ),
    .X(net2459));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1836 (.A(net910),
    .X(net2460));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1837 (.A(_0444_),
    .X(net2461));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1838 (.A(\gpio_configure[7][9] ),
    .X(net2462));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1839 (.A(net689),
    .X(net2463));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold184 (.A(net2141),
    .X(net808));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1840 (.A(\gpio_configure[30][2] ),
    .X(net2464));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1841 (.A(net986),
    .X(net2465));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1842 (.A(\gpio_configure[22][3] ),
    .X(net2466));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1843 (.A(net924),
    .X(net2467));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1844 (.A(_0628_),
    .X(net2468));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1845 (.A(\gpio_configure[23][2] ),
    .X(net2469));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1846 (.A(net946),
    .X(net2470));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1847 (.A(_0635_),
    .X(net2471));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1848 (.A(\gpio_configure[11][10] ),
    .X(net2472));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1849 (.A(net1130),
    .X(net2473));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold185 (.A(net2108),
    .X(net809));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1850 (.A(_0224_),
    .X(net2474));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1851 (.A(net1131),
    .X(net2475));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1852 (.A(\gpio_configure[1][10] ),
    .X(net2476));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1853 (.A(net1080),
    .X(net2477));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1854 (.A(_0150_),
    .X(net2478));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1855 (.A(net1081),
    .X(net2479));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1856 (.A(\gpio_configure[16][3] ),
    .X(net2480));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1857 (.A(net966),
    .X(net2481));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1858 (.A(_0580_),
    .X(net2482));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1859 (.A(net967),
    .X(net2483));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold186 (.A(net2110),
    .X(net810));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1860 (.A(\gpio_configure[0][3] ),
    .X(net2484));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1861 (.A(net970),
    .X(net2485));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1862 (.A(_0452_),
    .X(net2486));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1863 (.A(net971),
    .X(net2487));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1864 (.A(\gpio_configure[30][3] ),
    .X(net2488));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1865 (.A(net974),
    .X(net2489));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1866 (.A(\gpio_configure[26][2] ),
    .X(net2490));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1867 (.A(net1050),
    .X(net2491));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1868 (.A(\gpio_configure[21][6] ),
    .X(net2492));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1869 (.A(net744),
    .X(net2493));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold187 (.A(\gpio_configure[26][5] ),
    .X(net811));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1870 (.A(_0623_),
    .X(net2494));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1871 (.A(\gpio_configure[20][6] ),
    .X(net2495));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1872 (.A(net746),
    .X(net2496));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1873 (.A(_0615_),
    .X(net2497));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1874 (.A(\gpio_configure[22][1] ),
    .X(net2498));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1875 (.A(net687),
    .X(net2499));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1876 (.A(_0626_),
    .X(net2500));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1877 (.A(\gpio_configure[18][2] ),
    .X(net2501));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1878 (.A(net1122),
    .X(net2502));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1879 (.A(_0595_),
    .X(net2503));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold188 (.A(net2073),
    .X(net812));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1880 (.A(\gpio_configure[21][10] ),
    .X(net2504));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1881 (.A(net1072),
    .X(net2505));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1882 (.A(_0364_),
    .X(net2506));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1883 (.A(\gpio_configure[21][2] ),
    .X(net2507));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1884 (.A(net934),
    .X(net2508));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1885 (.A(_0619_),
    .X(net2509));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1886 (.A(\gpio_configure[3][10] ),
    .X(net2510));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1887 (.A(net1136),
    .X(net2511));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1888 (.A(\mgmt_gpio_data_buf[11] ),
    .X(net2512));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1889 (.A(net1028),
    .X(net2513));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold189 (.A(net2075),
    .X(net813));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1890 (.A(_0138_),
    .X(net2514));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1891 (.A(\clk2_output_dest[1] ),
    .X(net2515));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1892 (.A(net972),
    .X(net2516));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1893 (.A(_0431_),
    .X(net2517));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1894 (.A(\gpio_configure[12][3] ),
    .X(net2518));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1895 (.A(net952),
    .X(net2519));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1896 (.A(_0548_),
    .X(net2520));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1897 (.A(net953),
    .X(net2521));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1898 (.A(\gpio_configure[5][2] ),
    .X(net2522));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1899 (.A(net1056),
    .X(net2523));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold19 (.A(net2206),
    .X(net643));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold190 (.A(net2077),
    .X(net814));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1900 (.A(_0491_),
    .X(net2524));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1901 (.A(\gpio_configure[9][3] ),
    .X(net2525));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1902 (.A(net916),
    .X(net2526));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1903 (.A(_0524_),
    .X(net2527));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1904 (.A(net917),
    .X(net2528));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1905 (.A(\gpio_configure[33][6] ),
    .X(net2529));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1906 (.A(net1997),
    .X(net2530));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1907 (.A(_0719_),
    .X(net2531));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1908 (.A(\gpio_configure[17][3] ),
    .X(net2532));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1909 (.A(net990),
    .X(net2533));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold191 (.A(net2062),
    .X(net815));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1910 (.A(_0588_),
    .X(net2534));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1911 (.A(net268),
    .X(net2535));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1912 (.A(net1144),
    .X(net2536));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1913 (.A(_0401_),
    .X(net2537));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1914 (.A(\gpio_configure[36][6] ),
    .X(net2538));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1915 (.A(net738),
    .X(net2539));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1916 (.A(_0743_),
    .X(net2540));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1917 (.A(\mgmt_gpio_data_buf[14] ),
    .X(net2541));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1918 (.A(net748),
    .X(net2542));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1919 (.A(_0141_),
    .X(net2543));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold192 (.A(net2064),
    .X(net816));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1920 (.A(net262),
    .X(net2544));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1921 (.A(net1169),
    .X(net2545));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1922 (.A(_0396_),
    .X(net2546));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1923 (.A(net270),
    .X(net2547));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1924 (.A(net1148),
    .X(net2548));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1925 (.A(_0103_),
    .X(net2549));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1926 (.A(\gpio_configure[24][3] ),
    .X(net2550));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1927 (.A(net2010),
    .X(net2551));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1928 (.A(_0644_),
    .X(net2552));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1929 (.A(net273),
    .X(net2553));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold193 (.A(net2046),
    .X(net817));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1930 (.A(net978),
    .X(net2554));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1931 (.A(_0106_),
    .X(net2555));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1932 (.A(\gpio_configure[21][11] ),
    .X(net2556));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1933 (.A(net1030),
    .X(net2557));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1934 (.A(_0365_),
    .X(net2558));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1935 (.A(net298),
    .X(net2559));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1936 (.A(net1014),
    .X(net2560));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1937 (.A(_0417_),
    .X(net2561));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1938 (.A(\gpio_configure[15][3] ),
    .X(net2562));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1939 (.A(net984),
    .X(net2563));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold194 (.A(net2048),
    .X(net818));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1940 (.A(_0572_),
    .X(net2564));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1941 (.A(\gpio_configure[28][11] ),
    .X(net2565));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1942 (.A(net1040),
    .X(net2566));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1943 (.A(\gpio_configure[21][3] ),
    .X(net2567));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1944 (.A(net1052),
    .X(net2568));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1945 (.A(_0620_),
    .X(net2569));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1946 (.A(\gpio_configure[25][11] ),
    .X(net2570));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1947 (.A(net1090),
    .X(net2571));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1948 (.A(_0068_),
    .X(net2572));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1949 (.A(\gpio_configure[14][11] ),
    .X(net2573));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold195 (.A(net2180),
    .X(net819));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1950 (.A(net1100),
    .X(net2574));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1951 (.A(_0295_),
    .X(net2575));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1952 (.A(net1101),
    .X(net2576));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1953 (.A(\gpio_configure[10][11] ),
    .X(net2577));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1954 (.A(net1070),
    .X(net2578));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1955 (.A(_0220_),
    .X(net2579));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1956 (.A(net1071),
    .X(net2580));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1957 (.A(\gpio_configure[18][11] ),
    .X(net2581));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1958 (.A(net1048),
    .X(net2582));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1959 (.A(_0335_),
    .X(net2583));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold196 (.A(net2182),
    .X(net820));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1960 (.A(\gpio_configure[10][2] ),
    .X(net2584));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1961 (.A(net1177),
    .X(net2585));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1962 (.A(_0531_),
    .X(net2586));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1963 (.A(net1178),
    .X(net2587));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1964 (.A(\gpio_configure[16][2] ),
    .X(net2588));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1965 (.A(net1142),
    .X(net2589));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1966 (.A(_0579_),
    .X(net2590));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1967 (.A(net1143),
    .X(net2591));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1968 (.A(\gpio_configure[11][11] ),
    .X(net2592));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1969 (.A(net1046),
    .X(net2593));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold197 (.A(\gpio_configure[1][2] ),
    .X(net821));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1970 (.A(_0225_),
    .X(net2594));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1971 (.A(net1047),
    .X(net2595));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1972 (.A(\gpio_configure[9][11] ),
    .X(net2596));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1973 (.A(net938),
    .X(net2597));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1974 (.A(\gpio_configure[6][11] ),
    .X(net2598));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1975 (.A(net1074),
    .X(net2599));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1976 (.A(\gpio_configure[0][10] ),
    .X(net2600));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1977 (.A(net1112),
    .X(net2601));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1978 (.A(_0145_),
    .X(net2602));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1979 (.A(\gpio_configure[15][11] ),
    .X(net2603));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold198 (.A(net2095),
    .X(net822));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1980 (.A(net1076),
    .X(net2604));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1981 (.A(_0305_),
    .X(net2605));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1982 (.A(net1077),
    .X(net2606));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1983 (.A(\gpio_configure[20][11] ),
    .X(net2607));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1984 (.A(net1058),
    .X(net2608));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1985 (.A(_0355_),
    .X(net2609));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1986 (.A(\gpio_configure[29][11] ),
    .X(net2610));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1987 (.A(net994),
    .X(net2611));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1988 (.A(\gpio_configure[7][10] ),
    .X(net2612));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1989 (.A(net1196),
    .X(net2613));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold199 (.A(net2161),
    .X(net823));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1990 (.A(\gpio_configure[17][2] ),
    .X(net2614));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1991 (.A(net1173),
    .X(net2615));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1992 (.A(_0587_),
    .X(net2616));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1993 (.A(\gpio_configure[17][11] ),
    .X(net2617));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1994 (.A(net1102),
    .X(net2618));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1995 (.A(_0325_),
    .X(net2619));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1996 (.A(net1103),
    .X(net2620));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1997 (.A(\gpio_configure[8][10] ),
    .X(net2621));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1998 (.A(net1128),
    .X(net2622));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold1999 (.A(\gpio_configure[19][3] ),
    .X(net2623));
 sky130_fd_sc_hd__buf_8 hold2 (.A(net2016),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 hold20 (.A(net2208),
    .X(net644));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold200 (.A(net2163),
    .X(net824));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2000 (.A(net1064),
    .X(net2624));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2001 (.A(_0604_),
    .X(net2625));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2002 (.A(\mgmt_gpio_data_buf[22] ),
    .X(net2626));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2003 (.A(net759),
    .X(net2627));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2004 (.A(_0280_),
    .X(net2628));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2005 (.A(\gpio_configure[32][2] ),
    .X(net2629));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2006 (.A(net1175),
    .X(net2630));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2007 (.A(net278),
    .X(net2631));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2008 (.A(net1198),
    .X(net2632));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2009 (.A(_0407_),
    .X(net2633));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold201 (.A(net2058),
    .X(net825));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2010 (.A(\gpio_configure[4][10] ),
    .X(net2634));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2011 (.A(net1220),
    .X(net2635));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2012 (.A(net287),
    .X(net2636));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2013 (.A(net1118),
    .X(net2637));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2014 (.A(_0111_),
    .X(net2638));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2015 (.A(\gpio_configure[18][3] ),
    .X(net2639));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2016 (.A(net1054),
    .X(net2640));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2017 (.A(_0596_),
    .X(net2641));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2018 (.A(\gpio_configure[12][11] ),
    .X(net2642));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2019 (.A(net1062),
    .X(net2643));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold202 (.A(net2060),
    .X(net826));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2020 (.A(_0230_),
    .X(net2644));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2021 (.A(\gpio_configure[8][2] ),
    .X(net2645));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2022 (.A(net1183),
    .X(net2646));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2023 (.A(\gpio_configure[36][11] ),
    .X(net2647));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2024 (.A(net1134),
    .X(net2648));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2025 (.A(_0300_),
    .X(net2649));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2026 (.A(\gpio_configure[16][10] ),
    .X(net2650));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2027 (.A(net1232),
    .X(net2651));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2028 (.A(_0314_),
    .X(net2652));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2029 (.A(net1233),
    .X(net2653));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold203 (.A(net2146),
    .X(net827));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2030 (.A(\gpio_configure[22][11] ),
    .X(net2654));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2031 (.A(net1066),
    .X(net2655));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2032 (.A(_0370_),
    .X(net2656));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2033 (.A(\gpio_configure[37][11] ),
    .X(net2657));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2034 (.A(net1110),
    .X(net2658));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2035 (.A(_0290_),
    .X(net2659));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2036 (.A(\wbbd_data[0] ),
    .X(net2660));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2037 (.A(net1086),
    .X(net2661));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2038 (.A(_1461_),
    .X(net2662));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2039 (.A(net1087),
    .X(net2663));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold204 (.A(net2148),
    .X(net828));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2040 (.A(net500),
    .X(net2664));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2041 (.A(_0561_),
    .X(net2665));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2042 (.A(serial_bb_resetn),
    .X(net2666));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2043 (.A(net1202),
    .X(net2667));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2044 (.A(_0422_),
    .X(net2668));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2045 (.A(\gpio_configure[13][11] ),
    .X(net2669));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2046 (.A(net1106),
    .X(net2670));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2047 (.A(_0285_),
    .X(net2671));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2048 (.A(\gpio_configure[35][11] ),
    .X(net2672));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2049 (.A(net1114),
    .X(net2673));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold205 (.A(net2176),
    .X(net829));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2050 (.A(_0310_),
    .X(net2674));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2051 (.A(\gpio_configure[26][11] ),
    .X(net2675));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2052 (.A(net1008),
    .X(net2676));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2053 (.A(\gpio_configure[5][3] ),
    .X(net2677));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2054 (.A(net1189),
    .X(net2678));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2055 (.A(_0492_),
    .X(net2679));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2056 (.A(\gpio_configure[34][11] ),
    .X(net2680));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2057 (.A(net1132),
    .X(net2681));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2058 (.A(_0320_),
    .X(net2682));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2059 (.A(\gpio_configure[21][0] ),
    .X(net2683));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold206 (.A(net2178),
    .X(net830));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2060 (.A(net1246),
    .X(net2684));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2061 (.A(_0617_),
    .X(net2685));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2062 (.A(\mgmt_gpio_data[2] ),
    .X(net2686));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2063 (.A(net1306),
    .X(net2687));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2064 (.A(_0129_),
    .X(net2688));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2065 (.A(\gpio_configure[31][1] ),
    .X(net2689));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2066 (.A(net1166),
    .X(net2690));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2067 (.A(_0698_),
    .X(net2691));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2068 (.A(\hkspi.odata[4] ),
    .X(net2692));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2069 (.A(net706),
    .X(net2693));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold207 (.A(net2169),
    .X(net831));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2070 (.A(_1465_),
    .X(net2694));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2071 (.A(net791),
    .X(net2695));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2072 (.A(net707),
    .X(net2696));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2073 (.A(_0661_),
    .X(net2697));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2074 (.A(net721),
    .X(net2698));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2075 (.A(\gpio_configure[31][4] ),
    .X(net2699));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2076 (.A(net734),
    .X(net2700));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2077 (.A(_0701_),
    .X(net2701));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2078 (.A(\clk1_output_dest[1] ),
    .X(net2702));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2079 (.A(net732),
    .X(net2703));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold208 (.A(net2171),
    .X(net832));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2080 (.A(_0429_),
    .X(net2704));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2081 (.A(\mgmt_gpio_data[18] ),
    .X(net2705));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2082 (.A(net1338),
    .X(net2706));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2083 (.A(_0259_),
    .X(net2707));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2084 (.A(\mgmt_gpio_data[28] ),
    .X(net2708));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2085 (.A(net718),
    .X(net2709));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2086 (.A(_0270_),
    .X(net2710));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2087 (.A(net284),
    .X(net2711));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2088 (.A(net1247),
    .X(net2712));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2089 (.A(_0412_),
    .X(net2713));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold209 (.A(net2136),
    .X(net833));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2090 (.A(net292),
    .X(net2714));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2091 (.A(net1252),
    .X(net2715));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2092 (.A(_0116_),
    .X(net2716));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2093 (.A(\mgmt_gpio_data[19] ),
    .X(net2717));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2094 (.A(net1399),
    .X(net2718));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2095 (.A(_0260_),
    .X(net2719));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2096 (.A(\gpio_configure[25][12] ),
    .X(net2720));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2097 (.A(net767),
    .X(net2721));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2098 (.A(_0069_),
    .X(net2722));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2099 (.A(net275),
    .X(net2723));
 sky130_fd_sc_hd__buf_4 hold21 (.A(_0857_),
    .X(net645));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold210 (.A(net2138),
    .X(net834));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2100 (.A(net1279),
    .X(net2724));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2101 (.A(_0108_),
    .X(net2725));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2102 (.A(\gpio_configure[20][4] ),
    .X(net2726));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2103 (.A(net771),
    .X(net2727));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2104 (.A(_0613_),
    .X(net2728));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2105 (.A(\gpio_configure[17][12] ),
    .X(net2729));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2106 (.A(net782),
    .X(net2730));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2107 (.A(_0326_),
    .X(net2731));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2108 (.A(net783),
    .X(net2732));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2109 (.A(\gpio_configure[9][4] ),
    .X(net2733));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold211 (.A(net2153),
    .X(net835));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2110 (.A(net763),
    .X(net2734));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2111 (.A(_0525_),
    .X(net2735));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2112 (.A(net764),
    .X(net2736));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2113 (.A(\gpio_configure[25][0] ),
    .X(net2737));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2114 (.A(net1098),
    .X(net2738));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2115 (.A(\mgmt_gpio_data[10] ),
    .X(net2739));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2116 (.A(net1423),
    .X(net2740));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2117 (.A(_0121_),
    .X(net2741));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2118 (.A(\mgmt_gpio_data_buf[16] ),
    .X(net2742));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2119 (.A(net1993),
    .X(net2743));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold212 (.A(net2155),
    .X(net836));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2120 (.A(_0274_),
    .X(net2744));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2121 (.A(trap_output_dest),
    .X(net2745));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2122 (.A(net1092),
    .X(net2746));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2123 (.A(_0432_),
    .X(net2747));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2124 (.A(\gpio_configure[28][4] ),
    .X(net2748));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2125 (.A(net786),
    .X(net2749));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2126 (.A(\gpio_configure[14][12] ),
    .X(net2750));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2127 (.A(net773),
    .X(net2751));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2128 (.A(_0296_),
    .X(net2752));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2129 (.A(net774),
    .X(net2753));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold213 (.A(\gpio_configure[25][2] ),
    .X(net837));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2130 (.A(\mgmt_gpio_data[21] ),
    .X(net2754));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2131 (.A(net1449),
    .X(net2755));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2132 (.A(_0262_),
    .X(net2756));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2133 (.A(\mgmt_gpio_data_buf[8] ),
    .X(net2757));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2134 (.A(net1162),
    .X(net2758));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2135 (.A(_0135_),
    .X(net2759));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2136 (.A(\gpio_configure[37][12] ),
    .X(net2760));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2137 (.A(net2009),
    .X(net2761));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2138 (.A(_0291_),
    .X(net2762));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2139 (.A(\gpio_configure[35][4] ),
    .X(net2763));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold214 (.A(net2117),
    .X(net838));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2140 (.A(net769),
    .X(net2764));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2141 (.A(_0733_),
    .X(net2765));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2142 (.A(\gpio_configure[14][4] ),
    .X(net2766));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2143 (.A(net788),
    .X(net2767));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2144 (.A(_0565_),
    .X(net2768));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2145 (.A(net789),
    .X(net2769));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2146 (.A(\gpio_configure[36][12] ),
    .X(net2770));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2147 (.A(net2012),
    .X(net2771));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2148 (.A(_0301_),
    .X(net2772));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2149 (.A(\gpio_configure[21][4] ),
    .X(net2773));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold215 (.A(net2187),
    .X(net839));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2150 (.A(net765),
    .X(net2774));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2151 (.A(_0621_),
    .X(net2775));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2152 (.A(\mgmt_gpio_data[3] ),
    .X(net2776));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2153 (.A(net1441),
    .X(net2777));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2154 (.A(_0130_),
    .X(net2778));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2155 (.A(\gpio_configure[12][12] ),
    .X(net2779));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2156 (.A(net784),
    .X(net2780));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2157 (.A(_0231_),
    .X(net2781));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2158 (.A(\mgmt_gpio_data_buf[20] ),
    .X(net2782));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2159 (.A(net793),
    .X(net2783));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold216 (.A(net2189),
    .X(net840));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2160 (.A(_0278_),
    .X(net2784));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2161 (.A(\mgmt_gpio_data[14] ),
    .X(net2785));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2162 (.A(net1034),
    .X(net2786));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2163 (.A(_0125_),
    .X(net2787));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2164 (.A(\mgmt_gpio_data[11] ),
    .X(net2788));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2165 (.A(net1492),
    .X(net2789));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2166 (.A(_0122_),
    .X(net2790));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2167 (.A(net291),
    .X(net2791));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2168 (.A(net1471),
    .X(net2792));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2169 (.A(_0115_),
    .X(net2793));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold217 (.A(net2143),
    .X(net841));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2170 (.A(\gpio_configure[10][7] ),
    .X(net2794));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2171 (.A(net1018),
    .X(net2795));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2172 (.A(_0536_),
    .X(net2796));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2173 (.A(net1019),
    .X(net2797));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2174 (.A(\gpio_configure[4][7] ),
    .X(net2798));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2175 (.A(net1108),
    .X(net2799));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2176 (.A(\gpio_configure[6][7] ),
    .X(net2800));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2177 (.A(net1012),
    .X(net2801));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2178 (.A(\mgmt_gpio_data[34] ),
    .X(net2802));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2179 (.A(net1509),
    .X(net2803));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold218 (.A(net2145),
    .X(net842));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2180 (.A(\gpio_configure[1][5] ),
    .X(net2804));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2181 (.A(net1513),
    .X(net2805));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2182 (.A(\mgmt_gpio_data_buf[7] ),
    .X(net2806));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2183 (.A(net1060),
    .X(net2807));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2184 (.A(_0448_),
    .X(net2808));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2185 (.A(\gpio_configure[1][7] ),
    .X(net2809));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2186 (.A(net1016),
    .X(net2810));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2187 (.A(\mgmt_gpio_data[22] ),
    .X(net2811));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2188 (.A(net1104),
    .X(net2812));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2189 (.A(_0263_),
    .X(net2813));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold219 (.A(net2190),
    .X(net843));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2190 (.A(\gpio_configure[11][7] ),
    .X(net2814));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2191 (.A(net1120),
    .X(net2815));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2192 (.A(_0544_),
    .X(net2816));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2193 (.A(\gpio_configure[30][0] ),
    .X(net2817));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2194 (.A(net1238),
    .X(net2818));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2195 (.A(\gpio_configure[29][7] ),
    .X(net2819));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2196 (.A(net1068),
    .X(net2820));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2197 (.A(_0688_),
    .X(net2821));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2198 (.A(\gpio_configure[8][7] ),
    .X(net2822));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2199 (.A(net1084),
    .X(net2823));
 sky130_fd_sc_hd__clkbuf_2 hold22 (.A(net418),
    .X(net646));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold220 (.A(net2192),
    .X(net844));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2200 (.A(\gpio_configure[26][7] ),
    .X(net2824));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2201 (.A(net1116),
    .X(net2825));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2202 (.A(\gpio_configure[2][7] ),
    .X(net2826));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2203 (.A(net1082),
    .X(net2827));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2204 (.A(_0472_),
    .X(net2828));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2205 (.A(net274),
    .X(net2829));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2206 (.A(net1502),
    .X(net2830));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2207 (.A(_0107_),
    .X(net2831));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2208 (.A(\gpio_configure[3][7] ),
    .X(net2832));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2209 (.A(net1138),
    .X(net2833));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold221 (.A(net2050),
    .X(net845));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2210 (.A(_0480_),
    .X(net2834));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2211 (.A(\gpio_configure[23][7] ),
    .X(net2835));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2212 (.A(net1167),
    .X(net2836));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2213 (.A(_0640_),
    .X(net2837));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2214 (.A(\gpio_configure[6][5] ),
    .X(net2838));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2215 (.A(net1515),
    .X(net2839));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2216 (.A(\gpio_configure[28][0] ),
    .X(net2840));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2217 (.A(net1267),
    .X(net2841));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2218 (.A(\gpio_configure[0][7] ),
    .X(net2842));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2219 (.A(net1146),
    .X(net2843));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold222 (.A(net2052),
    .X(net846));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2220 (.A(_0456_),
    .X(net2844));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2221 (.A(net1147),
    .X(net2845));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2222 (.A(\hkspi.addr[7] ),
    .X(net2846));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2223 (.A(_0834_),
    .X(net2847));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2224 (.A(_0837_),
    .X(net2848));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2225 (.A(_0842_),
    .X(net2849));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2226 (.A(_0562_),
    .X(net2850));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2227 (.A(net1155),
    .X(net2851));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2228 (.A(\gpio_configure[5][7] ),
    .X(net2852));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2229 (.A(net1194),
    .X(net2853));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold223 (.A(net2183),
    .X(net847));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2230 (.A(_0496_),
    .X(net2854));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2231 (.A(\gpio_configure[22][7] ),
    .X(net2855));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2232 (.A(net1126),
    .X(net2856));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2233 (.A(_0632_),
    .X(net2857));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2234 (.A(\gpio_configure[32][1] ),
    .X(net2858));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2235 (.A(net1164),
    .X(net2859));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2236 (.A(\gpio_configure[15][7] ),
    .X(net2860));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2237 (.A(net1078),
    .X(net2861));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2238 (.A(_0576_),
    .X(net2862));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2239 (.A(\gpio_configure[8][1] ),
    .X(net2863));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold224 (.A(net2185),
    .X(net848));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2240 (.A(net1185),
    .X(net2864));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2241 (.A(\gpio_configure[27][7] ),
    .X(net2865));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2242 (.A(net1150),
    .X(net2866));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2243 (.A(_0672_),
    .X(net2867));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2244 (.A(\gpio_configure[2][1] ),
    .X(net2868));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2245 (.A(net1160),
    .X(net2869));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2246 (.A(_0466_),
    .X(net2870));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2247 (.A(\gpio_configure[14][7] ),
    .X(net2871));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2248 (.A(net1234),
    .X(net2872));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2249 (.A(net296),
    .X(net2873));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold225 (.A(net2127),
    .X(net849));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2250 (.A(net1096),
    .X(net2874));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2251 (.A(\gpio_configure[15][5] ),
    .X(net2875));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2252 (.A(net1527),
    .X(net2876));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2253 (.A(_0574_),
    .X(net2877));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2254 (.A(\gpio_configure[4][1] ),
    .X(net2878));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2255 (.A(net1228),
    .X(net2879));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2256 (.A(\gpio_configure[6][1] ),
    .X(net2880));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2257 (.A(net1156),
    .X(net2881));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2258 (.A(\gpio_configure[32][7] ),
    .X(net2882));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2259 (.A(net1158),
    .X(net2883));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold226 (.A(net2129),
    .X(net850));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2260 (.A(\gpio_configure[9][7] ),
    .X(net2884));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2261 (.A(net1214),
    .X(net2885));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2262 (.A(\gpio_configure[7][7] ),
    .X(net2886));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2263 (.A(net1222),
    .X(net2887));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2264 (.A(_0512_),
    .X(net2888));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2265 (.A(net1223),
    .X(net2889));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2266 (.A(\gpio_configure[25][7] ),
    .X(net2890));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2267 (.A(net1179),
    .X(net2891));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2268 (.A(\gpio_configure[32][4] ),
    .X(net2892));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2269 (.A(net716),
    .X(net2893));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold227 (.A(net2204),
    .X(net851));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2270 (.A(\gpio_configure[24][1] ),
    .X(net2894));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2271 (.A(net1192),
    .X(net2895));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2272 (.A(_0642_),
    .X(net2896));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2273 (.A(\gpio_configure[13][7] ),
    .X(net2897));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2274 (.A(net1206),
    .X(net2898));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2275 (.A(_0560_),
    .X(net2899));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2276 (.A(\gpio_configure[36][7] ),
    .X(net2900));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2277 (.A(net1140),
    .X(net2901));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2278 (.A(\gpio_configure[21][7] ),
    .X(net2902));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2279 (.A(net1181),
    .X(net2903));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold228 (.A(_0654_),
    .X(net852));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2280 (.A(_0624_),
    .X(net2904));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2281 (.A(\gpio_configure[1][4] ),
    .X(net2905));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2282 (.A(net2005),
    .X(net2906));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2283 (.A(\gpio_configure[18][7] ),
    .X(net2907));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2284 (.A(net1204),
    .X(net2908));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2285 (.A(_0600_),
    .X(net2909));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2286 (.A(\gpio_configure[8][4] ),
    .X(net2910));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2287 (.A(net710),
    .X(net2911));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2288 (.A(\gpio_configure[17][7] ),
    .X(net2912));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2289 (.A(net1224),
    .X(net2913));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold229 (.A(net2165),
    .X(net853));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2290 (.A(_0592_),
    .X(net2914));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2291 (.A(\gpio_configure[16][7] ),
    .X(net2915));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2292 (.A(net1226),
    .X(net2916));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2293 (.A(\mgmt_gpio_data_buf[1] ),
    .X(net2917));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2294 (.A(net1124),
    .X(net2918));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2295 (.A(_0442_),
    .X(net2919));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2296 (.A(\gpio_configure[16][5] ),
    .X(net2920));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2297 (.A(net1533),
    .X(net2921));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2298 (.A(\gpio_configure[5][5] ),
    .X(net2922));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2299 (.A(net1525),
    .X(net2923));
 sky130_fd_sc_hd__buf_4 hold23 (.A(_2625_),
    .X(net647));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold230 (.A(net2167),
    .X(net854));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2300 (.A(_0494_),
    .X(net2924));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2301 (.A(\gpio_configure[28][7] ),
    .X(net2925));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2302 (.A(net1187),
    .X(net2926));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2303 (.A(\gpio_configure[0][5] ),
    .X(net2927));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2304 (.A(net1547),
    .X(net2928));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2305 (.A(_0454_),
    .X(net2929));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2306 (.A(\gpio_configure[33][7] ),
    .X(net2930));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2307 (.A(net1208),
    .X(net2931));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2308 (.A(_0720_),
    .X(net2932));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2309 (.A(\mgmt_gpio_data[31] ),
    .X(net2933));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold231 (.A(net2243),
    .X(net855));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2310 (.A(net1171),
    .X(net2934));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2311 (.A(wbbd_busy),
    .X(net2935));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2312 (.A(net524),
    .X(net2936));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2313 (.A(_0851_),
    .X(net2937));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2314 (.A(_0506_),
    .X(net2938));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2315 (.A(net1211),
    .X(net2939));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2316 (.A(\gpio_configure[27][4] ),
    .X(net2940));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2317 (.A(net726),
    .X(net2941));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2318 (.A(\mgmt_gpio_data_buf[15] ),
    .X(net2942));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2319 (.A(net1236),
    .X(net2943));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold232 (.A(_0652_),
    .X(net856));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2320 (.A(_0142_),
    .X(net2944));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2321 (.A(\gpio_configure[5][1] ),
    .X(net2945));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2322 (.A(net1200),
    .X(net2946));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2323 (.A(\gpio_configure[2][10] ),
    .X(net2947));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2324 (.A(net1519),
    .X(net2948));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2325 (.A(\gpio_configure[5][11] ),
    .X(net2949));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2326 (.A(net1555),
    .X(net2950));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2327 (.A(\gpio_configure[3][1] ),
    .X(net2951));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2328 (.A(net1212),
    .X(net2952));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2329 (.A(\gpio_configure[13][5] ),
    .X(net2953));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold233 (.A(net2301),
    .X(net857));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2330 (.A(net1589),
    .X(net2954));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2331 (.A(\gpio_configure[5][4] ),
    .X(net2955));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2332 (.A(net722),
    .X(net2956));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2333 (.A(\gpio_configure[3][4] ),
    .X(net2957));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2334 (.A(net712),
    .X(net2958));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2335 (.A(\gpio_configure[24][11] ),
    .X(net2959));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2336 (.A(net1537),
    .X(net2960));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2337 (.A(_0250_),
    .X(net2961));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2338 (.A(\gpio_configure[0][1] ),
    .X(net2962));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2339 (.A(net1216),
    .X(net2963));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold234 (.A(net2303),
    .X(net858));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2340 (.A(_0450_),
    .X(net2964));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2341 (.A(\gpio_configure[17][5] ),
    .X(net2965));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2342 (.A(net1603),
    .X(net2966));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2343 (.A(_0590_),
    .X(net2967));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2344 (.A(\gpio_configure[2][5] ),
    .X(net2968));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2345 (.A(net1523),
    .X(net2969));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2346 (.A(\gpio_configure[31][11] ),
    .X(net2970));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2347 (.A(net1549),
    .X(net2971));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2348 (.A(\gpio_configure[33][11] ),
    .X(net2972));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2349 (.A(net1551),
    .X(net2973));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold235 (.A(net2226),
    .X(net859));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2350 (.A(\gpio_configure[0][4] ),
    .X(net2974));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2351 (.A(net724),
    .X(net2975));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2352 (.A(_0453_),
    .X(net2976));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2353 (.A(\gpio_configure[28][2] ),
    .X(net2977));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2354 (.A(net1559),
    .X(net2978));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2355 (.A(\gpio_configure[10][5] ),
    .X(net2979));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2356 (.A(net1521),
    .X(net2980));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2357 (.A(\gpio_configure[11][9] ),
    .X(net2981));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2358 (.A(net1253),
    .X(net2982));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2359 (.A(\gpio_configure[7][4] ),
    .X(net2983));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold236 (.A(net2228),
    .X(net860));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2360 (.A(net730),
    .X(net2984));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2361 (.A(_0509_),
    .X(net2985));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2362 (.A(\gpio_configure[32][11] ),
    .X(net2986));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2363 (.A(net1541),
    .X(net2987));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2364 (.A(\gpio_configure[22][10] ),
    .X(net2988));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2365 (.A(net1571),
    .X(net2989));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2366 (.A(_0369_),
    .X(net2990));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2367 (.A(\gpio_configure[9][10] ),
    .X(net2991));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2368 (.A(net1585),
    .X(net2992));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2369 (.A(\gpio_configure[32][5] ),
    .X(net2993));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold237 (.A(net2363),
    .X(net861));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2370 (.A(net1553),
    .X(net2994));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2371 (.A(\gpio_configure[22][9] ),
    .X(net2995));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2372 (.A(net1248),
    .X(net2996));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2373 (.A(_0368_),
    .X(net2997));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2374 (.A(\gpio_configure[10][10] ),
    .X(net2998));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2375 (.A(net1531),
    .X(net2999));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2376 (.A(\gpio_configure[36][10] ),
    .X(net3000));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2377 (.A(net1577),
    .X(net3001));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2378 (.A(\gpio_configure[24][7] ),
    .X(net3002));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2379 (.A(net1230),
    .X(net3003));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold238 (.A(net2365),
    .X(net862));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2380 (.A(_0648_),
    .X(net3004));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2381 (.A(\gpio_configure[12][5] ),
    .X(net3005));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2382 (.A(net1619),
    .X(net3006));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2383 (.A(\gpio_configure[3][5] ),
    .X(net3007));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2384 (.A(net1545),
    .X(net3008));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2385 (.A(\gpio_configure[12][9] ),
    .X(net3009));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2386 (.A(net1240),
    .X(net3010));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2387 (.A(\gpio_configure[30][11] ),
    .X(net3011));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2388 (.A(net1543),
    .X(net3012));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2389 (.A(\gpio_configure[4][11] ),
    .X(net3013));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold239 (.A(net2213),
    .X(net863));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2390 (.A(net1569),
    .X(net3014));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2391 (.A(\gpio_configure[7][11] ),
    .X(net3015));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2392 (.A(net1539),
    .X(net3016));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2393 (.A(\gpio_configure[19][10] ),
    .X(net3017));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2394 (.A(net1535),
    .X(net3018));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2395 (.A(_0344_),
    .X(net3019));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2396 (.A(\gpio_configure[14][5] ),
    .X(net3020));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2397 (.A(net1609),
    .X(net3021));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2398 (.A(\mgmt_gpio_data_buf[23] ),
    .X(net3022));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2399 (.A(net1257),
    .X(net3023));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold24 (.A(net2121),
    .X(net648));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold240 (.A(net2215),
    .X(net864));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2400 (.A(_0281_),
    .X(net3024));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2401 (.A(\gpio_configure[16][4] ),
    .X(net3025));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2402 (.A(net728),
    .X(net3026));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2403 (.A(\gpio_configure[1][11] ),
    .X(net3027));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2404 (.A(net1623),
    .X(net3028));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2405 (.A(_0151_),
    .X(net3029));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2406 (.A(\gpio_configure[20][2] ),
    .X(net3030));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2407 (.A(net1567),
    .X(net3031));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2408 (.A(_0611_),
    .X(net3032));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2409 (.A(\gpio_configure[34][1] ),
    .X(net3033));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold241 (.A(net2194),
    .X(net865));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2410 (.A(net1242),
    .X(net3034));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2411 (.A(_0722_),
    .X(net3035));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2412 (.A(\gpio_configure[14][10] ),
    .X(net3036));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2413 (.A(net1599),
    .X(net3037));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2414 (.A(\gpio_configure[34][10] ),
    .X(net3038));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2415 (.A(net1581),
    .X(net3039));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2416 (.A(\gpio_configure[35][10] ),
    .X(net3040));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2417 (.A(net1617),
    .X(net3041));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2418 (.A(\gpio_configure[16][11] ),
    .X(net3042));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2419 (.A(net1625),
    .X(net3043));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold242 (.A(net2196),
    .X(net866));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2420 (.A(\gpio_configure[37][10] ),
    .X(net3044));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2421 (.A(net1565),
    .X(net3045));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2422 (.A(\gpio_configure[8][5] ),
    .X(net3046));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2423 (.A(net1627),
    .X(net3047));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2424 (.A(\gpio_configure[1][6] ),
    .X(net3048));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2425 (.A(net1342),
    .X(net3049));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2426 (.A(\mgmt_gpio_data[33] ),
    .X(net3050));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2427 (.A(net1308),
    .X(net3051));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2428 (.A(\gpio_configure[20][10] ),
    .X(net3052));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2429 (.A(net1561),
    .X(net3053));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold243 (.A(net2245),
    .X(net867));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2430 (.A(_0354_),
    .X(net3054));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2431 (.A(\gpio_configure[8][11] ),
    .X(net3055));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2432 (.A(net1575),
    .X(net3056));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2433 (.A(net255),
    .X(net3057));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2434 (.A(net1563),
    .X(net3058));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2435 (.A(_0402_),
    .X(net3059));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2436 (.A(\gpio_configure[17][10] ),
    .X(net3060));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2437 (.A(net1611),
    .X(net3061));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2438 (.A(net277),
    .X(net3062));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2439 (.A(net1269),
    .X(net3063));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold244 (.A(net2247),
    .X(net868));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2440 (.A(_0406_),
    .X(net3064));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2441 (.A(\gpio_configure[4][5] ),
    .X(net3065));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2442 (.A(net1621),
    .X(net3066));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2443 (.A(\gpio_configure[10][6] ),
    .X(net3067));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2444 (.A(net1356),
    .X(net3068));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2445 (.A(_0535_),
    .X(net3069));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2446 (.A(\gpio_configure[14][2] ),
    .X(net3070));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2447 (.A(net1557),
    .X(net3071));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2448 (.A(\gpio_configure[36][9] ),
    .X(net3072));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2449 (.A(net1277),
    .X(net3073));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold245 (.A(net2290),
    .X(net869));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2450 (.A(\gpio_configure[4][4] ),
    .X(net3074));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2451 (.A(net761),
    .X(net3075));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2452 (.A(serial_bb_enable),
    .X(net3076));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2453 (.A(net1273),
    .X(net3077));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2454 (.A(_0425_),
    .X(net3078));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2455 (.A(\gpio_configure[11][5] ),
    .X(net3079));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2456 (.A(net1601),
    .X(net3080));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2457 (.A(\gpio_configure[3][11] ),
    .X(net3081));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2458 (.A(net1597),
    .X(net3082));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2459 (.A(net286),
    .X(net3083));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold246 (.A(net2292),
    .X(net870));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2460 (.A(net1280),
    .X(net3084));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2461 (.A(_0118_),
    .X(net3085));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2462 (.A(\gpio_configure[12][10] ),
    .X(net3086));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2463 (.A(net1605),
    .X(net3087));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2464 (.A(serial_bb_load),
    .X(net3088));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2465 (.A(net1639),
    .X(net3089));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2466 (.A(_0421_),
    .X(net3090));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2467 (.A(\gpio_configure[3][9] ),
    .X(net3091));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2468 (.A(net1286),
    .X(net3092));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2469 (.A(\gpio_configure[1][1] ),
    .X(net3093));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold247 (.A(net2251),
    .X(net871));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2470 (.A(net1255),
    .X(net3094));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2471 (.A(net280),
    .X(net3095));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2472 (.A(net1288),
    .X(net3096));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2473 (.A(\gpio_configure[13][10] ),
    .X(net3097));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2474 (.A(net1607),
    .X(net3098));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2475 (.A(\gpio_configure[29][10] ),
    .X(net3099));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2476 (.A(net1529),
    .X(net3100));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2477 (.A(net279),
    .X(net3101));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2478 (.A(net1629),
    .X(net3102));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2479 (.A(\gpio_configure[0][9] ),
    .X(net3103));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold248 (.A(net2253),
    .X(net872));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2480 (.A(net1282),
    .X(net3104));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2481 (.A(_0144_),
    .X(net3105));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2482 (.A(net261),
    .X(net3106));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2483 (.A(net1302),
    .X(net3107));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2484 (.A(_0395_),
    .X(net3108));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2485 (.A(\mgmt_gpio_data[35] ),
    .X(net3109));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2486 (.A(net1573),
    .X(net3110));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2487 (.A(\gpio_configure[35][9] ),
    .X(net3111));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2488 (.A(net1259),
    .X(net3112));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2489 (.A(\gpio_configure[25][10] ),
    .X(net3113));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold249 (.A(net2248),
    .X(net873));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2490 (.A(net1587),
    .X(net3114));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2491 (.A(_0067_),
    .X(net3115));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2492 (.A(\gpio_configure[5][9] ),
    .X(net3116));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2493 (.A(net1320),
    .X(net3117));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2494 (.A(net259),
    .X(net3118));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2495 (.A(net1300),
    .X(net3119));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2496 (.A(_0393_),
    .X(net3120));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2497 (.A(\gpio_configure[34][9] ),
    .X(net3121));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2498 (.A(net1294),
    .X(net3122));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2499 (.A(\gpio_configure[0][11] ),
    .X(net3123));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold25 (.A(net2133),
    .X(net649));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold250 (.A(net2250),
    .X(net874));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2500 (.A(net1595),
    .X(net3124));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2501 (.A(_0146_),
    .X(net3125));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2502 (.A(net271),
    .X(net3126));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2503 (.A(net1583),
    .X(net3127));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2504 (.A(\gpio_configure[15][1] ),
    .X(net3128));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2505 (.A(net1348),
    .X(net3129));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2506 (.A(\gpio_configure[17][9] ),
    .X(net3130));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2507 (.A(net1265),
    .X(net3131));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2508 (.A(net263),
    .X(net3132));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2509 (.A(net1579),
    .X(net3133));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold251 (.A(net2304),
    .X(net875));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2510 (.A(_0397_),
    .X(net3134));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2511 (.A(\gpio_configure[4][9] ),
    .X(net3135));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2512 (.A(net1292),
    .X(net3136));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2513 (.A(\gpio_configure[16][1] ),
    .X(net3137));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2514 (.A(net1296),
    .X(net3138));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2515 (.A(\gpio_configure[8][6] ),
    .X(net3139));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2516 (.A(net1407),
    .X(net3140));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2517 (.A(\gpio_configure[2][4] ),
    .X(net3141));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2518 (.A(net752),
    .X(net3142));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2519 (.A(\gpio_configure[16][9] ),
    .X(net3143));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold252 (.A(net2306),
    .X(net876));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2520 (.A(net1318),
    .X(net3144));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2521 (.A(\gpio_configure[10][1] ),
    .X(net3145));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2522 (.A(net1310),
    .X(net3146));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2523 (.A(\gpio_configure[8][9] ),
    .X(net3147));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2524 (.A(net1290),
    .X(net3148));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2525 (.A(\gpio_configure[17][6] ),
    .X(net3149));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2526 (.A(net1433),
    .X(net3150));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2527 (.A(_0591_),
    .X(net3151));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2528 (.A(\gpio_configure[31][12] ),
    .X(net3152));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2529 (.A(net750),
    .X(net3153));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold253 (.A(net2261),
    .X(net877));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2530 (.A(net267),
    .X(net3154));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2531 (.A(net1298),
    .X(net3155));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2532 (.A(_0400_),
    .X(net3156));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2533 (.A(\gpio_configure[33][9] ),
    .X(net3157));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2534 (.A(net1314),
    .X(net3158));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2535 (.A(\gpio_configure[26][6] ),
    .X(net3159));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2536 (.A(net1425),
    .X(net3160));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2537 (.A(\gpio_configure[15][10] ),
    .X(net3161));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2538 (.A(net1615),
    .X(net3162));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2539 (.A(\gpio_configure[31][9] ),
    .X(net3163));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold254 (.A(net2263),
    .X(net878));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2540 (.A(net1328),
    .X(net3164));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2541 (.A(\gpio_configure[15][6] ),
    .X(net3165));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2542 (.A(net1419),
    .X(net3166));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2543 (.A(net294),
    .X(net3167));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2544 (.A(net1284),
    .X(net3168));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2545 (.A(\mgmt_gpio_data_buf[6] ),
    .X(net3169));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2546 (.A(net1379),
    .X(net3170));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2547 (.A(_0447_),
    .X(net3171));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2548 (.A(\mgmt_gpio_data_buf[4] ),
    .X(net3172));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2549 (.A(net775),
    .X(net3173));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold255 (.A(net2237),
    .X(net879));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2550 (.A(_0445_),
    .X(net3174));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2551 (.A(\gpio_configure[37][6] ),
    .X(net3175));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2552 (.A(net1451),
    .X(net3176));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2553 (.A(\gpio_configure[3][6] ),
    .X(net3177));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2554 (.A(net1415),
    .X(net3178));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2555 (.A(\gpio_configure[27][6] ),
    .X(net3179));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2556 (.A(net1401),
    .X(net3180));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2557 (.A(\gpio_configure[22][6] ),
    .X(net3181));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2558 (.A(net1413),
    .X(net3182));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2559 (.A(\gpio_configure[9][5] ),
    .X(net3183));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold256 (.A(net2239),
    .X(net880));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2560 (.A(net1671),
    .X(net3184));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2561 (.A(irq_2_inputsrc),
    .X(net3185));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2562 (.A(net1326),
    .X(net3186));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2563 (.A(_0434_),
    .X(net3187));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2564 (.A(\gpio_configure[6][6] ),
    .X(net3188));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2565 (.A(net1445),
    .X(net3189));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2566 (.A(\gpio_configure[13][6] ),
    .X(net3190));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2567 (.A(net1417),
    .X(net3191));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2568 (.A(\gpio_configure[32][6] ),
    .X(net3192));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2569 (.A(net1455),
    .X(net3193));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold257 (.A(net2267),
    .X(net881));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2570 (.A(\gpio_configure[24][5] ),
    .X(net3194));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2571 (.A(net1681),
    .X(net3195));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2572 (.A(_0646_),
    .X(net3196));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2573 (.A(\gpio_configure[0][6] ),
    .X(net3197));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2574 (.A(net1463),
    .X(net3198));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2575 (.A(_0455_),
    .X(net3199));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2576 (.A(\gpio_configure[34][6] ),
    .X(net3200));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2577 (.A(net1427),
    .X(net3201));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2578 (.A(_0727_),
    .X(net3202));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2579 (.A(\gpio_configure[19][6] ),
    .X(net3203));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold258 (.A(net2269),
    .X(net882));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2580 (.A(net1429),
    .X(net3204));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2581 (.A(_0607_),
    .X(net3205));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2582 (.A(\gpio_configure[14][6] ),
    .X(net3206));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2583 (.A(net1437),
    .X(net3207));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2584 (.A(net288),
    .X(net3208));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2585 (.A(net1591),
    .X(net3209));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2586 (.A(\gpio_configure[4][6] ),
    .X(net3210));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2587 (.A(net1488),
    .X(net3211));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2588 (.A(\gpio_configure[18][1] ),
    .X(net3212));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2589 (.A(net1336),
    .X(net3213));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold259 (.A(net2240),
    .X(net883));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2590 (.A(_0594_),
    .X(net3214));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2591 (.A(\gpio_configure[4][0] ),
    .X(net3215));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2592 (.A(net1683),
    .X(net3216));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2593 (.A(\gpio_configure[2][6] ),
    .X(net3217));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2594 (.A(net1431),
    .X(net3218));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2595 (.A(\gpio_configure[17][1] ),
    .X(net3219));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2596 (.A(net1393),
    .X(net3220));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2597 (.A(_0586_),
    .X(net3221));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2598 (.A(\gpio_configure[29][1] ),
    .X(net3222));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2599 (.A(net1631),
    .X(net3223));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold26 (.A(net2135),
    .X(net650));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold260 (.A(net2242),
    .X(net884));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2600 (.A(_0682_),
    .X(net3224));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2601 (.A(net283),
    .X(net3225));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2602 (.A(net1469),
    .X(net3226));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2603 (.A(\gpio_configure[25][1] ),
    .X(net3227));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2604 (.A(net1636),
    .X(net3228));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2605 (.A(\gpio_configure[18][6] ),
    .X(net3229));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2606 (.A(net1474),
    .X(net3230));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2607 (.A(_0599_),
    .X(net3231));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2608 (.A(\gpio_configure[29][4] ),
    .X(net3232));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2609 (.A(net1244),
    .X(net3233));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold261 (.A(net2257),
    .X(net885));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2610 (.A(\gpio_configure[7][6] ),
    .X(net3234));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2611 (.A(net1500),
    .X(net3235));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2612 (.A(_0511_),
    .X(net3236));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2613 (.A(\gpio_configure[16][6] ),
    .X(net3237));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2614 (.A(net1496),
    .X(net3238));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2615 (.A(\gpio_configure[9][6] ),
    .X(net3239));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2616 (.A(net1478),
    .X(net3240));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2617 (.A(\gpio_configure[24][6] ),
    .X(net3241));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2618 (.A(net1494),
    .X(net3242));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2619 (.A(_0647_),
    .X(net3243));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold262 (.A(net2259),
    .X(net886));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2620 (.A(\gpio_configure[11][6] ),
    .X(net3244));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2621 (.A(net1507),
    .X(net3245));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2622 (.A(\mgmt_gpio_data[8] ),
    .X(net3246));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2623 (.A(net1503),
    .X(net3247));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2624 (.A(_0119_),
    .X(net3248));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2625 (.A(\gpio_configure[5][6] ),
    .X(net3249));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2626 (.A(net1465),
    .X(net3250));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2627 (.A(\mgmt_gpio_data_buf[12] ),
    .X(net3251));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2628 (.A(net1271),
    .X(net3252));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2629 (.A(_0139_),
    .X(net3253));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold263 (.A(net2223),
    .X(net887));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2630 (.A(serial_bb_data_2),
    .X(net3254));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2631 (.A(net1490),
    .X(net3255));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2632 (.A(_0424_),
    .X(net3256));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2633 (.A(\mgmt_gpio_data[36] ),
    .X(net3257));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2634 (.A(net1250),
    .X(net3258));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2635 (.A(\gpio_configure[12][6] ),
    .X(net3259));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2636 (.A(net1486),
    .X(net3260));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2637 (.A(\gpio_configure[36][4] ),
    .X(net3261));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2638 (.A(net1263),
    .X(net3262));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2639 (.A(\gpio_configure[13][4] ),
    .X(net3263));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold264 (.A(net2225),
    .X(net888));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2640 (.A(net1261),
    .X(net3264));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2641 (.A(\gpio_configure[12][4] ),
    .X(net3265));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2642 (.A(net1334),
    .X(net3266));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2643 (.A(\gpio_configure[33][4] ),
    .X(net3267));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2644 (.A(net1304),
    .X(net3268));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2645 (.A(_0717_),
    .X(net3269));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2646 (.A(\gpio_configure[37][4] ),
    .X(net3270));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2647 (.A(net1275),
    .X(net3271));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2648 (.A(\gpio_configure[34][4] ),
    .X(net3272));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2649 (.A(net1312),
    .X(net3273));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold265 (.A(net2220),
    .X(net889));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2650 (.A(_0725_),
    .X(net3274));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2651 (.A(\mgmt_gpio_data[23] ),
    .X(net3275));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2652 (.A(net1511),
    .X(net3276));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2653 (.A(_0264_),
    .X(net3277));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2654 (.A(\gpio_configure[22][4] ),
    .X(net3278));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2655 (.A(net1316),
    .X(net3279));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2656 (.A(\gpio_configure[2][12] ),
    .X(net3280));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2657 (.A(net1377),
    .X(net3281));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2658 (.A(\gpio_configure[21][1] ),
    .X(net3282));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2659 (.A(net1730),
    .X(net3283));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold266 (.A(net2222),
    .X(net890));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2660 (.A(_0618_),
    .X(net3284));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2661 (.A(\gpio_configure[30][4] ),
    .X(net3285));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2662 (.A(net1358),
    .X(net3286));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2663 (.A(\gpio_configure[15][4] ),
    .X(net3287));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2664 (.A(net1352),
    .X(net3288));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2665 (.A(\gpio_configure[11][4] ),
    .X(net3289));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2666 (.A(net1330),
    .X(net3290));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2667 (.A(\gpio_configure[10][12] ),
    .X(net3291));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2668 (.A(net1371),
    .X(net3292));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2669 (.A(\gpio_configure[9][12] ),
    .X(net3293));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold267 (.A(net2197),
    .X(net891));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2670 (.A(net1389),
    .X(net3294));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2671 (.A(\gpio_configure[24][4] ),
    .X(net3295));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2672 (.A(net1366),
    .X(net3296));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2673 (.A(_0645_),
    .X(net3297));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2674 (.A(\gpio_configure[23][4] ),
    .X(net3298));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2675 (.A(net1364),
    .X(net3299));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2676 (.A(_0637_),
    .X(net3300));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2677 (.A(\mgmt_gpio_data[1] ),
    .X(net3301));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2678 (.A(net1505),
    .X(net3302));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2679 (.A(_0128_),
    .X(net3303));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold268 (.A(net2199),
    .X(net892));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2680 (.A(\gpio_configure[17][4] ),
    .X(net3304));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2681 (.A(net1391),
    .X(net3305));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2682 (.A(_0589_),
    .X(net3306));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2683 (.A(\mgmt_gpio_data[15] ),
    .X(net3307));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2684 (.A(net1517),
    .X(net3308));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2685 (.A(_0126_),
    .X(net3309));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2686 (.A(\mgmt_gpio_data[7] ),
    .X(net3310));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2687 (.A(net1498),
    .X(net3311));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2688 (.A(_0134_),
    .X(net3312));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2689 (.A(\gpio_configure[21][12] ),
    .X(net3313));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold269 (.A(net2310),
    .X(net893));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2690 (.A(net1387),
    .X(net3314));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2691 (.A(_0366_),
    .X(net3315));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2692 (.A(\gpio_configure[18][4] ),
    .X(net3316));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2693 (.A(net1385),
    .X(net3317));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2694 (.A(_0597_),
    .X(net3318));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2695 (.A(\gpio_configure[25][4] ),
    .X(net3319));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2696 (.A(net1405),
    .X(net3320));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2697 (.A(net295),
    .X(net3321));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2698 (.A(net1593),
    .X(net3322));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2699 (.A(\gpio_configure[27][12] ),
    .X(net3323));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold27 (.A(\gpio_configure[20][7] ),
    .X(net651));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold270 (.A(net2312),
    .X(net894));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2700 (.A(net1332),
    .X(net3324));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2701 (.A(\gpio_configure[15][12] ),
    .X(net3325));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2702 (.A(net1421),
    .X(net3326));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2703 (.A(\gpio_configure[27][8] ),
    .X(net3327));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2704 (.A(net1763),
    .X(net3328));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2705 (.A(\gpio_configure[19][4] ),
    .X(net3329));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2706 (.A(net1381),
    .X(net3330));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2707 (.A(_0605_),
    .X(net3331));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2708 (.A(\gpio_configure[28][12] ),
    .X(net3332));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2709 (.A(net1443),
    .X(net3333));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold271 (.A(net2172),
    .X(net895));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2710 (.A(\gpio_configure[18][12] ),
    .X(net3334));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2711 (.A(net1457),
    .X(net3335));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2712 (.A(_0336_),
    .X(net3336));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2713 (.A(\gpio_configure[32][12] ),
    .X(net3337));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2714 (.A(net1453),
    .X(net3338));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2715 (.A(\gpio_configure[27][9] ),
    .X(net3339));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2716 (.A(net1749),
    .X(net3340));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2717 (.A(\gpio_configure[7][0] ),
    .X(net3341));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2718 (.A(net1641),
    .X(net3342));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2719 (.A(_0505_),
    .X(net3343));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold272 (.A(net2174),
    .X(net896));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2720 (.A(\gpio_configure[22][12] ),
    .X(net3344));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2721 (.A(net1447),
    .X(net3345));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2722 (.A(_0371_),
    .X(net3346));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2723 (.A(\gpio_configure[23][12] ),
    .X(net3347));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2724 (.A(net1435),
    .X(net3348));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2725 (.A(_0241_),
    .X(net3349));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2726 (.A(\gpio_configure[6][12] ),
    .X(net3350));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2727 (.A(net1467),
    .X(net3351));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2728 (.A(\gpio_configure[20][12] ),
    .X(net3352));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2729 (.A(net1461),
    .X(net3353));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold273 (.A(net2271),
    .X(net897));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2730 (.A(_0356_),
    .X(net3354));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2731 (.A(\gpio_configure[1][12] ),
    .X(net3355));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2732 (.A(net1472),
    .X(net3356));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2733 (.A(_0152_),
    .X(net3357));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2734 (.A(\gpio_configure[0][0] ),
    .X(net3358));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2735 (.A(net1661),
    .X(net3359));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2736 (.A(_0449_),
    .X(net3360));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2737 (.A(\gpio_configure[5][0] ),
    .X(net3361));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2738 (.A(net1659),
    .X(net3362));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2739 (.A(\gpio_configure[26][12] ),
    .X(net3363));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold274 (.A(net2273),
    .X(net898));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2740 (.A(net1459),
    .X(net3364));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2741 (.A(\gpio_configure[3][0] ),
    .X(net3365));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2742 (.A(net1653),
    .X(net3366));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2743 (.A(\gpio_configure[10][0] ),
    .X(net3367));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2744 (.A(net1637),
    .X(net3368));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2745 (.A(\gpio_configure[19][12] ),
    .X(net3369));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2746 (.A(net1439),
    .X(net3370));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2747 (.A(_0346_),
    .X(net3371));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2748 (.A(\mgmt_gpio_data_buf[0] ),
    .X(net3372));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2749 (.A(net1675),
    .X(net3373));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold275 (.A(net2230),
    .X(net899));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2750 (.A(_0441_),
    .X(net3374));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2751 (.A(net289),
    .X(net3375));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2752 (.A(net1368),
    .X(net3376));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2753 (.A(\mgmt_gpio_data[5] ),
    .X(net3377));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2754 (.A(net1841),
    .X(net3378));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2755 (.A(_0132_),
    .X(net3379));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2756 (.A(\gpio_configure[2][0] ),
    .X(net3380));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2757 (.A(net1634),
    .X(net3381));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2758 (.A(\gpio_configure[13][12] ),
    .X(net3382));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2759 (.A(net1476),
    .X(net3383));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold276 (.A(net2232),
    .X(net900));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2760 (.A(\gpio_configure[34][12] ),
    .X(net3384));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2761 (.A(net1482),
    .X(net3385));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2762 (.A(net326),
    .X(net3386));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2763 (.A(net1960),
    .X(net3387));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2764 (.A(net1777),
    .X(net3388));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2765 (.A(\gpio_configure[29][12] ),
    .X(net3389));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2766 (.A(net1480),
    .X(net3390));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2767 (.A(net340),
    .X(net3391));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2768 (.A(net1963),
    .X(net3392));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2769 (.A(net1785),
    .X(net3393));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold277 (.A(net2342),
    .X(net901));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2770 (.A(\gpio_configure[2][8] ),
    .X(net3394));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2771 (.A(net1649),
    .X(net3395));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2772 (.A(\gpio_configure[15][8] ),
    .X(net3396));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2773 (.A(net1679),
    .X(net3397));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2774 (.A(\gpio_configure[19][8] ),
    .X(net3398));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2775 (.A(net1677),
    .X(net3399));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2776 (.A(_0342_),
    .X(net3400));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2777 (.A(\gpio_configure[35][12] ),
    .X(net3401));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2778 (.A(net1484),
    .X(net3402));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2779 (.A(\gpio_configure[9][8] ),
    .X(net3403));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold278 (.A(net2344),
    .X(net902));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2780 (.A(net1643),
    .X(net3404));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2781 (.A(net320),
    .X(net3405));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2782 (.A(net1967),
    .X(net3406));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2783 (.A(net1793),
    .X(net3407));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2784 (.A(net325),
    .X(net3408));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2785 (.A(net1961),
    .X(net3409));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2786 (.A(net334),
    .X(net3410));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2787 (.A(net1968),
    .X(net3411));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2788 (.A(net1789),
    .X(net3412));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2789 (.A(net321),
    .X(net3413));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold279 (.A(\wbbd_addr[5] ),
    .X(net903));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2790 (.A(net1970),
    .X(net3414));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2791 (.A(net1799),
    .X(net3415));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2792 (.A(\gpio_configure[20][8] ),
    .X(net3416));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2793 (.A(net1684),
    .X(net3417));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2794 (.A(_0352_),
    .X(net3418));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2795 (.A(net323),
    .X(net3419));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2796 (.A(net1962),
    .X(net3420));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2797 (.A(net1783),
    .X(net3421));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2798 (.A(\gpio_configure[13][8] ),
    .X(net3422));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2799 (.A(net1686),
    .X(net3423));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold28 (.A(net2102),
    .X(net652));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold280 (.A(net2451),
    .X(net904));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2800 (.A(net343),
    .X(net3424));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2801 (.A(net1971),
    .X(net3425));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2802 (.A(net1797),
    .X(net3426));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2803 (.A(\gpio_configure[35][8] ),
    .X(net3427));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2804 (.A(net1698),
    .X(net3428));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2805 (.A(net339),
    .X(net3429));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2806 (.A(net1964),
    .X(net3430));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2807 (.A(net1787),
    .X(net3431));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2808 (.A(net327),
    .X(net3432));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2809 (.A(net1959),
    .X(net3433));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold281 (.A(_0868_),
    .X(net905));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2810 (.A(net1775),
    .X(net3434));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2811 (.A(\gpio_configure[1][0] ),
    .X(net3435));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2812 (.A(net1690),
    .X(net3436));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2813 (.A(\gpio_configure[37][8] ),
    .X(net3437));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2814 (.A(net1700),
    .X(net3438));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2815 (.A(net313),
    .X(net3439));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2816 (.A(net1976),
    .X(net3440));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2817 (.A(net1813),
    .X(net3441));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2818 (.A(net312),
    .X(net3442));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2819 (.A(net1966),
    .X(net3443));
 sky130_fd_sc_hd__buf_2 hold282 (.A(net386),
    .X(net906));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2820 (.A(net1791),
    .X(net3444));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2821 (.A(\gpio_configure[10][8] ),
    .X(net3445));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2822 (.A(net1688),
    .X(net3446));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2823 (.A(net330),
    .X(net3447));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2824 (.A(net1977),
    .X(net3448));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2825 (.A(\mgmt_gpio_data[25] ),
    .X(net3449));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2826 (.A(net1632),
    .X(net3450));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2827 (.A(net322),
    .X(net3451));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2828 (.A(net1972),
    .X(net3452));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2829 (.A(\gpio_configure[20][0] ),
    .X(net3453));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold283 (.A(net2294),
    .X(net907));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2830 (.A(net1706),
    .X(net3454));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2831 (.A(_0609_),
    .X(net3455));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2832 (.A(\gpio_configure[12][8] ),
    .X(net3456));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2833 (.A(net1694),
    .X(net3457));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2834 (.A(\mgmt_gpio_data_buf[17] ),
    .X(net3458));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2835 (.A(net1647),
    .X(net3459));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2836 (.A(_0275_),
    .X(net3460));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2837 (.A(net314),
    .X(net3461));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2838 (.A(net1973),
    .X(net3462));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2839 (.A(net331),
    .X(net3463));
 sky130_fd_sc_hd__buf_6 hold284 (.A(net2388),
    .X(net908));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2840 (.A(net1984),
    .X(net3464));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2841 (.A(\gpio_configure[25][8] ),
    .X(net3465));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2842 (.A(net1692),
    .X(net3466));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2843 (.A(_0065_),
    .X(net3467));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2844 (.A(\mgmt_gpio_data[4] ),
    .X(net3468));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2845 (.A(net1218),
    .X(net3469));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2846 (.A(_0131_),
    .X(net3470));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2847 (.A(net316),
    .X(net3471));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2848 (.A(net1975),
    .X(net3472));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2849 (.A(net337),
    .X(net3473));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold285 (.A(net2390),
    .X(net909));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2850 (.A(net1965),
    .X(net3474));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2851 (.A(net1781),
    .X(net3475));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2852 (.A(net319),
    .X(net3476));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2853 (.A(net1981),
    .X(net3477));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2854 (.A(\mgmt_gpio_data[6] ),
    .X(net3478));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2855 (.A(net1669),
    .X(net3479));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2856 (.A(_0133_),
    .X(net3480));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2857 (.A(\gpio_configure[17][0] ),
    .X(net3481));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2858 (.A(net1726),
    .X(net3482));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2859 (.A(_0585_),
    .X(net3483));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold286 (.A(net2459),
    .X(net910));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2860 (.A(net336),
    .X(net3484));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2861 (.A(net1980),
    .X(net3485));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2862 (.A(net341),
    .X(net3486));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2863 (.A(net1974),
    .X(net3487));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2864 (.A(\gpio_configure[34][8] ),
    .X(net3488));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2865 (.A(net1696),
    .X(net3489));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2866 (.A(\gpio_configure[17][8] ),
    .X(net3490));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2867 (.A(net1710),
    .X(net3491));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2868 (.A(net335),
    .X(net3492));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2869 (.A(net1983),
    .X(net3493));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold287 (.A(net2461),
    .X(net911));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2870 (.A(net315),
    .X(net3494));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2871 (.A(net1982),
    .X(net3495));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2872 (.A(\gpio_configure[29][8] ),
    .X(net3496));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2873 (.A(net1718),
    .X(net3497));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2874 (.A(\gpio_configure[36][8] ),
    .X(net3498));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2875 (.A(net1722),
    .X(net3499));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2876 (.A(net342),
    .X(net3500));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2877 (.A(net1979),
    .X(net3501));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2878 (.A(\gpio_configure[30][1] ),
    .X(net3502));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2879 (.A(net1665),
    .X(net3503));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold288 (.A(net2329),
    .X(net912));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2880 (.A(\gpio_configure[27][0] ),
    .X(net3504));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2881 (.A(net1728),
    .X(net3505));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2882 (.A(net317),
    .X(net3506));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2883 (.A(net1969),
    .X(net3507));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2884 (.A(\gpio_configure[23][1] ),
    .X(net3508));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2885 (.A(net1645),
    .X(net3509));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2886 (.A(_0634_),
    .X(net3510));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2887 (.A(\gpio_configure[26][1] ),
    .X(net3511));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2888 (.A(net1667),
    .X(net3512));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2889 (.A(\clk2_output_dest[0] ),
    .X(net3513));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold289 (.A(net2331),
    .X(net913));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2890 (.A(net1663),
    .X(net3514));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2891 (.A(_0430_),
    .X(net3515));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2892 (.A(\gpio_configure[22][8] ),
    .X(net3516));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2893 (.A(net1720),
    .X(net3517));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2894 (.A(_0367_),
    .X(net3518));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2895 (.A(net329),
    .X(net3519));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2896 (.A(net1985),
    .X(net3520));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2897 (.A(\mgmt_gpio_data_buf[9] ),
    .X(net3521));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2898 (.A(net1651),
    .X(net3522));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2899 (.A(_0136_),
    .X(net3523));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold29 (.A(net2157),
    .X(net653));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold290 (.A(net2280),
    .X(net914));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2900 (.A(net318),
    .X(net3524));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2901 (.A(net1978),
    .X(net3525));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2902 (.A(\gpio_configure[14][8] ),
    .X(net3526));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2903 (.A(net1704),
    .X(net3527));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2904 (.A(\gpio_configure[33][1] ),
    .X(net3528));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2905 (.A(net1657),
    .X(net3529));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2906 (.A(_0714_),
    .X(net3530));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2907 (.A(\gpio_configure[35][1] ),
    .X(net3531));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2908 (.A(net1655),
    .X(net3532));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2909 (.A(\gpio_configure[15][0] ),
    .X(net3533));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold291 (.A(net2282),
    .X(net915));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2910 (.A(net1757),
    .X(net3534));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2911 (.A(net338),
    .X(net3535));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2912 (.A(net1987),
    .X(net3536));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2913 (.A(net333),
    .X(net3537));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2914 (.A(net1986),
    .X(net3538));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2915 (.A(net328),
    .X(net3539));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2916 (.A(net1988),
    .X(net3540));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2917 (.A(\gpio_configure[2][9] ),
    .X(net3541));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2918 (.A(net1708),
    .X(net3542));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2919 (.A(\gpio_configure[36][1] ),
    .X(net3543));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold292 (.A(net2525),
    .X(net916));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2920 (.A(net1673),
    .X(net3544));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2921 (.A(\gpio_configure[19][1] ),
    .X(net3545));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2922 (.A(net1714),
    .X(net3546));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2923 (.A(_0602_),
    .X(net3547));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2924 (.A(net324),
    .X(net3548));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2925 (.A(net1989),
    .X(net3549));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2926 (.A(\gpio_configure[23][9] ),
    .X(net3550));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2927 (.A(net1702),
    .X(net3551));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2928 (.A(_0238_),
    .X(net3552));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2929 (.A(\gpio_configure[13][9] ),
    .X(net3553));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold293 (.A(net2527),
    .X(net917));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2930 (.A(net1712),
    .X(net3554));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2931 (.A(\gpio_configure[12][1] ),
    .X(net3555));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2932 (.A(net1724),
    .X(net3556));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2933 (.A(\gpio_configure[9][9] ),
    .X(net3557));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2934 (.A(net1716),
    .X(net3558));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2935 (.A(\gpio_configure[28][9] ),
    .X(net3559));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2936 (.A(net1737),
    .X(net3560));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2937 (.A(\gpio_configure[7][12] ),
    .X(net3561));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2938 (.A(net1322),
    .X(net3562));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2939 (.A(irq_spi),
    .X(net3563));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold294 (.A(net2395),
    .X(net918));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2940 (.A(net1866),
    .X(net3564));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2941 (.A(\gpio_configure[24][12] ),
    .X(net3565));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2942 (.A(net1324),
    .X(net3566));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2943 (.A(_0251_),
    .X(net3567));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2944 (.A(\mgmt_gpio_data[16] ),
    .X(net3568));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2945 (.A(net1931),
    .X(net3569));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2946 (.A(_0257_),
    .X(net3570));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2947 (.A(\gpio_configure[27][1] ),
    .X(net3571));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2948 (.A(net1733),
    .X(net3572));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2949 (.A(\gpio_configure[23][0] ),
    .X(net3573));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold295 (.A(_0460_),
    .X(net919));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2950 (.A(net1863),
    .X(net3574));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2951 (.A(_0633_),
    .X(net3575));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2952 (.A(\mgmt_gpio_data[20] ),
    .X(net3576));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2953 (.A(net1769),
    .X(net3577));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2954 (.A(_0261_),
    .X(net3578));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2955 (.A(\gpio_configure[6][4] ),
    .X(net3579));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2956 (.A(net1340),
    .X(net3580));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2957 (.A(\gpio_configure[29][0] ),
    .X(net3581));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2958 (.A(net1862),
    .X(net3582));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2959 (.A(_0681_),
    .X(net3583));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold296 (.A(net2371),
    .X(net920));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2960 (.A(\gpio_configure[28][1] ),
    .X(net3584));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2961 (.A(net1743),
    .X(net3585));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2962 (.A(\gpio_configure[32][9] ),
    .X(net3586));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2963 (.A(net1741),
    .X(net3587));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2964 (.A(\gpio_configure[11][0] ),
    .X(net3588));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2965 (.A(net1857),
    .X(net3589));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2966 (.A(_0537_),
    .X(net3590));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2967 (.A(\mgmt_gpio_data[12] ),
    .X(net3591));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2968 (.A(net1613),
    .X(net3592));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2969 (.A(_0123_),
    .X(net3593));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold297 (.A(net2373),
    .X(net921));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2970 (.A(\gpio_configure[1][9] ),
    .X(net3594));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2971 (.A(net1761),
    .X(net3595));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2972 (.A(_0149_),
    .X(net3596));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2973 (.A(\gpio_configure[15][9] ),
    .X(net3597));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2974 (.A(net1753),
    .X(net3598));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2975 (.A(\gpio_configure[21][9] ),
    .X(net3599));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2976 (.A(net1745),
    .X(net3600));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2977 (.A(_0363_),
    .X(net3601));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2978 (.A(\gpio_configure[20][9] ),
    .X(net3602));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2979 (.A(net1751),
    .X(net3603));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold298 (.A(net2217),
    .X(net922));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2980 (.A(_0353_),
    .X(net3604));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2981 (.A(\gpio_configure[18][9] ),
    .X(net3605));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2982 (.A(net1747),
    .X(net3606));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2983 (.A(_0333_),
    .X(net3607));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2984 (.A(\gpio_configure[25][9] ),
    .X(net3608));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2985 (.A(net1771),
    .X(net3609));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2986 (.A(_0066_),
    .X(net3610));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2987 (.A(\gpio_configure[14][9] ),
    .X(net3611));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2988 (.A(net1767),
    .X(net3612));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2989 (.A(\gpio_configure[4][12] ),
    .X(net3613));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold299 (.A(net2219),
    .X(net923));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2990 (.A(net1346),
    .X(net3614));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2991 (.A(\gpio_configure[9][1] ),
    .X(net3615));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2992 (.A(net1735),
    .X(net3616));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2993 (.A(\gpio_configure[19][9] ),
    .X(net3617));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2994 (.A(net1731),
    .X(net3618));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2995 (.A(_0343_),
    .X(net3619));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2996 (.A(\gpio_configure[10][4] ),
    .X(net3620));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2997 (.A(net1350),
    .X(net3621));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2998 (.A(hkspi_disable),
    .X(net3622));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold2999 (.A(net1869),
    .X(net3623));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3 (.A(net2019),
    .X(net627));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold30 (.A(net2159),
    .X(net654));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold300 (.A(net2466),
    .X(net924));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3000 (.A(_0427_),
    .X(net3624));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3001 (.A(\mgmt_gpio_data[24] ),
    .X(net3625));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3002 (.A(net1851),
    .X(net3626));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3003 (.A(\gpio_configure[20][1] ),
    .X(net3627));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3004 (.A(net1739),
    .X(net3628));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3005 (.A(_0610_),
    .X(net3629));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3006 (.A(\gpio_configure[6][9] ),
    .X(net3630));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3007 (.A(net1759),
    .X(net3631));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3008 (.A(net272),
    .X(net3632));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3009 (.A(net1354),
    .X(net3633));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold301 (.A(net2468),
    .X(net925));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3010 (.A(\gpio_configure[30][12] ),
    .X(net3634));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3011 (.A(net1397),
    .X(net3635));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3012 (.A(\gpio_configure[33][12] ),
    .X(net3636));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3013 (.A(net1403),
    .X(net3637));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3014 (.A(\mgmt_gpio_data[17] ),
    .X(net3638));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3015 (.A(net1843),
    .X(net3639));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3016 (.A(net264),
    .X(net3640));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3017 (.A(net1362),
    .X(net3641));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3018 (.A(_0398_),
    .X(net3642));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3019 (.A(\gpio_configure[10][9] ),
    .X(net3643));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold302 (.A(net2385),
    .X(net926));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3020 (.A(net1755),
    .X(net3644));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3021 (.A(\gpio_configure[29][9] ),
    .X(net3645));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3022 (.A(net1765),
    .X(net3646));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3023 (.A(\gpio_configure[8][12] ),
    .X(net3647));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3024 (.A(net1373),
    .X(net3648));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3025 (.A(net256),
    .X(net3649));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3026 (.A(net1375),
    .X(net3650));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3027 (.A(_0403_),
    .X(net3651));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3028 (.A(net260),
    .X(net3652));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3029 (.A(net1924),
    .X(net3653));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold303 (.A(net2387),
    .X(net927));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3030 (.A(_0394_),
    .X(net3654));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3031 (.A(net281),
    .X(net3655));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3032 (.A(net1411),
    .X(net3656));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3033 (.A(\gpio_configure[6][0] ),
    .X(net3657));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3034 (.A(net1847),
    .X(net3658));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3035 (.A(\gpio_configure[37][9] ),
    .X(net3659));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3036 (.A(net1773),
    .X(net3660));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3037 (.A(serial_bb_clock),
    .X(net3661));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3038 (.A(net1360),
    .X(net3662));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3039 (.A(_0420_),
    .X(net3663));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold304 (.A(net2444),
    .X(net928));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3040 (.A(\gpio_configure[0][12] ),
    .X(net3664));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3041 (.A(net1383),
    .X(net3665));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3042 (.A(_0147_),
    .X(net3666));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3043 (.A(\gpio_configure[5][12] ),
    .X(net3667));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3044 (.A(net1409),
    .X(net3668));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3045 (.A(irq_1_inputsrc),
    .X(net3669));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3046 (.A(net1914),
    .X(net3670));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3047 (.A(_0433_),
    .X(net3671));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3048 (.A(\gpio_configure[11][12] ),
    .X(net3672));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3049 (.A(net1344),
    .X(net3673));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold305 (.A(net2446),
    .X(net929));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3050 (.A(net266),
    .X(net3674));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3051 (.A(net1853),
    .X(net3675));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3052 (.A(_0399_),
    .X(net3676));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3053 (.A(\gpio_configure[3][12] ),
    .X(net3677));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3054 (.A(net1369),
    .X(net3678));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3055 (.A(\gpio_configure[16][12] ),
    .X(net3679));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3056 (.A(net1395),
    .X(net3680));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3057 (.A(\gpio_configure[26][9] ),
    .X(net3681));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3058 (.A(net1795),
    .X(net3682));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3059 (.A(\mgmt_gpio_data[0] ),
    .X(net3683));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold306 (.A(net2339),
    .X(net930));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3060 (.A(net1845),
    .X(net3684));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3061 (.A(_0127_),
    .X(net3685));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3062 (.A(\mgmt_gpio_data[32] ),
    .X(net3686));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3063 (.A(net1937),
    .X(net3687));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3064 (.A(\gpio_configure[18][8] ),
    .X(net3688));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3065 (.A(net1878),
    .X(net3689));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3066 (.A(_0332_),
    .X(net3690));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3067 (.A(\mgmt_gpio_data[9] ),
    .X(net3691));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3068 (.A(net1849),
    .X(net3692));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3069 (.A(\gpio_configure[26][8] ),
    .X(net3693));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold307 (.A(net2341),
    .X(net931));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3070 (.A(net1884),
    .X(net3694));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3071 (.A(reset_reg),
    .X(net3695));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3072 (.A(net1941),
    .X(net3696));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3073 (.A(_0418_),
    .X(net3697));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3074 (.A(\gpio_configure[22][0] ),
    .X(net3698));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3075 (.A(net1860),
    .X(net3699));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3076 (.A(\gpio_configure[12][0] ),
    .X(net3700));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3077 (.A(net1886),
    .X(net3701));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3078 (.A(\gpio_configure[13][0] ),
    .X(net3702));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3079 (.A(net1855),
    .X(net3703));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold308 (.A(net2409),
    .X(net932));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3080 (.A(net332),
    .X(net3704));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3081 (.A(net1990),
    .X(net3705));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3082 (.A(\gpio_configure[31][0] ),
    .X(net3706));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3083 (.A(net1864),
    .X(net3707));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3084 (.A(\gpio_configure[36][0] ),
    .X(net3708));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3085 (.A(net1870),
    .X(net3709));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3086 (.A(\gpio_configure[7][8] ),
    .X(net3710));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3087 (.A(net1918),
    .X(net3711));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3088 (.A(\gpio_configure[37][0] ),
    .X(net3712));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3089 (.A(net1858),
    .X(net3713));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold309 (.A(net2411),
    .X(net933));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3090 (.A(\gpio_configure[21][8] ),
    .X(net3714));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3091 (.A(net1910),
    .X(net3715));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3092 (.A(_0362_),
    .X(net3716));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3093 (.A(\gpio_configure[26][0] ),
    .X(net3717));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3094 (.A(net1872),
    .X(net3718));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3095 (.A(\gpio_configure[33][0] ),
    .X(net3719));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3096 (.A(net1874),
    .X(net3720));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3097 (.A(_0713_),
    .X(net3721));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3098 (.A(\gpio_configure[5][8] ),
    .X(net3722));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3099 (.A(net1892),
    .X(net3723));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold31 (.A(net2150),
    .X(net655));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold310 (.A(net2507),
    .X(net934));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3100 (.A(\gpio_configure[33][8] ),
    .X(net3724));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3101 (.A(net1902),
    .X(net3725));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3102 (.A(\gpio_configure[11][8] ),
    .X(net3726));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3103 (.A(net1922),
    .X(net3727));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3104 (.A(\gpio_configure[28][8] ),
    .X(net3728));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3105 (.A(net1906),
    .X(net3729));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3106 (.A(\gpio_configure[8][8] ),
    .X(net3730));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3107 (.A(net1951),
    .X(net3731));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3108 (.A(\gpio_configure[34][0] ),
    .X(net3732));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3109 (.A(net1876),
    .X(net3733));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold311 (.A(net2509),
    .X(net935));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3110 (.A(_0721_),
    .X(net3734));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3111 (.A(\gpio_configure[32][8] ),
    .X(net3735));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3112 (.A(net1896),
    .X(net3736));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3113 (.A(\gpio_configure[1][8] ),
    .X(net3737));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3114 (.A(net1900),
    .X(net3738));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3115 (.A(_0148_),
    .X(net3739));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3116 (.A(\gpio_configure[19][0] ),
    .X(net3740));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3117 (.A(net1882),
    .X(net3741));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3118 (.A(_0601_),
    .X(net3742));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3119 (.A(\gpio_configure[18][0] ),
    .X(net3743));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold312 (.A(net2326),
    .X(net936));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3120 (.A(net1890),
    .X(net3744));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3121 (.A(_0593_),
    .X(net3745));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3122 (.A(\gpio_configure[0][8] ),
    .X(net3746));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3123 (.A(net1945),
    .X(net3747));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3124 (.A(_0143_),
    .X(net3748));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3125 (.A(net265),
    .X(net3749));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3126 (.A(net1926),
    .X(net3750));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3127 (.A(_0392_),
    .X(net3751));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3128 (.A(\gpio_configure[16][8] ),
    .X(net3752));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3129 (.A(net1957),
    .X(net3753));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold313 (.A(net2328),
    .X(net937));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3130 (.A(serial_xfer),
    .X(net3754));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3131 (.A(net1929),
    .X(net3755));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3132 (.A(_2588_),
    .X(net3756));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3133 (.A(net285),
    .X(net3757));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3134 (.A(net1933),
    .X(net3758));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3135 (.A(_0117_),
    .X(net3759));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3136 (.A(\gpio_configure[24][8] ),
    .X(net3760));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3137 (.A(net1904),
    .X(net3761));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3138 (.A(_0247_),
    .X(net3762));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3139 (.A(\gpio_configure[31][8] ),
    .X(net3763));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold314 (.A(net2596),
    .X(net938));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3140 (.A(net1898),
    .X(net3764));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3141 (.A(\gpio_configure[23][8] ),
    .X(net3765));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3142 (.A(net1888),
    .X(net3766));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3143 (.A(_0237_),
    .X(net3767));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3144 (.A(\gpio_configure[9][0] ),
    .X(net3768));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3145 (.A(net1912),
    .X(net3769));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3146 (.A(\gpio_configure[6][8] ),
    .X(net3770));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3147 (.A(net1916),
    .X(net3771));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3148 (.A(\gpio_configure[35][0] ),
    .X(net3772));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3149 (.A(net1880),
    .X(net3773));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold315 (.A(_0215_),
    .X(net939));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3150 (.A(\gpio_configure[30][8] ),
    .X(net3774));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3151 (.A(net1908),
    .X(net3775));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3152 (.A(\gpio_configure[24][0] ),
    .X(net3776));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3153 (.A(net1894),
    .X(net3777));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3154 (.A(_0641_),
    .X(net3778));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3155 (.A(\gpio_configure[3][8] ),
    .X(net3779));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3156 (.A(net1949),
    .X(net3780));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3157 (.A(net258),
    .X(net3781));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3158 (.A(net1928),
    .X(net3782));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3159 (.A(_0413_),
    .X(net3783));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold316 (.A(net2354),
    .X(net940));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3160 (.A(\gpio_configure[4][8] ),
    .X(net3784));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3161 (.A(net1920),
    .X(net3785));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3162 (.A(\gpio_configure[32][0] ),
    .X(net3786));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3163 (.A(net1935),
    .X(net3787));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3164 (.A(\gpio_configure[8][0] ),
    .X(net3788));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3165 (.A(net1939),
    .X(net3789));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3166 (.A(net293),
    .X(net3790));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3167 (.A(net1943),
    .X(net3791));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3168 (.A(net276),
    .X(net3792));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3169 (.A(net1955),
    .X(net3793));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold317 (.A(net2356),
    .X(net941));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3170 (.A(net269),
    .X(net3794));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3171 (.A(net1947),
    .X(net3795));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3172 (.A(\gpio_configure[16][0] ),
    .X(net3796));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3173 (.A(net1953),
    .X(net3797));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3174 (.A(\hkspi.ldata[6] ),
    .X(net3798));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3175 (.A(_0390_),
    .X(net3799));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3176 (.A(\hkspi.ldata[1] ),
    .X(net3800));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3177 (.A(_0385_),
    .X(net3801));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3178 (.A(\hkspi.ldata[0] ),
    .X(net3802));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3179 (.A(\hkspi.ldata[3] ),
    .X(net3803));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold318 (.A(\gpio_configure[32][10] ),
    .X(net942));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3180 (.A(_0387_),
    .X(net3804));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3181 (.A(\wbbd_state[5] ),
    .X(net3805));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3182 (.A(\hkspi.ldata[5] ),
    .X(net3806));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3183 (.A(_0389_),
    .X(net3807));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3184 (.A(\wbbd_state[2] ),
    .X(net3808));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3185 (.A(\wbbd_state[3] ),
    .X(net3809));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3186 (.A(\wbbd_state[1] ),
    .X(net3810));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3187 (.A(_3366_),
    .X(net3811));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3188 (.A(\hkspi.ldata[2] ),
    .X(net3812));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3189 (.A(\wbbd_state[7] ),
    .X(net3813));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold319 (.A(net2299),
    .X(net943));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3190 (.A(\serial_data_staging_2[9] ),
    .X(net3814));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3191 (.A(_0793_),
    .X(net3815));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3192 (.A(\wbbd_data[6] ),
    .X(net3816));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3193 (.A(\serial_data_staging_2[1] ),
    .X(net3817));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3194 (.A(_0785_),
    .X(net3818));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3195 (.A(\serial_data_staging_1[8] ),
    .X(net3819));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3196 (.A(_0779_),
    .X(net3820));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3197 (.A(\wbbd_data[2] ),
    .X(net3821));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3198 (.A(\wbbd_data[4] ),
    .X(net3822));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3199 (.A(\serial_data_staging_1[4] ),
    .X(net3823));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold32 (.A(net2152),
    .X(net656));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold320 (.A(net2276),
    .X(net944));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3200 (.A(_0775_),
    .X(net3824));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3201 (.A(\serial_data_staging_2[10] ),
    .X(net3825));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3202 (.A(\serial_data_staging_2[3] ),
    .X(net3826));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3203 (.A(_0787_),
    .X(net3827));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3204 (.A(\serial_data_staging_2[11] ),
    .X(net3828));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3205 (.A(\serial_data_staging_2[2] ),
    .X(net3829));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3206 (.A(\wbbd_data[7] ),
    .X(net3830));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3207 (.A(\serial_data_staging_1[3] ),
    .X(net3831));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3208 (.A(_0774_),
    .X(net3832));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3209 (.A(\serial_data_staging_2[4] ),
    .X(net3833));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold321 (.A(net2278),
    .X(net945));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3210 (.A(\wbbd_state[6] ),
    .X(net3834));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3211 (.A(\serial_data_staging_2[6] ),
    .X(net3835));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3212 (.A(_0790_),
    .X(net3836));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3213 (.A(\serial_data_staging_2[0] ),
    .X(net3837));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3214 (.A(_0784_),
    .X(net3838));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3215 (.A(\serial_data_staging_1[10] ),
    .X(net3839));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3216 (.A(_0781_),
    .X(net3840));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3217 (.A(\serial_data_staging_1[9] ),
    .X(net3841));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3218 (.A(\serial_data_staging_1[0] ),
    .X(net3842));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3219 (.A(\serial_data_staging_1[1] ),
    .X(net3843));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold322 (.A(net2469),
    .X(net946));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3220 (.A(\serial_data_staging_1[5] ),
    .X(net3844));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3221 (.A(\wbbd_data[1] ),
    .X(net3845));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3222 (.A(\hkspi.pre_pass_thru_user ),
    .X(net3846));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3223 (.A(_0089_),
    .X(net3847));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3224 (.A(\hkspi.addr[6] ),
    .X(net3848));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3225 (.A(\hkspi.state[1] ),
    .X(net3849));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3226 (.A(\serial_data_staging_2[7] ),
    .X(net3850));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3227 (.A(\serial_data_staging_2[8] ),
    .X(net3851));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3228 (.A(\serial_data_staging_1[2] ),
    .X(net3852));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3229 (.A(serial_clock_pre),
    .X(net3853));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold323 (.A(net2471),
    .X(net947));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3230 (.A(\wbbd_state[4] ),
    .X(net3854));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3231 (.A(_0009_),
    .X(net3855));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3232 (.A(\wbbd_addr[5] ),
    .X(net3856));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3233 (.A(\wbbd_data[5] ),
    .X(net3857));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3234 (.A(\serial_data_staging_1[12] ),
    .X(net3858));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3235 (.A(_0783_),
    .X(net3859));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3236 (.A(\hkspi.state[4] ),
    .X(net3860));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3237 (.A(_0008_),
    .X(net3861));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3238 (.A(\serial_data_staging_1[11] ),
    .X(net3862));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3239 (.A(\serial_data_staging_2[5] ),
    .X(net3863));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold324 (.A(net2254),
    .X(net948));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3240 (.A(\wbbd_addr[6] ),
    .X(net3864));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3241 (.A(\serial_data_staging_2[12] ),
    .X(net3865));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3242 (.A(\serial_data_staging_1[6] ),
    .X(net3866));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3243 (.A(\wbbd_data[3] ),
    .X(net3867));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3244 (.A(\serial_data_staging_1[7] ),
    .X(net3868));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3245 (.A(serial_load_pre),
    .X(net3869));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3246 (.A(_0770_),
    .X(net3870));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3247 (.A(\hkspi.pass_thru_user ),
    .X(net3871));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3248 (.A(\hkspi.pre_pass_thru_mgmt ),
    .X(net3872));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3249 (.A(\hkspi.SDO ),
    .X(net3873));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold325 (.A(net2256),
    .X(net949));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3250 (.A(\hkspi.pass_thru_mgmt ),
    .X(net3874));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3251 (.A(\wbbd_state[0] ),
    .X(net3875));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3252 (.A(\wbbd_state[6] ),
    .X(net3876));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3253 (.A(serial_busy),
    .X(net3877));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3254 (.A(\hkspi.fixed[0] ),
    .X(net3878));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3255 (.A(_0081_),
    .X(net3879));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3256 (.A(\hkspi.fixed[2] ),
    .X(net3880));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3257 (.A(\hkspi.addr[3] ),
    .X(net3881));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3258 (.A(\hkspi.addr[4] ),
    .X(net3882));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3259 (.A(net311),
    .X(net3883));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold326 (.A(net2457),
    .X(net950));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3260 (.A(_0797_),
    .X(net3884));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3261 (.A(\hkspi.addr[2] ),
    .X(net3885));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3262 (.A(\hkspi.writemode ),
    .X(net3886));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3263 (.A(\hkspi.fixed[1] ),
    .X(net3887));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3264 (.A(\hkspi.pass_thru_mgmt_delay ),
    .X(net3888));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3265 (.A(\xfer_count[1] ),
    .X(net3889));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3266 (.A(\hkspi.count[1] ),
    .X(net3890));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3267 (.A(\hkspi.readmode ),
    .X(net3891));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3268 (.A(\hkspi.addr[0] ),
    .X(net3892));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3269 (.A(\wbbd_state[7] ),
    .X(net3893));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold327 (.A(_0156_),
    .X(net951));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3270 (.A(\xfer_count[0] ),
    .X(net3894));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3271 (.A(_1436_),
    .X(net3895));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3272 (.A(_0014_),
    .X(net3896));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3273 (.A(\pad_count_2[5] ),
    .X(net3897));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3274 (.A(\hkspi.count[0] ),
    .X(net3898));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3275 (.A(\hkspi.state[3] ),
    .X(net3899));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3276 (.A(\pad_count_2[4] ),
    .X(net3900));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3277 (.A(\pad_count_1[0] ),
    .X(net3901));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3278 (.A(\hkspi.state[2] ),
    .X(net3902));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3279 (.A(\hkspi.wrstb ),
    .X(net3903));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold328 (.A(net2518),
    .X(net952));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3280 (.A(\hkspi.addr[1] ),
    .X(net3904));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3281 (.A(\hkspi.rdstb ),
    .X(net3905));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3282 (.A(\gpio_configure[14][0] ),
    .X(net3906));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3283 (.A(\hkspi.state[3] ),
    .X(net3907));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3284 (.A(\hkspi.count[1] ),
    .X(net3908));
 sky130_fd_sc_hd__clkdlybuf4s50_2 hold3285 (.A(hkspi_disable),
    .X(net3909));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold329 (.A(net2520),
    .X(net953));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold33 (.A(net2295),
    .X(net657));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold330 (.A(net2421),
    .X(net954));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold331 (.A(_0660_),
    .X(net955));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold332 (.A(net2332),
    .X(net956));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold333 (.A(net2334),
    .X(net957));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold334 (.A(net2397),
    .X(net958));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold335 (.A(net2399),
    .X(net959));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold336 (.A(net2335),
    .X(net960));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold337 (.A(net2337),
    .X(net961));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold338 (.A(net2307),
    .X(net962));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold339 (.A(net2309),
    .X(net963));
 sky130_fd_sc_hd__buf_2 hold34 (.A(net2297),
    .X(net658));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold340 (.A(net2264),
    .X(net964));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold341 (.A(net2266),
    .X(net965));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold342 (.A(net2480),
    .X(net966));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold343 (.A(net2482),
    .X(net967));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold344 (.A(net2423),
    .X(net968));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold345 (.A(net2425),
    .X(net969));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold346 (.A(net2484),
    .X(net970));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold347 (.A(net2486),
    .X(net971));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold348 (.A(net2515),
    .X(net972));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold349 (.A(net2517),
    .X(net973));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold35 (.A(_0847_),
    .X(net659));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold350 (.A(net2488),
    .X(net974));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold351 (.A(_0692_),
    .X(net975));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold352 (.A(net2352),
    .X(net976));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold353 (.A(_0349_),
    .X(net977));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold354 (.A(net2553),
    .X(net978));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold355 (.A(net2555),
    .X(net979));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold356 (.A(\gpio_configure[27][10] ),
    .X(net980));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold357 (.A(net2211),
    .X(net981));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold358 (.A(net2316),
    .X(net982));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold359 (.A(net2318),
    .X(net983));
 sky130_fd_sc_hd__buf_12 hold36 (.A(net421),
    .X(net660));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold360 (.A(net2562),
    .X(net984));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold361 (.A(net2564),
    .X(net985));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold362 (.A(net2464),
    .X(net986));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold363 (.A(_0691_),
    .X(net987));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold364 (.A(net2418),
    .X(net988));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold365 (.A(net2420),
    .X(net989));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold366 (.A(net2532),
    .X(net990));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold367 (.A(net2534),
    .X(net991));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold368 (.A(net2426),
    .X(net992));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold369 (.A(net2428),
    .X(net993));
 sky130_fd_sc_hd__buf_4 hold37 (.A(_2631_),
    .X(net661));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold370 (.A(net2610),
    .X(net994));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold371 (.A(_0235_),
    .X(net995));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold372 (.A(net2435),
    .X(net996));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold373 (.A(net2437),
    .X(net997));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold374 (.A(net2274),
    .X(net998));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold375 (.A(_0254_),
    .X(net999));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold376 (.A(net2441),
    .X(net1000));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold377 (.A(net2443),
    .X(net1001));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold378 (.A(net2404),
    .X(net1002));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold379 (.A(net2406),
    .X(net1003));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold38 (.A(net2203),
    .X(net662));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold380 (.A(net2447),
    .X(net1004));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold381 (.A(_0708_),
    .X(net1005));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold382 (.A(net2366),
    .X(net1006));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold383 (.A(_0245_),
    .X(net1007));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold384 (.A(net2675),
    .X(net1008));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold385 (.A(_0255_),
    .X(net1009));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold386 (.A(net2401),
    .X(net1010));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold387 (.A(net2403),
    .X(net1011));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold388 (.A(net2800),
    .X(net1012));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold389 (.A(_0504_),
    .X(net1013));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold39 (.A(net2233),
    .X(net663));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold390 (.A(net2559),
    .X(net1014));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold391 (.A(net2561),
    .X(net1015));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold392 (.A(net2809),
    .X(net1016));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold393 (.A(_0464_),
    .X(net1017));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold394 (.A(net2794),
    .X(net1018));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold395 (.A(net2796),
    .X(net1019));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold396 (.A(\hkspi.addr[3] ),
    .X(net1020));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold397 (.A(_0838_),
    .X(net1021));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold398 (.A(_0839_),
    .X(net1022));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold399 (.A(_0840_),
    .X(net1023));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold4 (.A(net2024),
    .X(net628));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold40 (.A(net2235),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd1_1 hold400 (.A(_0860_),
    .X(net1024));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold401 (.A(net2552),
    .X(net1025));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold402 (.A(net2412),
    .X(net1026));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold403 (.A(net2414),
    .X(net1027));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold404 (.A(net2512),
    .X(net1028));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold405 (.A(net2514),
    .X(net1029));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold406 (.A(net2556),
    .X(net1030));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold407 (.A(net2558),
    .X(net1031));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold408 (.A(net2360),
    .X(net1032));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold409 (.A(net2362),
    .X(net1033));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold41 (.A(net2345),
    .X(net665));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold410 (.A(net2785),
    .X(net1034));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold411 (.A(net2787),
    .X(net1035));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold412 (.A(net2430),
    .X(net1036));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold413 (.A(net2432),
    .X(net1037));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold414 (.A(net2320),
    .X(net1038));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold415 (.A(net2322),
    .X(net1039));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold416 (.A(net2565),
    .X(net1040));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold417 (.A(_0382_),
    .X(net1041));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold418 (.A(net2407),
    .X(net1042));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold419 (.A(_0381_),
    .X(net1043));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold42 (.A(net2347),
    .X(net666));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold420 (.A(net2438),
    .X(net1044));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold421 (.A(net2440),
    .X(net1045));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold422 (.A(net2592),
    .X(net1046));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold423 (.A(net2594),
    .X(net1047));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold424 (.A(net2581),
    .X(net1048));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold425 (.A(net2583),
    .X(net1049));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold426 (.A(net2490),
    .X(net1050));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold427 (.A(_0659_),
    .X(net1051));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold428 (.A(net2567),
    .X(net1052));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold429 (.A(net2569),
    .X(net1053));
 sky130_fd_sc_hd__buf_12 hold43 (.A(net2349),
    .X(net667));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold430 (.A(net2639),
    .X(net1054));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold431 (.A(net2641),
    .X(net1055));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold432 (.A(net2522),
    .X(net1056));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold433 (.A(net2524),
    .X(net1057));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold434 (.A(net2607),
    .X(net1058));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold435 (.A(net2609),
    .X(net1059));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold436 (.A(net2806),
    .X(net1060));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold437 (.A(net2808),
    .X(net1061));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold438 (.A(net2642),
    .X(net1062));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold439 (.A(net2644),
    .X(net1063));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold44 (.A(net2394),
    .X(net668));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold440 (.A(net2623),
    .X(net1064));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold441 (.A(net2625),
    .X(net1065));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold442 (.A(net2654),
    .X(net1066));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold443 (.A(net2656),
    .X(net1067));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold444 (.A(net2819),
    .X(net1068));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold445 (.A(net2821),
    .X(net1069));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold446 (.A(net2577),
    .X(net1070));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold447 (.A(net2579),
    .X(net1071));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold448 (.A(net2504),
    .X(net1072));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold449 (.A(net2506),
    .X(net1073));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold45 (.A(net2039),
    .X(net669));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold450 (.A(net2598),
    .X(net1074));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold451 (.A(_0200_),
    .X(net1075));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold452 (.A(net2603),
    .X(net1076));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold453 (.A(net2605),
    .X(net1077));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold454 (.A(net2860),
    .X(net1078));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold455 (.A(net2862),
    .X(net1079));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold456 (.A(net2476),
    .X(net1080));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold457 (.A(net2478),
    .X(net1081));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold458 (.A(net2826),
    .X(net1082));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold459 (.A(net2828),
    .X(net1083));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold46 (.A(net2041),
    .X(net670));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold460 (.A(net2822),
    .X(net1084));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold461 (.A(_0520_),
    .X(net1085));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold462 (.A(net2660),
    .X(net1086));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold463 (.A(net2662),
    .X(net1087));
 sky130_fd_sc_hd__buf_12 hold464 (.A(net2664),
    .X(net1088));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold465 (.A(net2744),
    .X(net1089));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold466 (.A(net2570),
    .X(net1090));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold467 (.A(net2572),
    .X(net1091));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold468 (.A(net2745),
    .X(net1092));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold469 (.A(net2747),
    .X(net1093));
 sky130_fd_sc_hd__buf_12 hold47 (.A(net506),
    .X(net671));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold470 (.A(\gpio_configure[6][10] ),
    .X(net1094));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold471 (.A(net2455),
    .X(net1095));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold472 (.A(net2873),
    .X(net1096));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold473 (.A(_0415_),
    .X(net1097));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold474 (.A(net2737),
    .X(net1098));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold475 (.A(_0649_),
    .X(net1099));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold476 (.A(net2573),
    .X(net1100));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold477 (.A(net2575),
    .X(net1101));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold478 (.A(net2617),
    .X(net1102));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold479 (.A(net2619),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_16 hold48 (.A(net505),
    .X(net672));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold480 (.A(net2811),
    .X(net1104));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold481 (.A(net2813),
    .X(net1105));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold482 (.A(net2669),
    .X(net1106));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold483 (.A(net2671),
    .X(net1107));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold484 (.A(net2798),
    .X(net1108));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold485 (.A(_0488_),
    .X(net1109));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold486 (.A(net2657),
    .X(net1110));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold487 (.A(net2659),
    .X(net1111));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold488 (.A(net2600),
    .X(net1112));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold489 (.A(net2602),
    .X(net1113));
 sky130_fd_sc_hd__buf_6 hold49 (.A(_2607_),
    .X(net673));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold490 (.A(net2672),
    .X(net1114));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold491 (.A(net2674),
    .X(net1115));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold492 (.A(net2824),
    .X(net1116));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold493 (.A(_0664_),
    .X(net1117));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold494 (.A(net2636),
    .X(net1118));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold495 (.A(net2638),
    .X(net1119));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold496 (.A(net2814),
    .X(net1120));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold497 (.A(net2816),
    .X(net1121));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold498 (.A(net2501),
    .X(net1122));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold499 (.A(net2503),
    .X(net1123));
 sky130_fd_sc_hd__buf_12 hold5 (.A(net2026),
    .X(net629));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold50 (.A(net2370),
    .X(net674));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold500 (.A(net2917),
    .X(net1124));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold501 (.A(net2919),
    .X(net1125));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold502 (.A(net2855),
    .X(net1126));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold503 (.A(net2857),
    .X(net1127));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold504 (.A(net2621),
    .X(net1128));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold505 (.A(_0209_),
    .X(net1129));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold506 (.A(net2472),
    .X(net1130));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold507 (.A(net2474),
    .X(net1131));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold508 (.A(net2680),
    .X(net1132));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold509 (.A(net2682),
    .X(net1133));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold51 (.A(\hkspi.addr[6] ),
    .X(net675));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold510 (.A(net2647),
    .X(net1134));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold511 (.A(net2649),
    .X(net1135));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold512 (.A(net2510),
    .X(net1136));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold513 (.A(_0176_),
    .X(net1137));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold514 (.A(net2832),
    .X(net1138));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold515 (.A(net2834),
    .X(net1139));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold516 (.A(net2900),
    .X(net1140));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold517 (.A(_0744_),
    .X(net1141));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold518 (.A(net2588),
    .X(net1142));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold519 (.A(net2590),
    .X(net1143));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold52 (.A(net2847),
    .X(net676));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold520 (.A(net2535),
    .X(net1144));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold521 (.A(net2537),
    .X(net1145));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold522 (.A(net2842),
    .X(net1146));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold523 (.A(net2844),
    .X(net1147));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold524 (.A(net2547),
    .X(net1148));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold525 (.A(net2549),
    .X(net1149));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold526 (.A(net2865),
    .X(net1150));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold527 (.A(net2867),
    .X(net1151));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold528 (.A(\wbbd_addr[6] ),
    .X(net1152));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold529 (.A(_0836_),
    .X(net1153));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold53 (.A(_0858_),
    .X(net677));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold530 (.A(net2848),
    .X(net1154));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold531 (.A(net2850),
    .X(net1155));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold532 (.A(net2880),
    .X(net1156));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold533 (.A(_0498_),
    .X(net1157));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold534 (.A(net2882),
    .X(net1158));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold535 (.A(_0712_),
    .X(net1159));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold536 (.A(net2868),
    .X(net1160));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold537 (.A(net2870),
    .X(net1161));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold538 (.A(net2757),
    .X(net1162));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold539 (.A(net2759),
    .X(net1163));
 sky130_fd_sc_hd__buf_2 hold54 (.A(_0859_),
    .X(net678));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold540 (.A(net2858),
    .X(net1164));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold541 (.A(_0706_),
    .X(net1165));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold542 (.A(net2689),
    .X(net1166));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold543 (.A(net2835),
    .X(net1167));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold544 (.A(net2837),
    .X(net1168));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold545 (.A(net2544),
    .X(net1169));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold546 (.A(net2546),
    .X(net1170));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold547 (.A(net2933),
    .X(net1171));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold548 (.A(_0273_),
    .X(net1172));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold549 (.A(net2614),
    .X(net1173));
 sky130_fd_sc_hd__buf_4 hold55 (.A(net2114),
    .X(net679));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold550 (.A(net2616),
    .X(net1174));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold551 (.A(net2629),
    .X(net1175));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold552 (.A(_0707_),
    .X(net1176));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold553 (.A(net2584),
    .X(net1177));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold554 (.A(net2586),
    .X(net1178));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold555 (.A(net2890),
    .X(net1179));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold556 (.A(_0656_),
    .X(net1180));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold557 (.A(net2902),
    .X(net1181));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold558 (.A(net2904),
    .X(net1182));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold559 (.A(net2645),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_4 hold56 (.A(net354),
    .X(net680));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold560 (.A(_0515_),
    .X(net1184));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold561 (.A(net2863),
    .X(net1185));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold562 (.A(_0514_),
    .X(net1186));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold563 (.A(net2925),
    .X(net1187));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold564 (.A(_0680_),
    .X(net1188));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold565 (.A(net2677),
    .X(net1189));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold566 (.A(net2679),
    .X(net1190));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold567 (.A(net3906),
    .X(net1191));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold568 (.A(net2894),
    .X(net1192));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold569 (.A(net2896),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_4 hold57 (.A(_1558_),
    .X(net681));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold570 (.A(net2852),
    .X(net1194));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold571 (.A(net2854),
    .X(net1195));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold572 (.A(net2612),
    .X(net1196));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold573 (.A(_0204_),
    .X(net1197));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold574 (.A(net2631),
    .X(net1198));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold575 (.A(net2633),
    .X(net1199));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold576 (.A(net2945),
    .X(net1200));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold577 (.A(_0490_),
    .X(net1201));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold578 (.A(net2666),
    .X(net1202));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold579 (.A(net2668),
    .X(net1203));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold58 (.A(net2350),
    .X(net682));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold580 (.A(net2907),
    .X(net1204));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold581 (.A(net2909),
    .X(net1205));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold582 (.A(net2897),
    .X(net1206));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold583 (.A(net2899),
    .X(net1207));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold584 (.A(net2930),
    .X(net1208));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold585 (.A(net2932),
    .X(net1209));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold586 (.A(\gpio_configure[7][1] ),
    .X(net1210));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold587 (.A(net2938),
    .X(net1211));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold588 (.A(net2951),
    .X(net1212));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold589 (.A(_0474_),
    .X(net1213));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold59 (.A(net2283),
    .X(net683));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold590 (.A(net2884),
    .X(net1214));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold591 (.A(_0528_),
    .X(net1215));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold592 (.A(net2962),
    .X(net1216));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold593 (.A(net2964),
    .X(net1217));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold594 (.A(net3468),
    .X(net1218));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold595 (.A(net3470),
    .X(net1219));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold596 (.A(net2634),
    .X(net1220));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold597 (.A(_0189_),
    .X(net1221));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold598 (.A(net2886),
    .X(net1222));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold599 (.A(net2888),
    .X(net1223));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold6 (.A(net2029),
    .X(net630));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold60 (.A(net2285),
    .X(net684));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold600 (.A(net2912),
    .X(net1224));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold601 (.A(net2914),
    .X(net1225));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold602 (.A(net2915),
    .X(net1226));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold603 (.A(_0584_),
    .X(net1227));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold604 (.A(net2878),
    .X(net1228));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold605 (.A(_0482_),
    .X(net1229));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold606 (.A(net3002),
    .X(net1230));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold607 (.A(net3004),
    .X(net1231));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold608 (.A(net2650),
    .X(net1232));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold609 (.A(net2652),
    .X(net1233));
 sky130_fd_sc_hd__buf_12 hold61 (.A(net2287),
    .X(net685));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold610 (.A(net2871),
    .X(net1234));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold611 (.A(_0568_),
    .X(net1235));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold612 (.A(net2942),
    .X(net1236));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold613 (.A(net2944),
    .X(net1237));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold614 (.A(net2817),
    .X(net1238));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold615 (.A(_0689_),
    .X(net1239));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold616 (.A(net3009),
    .X(net1240));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold617 (.A(_0228_),
    .X(net1241));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold618 (.A(net3033),
    .X(net1242));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold619 (.A(net3035),
    .X(net1243));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold62 (.A(net2325),
    .X(net686));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold620 (.A(net3232),
    .X(net1244));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold621 (.A(_0685_),
    .X(net1245));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold622 (.A(net2683),
    .X(net1246));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold623 (.A(net2711),
    .X(net1247));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold624 (.A(net2995),
    .X(net1248));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold625 (.A(net2997),
    .X(net1249));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold626 (.A(net3257),
    .X(net1250));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold627 (.A(_0439_),
    .X(net1251));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold628 (.A(net2714),
    .X(net1252));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold629 (.A(net2981),
    .X(net1253));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold63 (.A(net2498),
    .X(net687));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold630 (.A(_0223_),
    .X(net1254));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold631 (.A(net3093),
    .X(net1255));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold632 (.A(_0458_),
    .X(net1256));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold633 (.A(net3022),
    .X(net1257));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold634 (.A(net3024),
    .X(net1258));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold635 (.A(net3111),
    .X(net1259));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold636 (.A(_0308_),
    .X(net1260));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold637 (.A(net3263),
    .X(net1261));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold638 (.A(_0557_),
    .X(net1262));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold639 (.A(net3261),
    .X(net1263));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold64 (.A(net2500),
    .X(net688));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold640 (.A(_0741_),
    .X(net1264));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold641 (.A(net3130),
    .X(net1265));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold642 (.A(_0323_),
    .X(net1266));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold643 (.A(net2840),
    .X(net1267));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold644 (.A(_0673_),
    .X(net1268));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold645 (.A(net3062),
    .X(net1269));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold646 (.A(net3064),
    .X(net1270));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold647 (.A(net3251),
    .X(net1271));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold648 (.A(net3253),
    .X(net1272));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold649 (.A(net3076),
    .X(net1273));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold65 (.A(net2462),
    .X(net689));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold650 (.A(net3078),
    .X(net1274));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold651 (.A(net3270),
    .X(net1275));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold652 (.A(_0749_),
    .X(net1276));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold653 (.A(net3072),
    .X(net1277));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold654 (.A(_0298_),
    .X(net1278));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold655 (.A(net2723),
    .X(net1279));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold656 (.A(net3083),
    .X(net1280));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold657 (.A(net3085),
    .X(net1281));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold658 (.A(net3103),
    .X(net1282));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold659 (.A(net3105),
    .X(net1283));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold66 (.A(_0203_),
    .X(net690));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold660 (.A(net3167),
    .X(net1284));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold661 (.A(_0102_),
    .X(net1285));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold662 (.A(net3091),
    .X(net1286));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold663 (.A(_0175_),
    .X(net1287));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold664 (.A(net3095),
    .X(net1288));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold665 (.A(_0110_),
    .X(net1289));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold666 (.A(net3147),
    .X(net1290));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold667 (.A(_0208_),
    .X(net1291));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold668 (.A(net3135),
    .X(net1292));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold669 (.A(_0188_),
    .X(net1293));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold67 (.A(net2382),
    .X(net691));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold670 (.A(net3121),
    .X(net1294));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold671 (.A(_0318_),
    .X(net1295));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold672 (.A(net3137),
    .X(net1296));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold673 (.A(_0578_),
    .X(net1297));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold674 (.A(net3154),
    .X(net1298));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold675 (.A(net3156),
    .X(net1299));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold676 (.A(net3118),
    .X(net1300));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold677 (.A(net3120),
    .X(net1301));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold678 (.A(net3106),
    .X(net1302));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold679 (.A(net3108),
    .X(net1303));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold68 (.A(net2384),
    .X(net692));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold680 (.A(net3267),
    .X(net1304));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold681 (.A(net3269),
    .X(net1305));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold682 (.A(net2686),
    .X(net1306));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold683 (.A(net2688),
    .X(net1307));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold684 (.A(net3050),
    .X(net1308));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold685 (.A(_0436_),
    .X(net1309));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold686 (.A(net3145),
    .X(net1310));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold687 (.A(_0530_),
    .X(net1311));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold688 (.A(net3272),
    .X(net1312));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold689 (.A(net3274),
    .X(net1313));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold69 (.A(net2087),
    .X(net693));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold690 (.A(net3157),
    .X(net1314));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold691 (.A(_0328_),
    .X(net1315));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold692 (.A(net3278),
    .X(net1316));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold693 (.A(_0629_),
    .X(net1317));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold694 (.A(net3143),
    .X(net1318));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold695 (.A(_0313_),
    .X(net1319));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold696 (.A(net3116),
    .X(net1320));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold697 (.A(_0193_),
    .X(net1321));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold698 (.A(net3561),
    .X(net1322));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold699 (.A(_0206_),
    .X(net1323));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold7 (.A(net2030),
    .X(net631));
 sky130_fd_sc_hd__buf_2 hold70 (.A(net2089),
    .X(net694));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold700 (.A(net3565),
    .X(net1324));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold701 (.A(net3567),
    .X(net1325));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold702 (.A(net3185),
    .X(net1326));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold703 (.A(net3187),
    .X(net1327));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold704 (.A(net3163),
    .X(net1328));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold705 (.A(_0348_),
    .X(net1329));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold706 (.A(net3289),
    .X(net1330));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold707 (.A(_0541_),
    .X(net1331));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold708 (.A(net3323),
    .X(net1332));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold709 (.A(_0246_),
    .X(net1333));
 sky130_fd_sc_hd__buf_2 hold71 (.A(_0866_),
    .X(net695));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold710 (.A(net3265),
    .X(net1334));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold711 (.A(_0549_),
    .X(net1335));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold712 (.A(net3212),
    .X(net1336));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold713 (.A(net3214),
    .X(net1337));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold714 (.A(net2705),
    .X(net1338));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold715 (.A(net2707),
    .X(net1339));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold716 (.A(net3579),
    .X(net1340));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold717 (.A(_0501_),
    .X(net1341));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold718 (.A(net3048),
    .X(net1342));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold719 (.A(_0463_),
    .X(net1343));
 sky130_fd_sc_hd__clkbuf_2 hold72 (.A(_0899_),
    .X(net696));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold720 (.A(net3672),
    .X(net1344));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold721 (.A(_0226_),
    .X(net1345));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold722 (.A(net3613),
    .X(net1346));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold723 (.A(_0191_),
    .X(net1347));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold724 (.A(net3128),
    .X(net1348));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold725 (.A(_0570_),
    .X(net1349));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold726 (.A(net3620),
    .X(net1350));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold727 (.A(_0533_),
    .X(net1351));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold728 (.A(net3287),
    .X(net1352));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold729 (.A(_0573_),
    .X(net1353));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold73 (.A(net2417),
    .X(net697));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold730 (.A(net3632),
    .X(net1354));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold731 (.A(_0105_),
    .X(net1355));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold732 (.A(net3067),
    .X(net1356));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold733 (.A(net3069),
    .X(net1357));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold734 (.A(net3285),
    .X(net1358));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold735 (.A(_0693_),
    .X(net1359));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold736 (.A(net3661),
    .X(net1360));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold737 (.A(net3663),
    .X(net1361));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold738 (.A(net3640),
    .X(net1362));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold739 (.A(net3642),
    .X(net1363));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold74 (.A(net2376),
    .X(net698));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold740 (.A(net3298),
    .X(net1364));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold741 (.A(net3300),
    .X(net1365));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold742 (.A(net3295),
    .X(net1366));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold743 (.A(net3297),
    .X(net1367));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold744 (.A(net3375),
    .X(net1368));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold745 (.A(net3677),
    .X(net1369));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold746 (.A(_0178_),
    .X(net1370));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold747 (.A(net3291),
    .X(net1371));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold748 (.A(_0221_),
    .X(net1372));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold749 (.A(net3647),
    .X(net1373));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold75 (.A(net2378),
    .X(net699));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold750 (.A(_0211_),
    .X(net1374));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold751 (.A(net3649),
    .X(net1375));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold752 (.A(net3651),
    .X(net1376));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold753 (.A(net3280),
    .X(net1377));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold754 (.A(_0157_),
    .X(net1378));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold755 (.A(net3169),
    .X(net1379));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold756 (.A(net3171),
    .X(net1380));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold757 (.A(net3329),
    .X(net1381));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold758 (.A(net3331),
    .X(net1382));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold759 (.A(net3664),
    .X(net1383));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold76 (.A(\gpio_configure[28][6] ),
    .X(net700));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold760 (.A(net3666),
    .X(net1384));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold761 (.A(net3316),
    .X(net1385));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold762 (.A(net3318),
    .X(net1386));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold763 (.A(net3313),
    .X(net1387));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold764 (.A(net3315),
    .X(net1388));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold765 (.A(net3293),
    .X(net1389));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold766 (.A(_0216_),
    .X(net1390));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold767 (.A(net3304),
    .X(net1391));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold768 (.A(net3306),
    .X(net1392));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold769 (.A(net3219),
    .X(net1393));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold77 (.A(net2288),
    .X(net701));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold770 (.A(net3221),
    .X(net1394));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold771 (.A(net3679),
    .X(net1395));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold772 (.A(_0316_),
    .X(net1396));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold773 (.A(net3634),
    .X(net1397));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold774 (.A(_0361_),
    .X(net1398));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold775 (.A(net2717),
    .X(net1399));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold776 (.A(net2719),
    .X(net1400));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold777 (.A(net3179),
    .X(net1401));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold778 (.A(_0671_),
    .X(net1402));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold779 (.A(net3636),
    .X(net1403));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold78 (.A(net2313),
    .X(net702));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold780 (.A(_0331_),
    .X(net1404));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold781 (.A(net3319),
    .X(net1405));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold782 (.A(_0653_),
    .X(net1406));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold783 (.A(net3139),
    .X(net1407));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold784 (.A(_0519_),
    .X(net1408));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold785 (.A(net3667),
    .X(net1409));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold786 (.A(_0196_),
    .X(net1410));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold787 (.A(net3655),
    .X(net1411));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold788 (.A(_0409_),
    .X(net1412));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold789 (.A(net3181),
    .X(net1413));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold79 (.A(net2315),
    .X(net703));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold790 (.A(_0631_),
    .X(net1414));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold791 (.A(net3177),
    .X(net1415));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold792 (.A(_0479_),
    .X(net1416));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold793 (.A(net3190),
    .X(net1417));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold794 (.A(_0559_),
    .X(net1418));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold795 (.A(net3165),
    .X(net1419));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold796 (.A(_0575_),
    .X(net1420));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold797 (.A(net3325),
    .X(net1421));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold798 (.A(_0306_),
    .X(net1422));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold799 (.A(net2739),
    .X(net1423));
 sky130_fd_sc_hd__buf_12 hold8 (.A(net2032),
    .X(net632));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold80 (.A(net2374),
    .X(net704));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold800 (.A(net2741),
    .X(net1424));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold801 (.A(net3159),
    .X(net1425));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold802 (.A(_0663_),
    .X(net1426));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold803 (.A(net3200),
    .X(net1427));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold804 (.A(net3202),
    .X(net1428));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold805 (.A(net3203),
    .X(net1429));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold806 (.A(net3205),
    .X(net1430));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold807 (.A(net3217),
    .X(net1431));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold808 (.A(_0471_),
    .X(net1432));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold809 (.A(net3149),
    .X(net1433));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold81 (.A(_0655_),
    .X(net705));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold810 (.A(net3151),
    .X(net1434));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold811 (.A(net3347),
    .X(net1435));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold812 (.A(net3349),
    .X(net1436));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold813 (.A(net3206),
    .X(net1437));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold814 (.A(_0567_),
    .X(net1438));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold815 (.A(net3369),
    .X(net1439));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold816 (.A(net3371),
    .X(net1440));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold817 (.A(net2776),
    .X(net1441));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold818 (.A(net2778),
    .X(net1442));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold819 (.A(net3332),
    .X(net1443));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold82 (.A(net2692),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold820 (.A(_0383_),
    .X(net1444));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold821 (.A(net3188),
    .X(net1445));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold822 (.A(_0503_),
    .X(net1446));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold823 (.A(net3344),
    .X(net1447));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold824 (.A(net3346),
    .X(net1448));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold825 (.A(net2754),
    .X(net1449));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold826 (.A(net2756),
    .X(net1450));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold827 (.A(net3175),
    .X(net1451));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold828 (.A(_0751_),
    .X(net1452));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold829 (.A(net3337),
    .X(net1453));
 sky130_fd_sc_hd__clkbuf_4 hold83 (.A(net2695),
    .X(net707));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold830 (.A(_0341_),
    .X(net1454));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold831 (.A(net3192),
    .X(net1455));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold832 (.A(_0711_),
    .X(net1456));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold833 (.A(net3334),
    .X(net1457));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold834 (.A(net3336),
    .X(net1458));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold835 (.A(net3363),
    .X(net1459));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold836 (.A(_0256_),
    .X(net1460));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold837 (.A(net3352),
    .X(net1461));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold838 (.A(net3354),
    .X(net1462));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold839 (.A(net3197),
    .X(net1463));
 sky130_fd_sc_hd__buf_12 hold84 (.A(net475),
    .X(net708));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold840 (.A(net3199),
    .X(net1464));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold841 (.A(net3249),
    .X(net1465));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold842 (.A(_0495_),
    .X(net1466));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold843 (.A(net3350),
    .X(net1467));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold844 (.A(_0201_),
    .X(net1468));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold845 (.A(net3225),
    .X(net1469));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold846 (.A(_0411_),
    .X(net1470));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold847 (.A(net2791),
    .X(net1471));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold848 (.A(net3355),
    .X(net1472));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold849 (.A(net3357),
    .X(net1473));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold85 (.A(_0461_),
    .X(net709));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold850 (.A(net3229),
    .X(net1474));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold851 (.A(net3231),
    .X(net1475));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold852 (.A(net3382),
    .X(net1476));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold853 (.A(_0286_),
    .X(net1477));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold854 (.A(net3239),
    .X(net1478));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold855 (.A(_0527_),
    .X(net1479));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold856 (.A(net3389),
    .X(net1480));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold857 (.A(_0236_),
    .X(net1481));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold858 (.A(net3384),
    .X(net1482));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold859 (.A(_0321_),
    .X(net1483));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold86 (.A(net2910),
    .X(net710));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold860 (.A(net3401),
    .X(net1484));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold861 (.A(_0311_),
    .X(net1485));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold862 (.A(net3259),
    .X(net1486));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold863 (.A(_0551_),
    .X(net1487));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold864 (.A(net3210),
    .X(net1488));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold865 (.A(_0487_),
    .X(net1489));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold866 (.A(net3254),
    .X(net1490));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold867 (.A(net3256),
    .X(net1491));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold868 (.A(net2788),
    .X(net1492));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold869 (.A(net2790),
    .X(net1493));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold87 (.A(_0517_),
    .X(net711));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold870 (.A(net3241),
    .X(net1494));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold871 (.A(net3243),
    .X(net1495));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold872 (.A(net3237),
    .X(net1496));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold873 (.A(_0583_),
    .X(net1497));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold874 (.A(net3310),
    .X(net1498));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold875 (.A(net3312),
    .X(net1499));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold876 (.A(net3234),
    .X(net1500));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold877 (.A(net3236),
    .X(net1501));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold878 (.A(net2829),
    .X(net1502));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold879 (.A(net3246),
    .X(net1503));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold88 (.A(net2957),
    .X(net712));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold880 (.A(net3248),
    .X(net1504));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold881 (.A(net3301),
    .X(net1505));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold882 (.A(net3303),
    .X(net1506));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold883 (.A(net3244),
    .X(net1507));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold884 (.A(_0543_),
    .X(net1508));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold885 (.A(net2802),
    .X(net1509));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold886 (.A(_0437_),
    .X(net1510));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold887 (.A(net3275),
    .X(net1511));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold888 (.A(net3277),
    .X(net1512));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold889 (.A(net2804),
    .X(net1513));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold89 (.A(_0477_),
    .X(net713));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold890 (.A(_0462_),
    .X(net1514));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold891 (.A(net2838),
    .X(net1515));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold892 (.A(_0502_),
    .X(net1516));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold893 (.A(net3307),
    .X(net1517));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold894 (.A(net3309),
    .X(net1518));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold895 (.A(net2947),
    .X(net1519));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold896 (.A(_0155_),
    .X(net1520));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold897 (.A(net2979),
    .X(net1521));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold898 (.A(_0534_),
    .X(net1522));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold899 (.A(net2968),
    .X(net1523));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold9 (.A(net2035),
    .X(net633));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold90 (.A(net2020),
    .X(net714));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold900 (.A(_0470_),
    .X(net1524));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold901 (.A(net2922),
    .X(net1525));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold902 (.A(net2924),
    .X(net1526));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold903 (.A(net2875),
    .X(net1527));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold904 (.A(net2877),
    .X(net1528));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold905 (.A(net3099),
    .X(net1529));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold906 (.A(_0234_),
    .X(net1530));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold907 (.A(net2998),
    .X(net1531));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold908 (.A(_0219_),
    .X(net1532));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold909 (.A(net2920),
    .X(net1533));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold91 (.A(net2022),
    .X(net715));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold910 (.A(_0582_),
    .X(net1534));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold911 (.A(net3017),
    .X(net1535));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold912 (.A(net3019),
    .X(net1536));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold913 (.A(net2959),
    .X(net1537));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold914 (.A(net2961),
    .X(net1538));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold915 (.A(net3015),
    .X(net1539));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold916 (.A(_0205_),
    .X(net1540));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold917 (.A(net2986),
    .X(net1541));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold918 (.A(_0340_),
    .X(net1542));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold919 (.A(net3011),
    .X(net1543));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold92 (.A(net2892),
    .X(net716));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold920 (.A(_0360_),
    .X(net1544));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold921 (.A(net3007),
    .X(net1545));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold922 (.A(_0478_),
    .X(net1546));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold923 (.A(net2927),
    .X(net1547));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold924 (.A(net2929),
    .X(net1548));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold925 (.A(net2970),
    .X(net1549));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold926 (.A(_0350_),
    .X(net1550));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold927 (.A(net2972),
    .X(net1551));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold928 (.A(_0330_),
    .X(net1552));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold929 (.A(net2993),
    .X(net1553));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold93 (.A(_0709_),
    .X(net717));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold930 (.A(_0710_),
    .X(net1554));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold931 (.A(net2949),
    .X(net1555));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold932 (.A(_0195_),
    .X(net1556));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold933 (.A(net3070),
    .X(net1557));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold934 (.A(_0563_),
    .X(net1558));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold935 (.A(net2977),
    .X(net1559));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold936 (.A(_0675_),
    .X(net1560));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold937 (.A(net3052),
    .X(net1561));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold938 (.A(net3054),
    .X(net1562));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold939 (.A(net3057),
    .X(net1563));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold94 (.A(net2708),
    .X(net718));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold940 (.A(net3059),
    .X(net1564));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold941 (.A(net3044),
    .X(net1565));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold942 (.A(_0289_),
    .X(net1566));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold943 (.A(net3030),
    .X(net1567));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold944 (.A(net3032),
    .X(net1568));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold945 (.A(net3013),
    .X(net1569));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold946 (.A(_0190_),
    .X(net1570));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold947 (.A(net2988),
    .X(net1571));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold948 (.A(net2990),
    .X(net1572));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold949 (.A(net3109),
    .X(net1573));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold95 (.A(net2710),
    .X(net719));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold950 (.A(_0438_),
    .X(net1574));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold951 (.A(net3055),
    .X(net1575));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold952 (.A(_0210_),
    .X(net1576));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold953 (.A(net3000),
    .X(net1577));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold954 (.A(_0299_),
    .X(net1578));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold955 (.A(net3132),
    .X(net1579));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold956 (.A(net3134),
    .X(net1580));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold957 (.A(net3038),
    .X(net1581));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold958 (.A(_0319_),
    .X(net1582));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold959 (.A(net3126),
    .X(net1583));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold96 (.A(\gpio_configure[26][4] ),
    .X(net720));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold960 (.A(_0104_),
    .X(net1584));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold961 (.A(net2991),
    .X(net1585));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold962 (.A(_0214_),
    .X(net1586));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold963 (.A(net3113),
    .X(net1587));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold964 (.A(net3115),
    .X(net1588));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold965 (.A(net2953),
    .X(net1589));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold966 (.A(_0558_),
    .X(net1590));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold967 (.A(net3208),
    .X(net1591));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold968 (.A(_0112_),
    .X(net1592));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold969 (.A(net3321),
    .X(net1593));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold97 (.A(net2697),
    .X(net721));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold970 (.A(_0414_),
    .X(net1594));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold971 (.A(net3123),
    .X(net1595));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold972 (.A(net3125),
    .X(net1596));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold973 (.A(net3081),
    .X(net1597));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold974 (.A(_0177_),
    .X(net1598));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold975 (.A(net3036),
    .X(net1599));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold976 (.A(_0294_),
    .X(net1600));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold977 (.A(net3079),
    .X(net1601));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold978 (.A(_0542_),
    .X(net1602));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold979 (.A(net2965),
    .X(net1603));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold98 (.A(net2955),
    .X(net722));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold980 (.A(net2967),
    .X(net1604));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold981 (.A(net3086),
    .X(net1605));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold982 (.A(_0229_),
    .X(net1606));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold983 (.A(net3097),
    .X(net1607));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold984 (.A(_0284_),
    .X(net1608));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold985 (.A(net3020),
    .X(net1609));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold986 (.A(_0566_),
    .X(net1610));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold987 (.A(net3060),
    .X(net1611));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold988 (.A(_0324_),
    .X(net1612));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold989 (.A(net3591),
    .X(net1613));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold99 (.A(_0493_),
    .X(net723));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold990 (.A(net3593),
    .X(net1614));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold991 (.A(net3161),
    .X(net1615));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold992 (.A(_0304_),
    .X(net1616));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold993 (.A(net3040),
    .X(net1617));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold994 (.A(_0309_),
    .X(net1618));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold995 (.A(net3005),
    .X(net1619));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold996 (.A(_0550_),
    .X(net1620));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold997 (.A(net3065),
    .X(net1621));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold998 (.A(_0486_),
    .X(net1622));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold999 (.A(net3027),
    .X(net1623));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(debug_mode),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(mask_rev_in[15]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(wb_adr_i[10]),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 input101 (.A(wb_adr_i[11]),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 input102 (.A(wb_adr_i[12]),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 input103 (.A(wb_adr_i[13]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(wb_adr_i[14]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(wb_adr_i[15]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(wb_adr_i[16]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(wb_adr_i[17]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(wb_adr_i[18]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(wb_adr_i[19]),
    .X(net109));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(mask_rev_in[16]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input110 (.A(wb_adr_i[1]),
    .X(net110));
 sky130_fd_sc_hd__buf_12 input111 (.A(wb_adr_i[20]),
    .X(net111));
 sky130_fd_sc_hd__buf_12 input112 (.A(wb_adr_i[21]),
    .X(net112));
 sky130_fd_sc_hd__buf_8 input113 (.A(wb_adr_i[22]),
    .X(net113));
 sky130_fd_sc_hd__buf_8 input114 (.A(wb_adr_i[23]),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 input115 (.A(wb_adr_i[24]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input116 (.A(wb_adr_i[25]),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(wb_adr_i[26]),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 input118 (.A(wb_adr_i[27]),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 input119 (.A(wb_adr_i[28]),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(mask_rev_in[17]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input120 (.A(wb_adr_i[29]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 input121 (.A(wb_adr_i[2]),
    .X(net121));
 sky130_fd_sc_hd__dlymetal6s2s_1 input122 (.A(wb_adr_i[30]),
    .X(net122));
 sky130_fd_sc_hd__dlymetal6s2s_1 input123 (.A(wb_adr_i[31]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 input124 (.A(wb_adr_i[3]),
    .X(net124));
 sky130_fd_sc_hd__buf_4 input125 (.A(wb_adr_i[4]),
    .X(net125));
 sky130_fd_sc_hd__dlymetal6s2s_1 input126 (.A(wb_adr_i[5]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 input127 (.A(wb_adr_i[6]),
    .X(net127));
 sky130_fd_sc_hd__buf_6 input128 (.A(wb_adr_i[7]),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 input129 (.A(wb_adr_i[8]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(mask_rev_in[18]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(wb_adr_i[9]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(wb_cyc_i),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(wb_dat_i[0]),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 input133 (.A(wb_dat_i[10]),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(wb_dat_i[11]),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 input135 (.A(wb_dat_i[12]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(wb_dat_i[13]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(wb_dat_i[14]),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 input138 (.A(wb_dat_i[15]),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 input139 (.A(wb_dat_i[16]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(mask_rev_in[19]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input140 (.A(wb_dat_i[17]),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 input141 (.A(wb_dat_i[18]),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 input142 (.A(wb_dat_i[19]),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 input143 (.A(wb_dat_i[1]),
    .X(net143));
 sky130_fd_sc_hd__dlymetal6s2s_1 input144 (.A(wb_dat_i[20]),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(wb_dat_i[21]),
    .X(net145));
 sky130_fd_sc_hd__dlymetal6s2s_1 input146 (.A(wb_dat_i[22]),
    .X(net146));
 sky130_fd_sc_hd__dlymetal6s2s_1 input147 (.A(wb_dat_i[23]),
    .X(net147));
 sky130_fd_sc_hd__dlymetal6s2s_1 input148 (.A(wb_dat_i[24]),
    .X(net148));
 sky130_fd_sc_hd__dlymetal6s2s_1 input149 (.A(wb_dat_i[25]),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input15 (.A(mask_rev_in[1]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input150 (.A(wb_dat_i[26]),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 input151 (.A(wb_dat_i[27]),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 input152 (.A(wb_dat_i[28]),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 input153 (.A(wb_dat_i[29]),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 input154 (.A(wb_dat_i[2]),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 input155 (.A(wb_dat_i[30]),
    .X(net155));
 sky130_fd_sc_hd__dlymetal6s2s_1 input156 (.A(wb_dat_i[31]),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 input157 (.A(wb_dat_i[3]),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 input158 (.A(wb_dat_i[4]),
    .X(net158));
 sky130_fd_sc_hd__dlymetal6s2s_1 input159 (.A(wb_dat_i[5]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(mask_rev_in[20]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input160 (.A(wb_dat_i[6]),
    .X(net160));
 sky130_fd_sc_hd__dlymetal6s2s_1 input161 (.A(wb_dat_i[7]),
    .X(net161));
 sky130_fd_sc_hd__dlymetal6s2s_1 input162 (.A(wb_dat_i[8]),
    .X(net162));
 sky130_fd_sc_hd__dlymetal6s2s_1 input163 (.A(wb_dat_i[9]),
    .X(net163));
 sky130_fd_sc_hd__buf_4 input164 (.A(wb_rstn_i),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 input165 (.A(wb_sel_i[0]),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 input166 (.A(wb_sel_i[1]),
    .X(net166));
 sky130_fd_sc_hd__dlymetal6s2s_1 input167 (.A(wb_sel_i[2]),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 input168 (.A(wb_sel_i[3]),
    .X(net168));
 sky130_fd_sc_hd__buf_4 input169 (.A(wb_stb_i),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(mask_rev_in[21]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input170 (.A(wb_we_i),
    .X(net170));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(mask_rev_in[22]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(mask_rev_in[23]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(debug_oeb),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(mask_rev_in[24]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(mask_rev_in[25]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(mask_rev_in[26]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(mask_rev_in[27]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(mask_rev_in[28]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(mask_rev_in[29]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(mask_rev_in[2]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(mask_rev_in[30]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(mask_rev_in[31]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(mask_rev_in[3]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(debug_out),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(mask_rev_in[4]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(mask_rev_in[5]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(mask_rev_in[6]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(mask_rev_in[7]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(mask_rev_in[8]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(mask_rev_in[9]),
    .X(net35));
 sky130_fd_sc_hd__buf_8 input36 (.A(mgmt_gpio_in[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(mgmt_gpio_in[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(mgmt_gpio_in[11]),
    .X(net38));
 sky130_fd_sc_hd__buf_6 input39 (.A(mgmt_gpio_in[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(mask_rev_in[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(mgmt_gpio_in[13]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(mgmt_gpio_in[14]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(mgmt_gpio_in[15]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(mgmt_gpio_in[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mgmt_gpio_in[17]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(mgmt_gpio_in[18]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(mgmt_gpio_in[19]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(mgmt_gpio_in[1]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(mgmt_gpio_in[20]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(mgmt_gpio_in[21]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(mask_rev_in[10]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(mgmt_gpio_in[22]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(mgmt_gpio_in[23]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(mgmt_gpio_in[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(mgmt_gpio_in[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(mgmt_gpio_in[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(mgmt_gpio_in[27]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(mgmt_gpio_in[28]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(mgmt_gpio_in[29]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(mgmt_gpio_in[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(mgmt_gpio_in[30]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(mask_rev_in[11]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input60 (.A(mgmt_gpio_in[31]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(mgmt_gpio_in[32]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(mgmt_gpio_in[33]),
    .X(net62));
 sky130_fd_sc_hd__buf_8 input63 (.A(mgmt_gpio_in[34]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(mgmt_gpio_in[35]),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input65 (.A(mgmt_gpio_in[36]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(mgmt_gpio_in[37]),
    .X(net66));
 sky130_fd_sc_hd__buf_12 input67 (.A(mgmt_gpio_in[3]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(mgmt_gpio_in[5]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(mgmt_gpio_in[6]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(mask_rev_in[12]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input70 (.A(mgmt_gpio_in[7]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(mgmt_gpio_in[8]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(mgmt_gpio_in[9]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(pad_flash_io0_di),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(pad_flash_io1_di),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(porb),
    .X(net75));
 sky130_fd_sc_hd__buf_12 input76 (.A(qspi_enabled),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(ser_tx),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(spi_csb),
    .X(net78));
 sky130_fd_sc_hd__buf_6 input79 (.A(spi_enabled),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(mask_rev_in[13]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(spi_sck),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(spi_sdo),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(spi_sdoenb),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(spimemio_flash_clk),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(spimemio_flash_csb),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(spimemio_flash_io0_do),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input86 (.A(spimemio_flash_io0_oeb),
    .X(net86));
 sky130_fd_sc_hd__buf_4 input87 (.A(spimemio_flash_io1_do),
    .X(net87));
 sky130_fd_sc_hd__buf_4 input88 (.A(spimemio_flash_io1_oeb),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(spimemio_flash_io2_do),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(mask_rev_in[14]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(spimemio_flash_io2_oeb),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(spimemio_flash_io3_do),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 input92 (.A(spimemio_flash_io3_oeb),
    .X(net92));
 sky130_fd_sc_hd__buf_6 input93 (.A(trap),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(uart_enabled),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(usr1_vcc_pwrgood),
    .X(net95));
 sky130_fd_sc_hd__buf_4 input96 (.A(usr1_vdd_pwrgood),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(usr2_vcc_pwrgood),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(usr2_vdd_pwrgood),
    .X(net98));
 sky130_fd_sc_hd__dlymetal6s2s_1 input99 (.A(wb_adr_i[0]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 max_cap351 (.A(_2593_),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 max_cap352 (.A(_2593_),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 max_cap362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 max_cap363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 max_cap395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_6 max_cap399 (.A(_1693_),
    .X(net399));
 sky130_fd_sc_hd__buf_6 max_cap400 (.A(_1681_),
    .X(net400));
 sky130_fd_sc_hd__buf_6 max_cap401 (.A(_1651_),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 max_cap402 (.A(_1645_),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 max_cap404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 max_cap405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_4 max_cap424 (.A(_1880_),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_8 max_cap426 (.A(_1753_),
    .X(net426));
 sky130_fd_sc_hd__buf_6 max_cap428 (.A(_1624_),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 max_cap449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 max_cap450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 max_cap451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_4 max_cap454 (.A(_1747_),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 max_cap455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 max_cap456 (.A(_1725_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 max_cap459 (.A(_1671_),
    .X(net459));
 sky130_fd_sc_hd__buf_6 max_cap460 (.A(_1639_),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 max_cap461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 max_cap464 (.A(_1537_),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 max_cap509 (.A(_0829_),
    .X(net509));
 sky130_fd_sc_hd__buf_8 max_cap530 (.A(_1892_),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_4 max_cap534 (.A(_1860_),
    .X(net534));
 sky130_fd_sc_hd__buf_2 max_cap537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_2 max_cap539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_2 max_cap541 (.A(_1719_),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 max_cap544 (.A(_1708_),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_2 max_cap545 (.A(_1708_),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 max_cap547 (.A(net549),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_2 max_cap548 (.A(_1706_),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_2 max_cap549 (.A(_1706_),
    .X(net549));
 sky130_fd_sc_hd__buf_6 max_cap550 (.A(_1612_),
    .X(net550));
 sky130_fd_sc_hd__buf_12 max_cap551 (.A(_1610_),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 max_cap553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 max_cap554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_2 max_cap555 (.A(_1608_),
    .X(net555));
 sky130_fd_sc_hd__buf_12 max_cap556 (.A(_1600_),
    .X(net556));
 sky130_fd_sc_hd__buf_8 max_cap557 (.A(_1586_),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_14_buff_inst (.A(mgmt_gpio_out_14_prebuff),
    .X(mgmt_gpio_out[14]));
 sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_15_buff_inst (.A(mgmt_gpio_out_15_prebuff),
    .X(mgmt_gpio_out[15]));
 sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_30_buff_inst (.A(mgmt_gpio_out_30_prebuff),
    .X(mgmt_gpio_out[30]));
 sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_31_buff_inst (.A(mgmt_gpio_out_31_prebuff),
    .X(mgmt_gpio_out[31]));
 sky130_fd_sc_hd__clkbuf_8 mgmt_gpio_9_buff_inst (.A(mgmt_gpio_out_9_prebuff),
    .X(mgmt_gpio_out[9]));
 sky130_fd_sc_hd__buf_12 output171 (.A(net171),
    .X(debug_in));
 sky130_fd_sc_hd__buf_12 output172 (.A(net172),
    .X(irq[0]));
 sky130_fd_sc_hd__buf_12 output173 (.A(net173),
    .X(irq[1]));
 sky130_fd_sc_hd__buf_12 output174 (.A(net174),
    .X(irq[2]));
 sky130_fd_sc_hd__buf_12 output175 (.A(net175),
    .X(mgmt_gpio_oeb[0]));
 sky130_fd_sc_hd__buf_12 output176 (.A(net176),
    .X(mgmt_gpio_oeb[10]));
 sky130_fd_sc_hd__buf_12 output177 (.A(net177),
    .X(mgmt_gpio_oeb[11]));
 sky130_fd_sc_hd__buf_12 output178 (.A(net178),
    .X(mgmt_gpio_oeb[12]));
 sky130_fd_sc_hd__buf_12 output179 (.A(net179),
    .X(mgmt_gpio_oeb[13]));
 sky130_fd_sc_hd__buf_12 output180 (.A(net180),
    .X(mgmt_gpio_oeb[14]));
 sky130_fd_sc_hd__buf_12 output181 (.A(net181),
    .X(mgmt_gpio_oeb[15]));
 sky130_fd_sc_hd__buf_12 output182 (.A(net182),
    .X(mgmt_gpio_oeb[16]));
 sky130_fd_sc_hd__buf_12 output183 (.A(net183),
    .X(mgmt_gpio_oeb[17]));
 sky130_fd_sc_hd__buf_12 output184 (.A(net184),
    .X(mgmt_gpio_oeb[18]));
 sky130_fd_sc_hd__buf_12 output185 (.A(net185),
    .X(mgmt_gpio_oeb[19]));
 sky130_fd_sc_hd__buf_12 output186 (.A(net186),
    .X(mgmt_gpio_oeb[1]));
 sky130_fd_sc_hd__buf_12 output187 (.A(net187),
    .X(mgmt_gpio_oeb[20]));
 sky130_fd_sc_hd__buf_12 output188 (.A(net188),
    .X(mgmt_gpio_oeb[21]));
 sky130_fd_sc_hd__buf_12 output189 (.A(net189),
    .X(mgmt_gpio_oeb[22]));
 sky130_fd_sc_hd__buf_12 output190 (.A(net190),
    .X(mgmt_gpio_oeb[23]));
 sky130_fd_sc_hd__buf_12 output191 (.A(net191),
    .X(mgmt_gpio_oeb[24]));
 sky130_fd_sc_hd__buf_12 output192 (.A(net192),
    .X(mgmt_gpio_oeb[25]));
 sky130_fd_sc_hd__buf_12 output193 (.A(net193),
    .X(mgmt_gpio_oeb[26]));
 sky130_fd_sc_hd__buf_12 output194 (.A(net194),
    .X(mgmt_gpio_oeb[27]));
 sky130_fd_sc_hd__buf_12 output195 (.A(net195),
    .X(mgmt_gpio_oeb[28]));
 sky130_fd_sc_hd__buf_12 output196 (.A(net196),
    .X(mgmt_gpio_oeb[29]));
 sky130_fd_sc_hd__buf_12 output197 (.A(net197),
    .X(mgmt_gpio_oeb[2]));
 sky130_fd_sc_hd__buf_12 output198 (.A(net198),
    .X(mgmt_gpio_oeb[30]));
 sky130_fd_sc_hd__buf_12 output199 (.A(net199),
    .X(mgmt_gpio_oeb[31]));
 sky130_fd_sc_hd__buf_12 output200 (.A(net200),
    .X(mgmt_gpio_oeb[32]));
 sky130_fd_sc_hd__buf_12 output201 (.A(net201),
    .X(mgmt_gpio_oeb[33]));
 sky130_fd_sc_hd__buf_12 output202 (.A(net202),
    .X(mgmt_gpio_oeb[34]));
 sky130_fd_sc_hd__buf_12 output203 (.A(net365),
    .X(mgmt_gpio_oeb[35]));
 sky130_fd_sc_hd__buf_12 output204 (.A(net204),
    .X(mgmt_gpio_oeb[36]));
 sky130_fd_sc_hd__buf_12 output205 (.A(net205),
    .X(mgmt_gpio_oeb[37]));
 sky130_fd_sc_hd__buf_12 output206 (.A(net206),
    .X(mgmt_gpio_oeb[3]));
 sky130_fd_sc_hd__buf_12 output207 (.A(net207),
    .X(mgmt_gpio_oeb[4]));
 sky130_fd_sc_hd__buf_12 output208 (.A(net208),
    .X(mgmt_gpio_oeb[5]));
 sky130_fd_sc_hd__buf_12 output209 (.A(net209),
    .X(mgmt_gpio_oeb[6]));
 sky130_fd_sc_hd__buf_12 output210 (.A(net210),
    .X(mgmt_gpio_oeb[7]));
 sky130_fd_sc_hd__buf_12 output211 (.A(net211),
    .X(mgmt_gpio_oeb[8]));
 sky130_fd_sc_hd__buf_12 output212 (.A(net212),
    .X(mgmt_gpio_oeb[9]));
 sky130_fd_sc_hd__buf_12 output213 (.A(net213),
    .X(mgmt_gpio_out[0]));
 sky130_fd_sc_hd__buf_12 output214 (.A(net214),
    .X(mgmt_gpio_out[10]));
 sky130_fd_sc_hd__buf_12 output215 (.A(net215),
    .X(mgmt_gpio_out[11]));
 sky130_fd_sc_hd__buf_12 output216 (.A(net216),
    .X(mgmt_gpio_out[12]));
 sky130_fd_sc_hd__buf_12 output217 (.A(net217),
    .X(mgmt_gpio_out[13]));
 sky130_fd_sc_hd__buf_12 output218 (.A(net218),
    .X(mgmt_gpio_out[16]));
 sky130_fd_sc_hd__buf_12 output219 (.A(net219),
    .X(mgmt_gpio_out[17]));
 sky130_fd_sc_hd__buf_12 output220 (.A(net220),
    .X(mgmt_gpio_out[18]));
 sky130_fd_sc_hd__buf_12 output221 (.A(net221),
    .X(mgmt_gpio_out[19]));
 sky130_fd_sc_hd__buf_12 output222 (.A(net222),
    .X(mgmt_gpio_out[1]));
 sky130_fd_sc_hd__buf_12 output223 (.A(net223),
    .X(mgmt_gpio_out[20]));
 sky130_fd_sc_hd__buf_12 output224 (.A(net224),
    .X(mgmt_gpio_out[21]));
 sky130_fd_sc_hd__buf_12 output225 (.A(net225),
    .X(mgmt_gpio_out[22]));
 sky130_fd_sc_hd__buf_12 output226 (.A(net226),
    .X(mgmt_gpio_out[23]));
 sky130_fd_sc_hd__buf_12 output227 (.A(net227),
    .X(mgmt_gpio_out[24]));
 sky130_fd_sc_hd__buf_12 output228 (.A(net228),
    .X(mgmt_gpio_out[25]));
 sky130_fd_sc_hd__buf_12 output229 (.A(net229),
    .X(mgmt_gpio_out[26]));
 sky130_fd_sc_hd__buf_12 output230 (.A(net230),
    .X(mgmt_gpio_out[27]));
 sky130_fd_sc_hd__buf_12 output231 (.A(net231),
    .X(mgmt_gpio_out[28]));
 sky130_fd_sc_hd__buf_12 output232 (.A(net232),
    .X(mgmt_gpio_out[29]));
 sky130_fd_sc_hd__buf_12 output233 (.A(net233),
    .X(mgmt_gpio_out[2]));
 sky130_fd_sc_hd__buf_12 output234 (.A(net234),
    .X(mgmt_gpio_out[32]));
 sky130_fd_sc_hd__buf_12 output235 (.A(net235),
    .X(mgmt_gpio_out[33]));
 sky130_fd_sc_hd__buf_12 output236 (.A(net236),
    .X(mgmt_gpio_out[34]));
 sky130_fd_sc_hd__buf_12 output237 (.A(net237),
    .X(mgmt_gpio_out[35]));
 sky130_fd_sc_hd__buf_12 output238 (.A(net238),
    .X(mgmt_gpio_out[36]));
 sky130_fd_sc_hd__buf_12 output239 (.A(net239),
    .X(mgmt_gpio_out[37]));
 sky130_fd_sc_hd__buf_12 output240 (.A(net240),
    .X(mgmt_gpio_out[3]));
 sky130_fd_sc_hd__buf_12 output241 (.A(net241),
    .X(mgmt_gpio_out[4]));
 sky130_fd_sc_hd__buf_12 output242 (.A(net242),
    .X(mgmt_gpio_out[5]));
 sky130_fd_sc_hd__buf_12 output243 (.A(net243),
    .X(mgmt_gpio_out[6]));
 sky130_fd_sc_hd__buf_12 output244 (.A(net244),
    .X(mgmt_gpio_out[7]));
 sky130_fd_sc_hd__buf_12 output245 (.A(net245),
    .X(mgmt_gpio_out[8]));
 sky130_fd_sc_hd__buf_12 output246 (.A(net246),
    .X(pad_flash_clk_oeb));
 sky130_fd_sc_hd__buf_12 output247 (.A(net247),
    .X(pad_flash_csb));
 sky130_fd_sc_hd__buf_12 output248 (.A(net248),
    .X(pad_flash_csb_oeb));
 sky130_fd_sc_hd__buf_12 output249 (.A(net249),
    .X(pad_flash_io0_do));
 sky130_fd_sc_hd__buf_12 output250 (.A(net250),
    .X(pad_flash_io0_ieb));
 sky130_fd_sc_hd__buf_12 output251 (.A(net251),
    .X(pad_flash_io0_oeb));
 sky130_fd_sc_hd__buf_12 output252 (.A(net252),
    .X(pad_flash_io1_do));
 sky130_fd_sc_hd__buf_12 output253 (.A(net253),
    .X(pad_flash_io1_ieb));
 sky130_fd_sc_hd__buf_12 output254 (.A(net254),
    .X(pad_flash_io1_oeb));
 sky130_fd_sc_hd__buf_12 output255 (.A(net255),
    .X(pll90_sel[0]));
 sky130_fd_sc_hd__buf_12 output256 (.A(net256),
    .X(pll90_sel[1]));
 sky130_fd_sc_hd__buf_12 output257 (.A(net257),
    .X(pll90_sel[2]));
 sky130_fd_sc_hd__buf_12 output258 (.A(net258),
    .X(pll_bypass));
 sky130_fd_sc_hd__buf_12 output259 (.A(net259),
    .X(pll_dco_ena));
 sky130_fd_sc_hd__buf_12 output260 (.A(net260),
    .X(pll_div[0]));
 sky130_fd_sc_hd__buf_12 output261 (.A(net261),
    .X(pll_div[1]));
 sky130_fd_sc_hd__buf_12 output262 (.A(net262),
    .X(pll_div[2]));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(pll_div[3]));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(pll_div[4]));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(pll_ena));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(pll_sel[0]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(pll_sel[1]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(pll_sel[2]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(pll_trim[0]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(pll_trim[10]));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(pll_trim[11]));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(pll_trim[12]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(pll_trim[13]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(pll_trim[14]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(pll_trim[15]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(pll_trim[16]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(pll_trim[17]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(pll_trim[18]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(pll_trim[19]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(pll_trim[1]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(pll_trim[20]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(pll_trim[21]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(pll_trim[22]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(pll_trim[23]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(pll_trim[24]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(pll_trim[25]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(pll_trim[2]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(pll_trim[3]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(pll_trim[4]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(pll_trim[5]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(pll_trim[6]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(pll_trim[7]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(pll_trim[8]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(pll_trim[9]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(pwr_ctrl_out[0]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(pwr_ctrl_out[1]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(pwr_ctrl_out[2]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(pwr_ctrl_out[3]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(reset));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(ser_rx));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(serial_clock));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(serial_data_1));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(serial_data_2));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(serial_load));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(serial_resetn));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(spi_sdi));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(spimemio_flash_io0_di));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(spimemio_flash_io1_di));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(spimemio_flash_io2_di));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(spimemio_flash_io3_di));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_6 output312 (.A(net3444),
    .X(net1792));
 sky130_fd_sc_hd__buf_6 output313 (.A(net3441),
    .X(net1814));
 sky130_fd_sc_hd__buf_6 output314 (.A(net1807),
    .X(net1808));
 sky130_fd_sc_hd__buf_6 output315 (.A(net1829),
    .X(net1830));
 sky130_fd_sc_hd__buf_6 output316 (.A(net1811),
    .X(net1812));
 sky130_fd_sc_hd__buf_6 output317 (.A(net1809),
    .X(net1810));
 sky130_fd_sc_hd__buf_6 output318 (.A(net1817),
    .X(net1818));
 sky130_fd_sc_hd__buf_6 output319 (.A(net1827),
    .X(net1828));
 sky130_fd_sc_hd__buf_6 output320 (.A(net3407),
    .X(net1794));
 sky130_fd_sc_hd__buf_6 output321 (.A(net3415),
    .X(net1800));
 sky130_fd_sc_hd__buf_6 output322 (.A(net1801),
    .X(net1802));
 sky130_fd_sc_hd__buf_6 output323 (.A(net3421),
    .X(net1784));
 sky130_fd_sc_hd__buf_6 output324 (.A(net1833),
    .X(net1834));
 sky130_fd_sc_hd__buf_6 output325 (.A(net1779),
    .X(net1780));
 sky130_fd_sc_hd__buf_6 output326 (.A(net3388),
    .X(net1778));
 sky130_fd_sc_hd__buf_6 output327 (.A(net3434),
    .X(net1776));
 sky130_fd_sc_hd__buf_6 output328 (.A(net1821),
    .X(net1822));
 sky130_fd_sc_hd__buf_6 output329 (.A(net1837),
    .X(net1838));
 sky130_fd_sc_hd__buf_6 output330 (.A(net1815),
    .X(net1816));
 sky130_fd_sc_hd__buf_6 output331 (.A(net1835),
    .X(net1836));
 sky130_fd_sc_hd__buf_6 output332 (.A(net1839),
    .X(net1840));
 sky130_fd_sc_hd__buf_6 output333 (.A(net1805),
    .X(net1806));
 sky130_fd_sc_hd__buf_6 output334 (.A(net3412),
    .X(net1790));
 sky130_fd_sc_hd__buf_6 output335 (.A(net1831),
    .X(net1832));
 sky130_fd_sc_hd__buf_6 output336 (.A(net1825),
    .X(net1826));
 sky130_fd_sc_hd__buf_6 output337 (.A(net3475),
    .X(net1782));
 sky130_fd_sc_hd__buf_6 output338 (.A(net1819),
    .X(net1820));
 sky130_fd_sc_hd__buf_6 output339 (.A(net3431),
    .X(net1788));
 sky130_fd_sc_hd__buf_6 output340 (.A(net3393),
    .X(net1786));
 sky130_fd_sc_hd__buf_6 output341 (.A(net1803),
    .X(net1804));
 sky130_fd_sc_hd__buf_6 output342 (.A(net1823),
    .X(net1824));
 sky130_fd_sc_hd__buf_6 output343 (.A(net3426),
    .X(net1798));
 sky130_fd_sc_hd__clkbuf_8 pad_flashh_clk_buff_inst (.A(pad_flash_clk_prebuff),
    .X(pad_flash_clk));
 sky130_fd_sc_hd__clkbuf_2 wire344 (.A(_1263_),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 wire345 (.A(_1220_),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 wire346 (.A(_3322_),
    .X(net346));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire347 (.A(_3240_),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 wire348 (.A(_3040_),
    .X(net348));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire349 (.A(_2731_),
    .X(net349));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire350 (.A(_2715_),
    .X(net350));
 sky130_fd_sc_hd__buf_2 wire364 (.A(_1598_),
    .X(net364));
 sky130_fd_sc_hd__buf_6 wire365 (.A(net203),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 wire393 (.A(_3011_),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 wire396 (.A(_1698_),
    .X(net396));
 sky130_fd_sc_hd__buf_2 wire406 (.A(_0888_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 wire427 (.A(_1636_),
    .X(net427));
 sky130_fd_sc_hd__buf_6 wire429 (.A(_1618_),
    .X(net429));
 sky130_fd_sc_hd__buf_2 wire452 (.A(_1829_),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 wire453 (.A(_1747_),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 wire462 (.A(_1538_),
    .X(net462));
 sky130_fd_sc_hd__buf_4 wire463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_6 wire507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_4 wire508 (.A(_1412_),
    .X(net508));
 sky130_fd_sc_hd__buf_2 wire529 (.A(_2075_),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_4 wire533 (.A(_1860_),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_4 wire536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_2 wire538 (.A(_1835_),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 wire540 (.A(_1719_),
    .X(net540));
 sky130_fd_sc_hd__buf_2 wire546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_4 wire559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 wire560 (.A(_1564_),
    .X(net560));
endmodule

