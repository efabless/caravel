magic
tech sky130A
magscale 1 2
timestamp 1636973449
<< nwell >>
rect -38 261 20002 827
<< pwell >>
rect 29 -17 63 17
rect 305 -17 339 17
rect 1409 -17 1443 17
rect 2512 -11 2536 11
rect 2697 -17 2731 17
rect 3801 -17 3835 17
rect 4905 -17 4939 17
rect 5273 -17 5307 17
rect 6377 -17 6411 17
rect 7481 -17 7515 17
rect 7849 -17 7883 17
rect 8953 -17 8987 17
rect 10057 -17 10091 17
rect 10425 -17 10459 17
rect 11529 -17 11563 17
rect 12633 -17 12667 17
rect 13001 -17 13035 17
rect 14105 -17 14139 17
rect 15209 -17 15243 17
rect 15577 -17 15611 17
rect 16681 -17 16715 17
rect 17785 -17 17819 17
rect 18153 -17 18187 17
rect 19257 -17 19291 17
rect 19624 -11 19648 11
rect 19901 -17 19935 17
<< obsli1 >>
rect 0 -17 19964 1105
<< obsm1 >>
rect 0 -48 19964 1136
<< metal2 >>
rect 170 -48 230 1136
rect 4170 -48 4230 1136
rect 8170 -48 8230 1136
rect 12170 -48 12230 1136
rect 16170 -48 16230 1136
<< obsm2 >>
rect 8482 711 8538 814
<< metal3 >>
rect 0 882 19964 982
rect 0 688 800 808
rect 0 302 19964 402
<< obsm3 >>
rect 880 715 8543 781
<< labels >>
rlabel metal3 s 0 688 800 808 6 HI
port 1 nsew signal output
rlabel metal3 s 0 302 19964 402 6 vccd2
port 2 nsew power input
rlabel metal2 s 170 -48 230 1136 6 vccd2
port 2 nsew power input
rlabel metal2 s 8170 -48 8230 1136 6 vccd2
port 2 nsew power input
rlabel metal2 s 16170 -48 16230 1136 6 vccd2
port 2 nsew power input
rlabel metal3 s 0 882 19964 982 6 vssd2
port 3 nsew ground input
rlabel metal2 s 4170 -48 4230 1136 6 vssd2
port 3 nsew ground input
rlabel metal2 s 12170 -48 12230 1136 6 vssd2
port 3 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 20000 1400
string LEFview TRUE
string GDS_FILE ../gds/mprj2_logic_high.gds
string GDS_END 27684
string GDS_START 19178
<< end >>

