magic
tech sky130A
magscale 1 2
timestamp 1637551221
<< viali >>
rect 2237 3145 2271 3179
rect 2697 3145 2731 3179
rect 3525 3145 3559 3179
rect 4445 3145 4479 3179
rect 5089 3145 5123 3179
rect 5365 3145 5399 3179
rect 5641 3145 5675 3179
rect 6009 3145 6043 3179
rect 6561 3145 6595 3179
rect 6837 3145 6871 3179
rect 7113 3145 7147 3179
rect 7389 3145 7423 3179
rect 7665 3145 7699 3179
rect 7941 3145 7975 3179
rect 8217 3145 8251 3179
rect 8493 3145 8527 3179
rect 8769 3145 8803 3179
rect 9137 3145 9171 3179
rect 9689 3145 9723 3179
rect 9965 3145 9999 3179
rect 10793 3145 10827 3179
rect 11345 3145 11379 3179
rect 12173 3145 12207 3179
rect 12725 3145 12759 3179
rect 13277 3145 13311 3179
rect 13553 3145 13587 3179
rect 13829 3145 13863 3179
rect 14381 3145 14415 3179
rect 15209 3145 15243 3179
rect 15761 3145 15795 3179
rect 16865 3145 16899 3179
rect 17693 3145 17727 3179
rect 18521 3145 18555 3179
rect 19441 3145 19475 3179
rect 20269 3145 20303 3179
rect 21373 3145 21407 3179
rect 22569 3145 22603 3179
rect 23673 3145 23707 3179
rect 24869 3145 24903 3179
rect 26249 3145 26283 3179
rect 27445 3145 27479 3179
rect 28549 3145 28583 3179
rect 29745 3145 29779 3179
rect 30849 3145 30883 3179
rect 31953 3145 31987 3179
rect 32873 3145 32907 3179
rect 33977 3145 34011 3179
rect 35173 3145 35207 3179
rect 36553 3145 36587 3179
rect 37749 3145 37783 3179
rect 38853 3145 38887 3179
rect 40049 3145 40083 3179
rect 41153 3145 41187 3179
rect 42625 3145 42659 3179
rect 43453 3145 43487 3179
rect 44281 3145 44315 3179
rect 45201 3145 45235 3179
rect 47777 3145 47811 3179
rect 48697 3145 48731 3179
rect 48973 3145 49007 3179
rect 49249 3145 49283 3179
rect 49525 3145 49559 3179
rect 49801 3145 49835 3179
rect 50353 3145 50387 3179
rect 50905 3145 50939 3179
rect 51181 3145 51215 3179
rect 51733 3145 51767 3179
rect 52285 3145 52319 3179
rect 52561 3145 52595 3179
rect 53205 3145 53239 3179
rect 53757 3145 53791 3179
rect 54033 3145 54067 3179
rect 54585 3145 54619 3179
rect 55137 3145 55171 3179
rect 55781 3145 55815 3179
rect 56609 3145 56643 3179
rect 57161 3145 57195 3179
rect 58081 3145 58115 3179
rect 58909 3145 58943 3179
rect 59737 3145 59771 3179
rect 60657 3145 60691 3179
rect 61209 3145 61243 3179
rect 62037 3145 62071 3179
rect 62589 3145 62623 3179
rect 63509 3145 63543 3179
rect 65165 3145 65199 3179
rect 66361 3145 66395 3179
rect 66637 3145 66671 3179
rect 67097 3145 67131 3179
rect 67373 3145 67407 3179
rect 67649 3145 67683 3179
rect 2973 3077 3007 3111
rect 17141 3077 17175 3111
rect 17969 3077 18003 3111
rect 19073 3077 19107 3111
rect 19993 3077 20027 3111
rect 21097 3077 21131 3111
rect 22293 3077 22327 3111
rect 23397 3077 23431 3111
rect 24225 3077 24259 3111
rect 25421 3077 25455 3111
rect 27169 3077 27203 3111
rect 28273 3077 28307 3111
rect 30021 3077 30055 3111
rect 31125 3077 31159 3111
rect 32321 3077 32355 3111
rect 33425 3077 33459 3111
rect 34529 3077 34563 3111
rect 36001 3077 36035 3111
rect 37473 3077 37507 3111
rect 38577 3077 38611 3111
rect 39681 3077 39715 3111
rect 40877 3077 40911 3111
rect 42901 3077 42935 3111
rect 44005 3077 44039 3111
rect 45477 3077 45511 3111
rect 50629 3077 50663 3111
rect 52009 3077 52043 3111
rect 53481 3077 53515 3111
rect 54309 3077 54343 3111
rect 54861 3077 54895 3111
rect 55505 3077 55539 3111
rect 57437 3077 57471 3111
rect 58357 3077 58391 3111
rect 59185 3077 59219 3111
rect 60013 3077 60047 3111
rect 60933 3077 60967 3111
rect 61761 3077 61795 3111
rect 62865 3077 62899 3111
rect 63785 3077 63819 3111
rect 64889 3077 64923 3111
rect 66085 3077 66119 3111
rect 3065 3009 3099 3043
rect 9413 3009 9447 3043
rect 10517 3009 10551 3043
rect 11069 3009 11103 3043
rect 11713 3009 11747 3043
rect 12449 3009 12483 3043
rect 13001 3009 13035 3043
rect 14933 3009 14967 3043
rect 15485 3009 15519 3043
rect 16037 3009 16071 3043
rect 17417 3009 17451 3043
rect 18245 3009 18279 3043
rect 19717 3009 19751 3043
rect 20821 3009 20855 3043
rect 22017 3009 22051 3043
rect 22845 3009 22879 3043
rect 23949 3009 23983 3043
rect 25145 3009 25179 3043
rect 26525 3009 26559 3043
rect 27721 3009 27755 3043
rect 28825 3009 28859 3043
rect 30297 3009 30331 3043
rect 31401 3009 31435 3043
rect 32597 3009 32631 3043
rect 33701 3009 33735 3043
rect 34897 3009 34931 3043
rect 36277 3009 36311 3043
rect 36829 3009 36863 3043
rect 38025 3009 38059 3043
rect 39129 3009 39163 3043
rect 40325 3009 40359 3043
rect 41429 3009 41463 3043
rect 42257 3009 42291 3043
rect 43177 3009 43211 3043
rect 44557 3009 44591 3043
rect 45753 3009 45787 3043
rect 48053 3009 48087 3043
rect 51457 3009 51491 3043
rect 52929 3009 52963 3043
rect 56333 3009 56367 3043
rect 56885 3009 56919 3043
rect 57713 3009 57747 3043
rect 58633 3009 58667 3043
rect 59461 3009 59495 3043
rect 60289 3009 60323 3043
rect 61485 3009 61519 3043
rect 62313 3009 62347 3043
rect 63233 3009 63267 3043
rect 64337 3009 64371 3043
rect 65441 3009 65475 3043
rect 65993 3009 66027 3043
rect 3617 2941 3651 2975
rect 4169 2941 4203 2975
rect 4721 2941 4755 2975
rect 10241 2941 10275 2975
rect 14657 2941 14691 2975
rect 16313 2941 16347 2975
rect 18797 2941 18831 2975
rect 20545 2941 20579 2975
rect 21649 2941 21683 2975
rect 23121 2941 23155 2975
rect 24593 2941 24627 2975
rect 25697 2941 25731 2975
rect 25973 2941 26007 2975
rect 26801 2941 26835 2975
rect 27997 2941 28031 2975
rect 29101 2941 29135 2975
rect 29377 2941 29411 2975
rect 30573 2941 30607 2975
rect 31677 2941 31711 2975
rect 33149 2941 33183 2975
rect 34253 2941 34287 2975
rect 35449 2941 35483 2975
rect 35725 2941 35759 2975
rect 37105 2941 37139 2975
rect 38301 2941 38335 2975
rect 39405 2941 39439 2975
rect 40601 2941 40635 2975
rect 41705 2941 41739 2975
rect 41981 2941 42015 2975
rect 43729 2941 43763 2975
rect 44833 2941 44867 2975
rect 56057 2941 56091 2975
rect 64061 2941 64095 2975
rect 64613 2941 64647 2975
rect 2789 2465 2823 2499
rect 3525 2465 3559 2499
rect 4169 2465 4203 2499
rect 5273 2465 5307 2499
rect 6285 2465 6319 2499
rect 11897 2465 11931 2499
rect 28825 2465 28859 2499
rect 36553 2465 36587 2499
rect 41705 2465 41739 2499
rect 44281 2465 44315 2499
rect 45293 2465 45327 2499
rect 45569 2465 45603 2499
rect 45845 2465 45879 2499
rect 46121 2465 46155 2499
rect 46397 2465 46431 2499
rect 46673 2465 46707 2499
rect 46949 2465 46983 2499
rect 47225 2465 47259 2499
rect 48053 2465 48087 2499
rect 48329 2465 48363 2499
rect 64981 2465 65015 2499
rect 65441 2465 65475 2499
rect 65993 2465 66027 2499
rect 66269 2465 66303 2499
rect 66545 2465 66579 2499
rect 3065 2397 3099 2431
rect 5549 2397 5583 2431
rect 6561 2397 6595 2431
rect 4445 2329 4479 2363
rect 4997 2329 5031 2363
rect 2513 2261 2547 2295
rect 3617 2261 3651 2295
rect 4721 2261 4755 2295
rect 5825 2261 5859 2295
rect 2145 2057 2179 2091
rect 3893 2057 3927 2091
rect 4169 2057 4203 2091
rect 6561 2057 6595 2091
rect 6837 2057 6871 2091
rect 4445 1989 4479 2023
rect 5825 1989 5859 2023
rect 2237 1921 2271 1955
rect 4721 1921 4755 1955
rect 6101 1921 6135 1955
rect 46121 1921 46155 1955
rect 2697 1853 2731 1887
rect 2789 1853 2823 1887
rect 3065 1853 3099 1887
rect 3341 1853 3375 1887
rect 3617 1853 3651 1887
rect 4997 1853 5031 1887
rect 5273 1853 5307 1887
rect 5549 1853 5583 1887
rect 7297 1853 7331 1887
rect 9873 1853 9907 1887
rect 12173 1853 12207 1887
rect 14105 1853 14139 1887
rect 16865 1853 16899 1887
rect 20269 1853 20303 1887
rect 22201 1853 22235 1887
rect 25053 1853 25087 1887
rect 29285 1853 29319 1887
rect 31493 1853 31527 1887
rect 32597 1853 32631 1887
rect 44373 1853 44407 1887
rect 45569 1853 45603 1887
rect 52285 1853 52319 1887
rect 27813 1377 27847 1411
rect 40417 1377 40451 1411
rect 46949 1377 46983 1411
rect 52285 1377 52319 1411
rect 2145 1309 2179 1343
rect 3065 1309 3099 1343
rect 4721 1309 4755 1343
rect 5549 1309 5583 1343
rect 5825 1309 5859 1343
rect 7205 1309 7239 1343
rect 7849 1309 7883 1343
rect 10149 1309 10183 1343
rect 11989 1309 12023 1343
rect 13553 1309 13587 1343
rect 14381 1309 14415 1343
rect 16313 1309 16347 1343
rect 17509 1309 17543 1343
rect 18337 1309 18371 1343
rect 19993 1309 20027 1343
rect 20821 1309 20855 1343
rect 21649 1309 21683 1343
rect 23029 1309 23063 1343
rect 24225 1309 24259 1343
rect 25605 1309 25639 1343
rect 26709 1309 26743 1343
rect 28089 1309 28123 1343
rect 29193 1309 29227 1343
rect 30389 1309 30423 1343
rect 31769 1309 31803 1343
rect 33149 1309 33183 1343
rect 33977 1309 34011 1343
rect 34897 1309 34931 1343
rect 35449 1309 35483 1343
rect 36553 1309 36587 1343
rect 37473 1309 37507 1343
rect 38301 1309 38335 1343
rect 39129 1309 39163 1343
rect 40693 1309 40727 1343
rect 41797 1309 41831 1343
rect 42901 1309 42935 1343
rect 44373 1309 44407 1343
rect 45201 1309 45235 1343
rect 46397 1309 46431 1343
rect 47777 1309 47811 1343
rect 48605 1309 48639 1343
rect 49709 1309 49743 1343
rect 50353 1309 50387 1343
rect 51181 1309 51215 1343
rect 52929 1309 52963 1343
rect 54033 1309 54067 1343
rect 55781 1309 55815 1343
rect 2513 1241 2547 1275
rect 4445 1241 4479 1275
rect 6101 1241 6135 1275
rect 6929 1241 6963 1275
rect 8125 1241 8159 1275
rect 8769 1241 8803 1275
rect 9413 1241 9447 1275
rect 10701 1241 10735 1275
rect 11253 1241 11287 1275
rect 12449 1241 12483 1275
rect 13277 1241 13311 1275
rect 14657 1241 14691 1275
rect 15209 1241 15243 1275
rect 17233 1241 17267 1275
rect 18613 1241 18647 1275
rect 19717 1241 19751 1275
rect 20545 1241 20579 1275
rect 21373 1241 21407 1275
rect 22477 1241 22511 1275
rect 23581 1241 23615 1275
rect 24593 1241 24627 1275
rect 25329 1241 25363 1275
rect 26433 1241 26467 1275
rect 27537 1241 27571 1275
rect 28917 1241 28951 1275
rect 29837 1241 29871 1275
rect 30665 1241 30699 1275
rect 31217 1241 31251 1275
rect 32873 1241 32907 1275
rect 33701 1241 33735 1275
rect 34529 1241 34563 1275
rect 36277 1241 36311 1275
rect 37105 1241 37139 1275
rect 38025 1241 38059 1275
rect 38853 1241 38887 1275
rect 40141 1241 40175 1275
rect 40969 1241 41003 1275
rect 41521 1241 41555 1275
rect 43545 1241 43579 1275
rect 45845 1241 45879 1275
rect 46673 1241 46707 1275
rect 47225 1241 47259 1275
rect 48329 1241 48363 1275
rect 49433 1241 49467 1275
rect 50629 1241 50663 1275
rect 52561 1241 52595 1275
rect 53481 1241 53515 1275
rect 54309 1241 54343 1275
rect 54861 1241 54895 1275
rect 56057 1241 56091 1275
rect 1869 1173 1903 1207
rect 2421 1173 2455 1207
rect 2789 1173 2823 1207
rect 3341 1173 3375 1207
rect 3617 1173 3651 1207
rect 4169 1173 4203 1207
rect 4997 1173 5031 1207
rect 5273 1173 5307 1207
rect 6653 1173 6687 1207
rect 7573 1173 7607 1207
rect 8493 1173 8527 1207
rect 9137 1173 9171 1207
rect 9689 1173 9723 1207
rect 10425 1173 10459 1207
rect 10977 1173 11011 1207
rect 11713 1173 11747 1207
rect 12725 1173 12759 1207
rect 13001 1173 13035 1207
rect 13829 1173 13863 1207
rect 14933 1173 14967 1207
rect 15485 1173 15519 1207
rect 15761 1173 15795 1207
rect 16037 1173 16071 1207
rect 16865 1173 16899 1207
rect 17785 1173 17819 1207
rect 18061 1173 18095 1207
rect 18889 1173 18923 1207
rect 19441 1173 19475 1207
rect 20269 1173 20303 1207
rect 21097 1173 21131 1207
rect 22017 1173 22051 1207
rect 22753 1173 22787 1207
rect 23305 1173 23339 1207
rect 23949 1173 23983 1207
rect 24869 1173 24903 1207
rect 25881 1173 25915 1207
rect 26157 1173 26191 1207
rect 27169 1173 27203 1207
rect 28365 1173 28399 1207
rect 28641 1173 28675 1207
rect 30113 1173 30147 1207
rect 30941 1173 30975 1207
rect 31493 1173 31527 1207
rect 32321 1173 32355 1207
rect 32597 1173 32631 1207
rect 33425 1173 33459 1207
rect 34253 1173 34287 1207
rect 35173 1173 35207 1207
rect 35725 1173 35759 1207
rect 36001 1173 36035 1207
rect 36829 1173 36863 1207
rect 37749 1173 37783 1207
rect 38577 1173 38611 1207
rect 39405 1173 39439 1207
rect 39681 1173 39715 1207
rect 41245 1173 41279 1207
rect 42073 1173 42107 1207
rect 42625 1173 42659 1207
rect 43177 1173 43211 1207
rect 43821 1173 43855 1207
rect 44097 1173 44131 1207
rect 44649 1173 44683 1207
rect 45477 1173 45511 1207
rect 46121 1173 46155 1207
rect 48053 1173 48087 1207
rect 48881 1173 48915 1207
rect 49157 1173 49191 1207
rect 49985 1173 50019 1207
rect 50905 1173 50939 1207
rect 51457 1173 51491 1207
rect 51733 1173 51767 1207
rect 52009 1173 52043 1207
rect 53205 1173 53239 1207
rect 53757 1173 53791 1207
rect 54585 1173 54619 1207
rect 55137 1173 55171 1207
rect 55505 1173 55539 1207
rect 56333 1173 56367 1207
<< metal1 >>
rect 658 3408 664 3460
rect 716 3448 722 3460
rect 6822 3448 6828 3460
rect 716 3420 6828 3448
rect 716 3408 722 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 5902 3380 5908 3392
rect 1728 3352 5908 3380
rect 1728 3340 1734 3352
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 25866 3380 25872 3392
rect 24912 3352 25872 3380
rect 24912 3340 24918 3352
rect 25866 3340 25872 3352
rect 25924 3340 25930 3392
rect 1288 3290 68816 3312
rect 1288 3238 13262 3290
rect 13314 3238 25262 3290
rect 25314 3238 37262 3290
rect 37314 3238 49262 3290
rect 49314 3238 61262 3290
rect 61314 3238 68816 3290
rect 1288 3216 68816 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 1452 3148 2237 3176
rect 1452 3136 1458 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 3326 3176 3332 3188
rect 2731 3148 3332 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 3602 3176 3608 3188
rect 3559 3148 3608 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4120 3148 4445 3176
rect 4120 3136 4126 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 4982 3136 4988 3188
rect 5040 3176 5046 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 5040 3148 5089 3176
rect 5040 3136 5046 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 5316 3148 5365 3176
rect 5316 3136 5322 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5868 3148 6009 3176
rect 5868 3136 5874 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 5997 3139 6055 3145
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6420 3148 6561 3176
rect 6420 3136 6426 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6696 3148 6837 3176
rect 6696 3136 6702 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6972 3148 7113 3176
rect 6972 3136 6978 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7374 3176 7380 3188
rect 7335 3148 7380 3176
rect 7101 3139 7159 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7524 3148 7665 3176
rect 7524 3136 7530 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 7800 3148 7941 3176
rect 7800 3136 7806 3148
rect 7929 3145 7941 3148
rect 7975 3145 7987 3179
rect 7929 3139 7987 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8076 3148 8217 3176
rect 8076 3136 8082 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8352 3148 8493 3176
rect 8352 3136 8358 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 8481 3139 8539 3145
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8628 3148 8769 3176
rect 8628 3136 8634 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 8757 3139 8815 3145
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8904 3148 9137 3176
rect 8904 3136 8910 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9125 3139 9183 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9824 3148 9965 3176
rect 9824 3136 9830 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 9953 3139 10011 3145
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 10560 3148 10793 3176
rect 10560 3136 10566 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 11112 3148 11345 3176
rect 11112 3136 11118 3148
rect 11333 3145 11345 3148
rect 11379 3145 11391 3179
rect 11333 3139 11391 3145
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11940 3148 12173 3176
rect 11940 3136 11946 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 12492 3148 12725 3176
rect 12492 3136 12498 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 12713 3139 12771 3145
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 13265 3179 13323 3185
rect 13265 3176 13277 3179
rect 13044 3148 13277 3176
rect 13044 3136 13050 3148
rect 13265 3145 13277 3148
rect 13311 3145 13323 3179
rect 13265 3139 13323 3145
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13504 3148 13553 3176
rect 13504 3136 13510 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13814 3176 13820 3188
rect 13775 3148 13820 3176
rect 13541 3139 13599 3145
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 14148 3148 14381 3176
rect 14148 3136 14154 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 14369 3139 14427 3145
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 15197 3179 15255 3185
rect 15197 3176 15209 3179
rect 14700 3148 15209 3176
rect 14700 3136 14706 3148
rect 15197 3145 15209 3148
rect 15243 3145 15255 3179
rect 15197 3139 15255 3145
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15344 3148 15761 3176
rect 15344 3136 15350 3148
rect 15749 3145 15761 3148
rect 15795 3145 15807 3179
rect 15749 3139 15807 3145
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16080 3148 16865 3176
rect 16080 3136 16086 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17000 3148 17693 3176
rect 17000 3136 17006 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 18509 3179 18567 3185
rect 18509 3176 18521 3179
rect 17828 3148 18521 3176
rect 17828 3136 17834 3148
rect 18509 3145 18521 3148
rect 18555 3145 18567 3179
rect 18509 3139 18567 3145
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 18656 3148 19441 3176
rect 18656 3136 18662 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 19576 3148 20269 3176
rect 19576 3136 19582 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 21361 3179 21419 3185
rect 21361 3176 21373 3179
rect 20496 3148 21373 3176
rect 20496 3136 20502 3148
rect 21361 3145 21373 3148
rect 21407 3145 21419 3179
rect 21361 3139 21419 3145
rect 21542 3136 21548 3188
rect 21600 3176 21606 3188
rect 22557 3179 22615 3185
rect 22557 3176 22569 3179
rect 21600 3148 22569 3176
rect 21600 3136 21606 3148
rect 22557 3145 22569 3148
rect 22603 3145 22615 3179
rect 22557 3139 22615 3145
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 23661 3179 23719 3185
rect 23661 3176 23673 3179
rect 22704 3148 23673 3176
rect 22704 3136 22710 3148
rect 23661 3145 23673 3148
rect 23707 3145 23719 3179
rect 23661 3139 23719 3145
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 23808 3148 24869 3176
rect 23808 3136 23814 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 25130 3136 25136 3188
rect 25188 3176 25194 3188
rect 26237 3179 26295 3185
rect 26237 3176 26249 3179
rect 25188 3148 26249 3176
rect 25188 3136 25194 3148
rect 26237 3145 26249 3148
rect 26283 3145 26295 3179
rect 26237 3139 26295 3145
rect 26326 3136 26332 3188
rect 26384 3176 26390 3188
rect 27433 3179 27491 3185
rect 27433 3176 27445 3179
rect 26384 3148 27445 3176
rect 26384 3136 26390 3148
rect 27433 3145 27445 3148
rect 27479 3145 27491 3179
rect 27433 3139 27491 3145
rect 27614 3136 27620 3188
rect 27672 3176 27678 3188
rect 28537 3179 28595 3185
rect 28537 3176 28549 3179
rect 27672 3148 28549 3176
rect 27672 3136 27678 3148
rect 28537 3145 28549 3148
rect 28583 3145 28595 3179
rect 28537 3139 28595 3145
rect 28718 3136 28724 3188
rect 28776 3176 28782 3188
rect 29733 3179 29791 3185
rect 29733 3176 29745 3179
rect 28776 3148 29745 3176
rect 28776 3136 28782 3148
rect 29733 3145 29745 3148
rect 29779 3145 29791 3179
rect 29733 3139 29791 3145
rect 29822 3136 29828 3188
rect 29880 3176 29886 3188
rect 30837 3179 30895 3185
rect 30837 3176 30849 3179
rect 29880 3148 30849 3176
rect 29880 3136 29886 3148
rect 30837 3145 30849 3148
rect 30883 3145 30895 3179
rect 30837 3139 30895 3145
rect 30926 3136 30932 3188
rect 30984 3176 30990 3188
rect 31941 3179 31999 3185
rect 31941 3176 31953 3179
rect 30984 3148 31953 3176
rect 30984 3136 30990 3148
rect 31941 3145 31953 3148
rect 31987 3145 31999 3179
rect 31941 3139 31999 3145
rect 32030 3136 32036 3188
rect 32088 3176 32094 3188
rect 32861 3179 32919 3185
rect 32861 3176 32873 3179
rect 32088 3148 32873 3176
rect 32088 3136 32094 3148
rect 32861 3145 32873 3148
rect 32907 3145 32919 3179
rect 32861 3139 32919 3145
rect 33134 3136 33140 3188
rect 33192 3176 33198 3188
rect 33965 3179 34023 3185
rect 33965 3176 33977 3179
rect 33192 3148 33977 3176
rect 33192 3136 33198 3148
rect 33965 3145 33977 3148
rect 34011 3145 34023 3179
rect 33965 3139 34023 3145
rect 34054 3136 34060 3188
rect 34112 3176 34118 3188
rect 35161 3179 35219 3185
rect 35161 3176 35173 3179
rect 34112 3148 35173 3176
rect 34112 3136 34118 3148
rect 35161 3145 35173 3148
rect 35207 3145 35219 3179
rect 35161 3139 35219 3145
rect 35342 3136 35348 3188
rect 35400 3176 35406 3188
rect 36541 3179 36599 3185
rect 36541 3176 36553 3179
rect 35400 3148 36553 3176
rect 35400 3136 35406 3148
rect 36541 3145 36553 3148
rect 36587 3145 36599 3179
rect 36541 3139 36599 3145
rect 36722 3136 36728 3188
rect 36780 3176 36786 3188
rect 37737 3179 37795 3185
rect 37737 3176 37749 3179
rect 36780 3148 37749 3176
rect 36780 3136 36786 3148
rect 37737 3145 37749 3148
rect 37783 3145 37795 3179
rect 37737 3139 37795 3145
rect 37826 3136 37832 3188
rect 37884 3176 37890 3188
rect 38841 3179 38899 3185
rect 38841 3176 38853 3179
rect 37884 3148 38853 3176
rect 37884 3136 37890 3148
rect 38841 3145 38853 3148
rect 38887 3145 38899 3179
rect 38841 3139 38899 3145
rect 38930 3136 38936 3188
rect 38988 3176 38994 3188
rect 40037 3179 40095 3185
rect 40037 3176 40049 3179
rect 38988 3148 40049 3176
rect 38988 3136 38994 3148
rect 40037 3145 40049 3148
rect 40083 3145 40095 3179
rect 40037 3139 40095 3145
rect 40126 3136 40132 3188
rect 40184 3176 40190 3188
rect 41141 3179 41199 3185
rect 41141 3176 41153 3179
rect 40184 3148 41153 3176
rect 40184 3136 40190 3148
rect 41141 3145 41153 3148
rect 41187 3145 41199 3179
rect 41141 3139 41199 3145
rect 41230 3136 41236 3188
rect 41288 3176 41294 3188
rect 41288 3148 41644 3176
rect 41288 3136 41294 3148
rect 2961 3111 3019 3117
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 4154 3108 4160 3120
rect 3007 3080 4160 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 10226 3068 10232 3120
rect 10284 3108 10290 3120
rect 10284 3080 10548 3108
rect 10284 3068 10290 3080
rect 290 3000 296 3052
rect 348 3040 354 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 348 3012 3065 3040
rect 348 3000 354 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 10520 3049 10548 3080
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 17129 3111 17187 3117
rect 17129 3108 17141 3111
rect 16632 3080 17141 3108
rect 16632 3068 16638 3080
rect 17129 3077 17141 3080
rect 17175 3077 17187 3111
rect 17129 3071 17187 3077
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 17957 3111 18015 3117
rect 17957 3108 17969 3111
rect 17276 3080 17969 3108
rect 17276 3068 17282 3080
rect 17957 3077 17969 3080
rect 18003 3077 18015 3111
rect 17957 3071 18015 3077
rect 18322 3068 18328 3120
rect 18380 3108 18386 3120
rect 19061 3111 19119 3117
rect 19061 3108 19073 3111
rect 18380 3080 19073 3108
rect 18380 3068 18386 3080
rect 19061 3077 19073 3080
rect 19107 3077 19119 3111
rect 19061 3071 19119 3077
rect 19150 3068 19156 3120
rect 19208 3108 19214 3120
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 19208 3080 19993 3108
rect 19208 3068 19214 3080
rect 19981 3077 19993 3080
rect 20027 3077 20039 3111
rect 19981 3071 20039 3077
rect 20162 3068 20168 3120
rect 20220 3108 20226 3120
rect 21085 3111 21143 3117
rect 21085 3108 21097 3111
rect 20220 3080 21097 3108
rect 20220 3068 20226 3080
rect 21085 3077 21097 3080
rect 21131 3077 21143 3111
rect 21085 3071 21143 3077
rect 21266 3068 21272 3120
rect 21324 3108 21330 3120
rect 22281 3111 22339 3117
rect 22281 3108 22293 3111
rect 21324 3080 22293 3108
rect 21324 3068 21330 3080
rect 22281 3077 22293 3080
rect 22327 3077 22339 3111
rect 22281 3071 22339 3077
rect 22370 3068 22376 3120
rect 22428 3108 22434 3120
rect 23385 3111 23443 3117
rect 23385 3108 23397 3111
rect 22428 3080 23397 3108
rect 22428 3068 22434 3080
rect 23385 3077 23397 3080
rect 23431 3077 23443 3111
rect 23385 3071 23443 3077
rect 23474 3068 23480 3120
rect 23532 3108 23538 3120
rect 24213 3111 24271 3117
rect 24213 3108 24225 3111
rect 23532 3080 24225 3108
rect 23532 3068 23538 3080
rect 24213 3077 24225 3080
rect 24259 3077 24271 3111
rect 24213 3071 24271 3077
rect 24302 3068 24308 3120
rect 24360 3108 24366 3120
rect 25409 3111 25467 3117
rect 25409 3108 25421 3111
rect 24360 3080 25421 3108
rect 24360 3068 24366 3080
rect 25409 3077 25421 3080
rect 25455 3077 25467 3111
rect 25409 3071 25467 3077
rect 25958 3068 25964 3120
rect 26016 3108 26022 3120
rect 27157 3111 27215 3117
rect 27157 3108 27169 3111
rect 26016 3080 27169 3108
rect 26016 3068 26022 3080
rect 27157 3077 27169 3080
rect 27203 3077 27215 3111
rect 27157 3071 27215 3077
rect 27246 3068 27252 3120
rect 27304 3108 27310 3120
rect 28261 3111 28319 3117
rect 28261 3108 28273 3111
rect 27304 3080 28273 3108
rect 27304 3068 27310 3080
rect 28261 3077 28273 3080
rect 28307 3077 28319 3111
rect 28261 3071 28319 3077
rect 28994 3068 29000 3120
rect 29052 3108 29058 3120
rect 30009 3111 30067 3117
rect 30009 3108 30021 3111
rect 29052 3080 30021 3108
rect 29052 3068 29058 3080
rect 30009 3077 30021 3080
rect 30055 3077 30067 3111
rect 30009 3071 30067 3077
rect 30098 3068 30104 3120
rect 30156 3108 30162 3120
rect 31113 3111 31171 3117
rect 31113 3108 31125 3111
rect 30156 3080 31125 3108
rect 30156 3068 30162 3080
rect 31113 3077 31125 3080
rect 31159 3077 31171 3111
rect 31113 3071 31171 3077
rect 31754 3068 31760 3120
rect 31812 3108 31818 3120
rect 32309 3111 32367 3117
rect 32309 3108 32321 3111
rect 31812 3080 32321 3108
rect 31812 3068 31818 3080
rect 32309 3077 32321 3080
rect 32355 3077 32367 3111
rect 32309 3071 32367 3077
rect 32398 3068 32404 3120
rect 32456 3108 32462 3120
rect 33413 3111 33471 3117
rect 33413 3108 33425 3111
rect 32456 3080 33425 3108
rect 32456 3068 32462 3080
rect 33413 3077 33425 3080
rect 33459 3077 33471 3111
rect 33413 3071 33471 3077
rect 33502 3068 33508 3120
rect 33560 3108 33566 3120
rect 34517 3111 34575 3117
rect 34517 3108 34529 3111
rect 33560 3080 34529 3108
rect 33560 3068 33566 3080
rect 34517 3077 34529 3080
rect 34563 3077 34575 3111
rect 34517 3071 34575 3077
rect 34790 3068 34796 3120
rect 34848 3108 34854 3120
rect 35989 3111 36047 3117
rect 35989 3108 36001 3111
rect 34848 3080 36001 3108
rect 34848 3068 34854 3080
rect 35989 3077 36001 3080
rect 36035 3077 36047 3111
rect 35989 3071 36047 3077
rect 36446 3068 36452 3120
rect 36504 3108 36510 3120
rect 37461 3111 37519 3117
rect 37461 3108 37473 3111
rect 36504 3080 37473 3108
rect 36504 3068 36510 3080
rect 37461 3077 37473 3080
rect 37507 3077 37519 3111
rect 37461 3071 37519 3077
rect 37550 3068 37556 3120
rect 37608 3108 37614 3120
rect 38565 3111 38623 3117
rect 38565 3108 38577 3111
rect 37608 3080 38577 3108
rect 37608 3068 37614 3080
rect 38565 3077 38577 3080
rect 38611 3077 38623 3111
rect 38565 3071 38623 3077
rect 38654 3068 38660 3120
rect 38712 3108 38718 3120
rect 39669 3111 39727 3117
rect 39669 3108 39681 3111
rect 38712 3080 39681 3108
rect 38712 3068 38718 3080
rect 39669 3077 39681 3080
rect 39715 3077 39727 3111
rect 39669 3071 39727 3077
rect 39758 3068 39764 3120
rect 39816 3108 39822 3120
rect 40865 3111 40923 3117
rect 40865 3108 40877 3111
rect 39816 3080 40877 3108
rect 39816 3068 39822 3080
rect 40865 3077 40877 3080
rect 40911 3077 40923 3111
rect 40865 3071 40923 3077
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9180 3012 9413 3040
rect 9180 3000 9186 3012
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10505 3003 10563 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11388 3012 11713 3040
rect 11388 3000 11394 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 12434 3040 12440 3052
rect 12395 3012 12440 3040
rect 11701 3003 11759 3009
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12768 3012 13001 3040
rect 12768 3000 12774 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14424 3012 14933 3040
rect 14424 3000 14430 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 15252 3012 15485 3040
rect 15252 3000 15258 3012
rect 15473 3009 15485 3012
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15620 3012 16037 3040
rect 15620 3000 15626 3012
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 16666 3000 16672 3052
rect 16724 3040 16730 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 16724 3012 17417 3040
rect 16724 3000 16730 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 17552 3012 18245 3040
rect 17552 3000 17558 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 18932 3012 19717 3040
rect 18932 3000 18938 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 19886 3000 19892 3052
rect 19944 3040 19950 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 19944 3012 20821 3040
rect 19944 3000 19950 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 20990 3000 20996 3052
rect 21048 3040 21054 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21048 3012 22017 3040
rect 21048 3000 21054 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22833 3043 22891 3049
rect 22833 3040 22845 3043
rect 22152 3012 22845 3040
rect 22152 3000 22158 3012
rect 22833 3009 22845 3012
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 22922 3000 22928 3052
rect 22980 3040 22986 3052
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 22980 3012 23949 3040
rect 22980 3000 22986 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24084 3012 25145 3040
rect 24084 3000 24090 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25498 3000 25504 3052
rect 25556 3040 25562 3052
rect 26513 3043 26571 3049
rect 26513 3040 26525 3043
rect 25556 3012 26525 3040
rect 25556 3000 25562 3012
rect 26513 3009 26525 3012
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 26602 3000 26608 3052
rect 26660 3040 26666 3052
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 26660 3012 27721 3040
rect 26660 3000 26666 3012
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 27798 3000 27804 3052
rect 27856 3040 27862 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 27856 3012 28825 3040
rect 27856 3000 27862 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 29270 3000 29276 3052
rect 29328 3040 29334 3052
rect 30285 3043 30343 3049
rect 30285 3040 30297 3043
rect 29328 3012 30297 3040
rect 29328 3000 29334 3012
rect 30285 3009 30297 3012
rect 30331 3009 30343 3043
rect 30285 3003 30343 3009
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 30432 3012 31401 3040
rect 30432 3000 30438 3012
rect 31389 3009 31401 3012
rect 31435 3009 31447 3043
rect 31389 3003 31447 3009
rect 31846 3000 31852 3052
rect 31904 3040 31910 3052
rect 32585 3043 32643 3049
rect 32585 3040 32597 3043
rect 31904 3012 32597 3040
rect 31904 3000 31910 3012
rect 32585 3009 32597 3012
rect 32631 3009 32643 3043
rect 32585 3003 32643 3009
rect 32674 3000 32680 3052
rect 32732 3040 32738 3052
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 32732 3012 33701 3040
rect 32732 3000 32738 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 33689 3003 33747 3009
rect 33778 3000 33784 3052
rect 33836 3040 33842 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 33836 3012 34897 3040
rect 33836 3000 33842 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 34885 3003 34943 3009
rect 35066 3000 35072 3052
rect 35124 3040 35130 3052
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 35124 3012 36277 3040
rect 35124 3000 35130 3012
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36817 3043 36875 3049
rect 36817 3040 36829 3043
rect 36265 3003 36323 3009
rect 36372 3012 36829 3040
rect 14 2932 20 2984
rect 72 2972 78 2984
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 72 2944 3617 2972
rect 72 2932 78 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 4154 2972 4160 2984
rect 4115 2944 4160 2972
rect 3605 2935 3663 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 4724 2904 4752 2935
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 10008 2944 10241 2972
rect 10008 2932 10014 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14645 2975 14703 2981
rect 14645 2972 14657 2975
rect 13964 2944 14657 2972
rect 13964 2932 13970 2944
rect 14645 2941 14657 2944
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 15746 2932 15752 2984
rect 15804 2972 15810 2984
rect 16301 2975 16359 2981
rect 16301 2972 16313 2975
rect 15804 2944 16313 2972
rect 15804 2932 15810 2944
rect 16301 2941 16313 2944
rect 16347 2941 16359 2975
rect 16301 2935 16359 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18012 2944 18797 2972
rect 18012 2932 18018 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 19610 2932 19616 2984
rect 19668 2972 19674 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 19668 2944 20545 2972
rect 19668 2932 19674 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 20772 2944 21649 2972
rect 20772 2932 20778 2944
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 21637 2935 21695 2941
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 23109 2975 23167 2981
rect 23109 2972 23121 2975
rect 22244 2944 23121 2972
rect 22244 2932 22250 2944
rect 23109 2941 23121 2944
rect 23155 2941 23167 2975
rect 23109 2935 23167 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 23624 2944 24593 2972
rect 23624 2932 23630 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 24912 2944 25697 2972
rect 24912 2932 24918 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 25685 2935 25743 2941
rect 25866 2932 25872 2984
rect 25924 2972 25930 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25924 2944 25973 2972
rect 25924 2932 25930 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 26789 2975 26847 2981
rect 26789 2972 26801 2975
rect 25961 2935 26019 2941
rect 26206 2944 26801 2972
rect 624 2876 4752 2904
rect 624 2864 630 2876
rect 25774 2864 25780 2916
rect 25832 2904 25838 2916
rect 26206 2904 26234 2944
rect 26789 2941 26801 2944
rect 26835 2941 26847 2975
rect 26789 2935 26847 2941
rect 26878 2932 26884 2984
rect 26936 2972 26942 2984
rect 27985 2975 28043 2981
rect 27985 2972 27997 2975
rect 26936 2944 27997 2972
rect 26936 2932 26942 2944
rect 27985 2941 27997 2944
rect 28031 2941 28043 2975
rect 27985 2935 28043 2941
rect 28074 2932 28080 2984
rect 28132 2972 28138 2984
rect 29089 2975 29147 2981
rect 29089 2972 29101 2975
rect 28132 2944 29101 2972
rect 28132 2932 28138 2944
rect 29089 2941 29101 2944
rect 29135 2941 29147 2975
rect 29089 2935 29147 2941
rect 29365 2975 29423 2981
rect 29365 2941 29377 2975
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 25832 2876 26234 2904
rect 25832 2864 25838 2876
rect 28166 2864 28172 2916
rect 28224 2904 28230 2916
rect 29380 2904 29408 2935
rect 29546 2932 29552 2984
rect 29604 2972 29610 2984
rect 30561 2975 30619 2981
rect 30561 2972 30573 2975
rect 29604 2944 30573 2972
rect 29604 2932 29610 2944
rect 30561 2941 30573 2944
rect 30607 2941 30619 2975
rect 30561 2935 30619 2941
rect 30650 2932 30656 2984
rect 30708 2972 30714 2984
rect 31665 2975 31723 2981
rect 31665 2972 31677 2975
rect 30708 2944 31677 2972
rect 30708 2932 30714 2944
rect 31665 2941 31677 2944
rect 31711 2941 31723 2975
rect 31665 2935 31723 2941
rect 32122 2932 32128 2984
rect 32180 2972 32186 2984
rect 33137 2975 33195 2981
rect 33137 2972 33149 2975
rect 32180 2944 33149 2972
rect 32180 2932 32186 2944
rect 33137 2941 33149 2944
rect 33183 2941 33195 2975
rect 33137 2935 33195 2941
rect 33226 2932 33232 2984
rect 33284 2972 33290 2984
rect 34241 2975 34299 2981
rect 34241 2972 34253 2975
rect 33284 2944 34253 2972
rect 33284 2932 33290 2944
rect 34241 2941 34253 2944
rect 34287 2941 34299 2975
rect 34241 2935 34299 2941
rect 34514 2932 34520 2984
rect 34572 2972 34578 2984
rect 35437 2975 35495 2981
rect 35437 2972 35449 2975
rect 34572 2944 35449 2972
rect 34572 2932 34578 2944
rect 35437 2941 35449 2944
rect 35483 2941 35495 2975
rect 35437 2935 35495 2941
rect 35713 2975 35771 2981
rect 35713 2941 35725 2975
rect 35759 2941 35771 2975
rect 35713 2935 35771 2941
rect 28224 2876 29408 2904
rect 28224 2864 28230 2876
rect 34606 2864 34612 2916
rect 34664 2904 34670 2916
rect 35728 2904 35756 2935
rect 35894 2932 35900 2984
rect 35952 2972 35958 2984
rect 36372 2972 36400 3012
rect 36817 3009 36829 3012
rect 36863 3009 36875 3043
rect 36817 3003 36875 3009
rect 36998 3000 37004 3052
rect 37056 3040 37062 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37056 3012 38025 3040
rect 37056 3000 37062 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 38102 3000 38108 3052
rect 38160 3040 38166 3052
rect 39117 3043 39175 3049
rect 39117 3040 39129 3043
rect 38160 3012 39129 3040
rect 38160 3000 38166 3012
rect 39117 3009 39129 3012
rect 39163 3009 39175 3043
rect 39117 3003 39175 3009
rect 39206 3000 39212 3052
rect 39264 3040 39270 3052
rect 40313 3043 40371 3049
rect 40313 3040 40325 3043
rect 39264 3012 40325 3040
rect 39264 3000 39270 3012
rect 40313 3009 40325 3012
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 40402 3000 40408 3052
rect 40460 3040 40466 3052
rect 41417 3043 41475 3049
rect 41417 3040 41429 3043
rect 40460 3012 41429 3040
rect 40460 3000 40466 3012
rect 41417 3009 41429 3012
rect 41463 3009 41475 3043
rect 41616 3040 41644 3148
rect 41690 3136 41696 3188
rect 41748 3176 41754 3188
rect 42613 3179 42671 3185
rect 42613 3176 42625 3179
rect 41748 3148 42625 3176
rect 41748 3136 41754 3148
rect 42613 3145 42625 3148
rect 42659 3145 42671 3179
rect 42613 3139 42671 3145
rect 42794 3136 42800 3188
rect 42852 3176 42858 3188
rect 43441 3179 43499 3185
rect 43441 3176 43453 3179
rect 42852 3148 43453 3176
rect 42852 3136 42858 3148
rect 43441 3145 43453 3148
rect 43487 3145 43499 3179
rect 43441 3139 43499 3145
rect 43530 3136 43536 3188
rect 43588 3176 43594 3188
rect 44269 3179 44327 3185
rect 44269 3176 44281 3179
rect 43588 3148 44281 3176
rect 43588 3136 43594 3148
rect 44269 3145 44281 3148
rect 44315 3145 44327 3179
rect 44269 3139 44327 3145
rect 44450 3136 44456 3188
rect 44508 3176 44514 3188
rect 45189 3179 45247 3185
rect 45189 3176 45201 3179
rect 44508 3148 45201 3176
rect 44508 3136 44514 3148
rect 45189 3145 45201 3148
rect 45235 3145 45247 3179
rect 45189 3139 45247 3145
rect 47486 3136 47492 3188
rect 47544 3176 47550 3188
rect 47765 3179 47823 3185
rect 47765 3176 47777 3179
rect 47544 3148 47777 3176
rect 47544 3136 47550 3148
rect 47765 3145 47777 3148
rect 47811 3145 47823 3179
rect 47765 3139 47823 3145
rect 48590 3136 48596 3188
rect 48648 3176 48654 3188
rect 48685 3179 48743 3185
rect 48685 3176 48697 3179
rect 48648 3148 48697 3176
rect 48648 3136 48654 3148
rect 48685 3145 48697 3148
rect 48731 3145 48743 3179
rect 48685 3139 48743 3145
rect 48866 3136 48872 3188
rect 48924 3176 48930 3188
rect 48961 3179 49019 3185
rect 48961 3176 48973 3179
rect 48924 3148 48973 3176
rect 48924 3136 48930 3148
rect 48961 3145 48973 3148
rect 49007 3145 49019 3179
rect 48961 3139 49019 3145
rect 49142 3136 49148 3188
rect 49200 3176 49206 3188
rect 49237 3179 49295 3185
rect 49237 3176 49249 3179
rect 49200 3148 49249 3176
rect 49200 3136 49206 3148
rect 49237 3145 49249 3148
rect 49283 3145 49295 3179
rect 49237 3139 49295 3145
rect 49418 3136 49424 3188
rect 49476 3176 49482 3188
rect 49513 3179 49571 3185
rect 49513 3176 49525 3179
rect 49476 3148 49525 3176
rect 49476 3136 49482 3148
rect 49513 3145 49525 3148
rect 49559 3145 49571 3179
rect 49513 3139 49571 3145
rect 49694 3136 49700 3188
rect 49752 3176 49758 3188
rect 49789 3179 49847 3185
rect 49789 3176 49801 3179
rect 49752 3148 49801 3176
rect 49752 3136 49758 3148
rect 49789 3145 49801 3148
rect 49835 3145 49847 3179
rect 49789 3139 49847 3145
rect 49970 3136 49976 3188
rect 50028 3176 50034 3188
rect 50341 3179 50399 3185
rect 50341 3176 50353 3179
rect 50028 3148 50353 3176
rect 50028 3136 50034 3148
rect 50341 3145 50353 3148
rect 50387 3145 50399 3179
rect 50341 3139 50399 3145
rect 50522 3136 50528 3188
rect 50580 3176 50586 3188
rect 50893 3179 50951 3185
rect 50893 3176 50905 3179
rect 50580 3148 50905 3176
rect 50580 3136 50586 3148
rect 50893 3145 50905 3148
rect 50939 3145 50951 3179
rect 50893 3139 50951 3145
rect 51074 3136 51080 3188
rect 51132 3176 51138 3188
rect 51169 3179 51227 3185
rect 51169 3176 51181 3179
rect 51132 3148 51181 3176
rect 51132 3136 51138 3148
rect 51169 3145 51181 3148
rect 51215 3145 51227 3179
rect 51169 3139 51227 3145
rect 51350 3136 51356 3188
rect 51408 3176 51414 3188
rect 51721 3179 51779 3185
rect 51721 3176 51733 3179
rect 51408 3148 51733 3176
rect 51408 3136 51414 3148
rect 51721 3145 51733 3148
rect 51767 3145 51779 3179
rect 51721 3139 51779 3145
rect 51902 3136 51908 3188
rect 51960 3176 51966 3188
rect 52273 3179 52331 3185
rect 52273 3176 52285 3179
rect 51960 3148 52285 3176
rect 51960 3136 51966 3148
rect 52273 3145 52285 3148
rect 52319 3145 52331 3179
rect 52273 3139 52331 3145
rect 52454 3136 52460 3188
rect 52512 3176 52518 3188
rect 52549 3179 52607 3185
rect 52549 3176 52561 3179
rect 52512 3148 52561 3176
rect 52512 3136 52518 3148
rect 52549 3145 52561 3148
rect 52595 3145 52607 3179
rect 52549 3139 52607 3145
rect 52730 3136 52736 3188
rect 52788 3176 52794 3188
rect 53193 3179 53251 3185
rect 53193 3176 53205 3179
rect 52788 3148 53205 3176
rect 52788 3136 52794 3148
rect 53193 3145 53205 3148
rect 53239 3145 53251 3179
rect 53193 3139 53251 3145
rect 53282 3136 53288 3188
rect 53340 3176 53346 3188
rect 53745 3179 53803 3185
rect 53745 3176 53757 3179
rect 53340 3148 53757 3176
rect 53340 3136 53346 3148
rect 53745 3145 53757 3148
rect 53791 3145 53803 3179
rect 53745 3139 53803 3145
rect 53834 3136 53840 3188
rect 53892 3176 53898 3188
rect 54021 3179 54079 3185
rect 54021 3176 54033 3179
rect 53892 3148 54033 3176
rect 53892 3136 53898 3148
rect 54021 3145 54033 3148
rect 54067 3145 54079 3179
rect 54021 3139 54079 3145
rect 54110 3136 54116 3188
rect 54168 3176 54174 3188
rect 54573 3179 54631 3185
rect 54573 3176 54585 3179
rect 54168 3148 54585 3176
rect 54168 3136 54174 3148
rect 54573 3145 54585 3148
rect 54619 3145 54631 3179
rect 54573 3139 54631 3145
rect 54662 3136 54668 3188
rect 54720 3176 54726 3188
rect 55125 3179 55183 3185
rect 55125 3176 55137 3179
rect 54720 3148 55137 3176
rect 54720 3136 54726 3148
rect 55125 3145 55137 3148
rect 55171 3145 55183 3179
rect 55125 3139 55183 3145
rect 55398 3136 55404 3188
rect 55456 3176 55462 3188
rect 55769 3179 55827 3185
rect 55769 3176 55781 3179
rect 55456 3148 55781 3176
rect 55456 3136 55462 3148
rect 55769 3145 55781 3148
rect 55815 3145 55827 3179
rect 55769 3139 55827 3145
rect 56042 3136 56048 3188
rect 56100 3176 56106 3188
rect 56597 3179 56655 3185
rect 56597 3176 56609 3179
rect 56100 3148 56609 3176
rect 56100 3136 56106 3148
rect 56597 3145 56609 3148
rect 56643 3145 56655 3179
rect 56597 3139 56655 3145
rect 56686 3136 56692 3188
rect 56744 3176 56750 3188
rect 57149 3179 57207 3185
rect 57149 3176 57161 3179
rect 56744 3148 57161 3176
rect 56744 3136 56750 3148
rect 57149 3145 57161 3148
rect 57195 3145 57207 3179
rect 57149 3139 57207 3145
rect 57514 3136 57520 3188
rect 57572 3176 57578 3188
rect 58069 3179 58127 3185
rect 58069 3176 58081 3179
rect 57572 3148 58081 3176
rect 57572 3136 57578 3148
rect 58069 3145 58081 3148
rect 58115 3145 58127 3179
rect 58069 3139 58127 3145
rect 58250 3136 58256 3188
rect 58308 3176 58314 3188
rect 58897 3179 58955 3185
rect 58897 3176 58909 3179
rect 58308 3148 58909 3176
rect 58308 3136 58314 3148
rect 58897 3145 58909 3148
rect 58943 3145 58955 3179
rect 58897 3139 58955 3145
rect 59078 3136 59084 3188
rect 59136 3176 59142 3188
rect 59725 3179 59783 3185
rect 59725 3176 59737 3179
rect 59136 3148 59737 3176
rect 59136 3136 59142 3148
rect 59725 3145 59737 3148
rect 59771 3145 59783 3179
rect 59725 3139 59783 3145
rect 59906 3136 59912 3188
rect 59964 3176 59970 3188
rect 60645 3179 60703 3185
rect 60645 3176 60657 3179
rect 59964 3148 60657 3176
rect 59964 3136 59970 3148
rect 60645 3145 60657 3148
rect 60691 3145 60703 3179
rect 60645 3139 60703 3145
rect 60734 3136 60740 3188
rect 60792 3176 60798 3188
rect 61197 3179 61255 3185
rect 61197 3176 61209 3179
rect 60792 3148 61209 3176
rect 60792 3136 60798 3148
rect 61197 3145 61209 3148
rect 61243 3145 61255 3179
rect 61197 3139 61255 3145
rect 61378 3136 61384 3188
rect 61436 3176 61442 3188
rect 62025 3179 62083 3185
rect 62025 3176 62037 3179
rect 61436 3148 62037 3176
rect 61436 3136 61442 3148
rect 62025 3145 62037 3148
rect 62071 3145 62083 3179
rect 62025 3139 62083 3145
rect 62114 3136 62120 3188
rect 62172 3176 62178 3188
rect 62577 3179 62635 3185
rect 62577 3176 62589 3179
rect 62172 3148 62589 3176
rect 62172 3136 62178 3148
rect 62577 3145 62589 3148
rect 62623 3145 62635 3179
rect 62577 3139 62635 3145
rect 62666 3136 62672 3188
rect 62724 3176 62730 3188
rect 63497 3179 63555 3185
rect 63497 3176 63509 3179
rect 62724 3148 63509 3176
rect 62724 3136 62730 3148
rect 63497 3145 63509 3148
rect 63543 3145 63555 3179
rect 63497 3139 63555 3145
rect 64322 3136 64328 3188
rect 64380 3176 64386 3188
rect 65153 3179 65211 3185
rect 65153 3176 65165 3179
rect 64380 3148 65165 3176
rect 64380 3136 64386 3148
rect 65153 3145 65165 3148
rect 65199 3145 65211 3179
rect 65153 3139 65211 3145
rect 65702 3136 65708 3188
rect 65760 3176 65766 3188
rect 66349 3179 66407 3185
rect 66349 3176 66361 3179
rect 65760 3148 66361 3176
rect 65760 3136 65766 3148
rect 66349 3145 66361 3148
rect 66395 3145 66407 3179
rect 66349 3139 66407 3145
rect 66530 3136 66536 3188
rect 66588 3176 66594 3188
rect 66625 3179 66683 3185
rect 66625 3176 66637 3179
rect 66588 3148 66637 3176
rect 66588 3136 66594 3148
rect 66625 3145 66637 3148
rect 66671 3145 66683 3179
rect 67082 3176 67088 3188
rect 67043 3148 67088 3176
rect 66625 3139 66683 3145
rect 67082 3136 67088 3148
rect 67140 3136 67146 3188
rect 67361 3179 67419 3185
rect 67361 3145 67373 3179
rect 67407 3176 67419 3179
rect 67450 3176 67456 3188
rect 67407 3148 67456 3176
rect 67407 3145 67419 3148
rect 67361 3139 67419 3145
rect 67450 3136 67456 3148
rect 67508 3136 67514 3188
rect 67634 3176 67640 3188
rect 67595 3148 67640 3176
rect 67634 3136 67640 3148
rect 67692 3136 67698 3188
rect 41966 3068 41972 3120
rect 42024 3108 42030 3120
rect 42889 3111 42947 3117
rect 42889 3108 42901 3111
rect 42024 3080 42901 3108
rect 42024 3068 42030 3080
rect 42889 3077 42901 3080
rect 42935 3077 42947 3111
rect 42889 3071 42947 3077
rect 43070 3068 43076 3120
rect 43128 3108 43134 3120
rect 43993 3111 44051 3117
rect 43993 3108 44005 3111
rect 43128 3080 44005 3108
rect 43128 3068 43134 3080
rect 43993 3077 44005 3080
rect 44039 3077 44051 3111
rect 43993 3071 44051 3077
rect 44726 3068 44732 3120
rect 44784 3108 44790 3120
rect 45465 3111 45523 3117
rect 45465 3108 45477 3111
rect 44784 3080 45477 3108
rect 44784 3068 44790 3080
rect 45465 3077 45477 3080
rect 45511 3077 45523 3111
rect 45465 3071 45523 3077
rect 50246 3068 50252 3120
rect 50304 3108 50310 3120
rect 50617 3111 50675 3117
rect 50617 3108 50629 3111
rect 50304 3080 50629 3108
rect 50304 3068 50310 3080
rect 50617 3077 50629 3080
rect 50663 3077 50675 3111
rect 50617 3071 50675 3077
rect 51626 3068 51632 3120
rect 51684 3108 51690 3120
rect 51997 3111 52055 3117
rect 51997 3108 52009 3111
rect 51684 3080 52009 3108
rect 51684 3068 51690 3080
rect 51997 3077 52009 3080
rect 52043 3077 52055 3111
rect 51997 3071 52055 3077
rect 53006 3068 53012 3120
rect 53064 3108 53070 3120
rect 53469 3111 53527 3117
rect 53469 3108 53481 3111
rect 53064 3080 53481 3108
rect 53064 3068 53070 3080
rect 53469 3077 53481 3080
rect 53515 3077 53527 3111
rect 53469 3071 53527 3077
rect 53926 3068 53932 3120
rect 53984 3108 53990 3120
rect 54297 3111 54355 3117
rect 54297 3108 54309 3111
rect 53984 3080 54309 3108
rect 53984 3068 53990 3080
rect 54297 3077 54309 3080
rect 54343 3077 54355 3111
rect 54297 3071 54355 3077
rect 54386 3068 54392 3120
rect 54444 3108 54450 3120
rect 54849 3111 54907 3117
rect 54849 3108 54861 3111
rect 54444 3080 54861 3108
rect 54444 3068 54450 3080
rect 54849 3077 54861 3080
rect 54895 3077 54907 3111
rect 54849 3071 54907 3077
rect 54938 3068 54944 3120
rect 54996 3108 55002 3120
rect 55493 3111 55551 3117
rect 55493 3108 55505 3111
rect 54996 3080 55505 3108
rect 54996 3068 55002 3080
rect 55493 3077 55505 3080
rect 55539 3077 55551 3111
rect 55493 3071 55551 3077
rect 56962 3068 56968 3120
rect 57020 3108 57026 3120
rect 57425 3111 57483 3117
rect 57425 3108 57437 3111
rect 57020 3080 57437 3108
rect 57020 3068 57026 3080
rect 57425 3077 57437 3080
rect 57471 3077 57483 3111
rect 57425 3071 57483 3077
rect 57974 3068 57980 3120
rect 58032 3108 58038 3120
rect 58345 3111 58403 3117
rect 58345 3108 58357 3111
rect 58032 3080 58357 3108
rect 58032 3068 58038 3080
rect 58345 3077 58357 3080
rect 58391 3077 58403 3111
rect 58345 3071 58403 3077
rect 58526 3068 58532 3120
rect 58584 3108 58590 3120
rect 59173 3111 59231 3117
rect 59173 3108 59185 3111
rect 58584 3080 59185 3108
rect 58584 3068 58590 3080
rect 59173 3077 59185 3080
rect 59219 3077 59231 3111
rect 59173 3071 59231 3077
rect 59354 3068 59360 3120
rect 59412 3108 59418 3120
rect 60001 3111 60059 3117
rect 60001 3108 60013 3111
rect 59412 3080 60013 3108
rect 59412 3068 59418 3080
rect 60001 3077 60013 3080
rect 60047 3077 60059 3111
rect 60001 3071 60059 3077
rect 60182 3068 60188 3120
rect 60240 3108 60246 3120
rect 60921 3111 60979 3117
rect 60921 3108 60933 3111
rect 60240 3080 60933 3108
rect 60240 3068 60246 3080
rect 60921 3077 60933 3080
rect 60967 3077 60979 3111
rect 60921 3071 60979 3077
rect 61010 3068 61016 3120
rect 61068 3108 61074 3120
rect 61749 3111 61807 3117
rect 61749 3108 61761 3111
rect 61068 3080 61761 3108
rect 61068 3068 61074 3080
rect 61749 3077 61761 3080
rect 61795 3077 61807 3111
rect 61749 3071 61807 3077
rect 62206 3068 62212 3120
rect 62264 3108 62270 3120
rect 62853 3111 62911 3117
rect 62853 3108 62865 3111
rect 62264 3080 62865 3108
rect 62264 3068 62270 3080
rect 62853 3077 62865 3080
rect 62899 3077 62911 3111
rect 62853 3071 62911 3077
rect 62942 3068 62948 3120
rect 63000 3108 63006 3120
rect 63773 3111 63831 3117
rect 63773 3108 63785 3111
rect 63000 3080 63785 3108
rect 63000 3068 63006 3080
rect 63773 3077 63785 3080
rect 63819 3077 63831 3111
rect 63773 3071 63831 3077
rect 64046 3068 64052 3120
rect 64104 3108 64110 3120
rect 64877 3111 64935 3117
rect 64877 3108 64889 3111
rect 64104 3080 64889 3108
rect 64104 3068 64110 3080
rect 64877 3077 64889 3080
rect 64923 3077 64935 3111
rect 64877 3071 64935 3077
rect 65242 3068 65248 3120
rect 65300 3108 65306 3120
rect 66073 3111 66131 3117
rect 66073 3108 66085 3111
rect 65300 3080 66085 3108
rect 65300 3068 65306 3080
rect 66073 3077 66085 3080
rect 66119 3077 66131 3111
rect 66073 3071 66131 3077
rect 42245 3043 42303 3049
rect 42245 3040 42257 3043
rect 41616 3012 42257 3040
rect 41417 3003 41475 3009
rect 42245 3009 42257 3012
rect 42291 3009 42303 3043
rect 42245 3003 42303 3009
rect 42334 3000 42340 3052
rect 42392 3040 42398 3052
rect 43165 3043 43223 3049
rect 43165 3040 43177 3043
rect 42392 3012 43177 3040
rect 42392 3000 42398 3012
rect 43165 3009 43177 3012
rect 43211 3009 43223 3043
rect 43165 3003 43223 3009
rect 43622 3000 43628 3052
rect 43680 3040 43686 3052
rect 44545 3043 44603 3049
rect 44545 3040 44557 3043
rect 43680 3012 44557 3040
rect 43680 3000 43686 3012
rect 44545 3009 44557 3012
rect 44591 3009 44603 3043
rect 44545 3003 44603 3009
rect 45002 3000 45008 3052
rect 45060 3040 45066 3052
rect 45741 3043 45799 3049
rect 45741 3040 45753 3043
rect 45060 3012 45753 3040
rect 45060 3000 45066 3012
rect 45741 3009 45753 3012
rect 45787 3009 45799 3043
rect 45741 3003 45799 3009
rect 47762 3000 47768 3052
rect 47820 3040 47826 3052
rect 48041 3043 48099 3049
rect 48041 3040 48053 3043
rect 47820 3012 48053 3040
rect 47820 3000 47826 3012
rect 48041 3009 48053 3012
rect 48087 3009 48099 3043
rect 48041 3003 48099 3009
rect 51166 3000 51172 3052
rect 51224 3040 51230 3052
rect 51445 3043 51503 3049
rect 51445 3040 51457 3043
rect 51224 3012 51457 3040
rect 51224 3000 51230 3012
rect 51445 3009 51457 3012
rect 51491 3009 51503 3043
rect 51445 3003 51503 3009
rect 52546 3000 52552 3052
rect 52604 3040 52610 3052
rect 52917 3043 52975 3049
rect 52917 3040 52929 3043
rect 52604 3012 52929 3040
rect 52604 3000 52610 3012
rect 52917 3009 52929 3012
rect 52963 3009 52975 3043
rect 52917 3003 52975 3009
rect 55766 3000 55772 3052
rect 55824 3040 55830 3052
rect 56321 3043 56379 3049
rect 56321 3040 56333 3043
rect 55824 3012 56333 3040
rect 55824 3000 55830 3012
rect 56321 3009 56333 3012
rect 56367 3009 56379 3043
rect 56321 3003 56379 3009
rect 56594 3000 56600 3052
rect 56652 3040 56658 3052
rect 56873 3043 56931 3049
rect 56873 3040 56885 3043
rect 56652 3012 56885 3040
rect 56652 3000 56658 3012
rect 56873 3009 56885 3012
rect 56919 3009 56931 3043
rect 56873 3003 56931 3009
rect 57146 3000 57152 3052
rect 57204 3040 57210 3052
rect 57701 3043 57759 3049
rect 57701 3040 57713 3043
rect 57204 3012 57713 3040
rect 57204 3000 57210 3012
rect 57701 3009 57713 3012
rect 57747 3009 57759 3043
rect 57701 3003 57759 3009
rect 58066 3000 58072 3052
rect 58124 3040 58130 3052
rect 58621 3043 58679 3049
rect 58621 3040 58633 3043
rect 58124 3012 58633 3040
rect 58124 3000 58130 3012
rect 58621 3009 58633 3012
rect 58667 3009 58679 3043
rect 58621 3003 58679 3009
rect 58802 3000 58808 3052
rect 58860 3040 58866 3052
rect 59449 3043 59507 3049
rect 59449 3040 59461 3043
rect 58860 3012 59461 3040
rect 58860 3000 58866 3012
rect 59449 3009 59461 3012
rect 59495 3009 59507 3043
rect 59449 3003 59507 3009
rect 59630 3000 59636 3052
rect 59688 3040 59694 3052
rect 60277 3043 60335 3049
rect 60277 3040 60289 3043
rect 59688 3012 60289 3040
rect 59688 3000 59694 3012
rect 60277 3009 60289 3012
rect 60323 3009 60335 3043
rect 60277 3003 60335 3009
rect 60826 3000 60832 3052
rect 60884 3040 60890 3052
rect 61473 3043 61531 3049
rect 61473 3040 61485 3043
rect 60884 3012 61485 3040
rect 60884 3000 60890 3012
rect 61473 3009 61485 3012
rect 61519 3009 61531 3043
rect 61473 3003 61531 3009
rect 61562 3000 61568 3052
rect 61620 3040 61626 3052
rect 62301 3043 62359 3049
rect 62301 3040 62313 3043
rect 61620 3012 62313 3040
rect 61620 3000 61626 3012
rect 62301 3009 62313 3012
rect 62347 3009 62359 3043
rect 62301 3003 62359 3009
rect 62390 3000 62396 3052
rect 62448 3040 62454 3052
rect 63221 3043 63279 3049
rect 63221 3040 63233 3043
rect 62448 3012 63233 3040
rect 62448 3000 62454 3012
rect 63221 3009 63233 3012
rect 63267 3009 63279 3043
rect 63221 3003 63279 3009
rect 63586 3000 63592 3052
rect 63644 3040 63650 3052
rect 64325 3043 64383 3049
rect 64325 3040 64337 3043
rect 63644 3012 64337 3040
rect 63644 3000 63650 3012
rect 64325 3009 64337 3012
rect 64371 3009 64383 3043
rect 64325 3003 64383 3009
rect 64690 3000 64696 3052
rect 64748 3040 64754 3052
rect 65429 3043 65487 3049
rect 65429 3040 65441 3043
rect 64748 3012 65441 3040
rect 64748 3000 64754 3012
rect 65429 3009 65441 3012
rect 65475 3009 65487 3043
rect 65429 3003 65487 3009
rect 65981 3043 66039 3049
rect 65981 3009 65993 3043
rect 66027 3040 66039 3043
rect 67910 3040 67916 3052
rect 66027 3012 67916 3040
rect 66027 3009 66039 3012
rect 65981 3003 66039 3009
rect 67910 3000 67916 3012
rect 67968 3000 67974 3052
rect 35952 2944 36400 2972
rect 37093 2975 37151 2981
rect 35952 2932 35958 2944
rect 37093 2941 37105 2975
rect 37139 2941 37151 2975
rect 37093 2935 37151 2941
rect 34664 2876 35756 2904
rect 34664 2864 34670 2876
rect 35986 2864 35992 2916
rect 36044 2904 36050 2916
rect 37108 2904 37136 2935
rect 37366 2932 37372 2984
rect 37424 2972 37430 2984
rect 38289 2975 38347 2981
rect 38289 2972 38301 2975
rect 37424 2944 38301 2972
rect 37424 2932 37430 2944
rect 38289 2941 38301 2944
rect 38335 2941 38347 2975
rect 38289 2935 38347 2941
rect 38378 2932 38384 2984
rect 38436 2972 38442 2984
rect 39393 2975 39451 2981
rect 39393 2972 39405 2975
rect 38436 2944 39405 2972
rect 38436 2932 38442 2944
rect 39393 2941 39405 2944
rect 39439 2941 39451 2975
rect 39393 2935 39451 2941
rect 39482 2932 39488 2984
rect 39540 2972 39546 2984
rect 40589 2975 40647 2981
rect 40589 2972 40601 2975
rect 39540 2944 40601 2972
rect 39540 2932 39546 2944
rect 40589 2941 40601 2944
rect 40635 2941 40647 2975
rect 40589 2935 40647 2941
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41693 2975 41751 2981
rect 41693 2972 41705 2975
rect 40736 2944 41705 2972
rect 40736 2932 40742 2944
rect 41693 2941 41705 2944
rect 41739 2941 41751 2975
rect 41693 2935 41751 2941
rect 41969 2975 42027 2981
rect 41969 2941 41981 2975
rect 42015 2941 42027 2975
rect 41969 2935 42027 2941
rect 36044 2876 37136 2904
rect 36044 2864 36050 2876
rect 40862 2864 40868 2916
rect 40920 2904 40926 2916
rect 41984 2904 42012 2935
rect 42886 2932 42892 2984
rect 42944 2972 42950 2984
rect 43717 2975 43775 2981
rect 43717 2972 43729 2975
rect 42944 2944 43729 2972
rect 42944 2932 42950 2944
rect 43717 2941 43729 2944
rect 43763 2941 43775 2975
rect 43717 2935 43775 2941
rect 43898 2932 43904 2984
rect 43956 2972 43962 2984
rect 44821 2975 44879 2981
rect 44821 2972 44833 2975
rect 43956 2944 44833 2972
rect 43956 2932 43962 2944
rect 44821 2941 44833 2944
rect 44867 2941 44879 2975
rect 44821 2935 44879 2941
rect 55490 2932 55496 2984
rect 55548 2972 55554 2984
rect 56045 2975 56103 2981
rect 56045 2972 56057 2975
rect 55548 2944 56057 2972
rect 55548 2932 55554 2944
rect 56045 2941 56057 2944
rect 56091 2941 56103 2975
rect 56045 2935 56103 2941
rect 63494 2932 63500 2984
rect 63552 2972 63558 2984
rect 64049 2975 64107 2981
rect 64049 2972 64061 2975
rect 63552 2944 64061 2972
rect 63552 2932 63558 2944
rect 64049 2941 64061 2944
rect 64095 2941 64107 2975
rect 64049 2935 64107 2941
rect 64601 2975 64659 2981
rect 64601 2941 64613 2975
rect 64647 2941 64659 2975
rect 64601 2935 64659 2941
rect 40920 2876 42012 2904
rect 40920 2864 40926 2876
rect 63770 2864 63776 2916
rect 63828 2904 63834 2916
rect 64616 2904 64644 2935
rect 63828 2876 64644 2904
rect 63828 2864 63834 2876
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 5626 2836 5632 2848
rect 992 2808 5632 2836
rect 992 2796 998 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 1288 2746 68816 2768
rect 1288 2694 7262 2746
rect 7314 2694 19262 2746
rect 19314 2694 31262 2746
rect 31314 2694 43262 2746
rect 43314 2694 55262 2746
rect 55314 2694 67262 2746
rect 67314 2694 68816 2746
rect 1288 2672 68816 2694
rect 2958 2524 2964 2576
rect 3016 2564 3022 2576
rect 3016 2536 4200 2564
rect 3016 2524 3022 2536
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2004 2468 2789 2496
rect 2004 2456 2010 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 3878 2496 3884 2508
rect 3559 2468 3884 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4172 2505 4200 2536
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 4488 2468 5273 2496
rect 4488 2456 4494 2468
rect 5261 2465 5273 2468
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 6086 2456 6092 2508
rect 6144 2496 6150 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 6144 2468 6285 2496
rect 6144 2456 6150 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11664 2468 11897 2496
rect 11664 2456 11670 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 28442 2456 28448 2508
rect 28500 2496 28506 2508
rect 28813 2499 28871 2505
rect 28813 2496 28825 2499
rect 28500 2468 28825 2496
rect 28500 2456 28506 2468
rect 28813 2465 28825 2468
rect 28859 2465 28871 2499
rect 28813 2459 28871 2465
rect 36170 2456 36176 2508
rect 36228 2496 36234 2508
rect 36541 2499 36599 2505
rect 36541 2496 36553 2499
rect 36228 2468 36553 2496
rect 36228 2456 36234 2468
rect 36541 2465 36553 2468
rect 36587 2465 36599 2499
rect 36541 2459 36599 2465
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 41693 2499 41751 2505
rect 41693 2496 41705 2499
rect 41472 2468 41705 2496
rect 41472 2456 41478 2468
rect 41693 2465 41705 2468
rect 41739 2465 41751 2499
rect 41693 2459 41751 2465
rect 44174 2456 44180 2508
rect 44232 2496 44238 2508
rect 44269 2499 44327 2505
rect 44269 2496 44281 2499
rect 44232 2468 44281 2496
rect 44232 2456 44238 2468
rect 44269 2465 44281 2468
rect 44315 2465 44327 2499
rect 45278 2496 45284 2508
rect 45239 2468 45284 2496
rect 44269 2459 44327 2465
rect 45278 2456 45284 2468
rect 45336 2456 45342 2508
rect 45554 2456 45560 2508
rect 45612 2496 45618 2508
rect 45830 2496 45836 2508
rect 45612 2468 45657 2496
rect 45791 2468 45836 2496
rect 45612 2456 45618 2468
rect 45830 2456 45836 2468
rect 45888 2456 45894 2508
rect 46106 2496 46112 2508
rect 46067 2468 46112 2496
rect 46106 2456 46112 2468
rect 46164 2456 46170 2508
rect 46382 2496 46388 2508
rect 46343 2468 46388 2496
rect 46382 2456 46388 2468
rect 46440 2456 46446 2508
rect 46658 2496 46664 2508
rect 46619 2468 46664 2496
rect 46658 2456 46664 2468
rect 46716 2456 46722 2508
rect 46934 2496 46940 2508
rect 46895 2468 46940 2496
rect 46934 2456 46940 2468
rect 46992 2456 46998 2508
rect 47210 2496 47216 2508
rect 47171 2468 47216 2496
rect 47210 2456 47216 2468
rect 47268 2456 47274 2508
rect 48038 2496 48044 2508
rect 47999 2468 48044 2496
rect 48038 2456 48044 2468
rect 48096 2456 48102 2508
rect 48314 2496 48320 2508
rect 48275 2468 48320 2496
rect 48314 2456 48320 2468
rect 48372 2456 48378 2508
rect 64874 2456 64880 2508
rect 64932 2496 64938 2508
rect 64969 2499 65027 2505
rect 64969 2496 64981 2499
rect 64932 2468 64981 2496
rect 64932 2456 64938 2468
rect 64969 2465 64981 2468
rect 65015 2465 65027 2499
rect 65426 2496 65432 2508
rect 65387 2468 65432 2496
rect 64969 2459 65027 2465
rect 65426 2456 65432 2468
rect 65484 2456 65490 2508
rect 65978 2496 65984 2508
rect 65939 2468 65984 2496
rect 65978 2456 65984 2468
rect 66036 2456 66042 2508
rect 66254 2496 66260 2508
rect 66215 2468 66260 2496
rect 66254 2456 66260 2468
rect 66312 2456 66318 2508
rect 66533 2499 66591 2505
rect 66533 2465 66545 2499
rect 66579 2496 66591 2499
rect 66806 2496 66812 2508
rect 66579 2468 66812 2496
rect 66579 2465 66591 2468
rect 66533 2459 66591 2465
rect 66806 2456 66812 2468
rect 66864 2456 66870 2508
rect 2498 2388 2504 2440
rect 2556 2428 2562 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2556 2400 3065 2428
rect 2556 2388 2562 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 3786 2388 3792 2440
rect 3844 2428 3850 2440
rect 3844 2400 4568 2428
rect 3844 2388 3850 2400
rect 2222 2320 2228 2372
rect 2280 2360 2286 2372
rect 3326 2360 3332 2372
rect 2280 2332 3332 2360
rect 2280 2320 2286 2332
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 3694 2320 3700 2372
rect 3752 2360 3758 2372
rect 3752 2332 3832 2360
rect 3752 2320 3758 2332
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 2501 2295 2559 2301
rect 2501 2292 2513 2295
rect 900 2264 2513 2292
rect 900 2252 906 2264
rect 2501 2261 2513 2264
rect 2547 2261 2559 2295
rect 2501 2255 2559 2261
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 3510 2292 3516 2304
rect 2832 2264 3516 2292
rect 2832 2252 2838 2264
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 3602 2252 3608 2304
rect 3660 2292 3666 2304
rect 3804 2292 3832 2332
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4433 2363 4491 2369
rect 4433 2360 4445 2363
rect 4028 2332 4445 2360
rect 4028 2320 4034 2332
rect 4433 2329 4445 2332
rect 4479 2329 4491 2363
rect 4540 2360 4568 2400
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4764 2400 5549 2428
rect 4764 2388 4770 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5868 2400 6561 2428
rect 5868 2388 5874 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 4985 2363 5043 2369
rect 4985 2360 4997 2363
rect 4540 2332 4997 2360
rect 4433 2323 4491 2329
rect 4985 2329 4997 2332
rect 5031 2329 5043 2363
rect 4985 2323 5043 2329
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 3660 2264 3705 2292
rect 3804 2264 4721 2292
rect 3660 2252 3666 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 5813 2295 5871 2301
rect 5813 2292 5825 2295
rect 5776 2264 5825 2292
rect 5776 2252 5782 2264
rect 5813 2261 5825 2264
rect 5859 2261 5871 2295
rect 5813 2255 5871 2261
rect 1288 2202 68816 2224
rect 1288 2150 13262 2202
rect 13314 2150 25262 2202
rect 25314 2150 37262 2202
rect 37314 2150 49262 2202
rect 49314 2150 61262 2202
rect 61314 2150 68816 2202
rect 1288 2128 68816 2150
rect 2133 2091 2191 2097
rect 2133 2057 2145 2091
rect 2179 2088 2191 2091
rect 2958 2088 2964 2100
rect 2179 2060 2964 2088
rect 2179 2057 2191 2060
rect 2133 2051 2191 2057
rect 2958 2048 2964 2060
rect 3016 2048 3022 2100
rect 3050 2048 3056 2100
rect 3108 2088 3114 2100
rect 3881 2091 3939 2097
rect 3881 2088 3893 2091
rect 3108 2060 3893 2088
rect 3108 2048 3114 2060
rect 3881 2057 3893 2060
rect 3927 2057 3939 2091
rect 3881 2051 3939 2057
rect 4157 2091 4215 2097
rect 4157 2057 4169 2091
rect 4203 2088 4215 2091
rect 4246 2088 4252 2100
rect 4203 2060 4252 2088
rect 4203 2057 4215 2060
rect 4157 2051 4215 2057
rect 4246 2048 4252 2060
rect 4304 2048 4310 2100
rect 4706 2048 4712 2100
rect 4764 2088 4770 2100
rect 6549 2091 6607 2097
rect 6549 2088 6561 2091
rect 4764 2060 6561 2088
rect 4764 2048 4770 2060
rect 6549 2057 6561 2060
rect 6595 2057 6607 2091
rect 6822 2088 6828 2100
rect 6783 2060 6828 2088
rect 6549 2051 6607 2057
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 2774 1980 2780 2032
rect 2832 2020 2838 2032
rect 4433 2023 4491 2029
rect 4433 2020 4445 2023
rect 2832 1992 4445 2020
rect 2832 1980 2838 1992
rect 4433 1989 4445 1992
rect 4479 1989 4491 2023
rect 4433 1983 4491 1989
rect 5534 1980 5540 2032
rect 5592 2020 5598 2032
rect 5813 2023 5871 2029
rect 5813 2020 5825 2023
rect 5592 1992 5825 2020
rect 5592 1980 5598 1992
rect 5813 1989 5825 1992
rect 5859 1989 5871 2023
rect 5813 1983 5871 1989
rect 1118 1912 1124 1964
rect 1176 1952 1182 1964
rect 2225 1955 2283 1961
rect 2225 1952 2237 1955
rect 1176 1924 2237 1952
rect 1176 1912 1182 1924
rect 2225 1921 2237 1924
rect 2271 1921 2283 1955
rect 2225 1915 2283 1921
rect 2332 1924 2820 1952
rect 1394 1776 1400 1828
rect 1452 1816 1458 1828
rect 2332 1816 2360 1924
rect 2792 1893 2820 1924
rect 2866 1912 2872 1964
rect 2924 1952 2930 1964
rect 4709 1955 4767 1961
rect 4709 1952 4721 1955
rect 2924 1924 4721 1952
rect 2924 1912 2930 1924
rect 4709 1921 4721 1924
rect 4755 1921 4767 1955
rect 4709 1915 4767 1921
rect 5350 1912 5356 1964
rect 5408 1952 5414 1964
rect 6089 1955 6147 1961
rect 6089 1952 6101 1955
rect 5408 1924 6101 1952
rect 5408 1912 5414 1924
rect 6089 1921 6101 1924
rect 6135 1921 6147 1955
rect 6089 1915 6147 1921
rect 45002 1912 45008 1964
rect 45060 1952 45066 1964
rect 46109 1955 46167 1961
rect 46109 1952 46121 1955
rect 45060 1924 46121 1952
rect 45060 1912 45066 1924
rect 46109 1921 46121 1924
rect 46155 1921 46167 1955
rect 46109 1915 46167 1921
rect 2685 1887 2743 1893
rect 2685 1853 2697 1887
rect 2731 1853 2743 1887
rect 2685 1847 2743 1853
rect 2777 1887 2835 1893
rect 2777 1853 2789 1887
rect 2823 1853 2835 1887
rect 3050 1884 3056 1896
rect 3011 1856 3056 1884
rect 2777 1847 2835 1853
rect 1452 1788 2360 1816
rect 1452 1776 1458 1788
rect 2700 1748 2728 1847
rect 3050 1844 3056 1856
rect 3108 1844 3114 1896
rect 3326 1884 3332 1896
rect 3287 1856 3332 1884
rect 3326 1844 3332 1856
rect 3384 1844 3390 1896
rect 3510 1844 3516 1896
rect 3568 1884 3574 1896
rect 3605 1887 3663 1893
rect 3605 1884 3617 1887
rect 3568 1856 3617 1884
rect 3568 1844 3574 1856
rect 3605 1853 3617 1856
rect 3651 1853 3663 1887
rect 3605 1847 3663 1853
rect 4985 1887 5043 1893
rect 4985 1853 4997 1887
rect 5031 1853 5043 1887
rect 4985 1847 5043 1853
rect 2958 1776 2964 1828
rect 3016 1816 3022 1828
rect 5000 1816 5028 1847
rect 5166 1844 5172 1896
rect 5224 1884 5230 1896
rect 5261 1887 5319 1893
rect 5261 1884 5273 1887
rect 5224 1856 5273 1884
rect 5224 1844 5230 1856
rect 5261 1853 5273 1856
rect 5307 1853 5319 1887
rect 5261 1847 5319 1853
rect 5537 1887 5595 1893
rect 5537 1853 5549 1887
rect 5583 1884 5595 1887
rect 5902 1884 5908 1896
rect 5583 1856 5908 1884
rect 5583 1853 5595 1856
rect 5537 1847 5595 1853
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 6914 1844 6920 1896
rect 6972 1884 6978 1896
rect 7285 1887 7343 1893
rect 7285 1884 7297 1887
rect 6972 1856 7297 1884
rect 6972 1844 6978 1856
rect 7285 1853 7297 1856
rect 7331 1853 7343 1887
rect 7285 1847 7343 1853
rect 9398 1844 9404 1896
rect 9456 1884 9462 1896
rect 9861 1887 9919 1893
rect 9861 1884 9873 1887
rect 9456 1856 9873 1884
rect 9456 1844 9462 1856
rect 9861 1853 9873 1856
rect 9907 1853 9919 1887
rect 9861 1847 9919 1853
rect 11606 1844 11612 1896
rect 11664 1884 11670 1896
rect 12161 1887 12219 1893
rect 12161 1884 12173 1887
rect 11664 1856 12173 1884
rect 11664 1844 11670 1856
rect 12161 1853 12173 1856
rect 12207 1853 12219 1887
rect 12161 1847 12219 1853
rect 13538 1844 13544 1896
rect 13596 1884 13602 1896
rect 14093 1887 14151 1893
rect 14093 1884 14105 1887
rect 13596 1856 14105 1884
rect 13596 1844 13602 1856
rect 14093 1853 14105 1856
rect 14139 1853 14151 1887
rect 14093 1847 14151 1853
rect 16114 1844 16120 1896
rect 16172 1884 16178 1896
rect 16853 1887 16911 1893
rect 16853 1884 16865 1887
rect 16172 1856 16865 1884
rect 16172 1844 16178 1856
rect 16853 1853 16865 1856
rect 16899 1853 16911 1887
rect 16853 1847 16911 1853
rect 19610 1844 19616 1896
rect 19668 1884 19674 1896
rect 20257 1887 20315 1893
rect 20257 1884 20269 1887
rect 19668 1856 20269 1884
rect 19668 1844 19674 1856
rect 20257 1853 20269 1856
rect 20303 1853 20315 1887
rect 20257 1847 20315 1853
rect 21542 1844 21548 1896
rect 21600 1884 21606 1896
rect 22189 1887 22247 1893
rect 22189 1884 22201 1887
rect 21600 1856 22201 1884
rect 21600 1844 21606 1856
rect 22189 1853 22201 1856
rect 22235 1853 22247 1887
rect 22189 1847 22247 1853
rect 24302 1844 24308 1896
rect 24360 1884 24366 1896
rect 25041 1887 25099 1893
rect 25041 1884 25053 1887
rect 24360 1856 25053 1884
rect 24360 1844 24366 1856
rect 25041 1853 25053 1856
rect 25087 1853 25099 1887
rect 25041 1847 25099 1853
rect 28442 1844 28448 1896
rect 28500 1884 28506 1896
rect 29273 1887 29331 1893
rect 29273 1884 29285 1887
rect 28500 1856 29285 1884
rect 28500 1844 28506 1856
rect 29273 1853 29285 1856
rect 29319 1853 29331 1887
rect 29273 1847 29331 1853
rect 30650 1844 30656 1896
rect 30708 1884 30714 1896
rect 31481 1887 31539 1893
rect 31481 1884 31493 1887
rect 30708 1856 31493 1884
rect 30708 1844 30714 1856
rect 31481 1853 31493 1856
rect 31527 1853 31539 1887
rect 31481 1847 31539 1853
rect 31754 1844 31760 1896
rect 31812 1884 31818 1896
rect 32585 1887 32643 1893
rect 32585 1884 32597 1887
rect 31812 1856 32597 1884
rect 31812 1844 31818 1856
rect 32585 1853 32597 1856
rect 32631 1853 32643 1887
rect 32585 1847 32643 1853
rect 43438 1844 43444 1896
rect 43496 1884 43502 1896
rect 44361 1887 44419 1893
rect 44361 1884 44373 1887
rect 43496 1856 44373 1884
rect 43496 1844 43502 1856
rect 44361 1853 44373 1856
rect 44407 1853 44419 1887
rect 44361 1847 44419 1853
rect 44450 1844 44456 1896
rect 44508 1884 44514 1896
rect 45557 1887 45615 1893
rect 45557 1884 45569 1887
rect 44508 1856 45569 1884
rect 44508 1844 44514 1856
rect 45557 1853 45569 1856
rect 45603 1853 45615 1887
rect 45557 1847 45615 1853
rect 51074 1844 51080 1896
rect 51132 1884 51138 1896
rect 52273 1887 52331 1893
rect 52273 1884 52285 1887
rect 51132 1856 52285 1884
rect 51132 1844 51138 1856
rect 52273 1853 52285 1856
rect 52319 1853 52331 1887
rect 52273 1847 52331 1853
rect 3016 1788 5028 1816
rect 3016 1776 3022 1788
rect 3878 1748 3884 1760
rect 2700 1720 3884 1748
rect 3878 1708 3884 1720
rect 3936 1708 3942 1760
rect 1288 1658 68816 1680
rect 1288 1606 7262 1658
rect 7314 1606 19262 1658
rect 19314 1606 31262 1658
rect 31314 1606 43262 1658
rect 43314 1606 55262 1658
rect 55314 1606 67262 1658
rect 67314 1606 68816 1658
rect 1288 1584 68816 1606
rect 2222 1368 2228 1420
rect 2280 1408 2286 1420
rect 2280 1380 2636 1408
rect 2280 1368 2286 1380
rect 2133 1343 2191 1349
rect 2133 1309 2145 1343
rect 2179 1340 2191 1343
rect 2406 1340 2412 1352
rect 2179 1312 2412 1340
rect 2179 1309 2191 1312
rect 2133 1303 2191 1309
rect 2406 1300 2412 1312
rect 2464 1300 2470 1352
rect 2608 1340 2636 1380
rect 3142 1368 3148 1420
rect 3200 1408 3206 1420
rect 3602 1408 3608 1420
rect 3200 1380 3608 1408
rect 3200 1368 3206 1380
rect 3602 1368 3608 1380
rect 3660 1368 3666 1420
rect 26510 1368 26516 1420
rect 26568 1408 26574 1420
rect 27801 1411 27859 1417
rect 27801 1408 27813 1411
rect 26568 1380 27813 1408
rect 26568 1368 26574 1380
rect 27801 1377 27813 1380
rect 27847 1377 27859 1411
rect 27801 1371 27859 1377
rect 27890 1368 27896 1420
rect 27948 1408 27954 1420
rect 27948 1380 28212 1408
rect 27948 1368 27954 1380
rect 3053 1343 3111 1349
rect 3053 1340 3065 1343
rect 2608 1312 3065 1340
rect 3053 1309 3065 1312
rect 3099 1309 3111 1343
rect 3053 1303 3111 1309
rect 3786 1300 3792 1352
rect 3844 1340 3850 1352
rect 4709 1343 4767 1349
rect 4709 1340 4721 1343
rect 3844 1312 4721 1340
rect 3844 1300 3850 1312
rect 4709 1309 4721 1312
rect 4755 1309 4767 1343
rect 4709 1303 4767 1309
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 5537 1343 5595 1349
rect 5537 1340 5549 1343
rect 5040 1312 5549 1340
rect 5040 1300 5046 1312
rect 5537 1309 5549 1312
rect 5583 1309 5595 1343
rect 5537 1303 5595 1309
rect 5626 1300 5632 1352
rect 5684 1340 5690 1352
rect 5813 1343 5871 1349
rect 5813 1340 5825 1343
rect 5684 1312 5825 1340
rect 5684 1300 5690 1312
rect 5813 1309 5825 1312
rect 5859 1309 5871 1343
rect 5813 1303 5871 1309
rect 6638 1300 6644 1352
rect 6696 1340 6702 1352
rect 7193 1343 7251 1349
rect 7193 1340 7205 1343
rect 6696 1312 7205 1340
rect 6696 1300 6702 1312
rect 7193 1309 7205 1312
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 7466 1300 7472 1352
rect 7524 1340 7530 1352
rect 7837 1343 7895 1349
rect 7837 1340 7849 1343
rect 7524 1312 7849 1340
rect 7524 1300 7530 1312
rect 7837 1309 7849 1312
rect 7883 1309 7895 1343
rect 7837 1303 7895 1309
rect 9674 1300 9680 1352
rect 9732 1340 9738 1352
rect 10137 1343 10195 1349
rect 10137 1340 10149 1343
rect 9732 1312 10149 1340
rect 9732 1300 9738 1312
rect 10137 1309 10149 1312
rect 10183 1309 10195 1343
rect 10137 1303 10195 1309
rect 11330 1300 11336 1352
rect 11388 1340 11394 1352
rect 11977 1343 12035 1349
rect 11977 1340 11989 1343
rect 11388 1312 11989 1340
rect 11388 1300 11394 1312
rect 11977 1309 11989 1312
rect 12023 1309 12035 1343
rect 11977 1303 12035 1309
rect 12986 1300 12992 1352
rect 13044 1340 13050 1352
rect 13541 1343 13599 1349
rect 13541 1340 13553 1343
rect 13044 1312 13553 1340
rect 13044 1300 13050 1312
rect 13541 1309 13553 1312
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 13814 1300 13820 1352
rect 13872 1340 13878 1352
rect 14369 1343 14427 1349
rect 14369 1340 14381 1343
rect 13872 1312 14381 1340
rect 13872 1300 13878 1312
rect 14369 1309 14381 1312
rect 14415 1309 14427 1343
rect 14369 1303 14427 1309
rect 15746 1300 15752 1352
rect 15804 1340 15810 1352
rect 16301 1343 16359 1349
rect 16301 1340 16313 1343
rect 15804 1312 16313 1340
rect 15804 1300 15810 1312
rect 16301 1309 16313 1312
rect 16347 1309 16359 1343
rect 16301 1303 16359 1309
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 17497 1343 17555 1349
rect 17497 1340 17509 1343
rect 16908 1312 17509 1340
rect 16908 1300 16914 1312
rect 17497 1309 17509 1312
rect 17543 1309 17555 1343
rect 17497 1303 17555 1309
rect 17678 1300 17684 1352
rect 17736 1340 17742 1352
rect 18325 1343 18383 1349
rect 18325 1340 18337 1343
rect 17736 1312 18337 1340
rect 17736 1300 17742 1312
rect 18325 1309 18337 1312
rect 18371 1309 18383 1343
rect 18325 1303 18383 1309
rect 19426 1300 19432 1352
rect 19484 1340 19490 1352
rect 19981 1343 20039 1349
rect 19981 1340 19993 1343
rect 19484 1312 19993 1340
rect 19484 1300 19490 1312
rect 19981 1309 19993 1312
rect 20027 1309 20039 1343
rect 19981 1303 20039 1309
rect 20162 1300 20168 1352
rect 20220 1340 20226 1352
rect 20809 1343 20867 1349
rect 20809 1340 20821 1343
rect 20220 1312 20821 1340
rect 20220 1300 20226 1312
rect 20809 1309 20821 1312
rect 20855 1309 20867 1343
rect 20809 1303 20867 1309
rect 20990 1300 20996 1352
rect 21048 1340 21054 1352
rect 21637 1343 21695 1349
rect 21637 1340 21649 1343
rect 21048 1312 21649 1340
rect 21048 1300 21054 1312
rect 21637 1309 21649 1312
rect 21683 1309 21695 1343
rect 21637 1303 21695 1309
rect 22370 1300 22376 1352
rect 22428 1340 22434 1352
rect 23017 1343 23075 1349
rect 23017 1340 23029 1343
rect 22428 1312 23029 1340
rect 22428 1300 22434 1312
rect 23017 1309 23029 1312
rect 23063 1309 23075 1343
rect 23017 1303 23075 1309
rect 23474 1300 23480 1352
rect 23532 1340 23538 1352
rect 24213 1343 24271 1349
rect 24213 1340 24225 1343
rect 23532 1312 24225 1340
rect 23532 1300 23538 1312
rect 24213 1309 24225 1312
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 24854 1300 24860 1352
rect 24912 1340 24918 1352
rect 25593 1343 25651 1349
rect 25593 1340 25605 1343
rect 24912 1312 25605 1340
rect 24912 1300 24918 1312
rect 25593 1309 25605 1312
rect 25639 1309 25651 1343
rect 25593 1303 25651 1309
rect 25958 1300 25964 1352
rect 26016 1340 26022 1352
rect 26697 1343 26755 1349
rect 26697 1340 26709 1343
rect 26016 1312 26709 1340
rect 26016 1300 26022 1312
rect 26697 1309 26709 1312
rect 26743 1309 26755 1343
rect 26697 1303 26755 1309
rect 27338 1300 27344 1352
rect 27396 1340 27402 1352
rect 28077 1343 28135 1349
rect 28077 1340 28089 1343
rect 27396 1312 28089 1340
rect 27396 1300 27402 1312
rect 28077 1309 28089 1312
rect 28123 1309 28135 1343
rect 28184 1340 28212 1380
rect 38930 1368 38936 1420
rect 38988 1408 38994 1420
rect 40405 1411 40463 1417
rect 40405 1408 40417 1411
rect 38988 1380 40417 1408
rect 38988 1368 38994 1380
rect 40405 1377 40417 1380
rect 40451 1377 40463 1411
rect 40405 1371 40463 1377
rect 41414 1368 41420 1420
rect 41472 1408 41478 1420
rect 41472 1380 42012 1408
rect 41472 1368 41478 1380
rect 29181 1343 29239 1349
rect 29181 1340 29193 1343
rect 28184 1312 29193 1340
rect 28077 1303 28135 1309
rect 29181 1309 29193 1312
rect 29227 1309 29239 1343
rect 29181 1303 29239 1309
rect 29546 1300 29552 1352
rect 29604 1340 29610 1352
rect 30377 1343 30435 1349
rect 30377 1340 30389 1343
rect 29604 1312 30389 1340
rect 29604 1300 29610 1312
rect 30377 1309 30389 1312
rect 30423 1309 30435 1343
rect 30377 1303 30435 1309
rect 30926 1300 30932 1352
rect 30984 1340 30990 1352
rect 31757 1343 31815 1349
rect 31757 1340 31769 1343
rect 30984 1312 31769 1340
rect 30984 1300 30990 1312
rect 31757 1309 31769 1312
rect 31803 1309 31815 1343
rect 31757 1303 31815 1309
rect 32306 1300 32312 1352
rect 32364 1340 32370 1352
rect 33137 1343 33195 1349
rect 33137 1340 33149 1343
rect 32364 1312 33149 1340
rect 32364 1300 32370 1312
rect 33137 1309 33149 1312
rect 33183 1309 33195 1343
rect 33137 1303 33195 1309
rect 33226 1300 33232 1352
rect 33284 1340 33290 1352
rect 33965 1343 34023 1349
rect 33965 1340 33977 1343
rect 33284 1312 33977 1340
rect 33284 1300 33290 1312
rect 33965 1309 33977 1312
rect 34011 1309 34023 1343
rect 33965 1303 34023 1309
rect 34054 1300 34060 1352
rect 34112 1340 34118 1352
rect 34885 1343 34943 1349
rect 34885 1340 34897 1343
rect 34112 1312 34897 1340
rect 34112 1300 34118 1312
rect 34885 1309 34897 1312
rect 34931 1309 34943 1343
rect 35437 1343 35495 1349
rect 35437 1340 35449 1343
rect 34885 1303 34943 1309
rect 34992 1312 35449 1340
rect 1946 1232 1952 1284
rect 2004 1272 2010 1284
rect 2501 1275 2559 1281
rect 2501 1272 2513 1275
rect 2004 1244 2513 1272
rect 2004 1232 2010 1244
rect 2501 1241 2513 1244
rect 2547 1241 2559 1275
rect 3234 1272 3240 1284
rect 2501 1235 2559 1241
rect 2700 1244 3240 1272
rect 1854 1204 1860 1216
rect 1815 1176 1860 1204
rect 1854 1164 1860 1176
rect 1912 1164 1918 1216
rect 2409 1207 2467 1213
rect 2409 1173 2421 1207
rect 2455 1204 2467 1207
rect 2700 1204 2728 1244
rect 3234 1232 3240 1244
rect 3292 1232 3298 1284
rect 3510 1232 3516 1284
rect 3568 1272 3574 1284
rect 4433 1275 4491 1281
rect 4433 1272 4445 1275
rect 3568 1244 4445 1272
rect 3568 1232 3574 1244
rect 4433 1241 4445 1244
rect 4479 1241 4491 1275
rect 4433 1235 4491 1241
rect 4522 1232 4528 1284
rect 4580 1272 4586 1284
rect 6089 1275 6147 1281
rect 6089 1272 6101 1275
rect 4580 1244 6101 1272
rect 4580 1232 4586 1244
rect 6089 1241 6101 1244
rect 6135 1241 6147 1275
rect 6089 1235 6147 1241
rect 6178 1232 6184 1284
rect 6236 1272 6242 1284
rect 6917 1275 6975 1281
rect 6917 1272 6929 1275
rect 6236 1244 6929 1272
rect 6236 1232 6242 1244
rect 6917 1241 6929 1244
rect 6963 1241 6975 1275
rect 6917 1235 6975 1241
rect 7742 1232 7748 1284
rect 7800 1272 7806 1284
rect 8113 1275 8171 1281
rect 8113 1272 8125 1275
rect 7800 1244 8125 1272
rect 7800 1232 7806 1244
rect 8113 1241 8125 1244
rect 8159 1241 8171 1275
rect 8113 1235 8171 1241
rect 8294 1232 8300 1284
rect 8352 1272 8358 1284
rect 8757 1275 8815 1281
rect 8757 1272 8769 1275
rect 8352 1244 8769 1272
rect 8352 1232 8358 1244
rect 8757 1241 8769 1244
rect 8803 1241 8815 1275
rect 8757 1235 8815 1241
rect 8846 1232 8852 1284
rect 8904 1272 8910 1284
rect 9401 1275 9459 1281
rect 9401 1272 9413 1275
rect 8904 1244 9413 1272
rect 8904 1232 8910 1244
rect 9401 1241 9413 1244
rect 9447 1241 9459 1275
rect 9401 1235 9459 1241
rect 10226 1232 10232 1284
rect 10284 1272 10290 1284
rect 10689 1275 10747 1281
rect 10689 1272 10701 1275
rect 10284 1244 10701 1272
rect 10284 1232 10290 1244
rect 10689 1241 10701 1244
rect 10735 1241 10747 1275
rect 10689 1235 10747 1241
rect 10778 1232 10784 1284
rect 10836 1272 10842 1284
rect 11241 1275 11299 1281
rect 11241 1272 11253 1275
rect 10836 1244 11253 1272
rect 10836 1232 10842 1244
rect 11241 1241 11253 1244
rect 11287 1241 11299 1275
rect 11241 1235 11299 1241
rect 11882 1232 11888 1284
rect 11940 1272 11946 1284
rect 12437 1275 12495 1281
rect 12437 1272 12449 1275
rect 11940 1244 12449 1272
rect 11940 1232 11946 1244
rect 12437 1241 12449 1244
rect 12483 1241 12495 1275
rect 12437 1235 12495 1241
rect 12802 1232 12808 1284
rect 12860 1272 12866 1284
rect 13265 1275 13323 1281
rect 13265 1272 13277 1275
rect 12860 1244 13277 1272
rect 12860 1232 12866 1244
rect 13265 1241 13277 1244
rect 13311 1241 13323 1275
rect 13265 1235 13323 1241
rect 14090 1232 14096 1284
rect 14148 1272 14154 1284
rect 14645 1275 14703 1281
rect 14645 1272 14657 1275
rect 14148 1244 14657 1272
rect 14148 1232 14154 1244
rect 14645 1241 14657 1244
rect 14691 1241 14703 1275
rect 14645 1235 14703 1241
rect 14734 1232 14740 1284
rect 14792 1272 14798 1284
rect 15197 1275 15255 1281
rect 15197 1272 15209 1275
rect 14792 1244 15209 1272
rect 14792 1232 14798 1244
rect 15197 1241 15209 1244
rect 15243 1241 15255 1275
rect 15197 1235 15255 1241
rect 15286 1232 15292 1284
rect 15344 1272 15350 1284
rect 15344 1244 15792 1272
rect 15344 1232 15350 1244
rect 2455 1176 2728 1204
rect 2455 1173 2467 1176
rect 2409 1167 2467 1173
rect 2774 1164 2780 1216
rect 2832 1204 2838 1216
rect 3326 1204 3332 1216
rect 2832 1176 2877 1204
rect 3287 1176 3332 1204
rect 2832 1164 2838 1176
rect 3326 1164 3332 1176
rect 3384 1164 3390 1216
rect 3418 1164 3424 1216
rect 3476 1204 3482 1216
rect 3605 1207 3663 1213
rect 3605 1204 3617 1207
rect 3476 1176 3617 1204
rect 3476 1164 3482 1176
rect 3605 1173 3617 1176
rect 3651 1173 3663 1207
rect 3605 1167 3663 1173
rect 3694 1164 3700 1216
rect 3752 1204 3758 1216
rect 4157 1207 4215 1213
rect 4157 1204 4169 1207
rect 3752 1176 4169 1204
rect 3752 1164 3758 1176
rect 4157 1173 4169 1176
rect 4203 1173 4215 1207
rect 4157 1167 4215 1173
rect 4246 1164 4252 1216
rect 4304 1204 4310 1216
rect 4985 1207 5043 1213
rect 4985 1204 4997 1207
rect 4304 1176 4997 1204
rect 4304 1164 4310 1176
rect 4985 1173 4997 1176
rect 5031 1173 5043 1207
rect 4985 1167 5043 1173
rect 5074 1164 5080 1216
rect 5132 1204 5138 1216
rect 5261 1207 5319 1213
rect 5261 1204 5273 1207
rect 5132 1176 5273 1204
rect 5132 1164 5138 1176
rect 5261 1173 5273 1176
rect 5307 1173 5319 1207
rect 5261 1167 5319 1173
rect 6362 1164 6368 1216
rect 6420 1204 6426 1216
rect 6641 1207 6699 1213
rect 6641 1204 6653 1207
rect 6420 1176 6653 1204
rect 6420 1164 6426 1176
rect 6641 1173 6653 1176
rect 6687 1173 6699 1207
rect 6641 1167 6699 1173
rect 7374 1164 7380 1216
rect 7432 1204 7438 1216
rect 7561 1207 7619 1213
rect 7561 1204 7573 1207
rect 7432 1176 7573 1204
rect 7432 1164 7438 1176
rect 7561 1173 7573 1176
rect 7607 1173 7619 1207
rect 7561 1167 7619 1173
rect 8018 1164 8024 1216
rect 8076 1204 8082 1216
rect 8481 1207 8539 1213
rect 8481 1204 8493 1207
rect 8076 1176 8493 1204
rect 8076 1164 8082 1176
rect 8481 1173 8493 1176
rect 8527 1173 8539 1207
rect 8481 1167 8539 1173
rect 8570 1164 8576 1216
rect 8628 1204 8634 1216
rect 9125 1207 9183 1213
rect 9125 1204 9137 1207
rect 8628 1176 9137 1204
rect 8628 1164 8634 1176
rect 9125 1173 9137 1176
rect 9171 1173 9183 1207
rect 9125 1167 9183 1173
rect 9214 1164 9220 1216
rect 9272 1204 9278 1216
rect 9677 1207 9735 1213
rect 9677 1204 9689 1207
rect 9272 1176 9689 1204
rect 9272 1164 9278 1176
rect 9677 1173 9689 1176
rect 9723 1173 9735 1207
rect 9677 1167 9735 1173
rect 9950 1164 9956 1216
rect 10008 1204 10014 1216
rect 10413 1207 10471 1213
rect 10413 1204 10425 1207
rect 10008 1176 10425 1204
rect 10008 1164 10014 1176
rect 10413 1173 10425 1176
rect 10459 1173 10471 1207
rect 10413 1167 10471 1173
rect 10502 1164 10508 1216
rect 10560 1204 10566 1216
rect 10965 1207 11023 1213
rect 10965 1204 10977 1207
rect 10560 1176 10977 1204
rect 10560 1164 10566 1176
rect 10965 1173 10977 1176
rect 11011 1173 11023 1207
rect 10965 1167 11023 1173
rect 11054 1164 11060 1216
rect 11112 1204 11118 1216
rect 11701 1207 11759 1213
rect 11701 1204 11713 1207
rect 11112 1176 11713 1204
rect 11112 1164 11118 1176
rect 11701 1173 11713 1176
rect 11747 1173 11759 1207
rect 11701 1167 11759 1173
rect 12158 1164 12164 1216
rect 12216 1204 12222 1216
rect 12713 1207 12771 1213
rect 12713 1204 12725 1207
rect 12216 1176 12725 1204
rect 12216 1164 12222 1176
rect 12713 1173 12725 1176
rect 12759 1173 12771 1207
rect 12713 1167 12771 1173
rect 12894 1164 12900 1216
rect 12952 1204 12958 1216
rect 12989 1207 13047 1213
rect 12989 1204 13001 1207
rect 12952 1176 13001 1204
rect 12952 1164 12958 1176
rect 12989 1173 13001 1176
rect 13035 1173 13047 1207
rect 12989 1167 13047 1173
rect 13446 1164 13452 1216
rect 13504 1204 13510 1216
rect 13817 1207 13875 1213
rect 13817 1204 13829 1207
rect 13504 1176 13829 1204
rect 13504 1164 13510 1176
rect 13817 1173 13829 1176
rect 13863 1173 13875 1207
rect 13817 1167 13875 1173
rect 14366 1164 14372 1216
rect 14424 1204 14430 1216
rect 14921 1207 14979 1213
rect 14921 1204 14933 1207
rect 14424 1176 14933 1204
rect 14424 1164 14430 1176
rect 14921 1173 14933 1176
rect 14967 1173 14979 1207
rect 14921 1167 14979 1173
rect 15010 1164 15016 1216
rect 15068 1204 15074 1216
rect 15764 1213 15792 1244
rect 16574 1232 16580 1284
rect 16632 1272 16638 1284
rect 17221 1275 17279 1281
rect 17221 1272 17233 1275
rect 16632 1244 17233 1272
rect 16632 1232 16638 1244
rect 17221 1241 17233 1244
rect 17267 1241 17279 1275
rect 17221 1235 17279 1241
rect 17402 1232 17408 1284
rect 17460 1272 17466 1284
rect 17460 1244 17908 1272
rect 17460 1232 17466 1244
rect 15473 1207 15531 1213
rect 15473 1204 15485 1207
rect 15068 1176 15485 1204
rect 15068 1164 15074 1176
rect 15473 1173 15485 1176
rect 15519 1173 15531 1207
rect 15473 1167 15531 1173
rect 15749 1207 15807 1213
rect 15749 1173 15761 1207
rect 15795 1173 15807 1207
rect 16022 1204 16028 1216
rect 15983 1176 16028 1204
rect 15749 1167 15807 1173
rect 16022 1164 16028 1176
rect 16080 1164 16086 1216
rect 16390 1164 16396 1216
rect 16448 1204 16454 1216
rect 16853 1207 16911 1213
rect 16853 1204 16865 1207
rect 16448 1176 16865 1204
rect 16448 1164 16454 1176
rect 16853 1173 16865 1176
rect 16899 1173 16911 1207
rect 16853 1167 16911 1173
rect 17126 1164 17132 1216
rect 17184 1204 17190 1216
rect 17773 1207 17831 1213
rect 17773 1204 17785 1207
rect 17184 1176 17785 1204
rect 17184 1164 17190 1176
rect 17773 1173 17785 1176
rect 17819 1173 17831 1207
rect 17880 1204 17908 1244
rect 17954 1232 17960 1284
rect 18012 1272 18018 1284
rect 18601 1275 18659 1281
rect 18601 1272 18613 1275
rect 18012 1244 18613 1272
rect 18012 1232 18018 1244
rect 18601 1241 18613 1244
rect 18647 1241 18659 1275
rect 18601 1235 18659 1241
rect 19058 1232 19064 1284
rect 19116 1272 19122 1284
rect 19705 1275 19763 1281
rect 19705 1272 19717 1275
rect 19116 1244 19717 1272
rect 19116 1232 19122 1244
rect 19705 1241 19717 1244
rect 19751 1241 19763 1275
rect 19705 1235 19763 1241
rect 19886 1232 19892 1284
rect 19944 1272 19950 1284
rect 20533 1275 20591 1281
rect 20533 1272 20545 1275
rect 19944 1244 20545 1272
rect 19944 1232 19950 1244
rect 20533 1241 20545 1244
rect 20579 1241 20591 1275
rect 20533 1235 20591 1241
rect 20714 1232 20720 1284
rect 20772 1272 20778 1284
rect 21361 1275 21419 1281
rect 21361 1272 21373 1275
rect 20772 1244 21373 1272
rect 20772 1232 20778 1244
rect 21361 1241 21373 1244
rect 21407 1241 21419 1275
rect 21361 1235 21419 1241
rect 21818 1232 21824 1284
rect 21876 1272 21882 1284
rect 22465 1275 22523 1281
rect 22465 1272 22477 1275
rect 21876 1244 22477 1272
rect 21876 1232 21882 1244
rect 22465 1241 22477 1244
rect 22511 1241 22523 1275
rect 22465 1235 22523 1241
rect 22646 1232 22652 1284
rect 22704 1272 22710 1284
rect 22704 1244 22876 1272
rect 22704 1232 22710 1244
rect 18049 1207 18107 1213
rect 18049 1204 18061 1207
rect 17880 1176 18061 1204
rect 17773 1167 17831 1173
rect 18049 1173 18061 1176
rect 18095 1173 18107 1207
rect 18049 1167 18107 1173
rect 18230 1164 18236 1216
rect 18288 1204 18294 1216
rect 18877 1207 18935 1213
rect 18877 1204 18889 1207
rect 18288 1176 18889 1204
rect 18288 1164 18294 1176
rect 18877 1173 18889 1176
rect 18923 1173 18935 1207
rect 18877 1167 18935 1173
rect 18966 1164 18972 1216
rect 19024 1204 19030 1216
rect 19429 1207 19487 1213
rect 19429 1204 19441 1207
rect 19024 1176 19441 1204
rect 19024 1164 19030 1176
rect 19429 1173 19441 1176
rect 19475 1173 19487 1207
rect 20254 1204 20260 1216
rect 20215 1176 20260 1204
rect 19429 1167 19487 1173
rect 20254 1164 20260 1176
rect 20312 1164 20318 1216
rect 20622 1164 20628 1216
rect 20680 1204 20686 1216
rect 21085 1207 21143 1213
rect 21085 1204 21097 1207
rect 20680 1176 21097 1204
rect 20680 1164 20686 1176
rect 21085 1173 21097 1176
rect 21131 1173 21143 1207
rect 21085 1167 21143 1173
rect 21266 1164 21272 1216
rect 21324 1204 21330 1216
rect 22005 1207 22063 1213
rect 22005 1204 22017 1207
rect 21324 1176 22017 1204
rect 21324 1164 21330 1176
rect 22005 1173 22017 1176
rect 22051 1173 22063 1207
rect 22005 1167 22063 1173
rect 22094 1164 22100 1216
rect 22152 1204 22158 1216
rect 22741 1207 22799 1213
rect 22741 1204 22753 1207
rect 22152 1176 22753 1204
rect 22152 1164 22158 1176
rect 22741 1173 22753 1176
rect 22787 1173 22799 1207
rect 22848 1204 22876 1244
rect 22922 1232 22928 1284
rect 22980 1272 22986 1284
rect 23569 1275 23627 1281
rect 23569 1272 23581 1275
rect 22980 1244 23581 1272
rect 22980 1232 22986 1244
rect 23569 1241 23581 1244
rect 23615 1241 23627 1275
rect 23569 1235 23627 1241
rect 23750 1232 23756 1284
rect 23808 1272 23814 1284
rect 24581 1275 24639 1281
rect 24581 1272 24593 1275
rect 23808 1244 24593 1272
rect 23808 1232 23814 1244
rect 24581 1241 24593 1244
rect 24627 1241 24639 1275
rect 24581 1235 24639 1241
rect 24670 1232 24676 1284
rect 24728 1272 24734 1284
rect 25317 1275 25375 1281
rect 25317 1272 25329 1275
rect 24728 1244 25329 1272
rect 24728 1232 24734 1244
rect 25317 1241 25329 1244
rect 25363 1241 25375 1275
rect 25317 1235 25375 1241
rect 25682 1232 25688 1284
rect 25740 1272 25746 1284
rect 26421 1275 26479 1281
rect 26421 1272 26433 1275
rect 25740 1244 26433 1272
rect 25740 1232 25746 1244
rect 26421 1241 26433 1244
rect 26467 1241 26479 1275
rect 26421 1235 26479 1241
rect 26786 1232 26792 1284
rect 26844 1272 26850 1284
rect 27525 1275 27583 1281
rect 27525 1272 27537 1275
rect 26844 1244 27537 1272
rect 26844 1232 26850 1244
rect 27525 1241 27537 1244
rect 27571 1241 27583 1275
rect 27525 1235 27583 1241
rect 27614 1232 27620 1284
rect 27672 1272 27678 1284
rect 27672 1244 27936 1272
rect 27672 1232 27678 1244
rect 23293 1207 23351 1213
rect 23293 1204 23305 1207
rect 22848 1176 23305 1204
rect 22741 1167 22799 1173
rect 23293 1173 23305 1176
rect 23339 1173 23351 1207
rect 23293 1167 23351 1173
rect 23382 1164 23388 1216
rect 23440 1204 23446 1216
rect 23937 1207 23995 1213
rect 23937 1204 23949 1207
rect 23440 1176 23949 1204
rect 23440 1164 23446 1176
rect 23937 1173 23949 1176
rect 23983 1173 23995 1207
rect 23937 1167 23995 1173
rect 24026 1164 24032 1216
rect 24084 1204 24090 1216
rect 24857 1207 24915 1213
rect 24857 1204 24869 1207
rect 24084 1176 24869 1204
rect 24084 1164 24090 1176
rect 24857 1173 24869 1176
rect 24903 1173 24915 1207
rect 24857 1167 24915 1173
rect 25130 1164 25136 1216
rect 25188 1204 25194 1216
rect 25869 1207 25927 1213
rect 25869 1204 25881 1207
rect 25188 1176 25881 1204
rect 25188 1164 25194 1176
rect 25869 1173 25881 1176
rect 25915 1173 25927 1207
rect 26142 1204 26148 1216
rect 26103 1176 26148 1204
rect 25869 1167 25927 1173
rect 26142 1164 26148 1176
rect 26200 1164 26206 1216
rect 26234 1164 26240 1216
rect 26292 1204 26298 1216
rect 27157 1207 27215 1213
rect 27157 1204 27169 1207
rect 26292 1176 27169 1204
rect 26292 1164 26298 1176
rect 27157 1173 27169 1176
rect 27203 1173 27215 1207
rect 27908 1204 27936 1244
rect 28166 1232 28172 1284
rect 28224 1272 28230 1284
rect 28905 1275 28963 1281
rect 28905 1272 28917 1275
rect 28224 1244 28917 1272
rect 28224 1232 28230 1244
rect 28905 1241 28917 1244
rect 28951 1241 28963 1275
rect 28905 1235 28963 1241
rect 28994 1232 29000 1284
rect 29052 1272 29058 1284
rect 29825 1275 29883 1281
rect 29825 1272 29837 1275
rect 29052 1244 29837 1272
rect 29052 1232 29058 1244
rect 29825 1241 29837 1244
rect 29871 1241 29883 1275
rect 29825 1235 29883 1241
rect 29914 1232 29920 1284
rect 29972 1272 29978 1284
rect 30653 1275 30711 1281
rect 30653 1272 30665 1275
rect 29972 1244 30665 1272
rect 29972 1232 29978 1244
rect 30653 1241 30665 1244
rect 30699 1241 30711 1275
rect 31205 1275 31263 1281
rect 31205 1272 31217 1275
rect 30653 1235 30711 1241
rect 30760 1244 31217 1272
rect 28353 1207 28411 1213
rect 28353 1204 28365 1207
rect 27908 1176 28365 1204
rect 27157 1167 27215 1173
rect 28353 1173 28365 1176
rect 28399 1173 28411 1207
rect 28626 1204 28632 1216
rect 28587 1176 28632 1204
rect 28353 1167 28411 1173
rect 28626 1164 28632 1176
rect 28684 1164 28690 1216
rect 28718 1164 28724 1216
rect 28776 1204 28782 1216
rect 30101 1207 30159 1213
rect 30101 1204 30113 1207
rect 28776 1176 30113 1204
rect 28776 1164 28782 1176
rect 30101 1173 30113 1176
rect 30147 1173 30159 1207
rect 30101 1167 30159 1173
rect 30374 1164 30380 1216
rect 30432 1204 30438 1216
rect 30760 1204 30788 1244
rect 31205 1241 31217 1244
rect 31251 1241 31263 1275
rect 31205 1235 31263 1241
rect 32030 1232 32036 1284
rect 32088 1272 32094 1284
rect 32861 1275 32919 1281
rect 32861 1272 32873 1275
rect 32088 1244 32873 1272
rect 32088 1232 32094 1244
rect 32861 1241 32873 1244
rect 32907 1241 32919 1275
rect 32861 1235 32919 1241
rect 32950 1232 32956 1284
rect 33008 1272 33014 1284
rect 33689 1275 33747 1281
rect 33689 1272 33701 1275
rect 33008 1244 33701 1272
rect 33008 1232 33014 1244
rect 33689 1241 33701 1244
rect 33735 1241 33747 1275
rect 33689 1235 33747 1241
rect 33778 1232 33784 1284
rect 33836 1272 33842 1284
rect 34517 1275 34575 1281
rect 34517 1272 34529 1275
rect 33836 1244 34529 1272
rect 33836 1232 33842 1244
rect 34517 1241 34529 1244
rect 34563 1241 34575 1275
rect 34517 1235 34575 1241
rect 34606 1232 34612 1284
rect 34664 1272 34670 1284
rect 34992 1272 35020 1312
rect 35437 1309 35449 1312
rect 35483 1309 35495 1343
rect 35437 1303 35495 1309
rect 35618 1300 35624 1352
rect 35676 1340 35682 1352
rect 36541 1343 36599 1349
rect 36541 1340 36553 1343
rect 35676 1312 36553 1340
rect 35676 1300 35682 1312
rect 36541 1309 36553 1312
rect 36587 1309 36599 1343
rect 36541 1303 36599 1309
rect 36630 1300 36636 1352
rect 36688 1340 36694 1352
rect 37461 1343 37519 1349
rect 37461 1340 37473 1343
rect 36688 1312 37473 1340
rect 36688 1300 36694 1312
rect 37461 1309 37473 1312
rect 37507 1309 37519 1343
rect 37461 1303 37519 1309
rect 37550 1300 37556 1352
rect 37608 1340 37614 1352
rect 38289 1343 38347 1349
rect 38289 1340 38301 1343
rect 37608 1312 38301 1340
rect 37608 1300 37614 1312
rect 38289 1309 38301 1312
rect 38335 1309 38347 1343
rect 38289 1303 38347 1309
rect 38378 1300 38384 1352
rect 38436 1340 38442 1352
rect 39117 1343 39175 1349
rect 39117 1340 39129 1343
rect 38436 1312 39129 1340
rect 38436 1300 38442 1312
rect 39117 1309 39129 1312
rect 39163 1309 39175 1343
rect 39117 1303 39175 1309
rect 39482 1300 39488 1352
rect 39540 1340 39546 1352
rect 40681 1343 40739 1349
rect 40681 1340 40693 1343
rect 39540 1312 40693 1340
rect 39540 1300 39546 1312
rect 40681 1309 40693 1312
rect 40727 1309 40739 1343
rect 40681 1303 40739 1309
rect 40770 1300 40776 1352
rect 40828 1340 40834 1352
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 40828 1312 41797 1340
rect 40828 1300 40834 1312
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41984 1340 42012 1380
rect 45830 1368 45836 1420
rect 45888 1408 45894 1420
rect 46937 1411 46995 1417
rect 46937 1408 46949 1411
rect 45888 1380 46949 1408
rect 45888 1368 45894 1380
rect 46937 1377 46949 1380
rect 46983 1377 46995 1411
rect 46937 1371 46995 1377
rect 47394 1368 47400 1420
rect 47452 1408 47458 1420
rect 47452 1380 47992 1408
rect 47452 1368 47458 1380
rect 42889 1343 42947 1349
rect 42889 1340 42901 1343
rect 41984 1312 42901 1340
rect 41785 1303 41843 1309
rect 42889 1309 42901 1312
rect 42935 1309 42947 1343
rect 42889 1303 42947 1309
rect 43070 1300 43076 1352
rect 43128 1340 43134 1352
rect 44361 1343 44419 1349
rect 44361 1340 44373 1343
rect 43128 1312 44373 1340
rect 43128 1300 43134 1312
rect 44361 1309 44373 1312
rect 44407 1309 44419 1343
rect 45189 1343 45247 1349
rect 45189 1340 45201 1343
rect 44361 1303 44419 1309
rect 44468 1312 45201 1340
rect 34664 1244 35020 1272
rect 34664 1232 34670 1244
rect 35342 1232 35348 1284
rect 35400 1272 35406 1284
rect 36265 1275 36323 1281
rect 36265 1272 36277 1275
rect 35400 1244 36277 1272
rect 35400 1232 35406 1244
rect 36265 1241 36277 1244
rect 36311 1241 36323 1275
rect 36265 1235 36323 1241
rect 36354 1232 36360 1284
rect 36412 1272 36418 1284
rect 37093 1275 37151 1281
rect 37093 1272 37105 1275
rect 36412 1244 37105 1272
rect 36412 1232 36418 1244
rect 37093 1241 37105 1244
rect 37139 1241 37151 1275
rect 37093 1235 37151 1241
rect 37366 1232 37372 1284
rect 37424 1272 37430 1284
rect 38013 1275 38071 1281
rect 38013 1272 38025 1275
rect 37424 1244 38025 1272
rect 37424 1232 37430 1244
rect 38013 1241 38025 1244
rect 38059 1241 38071 1275
rect 38013 1235 38071 1241
rect 38102 1232 38108 1284
rect 38160 1272 38166 1284
rect 38841 1275 38899 1281
rect 38841 1272 38853 1275
rect 38160 1244 38853 1272
rect 38160 1232 38166 1244
rect 38841 1241 38853 1244
rect 38887 1241 38899 1275
rect 38841 1235 38899 1241
rect 39206 1232 39212 1284
rect 39264 1272 39270 1284
rect 40129 1275 40187 1281
rect 40129 1272 40141 1275
rect 39264 1244 40141 1272
rect 39264 1232 39270 1244
rect 40129 1241 40141 1244
rect 40175 1241 40187 1275
rect 40957 1275 41015 1281
rect 40957 1272 40969 1275
rect 40129 1235 40187 1241
rect 40236 1244 40969 1272
rect 30432 1176 30788 1204
rect 30432 1164 30438 1176
rect 30834 1164 30840 1216
rect 30892 1204 30898 1216
rect 30929 1207 30987 1213
rect 30929 1204 30941 1207
rect 30892 1176 30941 1204
rect 30892 1164 30898 1176
rect 30929 1173 30941 1176
rect 30975 1173 30987 1207
rect 30929 1167 30987 1173
rect 31018 1164 31024 1216
rect 31076 1204 31082 1216
rect 31481 1207 31539 1213
rect 31481 1204 31493 1207
rect 31076 1176 31493 1204
rect 31076 1164 31082 1176
rect 31481 1173 31493 1176
rect 31527 1173 31539 1207
rect 31481 1167 31539 1173
rect 31570 1164 31576 1216
rect 31628 1204 31634 1216
rect 32309 1207 32367 1213
rect 32309 1204 32321 1207
rect 31628 1176 32321 1204
rect 31628 1164 31634 1176
rect 32309 1173 32321 1176
rect 32355 1173 32367 1207
rect 32309 1167 32367 1173
rect 32398 1164 32404 1216
rect 32456 1204 32462 1216
rect 32585 1207 32643 1213
rect 32585 1204 32597 1207
rect 32456 1176 32597 1204
rect 32456 1164 32462 1176
rect 32585 1173 32597 1176
rect 32631 1173 32643 1207
rect 32585 1167 32643 1173
rect 32674 1164 32680 1216
rect 32732 1204 32738 1216
rect 33413 1207 33471 1213
rect 33413 1204 33425 1207
rect 32732 1176 33425 1204
rect 32732 1164 32738 1176
rect 33413 1173 33425 1176
rect 33459 1173 33471 1207
rect 33413 1167 33471 1173
rect 33502 1164 33508 1216
rect 33560 1204 33566 1216
rect 34241 1207 34299 1213
rect 34241 1204 34253 1207
rect 33560 1176 34253 1204
rect 33560 1164 33566 1176
rect 34241 1173 34253 1176
rect 34287 1173 34299 1207
rect 34241 1167 34299 1173
rect 34330 1164 34336 1216
rect 34388 1204 34394 1216
rect 35161 1207 35219 1213
rect 35161 1204 35173 1207
rect 34388 1176 35173 1204
rect 34388 1164 34394 1176
rect 35161 1173 35173 1176
rect 35207 1173 35219 1207
rect 35710 1204 35716 1216
rect 35671 1176 35716 1204
rect 35161 1167 35219 1173
rect 35710 1164 35716 1176
rect 35768 1164 35774 1216
rect 35802 1164 35808 1216
rect 35860 1204 35866 1216
rect 35989 1207 36047 1213
rect 35989 1204 36001 1207
rect 35860 1176 36001 1204
rect 35860 1164 35866 1176
rect 35989 1173 36001 1176
rect 36035 1173 36047 1207
rect 35989 1167 36047 1173
rect 36078 1164 36084 1216
rect 36136 1204 36142 1216
rect 36817 1207 36875 1213
rect 36817 1204 36829 1207
rect 36136 1176 36829 1204
rect 36136 1164 36142 1176
rect 36817 1173 36829 1176
rect 36863 1173 36875 1207
rect 36817 1167 36875 1173
rect 36906 1164 36912 1216
rect 36964 1204 36970 1216
rect 37737 1207 37795 1213
rect 37737 1204 37749 1207
rect 36964 1176 37749 1204
rect 36964 1164 36970 1176
rect 37737 1173 37749 1176
rect 37783 1173 37795 1207
rect 37737 1167 37795 1173
rect 37826 1164 37832 1216
rect 37884 1204 37890 1216
rect 38565 1207 38623 1213
rect 38565 1204 38577 1207
rect 37884 1176 38577 1204
rect 37884 1164 37890 1176
rect 38565 1173 38577 1176
rect 38611 1173 38623 1207
rect 38565 1167 38623 1173
rect 38654 1164 38660 1216
rect 38712 1204 38718 1216
rect 39393 1207 39451 1213
rect 39393 1204 39405 1207
rect 38712 1176 39405 1204
rect 38712 1164 38718 1176
rect 39393 1173 39405 1176
rect 39439 1173 39451 1207
rect 39666 1204 39672 1216
rect 39627 1176 39672 1204
rect 39393 1167 39451 1173
rect 39666 1164 39672 1176
rect 39724 1164 39730 1216
rect 39758 1164 39764 1216
rect 39816 1204 39822 1216
rect 40236 1204 40264 1244
rect 40957 1241 40969 1244
rect 41003 1241 41015 1275
rect 41509 1275 41567 1281
rect 41509 1272 41521 1275
rect 40957 1235 41015 1241
rect 41064 1244 41521 1272
rect 39816 1176 40264 1204
rect 39816 1164 39822 1176
rect 40494 1164 40500 1216
rect 40552 1204 40558 1216
rect 41064 1204 41092 1244
rect 41509 1241 41521 1244
rect 41555 1241 41567 1275
rect 41509 1235 41567 1241
rect 42518 1232 42524 1284
rect 42576 1272 42582 1284
rect 43533 1275 43591 1281
rect 43533 1272 43545 1275
rect 42576 1244 43545 1272
rect 42576 1232 42582 1244
rect 43533 1241 43545 1244
rect 43579 1241 43591 1275
rect 43533 1235 43591 1241
rect 43622 1232 43628 1284
rect 43680 1272 43686 1284
rect 44468 1272 44496 1312
rect 45189 1309 45201 1312
rect 45235 1309 45247 1343
rect 45189 1303 45247 1309
rect 45278 1300 45284 1352
rect 45336 1340 45342 1352
rect 46385 1343 46443 1349
rect 46385 1340 46397 1343
rect 45336 1312 46397 1340
rect 45336 1300 45342 1312
rect 46385 1309 46397 1312
rect 46431 1309 46443 1343
rect 46385 1303 46443 1309
rect 46474 1300 46480 1352
rect 46532 1340 46538 1352
rect 47765 1343 47823 1349
rect 47765 1340 47777 1343
rect 46532 1312 47777 1340
rect 46532 1300 46538 1312
rect 47765 1309 47777 1312
rect 47811 1309 47823 1343
rect 47964 1340 47992 1380
rect 48866 1368 48872 1420
rect 48924 1408 48930 1420
rect 48924 1380 49832 1408
rect 48924 1368 48930 1380
rect 48593 1343 48651 1349
rect 48593 1340 48605 1343
rect 47964 1312 48605 1340
rect 47765 1303 47823 1309
rect 48593 1309 48605 1312
rect 48639 1309 48651 1343
rect 48593 1303 48651 1309
rect 48682 1300 48688 1352
rect 48740 1340 48746 1352
rect 49697 1343 49755 1349
rect 49697 1340 49709 1343
rect 48740 1312 49709 1340
rect 48740 1300 48746 1312
rect 49697 1309 49709 1312
rect 49743 1309 49755 1343
rect 49804 1340 49832 1380
rect 49878 1368 49884 1420
rect 49936 1408 49942 1420
rect 49936 1380 50568 1408
rect 49936 1368 49942 1380
rect 50341 1343 50399 1349
rect 50341 1340 50353 1343
rect 49804 1312 50353 1340
rect 49697 1303 49755 1309
rect 50341 1309 50353 1312
rect 50387 1309 50399 1343
rect 50540 1340 50568 1380
rect 50798 1368 50804 1420
rect 50856 1408 50862 1420
rect 52273 1411 52331 1417
rect 52273 1408 52285 1411
rect 50856 1380 52285 1408
rect 50856 1368 50862 1380
rect 52273 1377 52285 1380
rect 52319 1377 52331 1411
rect 52273 1371 52331 1377
rect 51169 1343 51227 1349
rect 51169 1340 51181 1343
rect 50540 1312 51181 1340
rect 50341 1303 50399 1309
rect 51169 1309 51181 1312
rect 51215 1309 51227 1343
rect 51169 1303 51227 1309
rect 51626 1300 51632 1352
rect 51684 1340 51690 1352
rect 52917 1343 52975 1349
rect 52917 1340 52929 1343
rect 51684 1312 52929 1340
rect 51684 1300 51690 1312
rect 52917 1309 52929 1312
rect 52963 1309 52975 1343
rect 52917 1303 52975 1309
rect 53006 1300 53012 1352
rect 53064 1340 53070 1352
rect 54021 1343 54079 1349
rect 54021 1340 54033 1343
rect 53064 1312 54033 1340
rect 53064 1300 53070 1312
rect 54021 1309 54033 1312
rect 54067 1309 54079 1343
rect 54021 1303 54079 1309
rect 54662 1300 54668 1352
rect 54720 1340 54726 1352
rect 55769 1343 55827 1349
rect 55769 1340 55781 1343
rect 54720 1312 55781 1340
rect 54720 1300 54726 1312
rect 55769 1309 55781 1312
rect 55815 1309 55827 1343
rect 55769 1303 55827 1309
rect 43680 1244 44496 1272
rect 43680 1232 43686 1244
rect 44726 1232 44732 1284
rect 44784 1272 44790 1284
rect 45833 1275 45891 1281
rect 45833 1272 45845 1275
rect 44784 1244 45845 1272
rect 44784 1232 44790 1244
rect 45833 1241 45845 1244
rect 45879 1241 45891 1275
rect 46661 1275 46719 1281
rect 46661 1272 46673 1275
rect 45833 1235 45891 1241
rect 45940 1244 46673 1272
rect 41230 1204 41236 1216
rect 40552 1176 41092 1204
rect 41191 1176 41236 1204
rect 40552 1164 40558 1176
rect 41230 1164 41236 1176
rect 41288 1164 41294 1216
rect 41322 1164 41328 1216
rect 41380 1204 41386 1216
rect 42061 1207 42119 1213
rect 42061 1204 42073 1207
rect 41380 1176 42073 1204
rect 41380 1164 41386 1176
rect 42061 1173 42073 1176
rect 42107 1173 42119 1207
rect 42610 1204 42616 1216
rect 42571 1176 42616 1204
rect 42061 1167 42119 1173
rect 42610 1164 42616 1176
rect 42668 1164 42674 1216
rect 42794 1164 42800 1216
rect 42852 1204 42858 1216
rect 43165 1207 43223 1213
rect 43165 1204 43177 1207
rect 42852 1176 43177 1204
rect 42852 1164 42858 1176
rect 43165 1173 43177 1176
rect 43211 1173 43223 1207
rect 43806 1204 43812 1216
rect 43767 1176 43812 1204
rect 43165 1167 43223 1173
rect 43806 1164 43812 1176
rect 43864 1164 43870 1216
rect 44082 1204 44088 1216
rect 44043 1176 44088 1204
rect 44082 1164 44088 1176
rect 44140 1164 44146 1216
rect 44634 1204 44640 1216
rect 44595 1176 44640 1204
rect 44634 1164 44640 1176
rect 44692 1164 44698 1216
rect 45462 1204 45468 1216
rect 45423 1176 45468 1204
rect 45462 1164 45468 1176
rect 45520 1164 45526 1216
rect 45554 1164 45560 1216
rect 45612 1204 45618 1216
rect 45940 1204 45968 1244
rect 46661 1241 46673 1244
rect 46707 1241 46719 1275
rect 47213 1275 47271 1281
rect 47213 1272 47225 1275
rect 46661 1235 46719 1241
rect 46860 1244 47225 1272
rect 46106 1204 46112 1216
rect 45612 1176 45968 1204
rect 46067 1176 46112 1204
rect 45612 1164 45618 1176
rect 46106 1164 46112 1176
rect 46164 1164 46170 1216
rect 46198 1164 46204 1216
rect 46256 1204 46262 1216
rect 46860 1204 46888 1244
rect 47213 1241 47225 1244
rect 47259 1241 47271 1275
rect 47213 1235 47271 1241
rect 47302 1232 47308 1284
rect 47360 1272 47366 1284
rect 48317 1275 48375 1281
rect 48317 1272 48329 1275
rect 47360 1244 48329 1272
rect 47360 1232 47366 1244
rect 48317 1241 48329 1244
rect 48363 1241 48375 1275
rect 48317 1235 48375 1241
rect 48406 1232 48412 1284
rect 48464 1272 48470 1284
rect 49421 1275 49479 1281
rect 49421 1272 49433 1275
rect 48464 1244 49433 1272
rect 48464 1232 48470 1244
rect 49421 1241 49433 1244
rect 49467 1241 49479 1275
rect 49421 1235 49479 1241
rect 49510 1232 49516 1284
rect 49568 1272 49574 1284
rect 50617 1275 50675 1281
rect 50617 1272 50629 1275
rect 49568 1244 50629 1272
rect 49568 1232 49574 1244
rect 50617 1241 50629 1244
rect 50663 1241 50675 1275
rect 50617 1235 50675 1241
rect 50724 1244 51120 1272
rect 46256 1176 46888 1204
rect 46256 1164 46262 1176
rect 46934 1164 46940 1216
rect 46992 1204 46998 1216
rect 48041 1207 48099 1213
rect 48041 1204 48053 1207
rect 46992 1176 48053 1204
rect 46992 1164 46998 1176
rect 48041 1173 48053 1176
rect 48087 1173 48099 1207
rect 48041 1167 48099 1173
rect 48130 1164 48136 1216
rect 48188 1204 48194 1216
rect 48869 1207 48927 1213
rect 48869 1204 48881 1207
rect 48188 1176 48881 1204
rect 48188 1164 48194 1176
rect 48869 1173 48881 1176
rect 48915 1173 48927 1207
rect 49142 1204 49148 1216
rect 49103 1176 49148 1204
rect 48869 1167 48927 1173
rect 49142 1164 49148 1176
rect 49200 1164 49206 1216
rect 49970 1204 49976 1216
rect 49931 1176 49976 1204
rect 49970 1164 49976 1176
rect 50028 1164 50034 1216
rect 50062 1164 50068 1216
rect 50120 1204 50126 1216
rect 50724 1204 50752 1244
rect 50890 1204 50896 1216
rect 50120 1176 50752 1204
rect 50851 1176 50896 1204
rect 50120 1164 50126 1176
rect 50890 1164 50896 1176
rect 50948 1164 50954 1216
rect 51092 1204 51120 1244
rect 51350 1232 51356 1284
rect 51408 1272 51414 1284
rect 52549 1275 52607 1281
rect 52549 1272 52561 1275
rect 51408 1244 52561 1272
rect 51408 1232 51414 1244
rect 52549 1241 52561 1244
rect 52595 1241 52607 1275
rect 52549 1235 52607 1241
rect 52638 1232 52644 1284
rect 52696 1272 52702 1284
rect 53469 1275 53527 1281
rect 53469 1272 53481 1275
rect 52696 1244 53481 1272
rect 52696 1232 52702 1244
rect 53469 1241 53481 1244
rect 53515 1241 53527 1275
rect 54297 1275 54355 1281
rect 54297 1272 54309 1275
rect 53469 1235 53527 1241
rect 53576 1244 54309 1272
rect 51445 1207 51503 1213
rect 51445 1204 51457 1207
rect 51092 1176 51457 1204
rect 51445 1173 51457 1176
rect 51491 1173 51503 1207
rect 51718 1204 51724 1216
rect 51679 1176 51724 1204
rect 51445 1167 51503 1173
rect 51718 1164 51724 1176
rect 51776 1164 51782 1216
rect 51810 1164 51816 1216
rect 51868 1204 51874 1216
rect 51997 1207 52055 1213
rect 51997 1204 52009 1207
rect 51868 1176 52009 1204
rect 51868 1164 51874 1176
rect 51997 1173 52009 1176
rect 52043 1173 52055 1207
rect 51997 1167 52055 1173
rect 52362 1164 52368 1216
rect 52420 1204 52426 1216
rect 53193 1207 53251 1213
rect 53193 1204 53205 1207
rect 52420 1176 53205 1204
rect 52420 1164 52426 1176
rect 53193 1173 53205 1176
rect 53239 1173 53251 1207
rect 53193 1167 53251 1173
rect 53282 1164 53288 1216
rect 53340 1204 53346 1216
rect 53576 1204 53604 1244
rect 54297 1241 54309 1244
rect 54343 1241 54355 1275
rect 54849 1275 54907 1281
rect 54849 1272 54861 1275
rect 54297 1235 54355 1241
rect 54404 1244 54861 1272
rect 53742 1204 53748 1216
rect 53340 1176 53604 1204
rect 53703 1176 53748 1204
rect 53340 1164 53346 1176
rect 53742 1164 53748 1176
rect 53800 1164 53806 1216
rect 53834 1164 53840 1216
rect 53892 1204 53898 1216
rect 54404 1204 54432 1244
rect 54849 1241 54861 1244
rect 54895 1241 54907 1275
rect 54849 1235 54907 1241
rect 54938 1232 54944 1284
rect 54996 1272 55002 1284
rect 56045 1275 56103 1281
rect 56045 1272 56057 1275
rect 54996 1244 56057 1272
rect 54996 1232 55002 1244
rect 56045 1241 56057 1244
rect 56091 1241 56103 1275
rect 56045 1235 56103 1241
rect 54570 1204 54576 1216
rect 53892 1176 54432 1204
rect 54531 1176 54576 1204
rect 53892 1164 53898 1176
rect 54570 1164 54576 1176
rect 54628 1164 54634 1216
rect 55122 1204 55128 1216
rect 55083 1176 55128 1204
rect 55122 1164 55128 1176
rect 55180 1164 55186 1216
rect 55490 1204 55496 1216
rect 55451 1176 55496 1204
rect 55490 1164 55496 1176
rect 55548 1164 55554 1216
rect 56318 1204 56324 1216
rect 56279 1176 56324 1204
rect 56318 1164 56324 1176
rect 56376 1164 56382 1216
rect 1288 1114 68816 1136
rect 1288 1062 13262 1114
rect 13314 1062 25262 1114
rect 25314 1062 37262 1114
rect 37314 1062 49262 1114
rect 49314 1062 61262 1114
rect 61314 1062 68816 1114
rect 1288 1040 68816 1062
rect 1854 960 1860 1012
rect 1912 1000 1918 1012
rect 4154 1000 4160 1012
rect 1912 972 4160 1000
rect 1912 960 1918 972
rect 4154 960 4160 972
rect 4212 960 4218 1012
rect 1210 892 1216 944
rect 1268 932 1274 944
rect 5718 932 5724 944
rect 1268 904 5724 932
rect 1268 892 1274 904
rect 5718 892 5724 904
rect 5776 892 5782 944
rect 42242 892 42248 944
rect 42300 932 42306 944
rect 44082 932 44088 944
rect 42300 904 44088 932
rect 42300 892 42306 904
rect 44082 892 44088 904
rect 44140 892 44146 944
rect 53834 892 53840 944
rect 53892 932 53898 944
rect 55122 932 55128 944
rect 53892 904 55128 932
rect 53892 892 53898 904
rect 55122 892 55128 904
rect 55180 892 55186 944
rect 14 824 20 876
rect 72 864 78 876
rect 2774 864 2780 876
rect 72 836 2780 864
rect 72 824 78 836
rect 2774 824 2780 836
rect 2832 824 2838 876
rect 41966 824 41972 876
rect 42024 864 42030 876
rect 43806 864 43812 876
rect 42024 836 43812 864
rect 42024 824 42030 836
rect 43806 824 43812 836
rect 43864 824 43870 876
rect 53282 824 53288 876
rect 53340 864 53346 876
rect 54570 864 54576 876
rect 53340 836 54576 864
rect 53340 824 53346 836
rect 54570 824 54576 836
rect 54628 824 54634 876
rect 290 756 296 808
rect 348 796 354 808
rect 3326 796 3332 808
rect 348 768 3332 796
rect 348 756 354 768
rect 3326 756 3332 768
rect 3384 756 3390 808
rect 29270 756 29276 808
rect 29328 796 29334 808
rect 30834 796 30840 808
rect 29328 768 30840 796
rect 29328 756 29334 768
rect 30834 756 30840 768
rect 30892 756 30898 808
rect 34790 756 34796 808
rect 34848 796 34854 808
rect 35710 796 35716 808
rect 34848 768 35716 796
rect 34848 756 34854 768
rect 35710 756 35716 768
rect 35768 756 35774 808
rect 41138 756 41144 808
rect 41196 796 41202 808
rect 42610 796 42616 808
rect 41196 768 42616 796
rect 41196 756 41202 768
rect 42610 756 42616 768
rect 42668 756 42674 808
rect 44174 756 44180 808
rect 44232 796 44238 808
rect 46106 796 46112 808
rect 44232 768 46112 796
rect 44232 756 44238 768
rect 46106 756 46112 768
rect 46164 756 46170 808
rect 48590 756 48596 808
rect 48648 796 48654 808
rect 49970 796 49976 808
rect 48648 768 49976 796
rect 48648 756 48654 768
rect 49970 756 49976 768
rect 50028 756 50034 808
rect 50522 756 50528 808
rect 50580 796 50586 808
rect 51810 796 51816 808
rect 50580 768 51816 796
rect 50580 756 50586 768
rect 51810 756 51816 768
rect 51868 756 51874 808
rect 54386 756 54392 808
rect 54444 796 54450 808
rect 56318 796 56324 808
rect 54444 768 56324 796
rect 54444 756 54450 768
rect 56318 756 56324 768
rect 56376 756 56382 808
rect 2774 688 2780 740
rect 2832 728 2838 740
rect 5074 728 5080 740
rect 2832 700 5080 728
rect 2832 688 2838 700
rect 5074 688 5080 700
rect 5132 688 5138 740
rect 12434 688 12440 740
rect 12492 728 12498 740
rect 12894 728 12900 740
rect 12492 700 12900 728
rect 12492 688 12498 700
rect 12894 688 12900 700
rect 12952 688 12958 740
rect 15470 688 15476 740
rect 15528 728 15534 740
rect 16022 728 16028 740
rect 15528 700 16028 728
rect 15528 688 15534 700
rect 16022 688 16028 700
rect 16080 688 16086 740
rect 18782 688 18788 740
rect 18840 728 18846 740
rect 20254 728 20260 740
rect 18840 700 20260 728
rect 18840 688 18846 700
rect 20254 688 20260 700
rect 20312 688 20318 740
rect 25406 688 25412 740
rect 25464 728 25470 740
rect 26142 728 26148 740
rect 25464 700 26148 728
rect 25464 688 25470 700
rect 26142 688 26148 700
rect 26200 688 26206 740
rect 27062 688 27068 740
rect 27120 728 27126 740
rect 28626 728 28632 740
rect 27120 700 28632 728
rect 27120 688 27126 700
rect 28626 688 28632 700
rect 28684 688 28690 740
rect 30098 688 30104 740
rect 30156 728 30162 740
rect 31018 728 31024 740
rect 30156 700 31024 728
rect 30156 688 30162 700
rect 31018 688 31024 700
rect 31076 688 31082 740
rect 31478 688 31484 740
rect 31536 728 31542 740
rect 32398 728 32404 740
rect 31536 700 32404 728
rect 31536 688 31542 700
rect 32398 688 32404 700
rect 32456 688 32462 740
rect 35066 688 35072 740
rect 35124 728 35130 740
rect 35802 728 35808 740
rect 35124 700 35808 728
rect 35124 688 35130 700
rect 35802 688 35808 700
rect 35860 688 35866 740
rect 38654 688 38660 740
rect 38712 728 38718 740
rect 39666 728 39672 740
rect 38712 700 39672 728
rect 38712 688 38718 700
rect 39666 688 39672 700
rect 39724 688 39730 740
rect 40034 688 40040 740
rect 40092 728 40098 740
rect 41230 728 41236 740
rect 40092 700 41236 728
rect 40092 688 40098 700
rect 41230 688 41236 700
rect 41288 688 41294 740
rect 41690 688 41696 740
rect 41748 728 41754 740
rect 42794 728 42800 740
rect 41748 700 42800 728
rect 41748 688 41754 700
rect 42794 688 42800 700
rect 42852 688 42858 740
rect 43898 688 43904 740
rect 43956 728 43962 740
rect 45462 728 45468 740
rect 43956 700 45468 728
rect 43956 688 43962 700
rect 45462 688 45468 700
rect 45520 688 45526 740
rect 47762 688 47768 740
rect 47820 728 47826 740
rect 49142 728 49148 740
rect 47820 700 49148 728
rect 47820 688 47826 700
rect 49142 688 49148 700
rect 49200 688 49206 740
rect 50246 688 50252 740
rect 50304 728 50310 740
rect 51718 728 51724 740
rect 50304 700 51724 728
rect 50304 688 50310 700
rect 51718 688 51724 700
rect 51776 688 51782 740
rect 54110 688 54116 740
rect 54168 728 54174 740
rect 55490 728 55496 740
rect 54168 700 55496 728
rect 54168 688 54174 700
rect 55490 688 55496 700
rect 55548 688 55554 740
rect 1762 620 1768 672
rect 1820 660 1826 672
rect 5166 660 5172 672
rect 1820 632 5172 660
rect 1820 620 1826 632
rect 5166 620 5172 632
rect 5224 620 5230 672
rect 42886 620 42892 672
rect 42944 660 42950 672
rect 44634 660 44640 672
rect 42944 632 44640 660
rect 42944 620 42950 632
rect 44634 620 44640 632
rect 44692 620 44698 672
rect 49510 552 49516 604
rect 49568 592 49574 604
rect 50890 592 50896 604
rect 49568 564 50896 592
rect 49568 552 49574 564
rect 50890 552 50896 564
rect 50948 552 50954 604
rect 52546 552 52552 604
rect 52604 592 52610 604
rect 53742 592 53748 604
rect 52604 564 53748 592
rect 52604 552 52610 564
rect 53742 552 53748 564
rect 53800 552 53806 604
<< via1 >>
rect 664 3408 716 3460
rect 6828 3408 6880 3460
rect 1676 3340 1728 3392
rect 5908 3340 5960 3392
rect 24860 3340 24912 3392
rect 25872 3340 25924 3392
rect 13262 3238 13314 3290
rect 25262 3238 25314 3290
rect 37262 3238 37314 3290
rect 49262 3238 49314 3290
rect 61262 3238 61314 3290
rect 1400 3136 1452 3188
rect 3332 3136 3384 3188
rect 3608 3136 3660 3188
rect 4068 3136 4120 3188
rect 4988 3136 5040 3188
rect 5264 3136 5316 3188
rect 5540 3136 5592 3188
rect 5816 3136 5868 3188
rect 6368 3136 6420 3188
rect 6644 3136 6696 3188
rect 6920 3136 6972 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 7472 3136 7524 3188
rect 7748 3136 7800 3188
rect 8024 3136 8076 3188
rect 8300 3136 8352 3188
rect 8576 3136 8628 3188
rect 8852 3136 8904 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 9772 3136 9824 3188
rect 10508 3136 10560 3188
rect 11060 3136 11112 3188
rect 11888 3136 11940 3188
rect 12440 3136 12492 3188
rect 12992 3136 13044 3188
rect 13452 3136 13504 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14096 3136 14148 3188
rect 14648 3136 14700 3188
rect 15292 3136 15344 3188
rect 16028 3136 16080 3188
rect 16948 3136 17000 3188
rect 17776 3136 17828 3188
rect 18604 3136 18656 3188
rect 19524 3136 19576 3188
rect 20444 3136 20496 3188
rect 21548 3136 21600 3188
rect 22652 3136 22704 3188
rect 23756 3136 23808 3188
rect 25136 3136 25188 3188
rect 26332 3136 26384 3188
rect 27620 3136 27672 3188
rect 28724 3136 28776 3188
rect 29828 3136 29880 3188
rect 30932 3136 30984 3188
rect 32036 3136 32088 3188
rect 33140 3136 33192 3188
rect 34060 3136 34112 3188
rect 35348 3136 35400 3188
rect 36728 3136 36780 3188
rect 37832 3136 37884 3188
rect 38936 3136 38988 3188
rect 40132 3136 40184 3188
rect 41236 3136 41288 3188
rect 4160 3068 4212 3120
rect 10232 3068 10284 3120
rect 296 3000 348 3052
rect 9128 3000 9180 3052
rect 16580 3068 16632 3120
rect 17224 3068 17276 3120
rect 18328 3068 18380 3120
rect 19156 3068 19208 3120
rect 20168 3068 20220 3120
rect 21272 3068 21324 3120
rect 22376 3068 22428 3120
rect 23480 3068 23532 3120
rect 24308 3068 24360 3120
rect 25964 3068 26016 3120
rect 27252 3068 27304 3120
rect 29000 3068 29052 3120
rect 30104 3068 30156 3120
rect 31760 3068 31812 3120
rect 32404 3068 32456 3120
rect 33508 3068 33560 3120
rect 34796 3068 34848 3120
rect 36452 3068 36504 3120
rect 37556 3068 37608 3120
rect 38660 3068 38712 3120
rect 39764 3068 39816 3120
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11336 3000 11388 3052
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 12716 3000 12768 3052
rect 14372 3000 14424 3052
rect 15200 3000 15252 3052
rect 15568 3000 15620 3052
rect 16672 3000 16724 3052
rect 17500 3000 17552 3052
rect 18880 3000 18932 3052
rect 19892 3000 19944 3052
rect 20996 3000 21048 3052
rect 22100 3000 22152 3052
rect 22928 3000 22980 3052
rect 24032 3000 24084 3052
rect 25504 3000 25556 3052
rect 26608 3000 26660 3052
rect 27804 3000 27856 3052
rect 29276 3000 29328 3052
rect 30380 3000 30432 3052
rect 31852 3000 31904 3052
rect 32680 3000 32732 3052
rect 33784 3000 33836 3052
rect 35072 3000 35124 3052
rect 20 2932 72 2984
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 572 2864 624 2916
rect 9956 2932 10008 2984
rect 13912 2932 13964 2984
rect 15752 2932 15804 2984
rect 17960 2932 18012 2984
rect 19616 2932 19668 2984
rect 20720 2932 20772 2984
rect 22192 2932 22244 2984
rect 23572 2932 23624 2984
rect 24860 2932 24912 2984
rect 25872 2932 25924 2984
rect 25780 2864 25832 2916
rect 26884 2932 26936 2984
rect 28080 2932 28132 2984
rect 28172 2864 28224 2916
rect 29552 2932 29604 2984
rect 30656 2932 30708 2984
rect 32128 2932 32180 2984
rect 33232 2932 33284 2984
rect 34520 2932 34572 2984
rect 34612 2864 34664 2916
rect 35900 2932 35952 2984
rect 37004 3000 37056 3052
rect 38108 3000 38160 3052
rect 39212 3000 39264 3052
rect 40408 3000 40460 3052
rect 41696 3136 41748 3188
rect 42800 3136 42852 3188
rect 43536 3136 43588 3188
rect 44456 3136 44508 3188
rect 47492 3136 47544 3188
rect 48596 3136 48648 3188
rect 48872 3136 48924 3188
rect 49148 3136 49200 3188
rect 49424 3136 49476 3188
rect 49700 3136 49752 3188
rect 49976 3136 50028 3188
rect 50528 3136 50580 3188
rect 51080 3136 51132 3188
rect 51356 3136 51408 3188
rect 51908 3136 51960 3188
rect 52460 3136 52512 3188
rect 52736 3136 52788 3188
rect 53288 3136 53340 3188
rect 53840 3136 53892 3188
rect 54116 3136 54168 3188
rect 54668 3136 54720 3188
rect 55404 3136 55456 3188
rect 56048 3136 56100 3188
rect 56692 3136 56744 3188
rect 57520 3136 57572 3188
rect 58256 3136 58308 3188
rect 59084 3136 59136 3188
rect 59912 3136 59964 3188
rect 60740 3136 60792 3188
rect 61384 3136 61436 3188
rect 62120 3136 62172 3188
rect 62672 3136 62724 3188
rect 64328 3136 64380 3188
rect 65708 3136 65760 3188
rect 66536 3136 66588 3188
rect 67088 3179 67140 3188
rect 67088 3145 67097 3179
rect 67097 3145 67131 3179
rect 67131 3145 67140 3179
rect 67088 3136 67140 3145
rect 67456 3136 67508 3188
rect 67640 3179 67692 3188
rect 67640 3145 67649 3179
rect 67649 3145 67683 3179
rect 67683 3145 67692 3179
rect 67640 3136 67692 3145
rect 41972 3068 42024 3120
rect 43076 3068 43128 3120
rect 44732 3068 44784 3120
rect 50252 3068 50304 3120
rect 51632 3068 51684 3120
rect 53012 3068 53064 3120
rect 53932 3068 53984 3120
rect 54392 3068 54444 3120
rect 54944 3068 54996 3120
rect 56968 3068 57020 3120
rect 57980 3068 58032 3120
rect 58532 3068 58584 3120
rect 59360 3068 59412 3120
rect 60188 3068 60240 3120
rect 61016 3068 61068 3120
rect 62212 3068 62264 3120
rect 62948 3068 63000 3120
rect 64052 3068 64104 3120
rect 65248 3068 65300 3120
rect 42340 3000 42392 3052
rect 43628 3000 43680 3052
rect 45008 3000 45060 3052
rect 47768 3000 47820 3052
rect 51172 3000 51224 3052
rect 52552 3000 52604 3052
rect 55772 3000 55824 3052
rect 56600 3000 56652 3052
rect 57152 3000 57204 3052
rect 58072 3000 58124 3052
rect 58808 3000 58860 3052
rect 59636 3000 59688 3052
rect 60832 3000 60884 3052
rect 61568 3000 61620 3052
rect 62396 3000 62448 3052
rect 63592 3000 63644 3052
rect 64696 3000 64748 3052
rect 67916 3000 67968 3052
rect 35992 2864 36044 2916
rect 37372 2932 37424 2984
rect 38384 2932 38436 2984
rect 39488 2932 39540 2984
rect 40684 2932 40736 2984
rect 40868 2864 40920 2916
rect 42892 2932 42944 2984
rect 43904 2932 43956 2984
rect 55496 2932 55548 2984
rect 63500 2932 63552 2984
rect 63776 2864 63828 2916
rect 940 2796 992 2848
rect 5632 2796 5684 2848
rect 7262 2694 7314 2746
rect 19262 2694 19314 2746
rect 31262 2694 31314 2746
rect 43262 2694 43314 2746
rect 55262 2694 55314 2746
rect 67262 2694 67314 2746
rect 2964 2524 3016 2576
rect 1952 2456 2004 2508
rect 3884 2456 3936 2508
rect 4436 2456 4488 2508
rect 6092 2456 6144 2508
rect 11612 2456 11664 2508
rect 28448 2456 28500 2508
rect 36176 2456 36228 2508
rect 41420 2456 41472 2508
rect 44180 2456 44232 2508
rect 45284 2499 45336 2508
rect 45284 2465 45293 2499
rect 45293 2465 45327 2499
rect 45327 2465 45336 2499
rect 45284 2456 45336 2465
rect 45560 2499 45612 2508
rect 45560 2465 45569 2499
rect 45569 2465 45603 2499
rect 45603 2465 45612 2499
rect 45836 2499 45888 2508
rect 45560 2456 45612 2465
rect 45836 2465 45845 2499
rect 45845 2465 45879 2499
rect 45879 2465 45888 2499
rect 45836 2456 45888 2465
rect 46112 2499 46164 2508
rect 46112 2465 46121 2499
rect 46121 2465 46155 2499
rect 46155 2465 46164 2499
rect 46112 2456 46164 2465
rect 46388 2499 46440 2508
rect 46388 2465 46397 2499
rect 46397 2465 46431 2499
rect 46431 2465 46440 2499
rect 46388 2456 46440 2465
rect 46664 2499 46716 2508
rect 46664 2465 46673 2499
rect 46673 2465 46707 2499
rect 46707 2465 46716 2499
rect 46664 2456 46716 2465
rect 46940 2499 46992 2508
rect 46940 2465 46949 2499
rect 46949 2465 46983 2499
rect 46983 2465 46992 2499
rect 46940 2456 46992 2465
rect 47216 2499 47268 2508
rect 47216 2465 47225 2499
rect 47225 2465 47259 2499
rect 47259 2465 47268 2499
rect 47216 2456 47268 2465
rect 48044 2499 48096 2508
rect 48044 2465 48053 2499
rect 48053 2465 48087 2499
rect 48087 2465 48096 2499
rect 48044 2456 48096 2465
rect 48320 2499 48372 2508
rect 48320 2465 48329 2499
rect 48329 2465 48363 2499
rect 48363 2465 48372 2499
rect 48320 2456 48372 2465
rect 64880 2456 64932 2508
rect 65432 2499 65484 2508
rect 65432 2465 65441 2499
rect 65441 2465 65475 2499
rect 65475 2465 65484 2499
rect 65432 2456 65484 2465
rect 65984 2499 66036 2508
rect 65984 2465 65993 2499
rect 65993 2465 66027 2499
rect 66027 2465 66036 2499
rect 65984 2456 66036 2465
rect 66260 2499 66312 2508
rect 66260 2465 66269 2499
rect 66269 2465 66303 2499
rect 66303 2465 66312 2499
rect 66260 2456 66312 2465
rect 66812 2456 66864 2508
rect 2504 2388 2556 2440
rect 3792 2388 3844 2440
rect 2228 2320 2280 2372
rect 3332 2320 3384 2372
rect 3700 2320 3752 2372
rect 848 2252 900 2304
rect 2780 2252 2832 2304
rect 3516 2252 3568 2304
rect 3608 2295 3660 2304
rect 3608 2261 3617 2295
rect 3617 2261 3651 2295
rect 3651 2261 3660 2295
rect 3976 2320 4028 2372
rect 4712 2388 4764 2440
rect 5816 2388 5868 2440
rect 3608 2252 3660 2261
rect 5724 2252 5776 2304
rect 13262 2150 13314 2202
rect 25262 2150 25314 2202
rect 37262 2150 37314 2202
rect 49262 2150 49314 2202
rect 61262 2150 61314 2202
rect 2964 2048 3016 2100
rect 3056 2048 3108 2100
rect 4252 2048 4304 2100
rect 4712 2048 4764 2100
rect 6828 2091 6880 2100
rect 6828 2057 6837 2091
rect 6837 2057 6871 2091
rect 6871 2057 6880 2091
rect 6828 2048 6880 2057
rect 2780 1980 2832 2032
rect 5540 1980 5592 2032
rect 1124 1912 1176 1964
rect 1400 1776 1452 1828
rect 2872 1912 2924 1964
rect 5356 1912 5408 1964
rect 45008 1912 45060 1964
rect 3056 1887 3108 1896
rect 3056 1853 3065 1887
rect 3065 1853 3099 1887
rect 3099 1853 3108 1887
rect 3056 1844 3108 1853
rect 3332 1887 3384 1896
rect 3332 1853 3341 1887
rect 3341 1853 3375 1887
rect 3375 1853 3384 1887
rect 3332 1844 3384 1853
rect 3516 1844 3568 1896
rect 2964 1776 3016 1828
rect 5172 1844 5224 1896
rect 5908 1844 5960 1896
rect 6920 1844 6972 1896
rect 9404 1844 9456 1896
rect 11612 1844 11664 1896
rect 13544 1844 13596 1896
rect 16120 1844 16172 1896
rect 19616 1844 19668 1896
rect 21548 1844 21600 1896
rect 24308 1844 24360 1896
rect 28448 1844 28500 1896
rect 30656 1844 30708 1896
rect 31760 1844 31812 1896
rect 43444 1844 43496 1896
rect 44456 1844 44508 1896
rect 51080 1844 51132 1896
rect 3884 1708 3936 1760
rect 7262 1606 7314 1658
rect 19262 1606 19314 1658
rect 31262 1606 31314 1658
rect 43262 1606 43314 1658
rect 55262 1606 55314 1658
rect 67262 1606 67314 1658
rect 2228 1368 2280 1420
rect 2412 1300 2464 1352
rect 3148 1368 3200 1420
rect 3608 1368 3660 1420
rect 26516 1368 26568 1420
rect 27896 1368 27948 1420
rect 3792 1300 3844 1352
rect 4988 1300 5040 1352
rect 5632 1300 5684 1352
rect 6644 1300 6696 1352
rect 7472 1300 7524 1352
rect 9680 1300 9732 1352
rect 11336 1300 11388 1352
rect 12992 1300 13044 1352
rect 13820 1300 13872 1352
rect 15752 1300 15804 1352
rect 16856 1300 16908 1352
rect 17684 1300 17736 1352
rect 19432 1300 19484 1352
rect 20168 1300 20220 1352
rect 20996 1300 21048 1352
rect 22376 1300 22428 1352
rect 23480 1300 23532 1352
rect 24860 1300 24912 1352
rect 25964 1300 26016 1352
rect 27344 1300 27396 1352
rect 38936 1368 38988 1420
rect 41420 1368 41472 1420
rect 29552 1300 29604 1352
rect 30932 1300 30984 1352
rect 32312 1300 32364 1352
rect 33232 1300 33284 1352
rect 34060 1300 34112 1352
rect 1952 1232 2004 1284
rect 1860 1207 1912 1216
rect 1860 1173 1869 1207
rect 1869 1173 1903 1207
rect 1903 1173 1912 1207
rect 1860 1164 1912 1173
rect 3240 1232 3292 1284
rect 3516 1232 3568 1284
rect 4528 1232 4580 1284
rect 6184 1232 6236 1284
rect 7748 1232 7800 1284
rect 8300 1232 8352 1284
rect 8852 1232 8904 1284
rect 10232 1232 10284 1284
rect 10784 1232 10836 1284
rect 11888 1232 11940 1284
rect 12808 1232 12860 1284
rect 14096 1232 14148 1284
rect 14740 1232 14792 1284
rect 15292 1232 15344 1284
rect 2780 1207 2832 1216
rect 2780 1173 2789 1207
rect 2789 1173 2823 1207
rect 2823 1173 2832 1207
rect 3332 1207 3384 1216
rect 2780 1164 2832 1173
rect 3332 1173 3341 1207
rect 3341 1173 3375 1207
rect 3375 1173 3384 1207
rect 3332 1164 3384 1173
rect 3424 1164 3476 1216
rect 3700 1164 3752 1216
rect 4252 1164 4304 1216
rect 5080 1164 5132 1216
rect 6368 1164 6420 1216
rect 7380 1164 7432 1216
rect 8024 1164 8076 1216
rect 8576 1164 8628 1216
rect 9220 1164 9272 1216
rect 9956 1164 10008 1216
rect 10508 1164 10560 1216
rect 11060 1164 11112 1216
rect 12164 1164 12216 1216
rect 12900 1164 12952 1216
rect 13452 1164 13504 1216
rect 14372 1164 14424 1216
rect 15016 1164 15068 1216
rect 16580 1232 16632 1284
rect 17408 1232 17460 1284
rect 16028 1207 16080 1216
rect 16028 1173 16037 1207
rect 16037 1173 16071 1207
rect 16071 1173 16080 1207
rect 16028 1164 16080 1173
rect 16396 1164 16448 1216
rect 17132 1164 17184 1216
rect 17960 1232 18012 1284
rect 19064 1232 19116 1284
rect 19892 1232 19944 1284
rect 20720 1232 20772 1284
rect 21824 1232 21876 1284
rect 22652 1232 22704 1284
rect 18236 1164 18288 1216
rect 18972 1164 19024 1216
rect 20260 1207 20312 1216
rect 20260 1173 20269 1207
rect 20269 1173 20303 1207
rect 20303 1173 20312 1207
rect 20260 1164 20312 1173
rect 20628 1164 20680 1216
rect 21272 1164 21324 1216
rect 22100 1164 22152 1216
rect 22928 1232 22980 1284
rect 23756 1232 23808 1284
rect 24676 1232 24728 1284
rect 25688 1232 25740 1284
rect 26792 1232 26844 1284
rect 27620 1232 27672 1284
rect 23388 1164 23440 1216
rect 24032 1164 24084 1216
rect 25136 1164 25188 1216
rect 26148 1207 26200 1216
rect 26148 1173 26157 1207
rect 26157 1173 26191 1207
rect 26191 1173 26200 1207
rect 26148 1164 26200 1173
rect 26240 1164 26292 1216
rect 28172 1232 28224 1284
rect 29000 1232 29052 1284
rect 29920 1232 29972 1284
rect 28632 1207 28684 1216
rect 28632 1173 28641 1207
rect 28641 1173 28675 1207
rect 28675 1173 28684 1207
rect 28632 1164 28684 1173
rect 28724 1164 28776 1216
rect 30380 1164 30432 1216
rect 32036 1232 32088 1284
rect 32956 1232 33008 1284
rect 33784 1232 33836 1284
rect 34612 1232 34664 1284
rect 35624 1300 35676 1352
rect 36636 1300 36688 1352
rect 37556 1300 37608 1352
rect 38384 1300 38436 1352
rect 39488 1300 39540 1352
rect 40776 1300 40828 1352
rect 45836 1368 45888 1420
rect 47400 1368 47452 1420
rect 43076 1300 43128 1352
rect 35348 1232 35400 1284
rect 36360 1232 36412 1284
rect 37372 1232 37424 1284
rect 38108 1232 38160 1284
rect 39212 1232 39264 1284
rect 30840 1164 30892 1216
rect 31024 1164 31076 1216
rect 31576 1164 31628 1216
rect 32404 1164 32456 1216
rect 32680 1164 32732 1216
rect 33508 1164 33560 1216
rect 34336 1164 34388 1216
rect 35716 1207 35768 1216
rect 35716 1173 35725 1207
rect 35725 1173 35759 1207
rect 35759 1173 35768 1207
rect 35716 1164 35768 1173
rect 35808 1164 35860 1216
rect 36084 1164 36136 1216
rect 36912 1164 36964 1216
rect 37832 1164 37884 1216
rect 38660 1164 38712 1216
rect 39672 1207 39724 1216
rect 39672 1173 39681 1207
rect 39681 1173 39715 1207
rect 39715 1173 39724 1207
rect 39672 1164 39724 1173
rect 39764 1164 39816 1216
rect 40500 1164 40552 1216
rect 42524 1232 42576 1284
rect 43628 1232 43680 1284
rect 45284 1300 45336 1352
rect 46480 1300 46532 1352
rect 48872 1368 48924 1420
rect 48688 1300 48740 1352
rect 49884 1368 49936 1420
rect 50804 1368 50856 1420
rect 51632 1300 51684 1352
rect 53012 1300 53064 1352
rect 54668 1300 54720 1352
rect 44732 1232 44784 1284
rect 41236 1207 41288 1216
rect 41236 1173 41245 1207
rect 41245 1173 41279 1207
rect 41279 1173 41288 1207
rect 41236 1164 41288 1173
rect 41328 1164 41380 1216
rect 42616 1207 42668 1216
rect 42616 1173 42625 1207
rect 42625 1173 42659 1207
rect 42659 1173 42668 1207
rect 42616 1164 42668 1173
rect 42800 1164 42852 1216
rect 43812 1207 43864 1216
rect 43812 1173 43821 1207
rect 43821 1173 43855 1207
rect 43855 1173 43864 1207
rect 43812 1164 43864 1173
rect 44088 1207 44140 1216
rect 44088 1173 44097 1207
rect 44097 1173 44131 1207
rect 44131 1173 44140 1207
rect 44088 1164 44140 1173
rect 44640 1207 44692 1216
rect 44640 1173 44649 1207
rect 44649 1173 44683 1207
rect 44683 1173 44692 1207
rect 44640 1164 44692 1173
rect 45468 1207 45520 1216
rect 45468 1173 45477 1207
rect 45477 1173 45511 1207
rect 45511 1173 45520 1207
rect 45468 1164 45520 1173
rect 45560 1164 45612 1216
rect 46112 1207 46164 1216
rect 46112 1173 46121 1207
rect 46121 1173 46155 1207
rect 46155 1173 46164 1207
rect 46112 1164 46164 1173
rect 46204 1164 46256 1216
rect 47308 1232 47360 1284
rect 48412 1232 48464 1284
rect 49516 1232 49568 1284
rect 46940 1164 46992 1216
rect 48136 1164 48188 1216
rect 49148 1207 49200 1216
rect 49148 1173 49157 1207
rect 49157 1173 49191 1207
rect 49191 1173 49200 1207
rect 49148 1164 49200 1173
rect 49976 1207 50028 1216
rect 49976 1173 49985 1207
rect 49985 1173 50019 1207
rect 50019 1173 50028 1207
rect 49976 1164 50028 1173
rect 50068 1164 50120 1216
rect 50896 1207 50948 1216
rect 50896 1173 50905 1207
rect 50905 1173 50939 1207
rect 50939 1173 50948 1207
rect 50896 1164 50948 1173
rect 51356 1232 51408 1284
rect 52644 1232 52696 1284
rect 51724 1207 51776 1216
rect 51724 1173 51733 1207
rect 51733 1173 51767 1207
rect 51767 1173 51776 1207
rect 51724 1164 51776 1173
rect 51816 1164 51868 1216
rect 52368 1164 52420 1216
rect 53288 1164 53340 1216
rect 53748 1207 53800 1216
rect 53748 1173 53757 1207
rect 53757 1173 53791 1207
rect 53791 1173 53800 1207
rect 53748 1164 53800 1173
rect 53840 1164 53892 1216
rect 54944 1232 54996 1284
rect 54576 1207 54628 1216
rect 54576 1173 54585 1207
rect 54585 1173 54619 1207
rect 54619 1173 54628 1207
rect 54576 1164 54628 1173
rect 55128 1207 55180 1216
rect 55128 1173 55137 1207
rect 55137 1173 55171 1207
rect 55171 1173 55180 1207
rect 55128 1164 55180 1173
rect 55496 1207 55548 1216
rect 55496 1173 55505 1207
rect 55505 1173 55539 1207
rect 55539 1173 55548 1207
rect 55496 1164 55548 1173
rect 56324 1207 56376 1216
rect 56324 1173 56333 1207
rect 56333 1173 56367 1207
rect 56367 1173 56376 1207
rect 56324 1164 56376 1173
rect 13262 1062 13314 1114
rect 25262 1062 25314 1114
rect 37262 1062 37314 1114
rect 49262 1062 49314 1114
rect 61262 1062 61314 1114
rect 1860 960 1912 1012
rect 4160 960 4212 1012
rect 1216 892 1268 944
rect 5724 892 5776 944
rect 42248 892 42300 944
rect 44088 892 44140 944
rect 53840 892 53892 944
rect 55128 892 55180 944
rect 20 824 72 876
rect 2780 824 2832 876
rect 41972 824 42024 876
rect 43812 824 43864 876
rect 53288 824 53340 876
rect 54576 824 54628 876
rect 296 756 348 808
rect 3332 756 3384 808
rect 29276 756 29328 808
rect 30840 756 30892 808
rect 34796 756 34848 808
rect 35716 756 35768 808
rect 41144 756 41196 808
rect 42616 756 42668 808
rect 44180 756 44232 808
rect 46112 756 46164 808
rect 48596 756 48648 808
rect 49976 756 50028 808
rect 50528 756 50580 808
rect 51816 756 51868 808
rect 54392 756 54444 808
rect 56324 756 56376 808
rect 2780 688 2832 740
rect 5080 688 5132 740
rect 12440 688 12492 740
rect 12900 688 12952 740
rect 15476 688 15528 740
rect 16028 688 16080 740
rect 18788 688 18840 740
rect 20260 688 20312 740
rect 25412 688 25464 740
rect 26148 688 26200 740
rect 27068 688 27120 740
rect 28632 688 28684 740
rect 30104 688 30156 740
rect 31024 688 31076 740
rect 31484 688 31536 740
rect 32404 688 32456 740
rect 35072 688 35124 740
rect 35808 688 35860 740
rect 38660 688 38712 740
rect 39672 688 39724 740
rect 40040 688 40092 740
rect 41236 688 41288 740
rect 41696 688 41748 740
rect 42800 688 42852 740
rect 43904 688 43956 740
rect 45468 688 45520 740
rect 47768 688 47820 740
rect 49148 688 49200 740
rect 50252 688 50304 740
rect 51724 688 51776 740
rect 54116 688 54168 740
rect 55496 688 55548 740
rect 1768 620 1820 672
rect 5172 620 5224 672
rect 42892 620 42944 672
rect 44640 620 44692 672
rect 49516 552 49568 604
rect 50896 552 50948 604
rect 52552 552 52604 604
rect 53748 552 53800 604
<< metal2 >>
rect 18 3800 74 4400
rect 294 3800 350 4400
rect 570 3800 626 4400
rect 846 3800 902 4400
rect 1122 3800 1178 4400
rect 1398 3800 1454 4400
rect 1674 3800 1730 4400
rect 1950 3800 2006 4400
rect 2226 3800 2282 4400
rect 2502 3800 2558 4400
rect 2778 3800 2834 4400
rect 3054 3800 3110 4400
rect 3330 3800 3386 4400
rect 3606 3800 3662 4400
rect 3882 3800 3938 4400
rect 4158 3800 4214 4400
rect 4434 3800 4490 4400
rect 4710 3800 4766 4400
rect 4986 3800 5042 4400
rect 5262 3800 5318 4400
rect 5538 3800 5594 4400
rect 5814 3800 5870 4400
rect 6090 3800 6146 4400
rect 6366 3800 6422 4400
rect 6642 3800 6698 4400
rect 6918 3800 6974 4400
rect 7194 3800 7250 4400
rect 7470 3800 7526 4400
rect 7746 3800 7802 4400
rect 8022 3800 8078 4400
rect 8298 3800 8354 4400
rect 8574 3800 8630 4400
rect 8850 3800 8906 4400
rect 9126 3800 9182 4400
rect 9402 3800 9458 4400
rect 9678 3800 9734 4400
rect 9954 3800 10010 4400
rect 10230 3800 10286 4400
rect 10506 3800 10562 4400
rect 10782 3800 10838 4400
rect 11058 3800 11114 4400
rect 11334 3800 11390 4400
rect 11610 3800 11666 4400
rect 11886 3800 11942 4400
rect 12162 3800 12218 4400
rect 12438 3800 12494 4400
rect 12714 3800 12770 4400
rect 12990 3800 13046 4400
rect 13266 3800 13322 4400
rect 13542 3800 13598 4400
rect 13818 3800 13874 4400
rect 14094 3800 14150 4400
rect 14370 3800 14426 4400
rect 14646 3800 14702 4400
rect 14922 3800 14978 4400
rect 15198 3800 15254 4400
rect 15474 3800 15530 4400
rect 15750 3800 15806 4400
rect 16026 3800 16082 4400
rect 16302 3800 16358 4400
rect 16578 3800 16634 4400
rect 16854 3800 16910 4400
rect 17130 3800 17186 4400
rect 17406 3800 17462 4400
rect 17682 3800 17738 4400
rect 17958 3800 18014 4400
rect 18234 3800 18290 4400
rect 18510 3800 18566 4400
rect 18786 3800 18842 4400
rect 19062 3800 19118 4400
rect 19338 3800 19394 4400
rect 19614 3800 19670 4400
rect 19890 3800 19946 4400
rect 20166 3800 20222 4400
rect 20442 3800 20498 4400
rect 20718 3800 20774 4400
rect 20994 3800 21050 4400
rect 21270 3800 21326 4400
rect 21546 3800 21602 4400
rect 21822 3800 21878 4400
rect 22098 3800 22154 4400
rect 22374 3800 22430 4400
rect 22650 3800 22706 4400
rect 22926 3800 22982 4400
rect 23202 3800 23258 4400
rect 23478 3800 23534 4400
rect 23754 3800 23810 4400
rect 24030 3800 24086 4400
rect 24306 3800 24362 4400
rect 24582 3800 24638 4400
rect 24858 3800 24914 4400
rect 25134 3800 25190 4400
rect 25410 3800 25466 4400
rect 25686 3800 25742 4400
rect 25962 3800 26018 4400
rect 26238 3800 26294 4400
rect 26514 3800 26570 4400
rect 26790 3800 26846 4400
rect 27066 3800 27122 4400
rect 27342 3800 27398 4400
rect 27618 3800 27674 4400
rect 27894 3800 27950 4400
rect 28170 3800 28226 4400
rect 28446 3800 28502 4400
rect 28722 3800 28778 4400
rect 28998 3800 29054 4400
rect 29274 3800 29330 4400
rect 29550 3800 29606 4400
rect 29826 3800 29882 4400
rect 30102 3800 30158 4400
rect 30378 3800 30434 4400
rect 30654 3800 30710 4400
rect 30930 3800 30986 4400
rect 31206 3800 31262 4400
rect 31482 3800 31538 4400
rect 31758 3800 31814 4400
rect 32034 3800 32090 4400
rect 32310 3800 32366 4400
rect 32586 3800 32642 4400
rect 32862 3800 32918 4400
rect 33138 3800 33194 4400
rect 33414 3800 33470 4400
rect 33690 3800 33746 4400
rect 33966 3800 34022 4400
rect 34242 3800 34298 4400
rect 34518 3800 34574 4400
rect 34794 3800 34850 4400
rect 35070 3800 35126 4400
rect 35346 3800 35402 4400
rect 35622 3800 35678 4400
rect 35898 3800 35954 4400
rect 36174 3800 36230 4400
rect 36450 3800 36506 4400
rect 36726 3800 36782 4400
rect 37002 3800 37058 4400
rect 37278 3800 37334 4400
rect 37554 3800 37610 4400
rect 37830 3800 37886 4400
rect 38106 3800 38162 4400
rect 38382 3800 38438 4400
rect 38658 3800 38714 4400
rect 38934 3800 38990 4400
rect 39210 3800 39266 4400
rect 39486 3800 39542 4400
rect 39762 3800 39818 4400
rect 40038 3800 40094 4400
rect 40314 3800 40370 4400
rect 40590 3800 40646 4400
rect 40866 3800 40922 4400
rect 41142 3800 41198 4400
rect 41418 3800 41474 4400
rect 41694 3800 41750 4400
rect 41970 3800 42026 4400
rect 42246 3800 42302 4400
rect 42522 3800 42578 4400
rect 42798 3800 42854 4400
rect 43074 3800 43130 4400
rect 43350 3800 43406 4400
rect 43626 3800 43682 4400
rect 43902 3800 43958 4400
rect 44178 3800 44234 4400
rect 44454 3800 44510 4400
rect 44730 3800 44786 4400
rect 45006 3800 45062 4400
rect 45282 3800 45338 4400
rect 45558 3800 45614 4400
rect 45834 3800 45890 4400
rect 46110 3800 46166 4400
rect 46386 3800 46442 4400
rect 46662 3800 46718 4400
rect 46938 3800 46994 4400
rect 47214 3800 47270 4400
rect 47490 3800 47546 4400
rect 47766 3800 47822 4400
rect 48042 3800 48098 4400
rect 48318 3800 48374 4400
rect 48594 3800 48650 4400
rect 48870 3800 48926 4400
rect 49146 3800 49202 4400
rect 49422 3800 49478 4400
rect 49698 3800 49754 4400
rect 49974 3800 50030 4400
rect 50250 3800 50306 4400
rect 50526 3800 50582 4400
rect 50802 3800 50858 4400
rect 51078 3800 51134 4400
rect 51354 3800 51410 4400
rect 51630 3800 51686 4400
rect 51906 3800 51962 4400
rect 52182 3800 52238 4400
rect 52458 3800 52514 4400
rect 52734 3800 52790 4400
rect 53010 3800 53066 4400
rect 53286 3800 53342 4400
rect 53562 3800 53618 4400
rect 53838 3800 53894 4400
rect 54114 3800 54170 4400
rect 54390 3800 54446 4400
rect 54666 3800 54722 4400
rect 54942 3800 54998 4400
rect 55218 3800 55274 4400
rect 55494 3800 55550 4400
rect 55770 3800 55826 4400
rect 56046 3800 56102 4400
rect 56322 3800 56378 4400
rect 56598 3800 56654 4400
rect 56874 3800 56930 4400
rect 57150 3800 57206 4400
rect 57426 3800 57482 4400
rect 57702 3800 57758 4400
rect 57978 3800 58034 4400
rect 58254 3800 58310 4400
rect 58530 3800 58586 4400
rect 58806 3800 58862 4400
rect 59082 3800 59138 4400
rect 59358 3800 59414 4400
rect 59634 3800 59690 4400
rect 59910 3800 59966 4400
rect 60186 3800 60242 4400
rect 60462 3800 60518 4400
rect 60738 3800 60794 4400
rect 61014 3800 61070 4400
rect 61290 3800 61346 4400
rect 61566 3800 61622 4400
rect 61842 3800 61898 4400
rect 62118 3800 62174 4400
rect 62394 3800 62450 4400
rect 62670 3800 62726 4400
rect 62946 3800 63002 4400
rect 63222 3800 63278 4400
rect 63498 3800 63554 4400
rect 63774 3800 63830 4400
rect 64050 3800 64106 4400
rect 64326 3800 64382 4400
rect 64602 3800 64658 4400
rect 64878 3800 64934 4400
rect 65154 3800 65210 4400
rect 65430 3800 65486 4400
rect 65706 3800 65762 4400
rect 65982 3800 66038 4400
rect 66258 3800 66314 4400
rect 66534 3800 66590 4400
rect 66810 3800 66866 4400
rect 67086 3800 67142 4400
rect 67362 3800 67418 4400
rect 67638 3800 67694 4400
rect 67914 3800 67970 4400
rect 32 2990 60 3800
rect 308 3058 336 3800
rect 296 3052 348 3058
rect 296 2994 348 3000
rect 20 2984 72 2990
rect 20 2926 72 2932
rect 584 2922 612 3800
rect 664 3460 716 3466
rect 664 3402 716 3408
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 676 1034 704 3402
rect 860 2310 888 3800
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 584 1006 704 1034
rect 20 876 72 882
rect 20 818 72 824
rect 32 600 60 818
rect 296 808 348 814
rect 296 750 348 756
rect 308 600 336 750
rect 584 600 612 1006
rect 952 626 980 2790
rect 1136 2122 1164 3800
rect 1412 3194 1440 3800
rect 1688 3482 1716 3800
rect 1688 3454 1808 3482
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1136 2094 1256 2122
rect 1124 1964 1176 1970
rect 1124 1906 1176 1912
rect 860 600 980 626
rect 1136 600 1164 1906
rect 1228 950 1256 2094
rect 1400 1828 1452 1834
rect 1400 1770 1452 1776
rect 1216 944 1268 950
rect 1216 886 1268 892
rect 1412 600 1440 1770
rect 1688 600 1716 3334
rect 1780 678 1808 3454
rect 1964 2514 1992 3800
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2240 2378 2268 3800
rect 2516 2446 2544 3800
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 2792 2310 2820 3800
rect 2962 3768 3018 3777
rect 2962 3703 3018 3712
rect 2976 2582 3004 3703
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 3068 2106 3096 3800
rect 3344 3194 3372 3800
rect 3620 3194 3648 3800
rect 3698 3360 3754 3369
rect 3698 3295 3754 3304
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3712 2378 3740 3295
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3804 2446 3832 3023
rect 3896 2514 3924 3800
rect 4066 3768 4122 3777
rect 4066 3703 4122 3712
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3988 2378 4016 3567
rect 4080 3194 4108 3703
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4172 3126 4200 3800
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4066 2544 4122 2553
rect 4172 2530 4200 2926
rect 4250 2816 4306 2825
rect 4250 2751 4306 2760
rect 4122 2502 4200 2530
rect 4066 2479 4122 2488
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 3056 2100 3108 2106
rect 3056 2042 3108 2048
rect 2780 2032 2832 2038
rect 2778 2000 2780 2009
rect 2832 2000 2834 2009
rect 2976 1986 3004 2042
rect 2778 1935 2834 1944
rect 2872 1964 2924 1970
rect 2976 1958 3188 1986
rect 2872 1906 2924 1912
rect 2884 1737 2912 1906
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 2964 1828 3016 1834
rect 2964 1770 3016 1776
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 2976 1465 3004 1770
rect 2962 1456 3018 1465
rect 2228 1420 2280 1426
rect 2962 1391 3018 1400
rect 2228 1362 2280 1368
rect 1952 1284 2004 1290
rect 1952 1226 2004 1232
rect 1860 1216 1912 1222
rect 1860 1158 1912 1164
rect 1872 1018 1900 1158
rect 1860 1012 1912 1018
rect 1860 954 1912 960
rect 1768 672 1820 678
rect 1768 614 1820 620
rect 1964 600 1992 1226
rect 2240 600 2268 1362
rect 2412 1352 2464 1358
rect 2412 1294 2464 1300
rect 2424 626 2452 1294
rect 2780 1216 2832 1222
rect 2780 1158 2832 1164
rect 2792 882 2820 1158
rect 2780 876 2832 882
rect 2780 818 2832 824
rect 2780 740 2832 746
rect 2780 682 2832 688
rect 2424 600 2544 626
rect 2792 600 2820 682
rect 3068 600 3096 1838
rect 3160 1426 3188 1958
rect 3344 1902 3372 2314
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3528 1902 3556 2246
rect 3620 2145 3648 2246
rect 3606 2136 3662 2145
rect 4264 2106 4292 2751
rect 4448 2514 4476 3800
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4724 2446 4752 3800
rect 5000 3194 5028 3800
rect 5276 3194 5304 3800
rect 5552 3194 5580 3800
rect 5828 3194 5856 3800
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 3606 2071 3662 2080
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3884 1760 3936 1766
rect 3884 1702 3936 1708
rect 3148 1420 3200 1426
rect 3148 1362 3200 1368
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 3516 1284 3568 1290
rect 3516 1226 3568 1232
rect 3252 626 3280 1226
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3424 1216 3476 1222
rect 3424 1158 3476 1164
rect 3344 814 3372 1158
rect 3332 808 3384 814
rect 3332 750 3384 756
rect 3436 649 3464 1158
rect 3528 921 3556 1226
rect 3514 912 3570 921
rect 3514 847 3570 856
rect 3422 640 3478 649
rect 3252 600 3372 626
rect 18 0 74 600
rect 294 0 350 600
rect 570 0 626 600
rect 846 598 980 600
rect 846 0 902 598
rect 1122 0 1178 600
rect 1398 0 1454 600
rect 1674 0 1730 600
rect 1950 0 2006 600
rect 2226 0 2282 600
rect 2424 598 2558 600
rect 2502 0 2558 598
rect 2778 0 2834 600
rect 3054 0 3110 600
rect 3252 598 3386 600
rect 3330 0 3386 598
rect 3620 600 3648 1362
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3700 1216 3752 1222
rect 3700 1158 3752 1164
rect 3712 1057 3740 1158
rect 3698 1048 3754 1057
rect 3698 983 3754 992
rect 3804 649 3832 1294
rect 3790 640 3846 649
rect 3422 575 3478 584
rect 3606 0 3662 600
rect 3896 600 3924 1702
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 4252 1216 4304 1222
rect 4080 1164 4252 1170
rect 4080 1158 4304 1164
rect 4080 1142 4292 1158
rect 4080 649 4108 1142
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 4066 640 4122 649
rect 3790 575 3846 584
rect 3882 0 3938 600
rect 4172 600 4200 954
rect 4540 626 4568 1226
rect 4448 600 4568 626
rect 4724 600 4752 2042
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5000 600 5028 1294
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5092 746 5120 1158
rect 5080 740 5132 746
rect 5080 682 5132 688
rect 5184 678 5212 1838
rect 5368 1034 5396 1906
rect 5276 1006 5396 1034
rect 5172 672 5224 678
rect 5172 614 5224 620
rect 5276 600 5304 1006
rect 5552 600 5580 1974
rect 5644 1358 5672 2790
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 5736 950 5764 2246
rect 5724 944 5776 950
rect 5724 886 5776 892
rect 5828 600 5856 2382
rect 5920 1902 5948 3334
rect 6104 2514 6132 3800
rect 6380 3194 6408 3800
rect 6656 3194 6684 3800
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6840 2106 6868 3402
rect 6932 3194 6960 3800
rect 7208 3448 7236 3800
rect 7208 3420 7420 3448
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7238 2746 7338 3312
rect 7392 3194 7420 3420
rect 7484 3194 7512 3800
rect 7760 3194 7788 3800
rect 8036 3194 8064 3800
rect 8312 3194 8340 3800
rect 8588 3194 8616 3800
rect 8864 3194 8892 3800
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9140 3058 9168 3800
rect 9416 3176 9444 3800
rect 9692 3346 9720 3800
rect 9692 3318 9812 3346
rect 9784 3194 9812 3318
rect 9680 3188 9732 3194
rect 9416 3148 9680 3176
rect 9680 3130 9732 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9968 2990 9996 3800
rect 10244 3126 10272 3800
rect 10520 3194 10548 3800
rect 10508 3188 10560 3194
rect 10796 3176 10824 3800
rect 11072 3194 11100 3800
rect 11060 3188 11112 3194
rect 10796 3148 11008 3176
rect 10508 3130 10560 3136
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10980 3040 11008 3148
rect 11060 3130 11112 3136
rect 11348 3058 11376 3800
rect 11060 3052 11112 3058
rect 10980 3012 11060 3040
rect 11060 2994 11112 3000
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 7238 2694 7262 2746
rect 7314 2694 7338 2746
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6920 1896 6972 1902
rect 6920 1838 6972 1844
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6184 1284 6236 1290
rect 6184 1226 6236 1232
rect 6196 626 6224 1226
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6104 600 6224 626
rect 6380 600 6408 1158
rect 6656 600 6684 1294
rect 6932 600 6960 1838
rect 7238 1658 7338 2694
rect 11624 2514 11652 3800
rect 11900 3194 11928 3800
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12176 3040 12204 3800
rect 12452 3194 12480 3800
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12728 3058 12756 3800
rect 13004 3194 13032 3800
rect 13280 3448 13308 3800
rect 13280 3420 13492 3448
rect 13238 3290 13338 3312
rect 13238 3238 13262 3290
rect 13314 3238 13338 3290
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 12440 3052 12492 3058
rect 12176 3012 12440 3040
rect 12440 2994 12492 3000
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 13238 2348 13338 3238
rect 13464 3194 13492 3420
rect 13452 3188 13504 3194
rect 13556 3176 13584 3800
rect 13832 3346 13860 3800
rect 13832 3318 13952 3346
rect 13820 3188 13872 3194
rect 13556 3148 13820 3176
rect 13452 3130 13504 3136
rect 13820 3130 13872 3136
rect 13924 2990 13952 3318
rect 14108 3194 14136 3800
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14384 3058 14412 3800
rect 14660 3194 14688 3800
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14936 3074 14964 3800
rect 15212 3176 15240 3800
rect 15292 3188 15344 3194
rect 15212 3148 15292 3176
rect 15292 3130 15344 3136
rect 14936 3058 15240 3074
rect 14372 3052 14424 3058
rect 14936 3052 15252 3058
rect 14936 3046 15200 3052
rect 14372 2994 14424 3000
rect 15488 3040 15516 3800
rect 15568 3052 15620 3058
rect 15488 3012 15568 3040
rect 15200 2994 15252 3000
rect 15568 2994 15620 3000
rect 15764 2990 15792 3800
rect 16040 3194 16068 3800
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16316 3108 16344 3800
rect 16592 3210 16620 3800
rect 16592 3182 16712 3210
rect 16580 3120 16632 3126
rect 16316 3080 16580 3108
rect 16580 3062 16632 3068
rect 16684 3058 16712 3182
rect 16868 3176 16896 3800
rect 16948 3188 17000 3194
rect 16868 3148 16948 3176
rect 16948 3130 17000 3136
rect 17144 3108 17172 3800
rect 17224 3120 17276 3126
rect 17144 3080 17224 3108
rect 17224 3062 17276 3068
rect 16672 3052 16724 3058
rect 17420 3040 17448 3800
rect 17696 3176 17724 3800
rect 17776 3188 17828 3194
rect 17696 3148 17776 3176
rect 17776 3130 17828 3136
rect 17500 3052 17552 3058
rect 17420 3012 17500 3040
rect 16672 2994 16724 3000
rect 17500 2994 17552 3000
rect 17972 2990 18000 3800
rect 18248 3108 18276 3800
rect 18524 3176 18552 3800
rect 18604 3188 18656 3194
rect 18524 3148 18604 3176
rect 18604 3130 18656 3136
rect 18328 3120 18380 3126
rect 18248 3080 18328 3108
rect 18328 3062 18380 3068
rect 18800 3074 18828 3800
rect 19076 3108 19104 3800
rect 19352 3482 19380 3800
rect 19352 3454 19564 3482
rect 19156 3120 19208 3126
rect 19076 3080 19156 3108
rect 18800 3058 18920 3074
rect 19156 3062 19208 3068
rect 18800 3052 18932 3058
rect 18800 3046 18880 3052
rect 18880 2994 18932 3000
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 13238 2292 13260 2348
rect 13316 2292 13338 2348
rect 13238 2202 13338 2292
rect 13238 2150 13262 2202
rect 13314 2150 13338 2202
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 7238 1606 7262 1658
rect 7314 1606 7338 1658
rect 7238 1268 7338 1606
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7238 1212 7260 1268
rect 7316 1212 7338 1268
rect 7238 1040 7338 1212
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 7392 626 7420 1158
rect 7208 600 7420 626
rect 7484 600 7512 1294
rect 7748 1284 7800 1290
rect 7748 1226 7800 1232
rect 8300 1284 8352 1290
rect 8300 1226 8352 1232
rect 8852 1284 8904 1290
rect 8852 1226 8904 1232
rect 7760 600 7788 1226
rect 8024 1216 8076 1222
rect 8024 1158 8076 1164
rect 8036 600 8064 1158
rect 8312 600 8340 1226
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 8588 600 8616 1158
rect 8864 600 8892 1226
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9232 626 9260 1158
rect 9140 600 9260 626
rect 9416 600 9444 1838
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 11336 1352 11388 1358
rect 11336 1294 11388 1300
rect 9692 600 9720 1294
rect 10232 1284 10284 1290
rect 10232 1226 10284 1232
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 9956 1216 10008 1222
rect 9956 1158 10008 1164
rect 9968 600 9996 1158
rect 10244 600 10272 1226
rect 10508 1216 10560 1222
rect 10508 1158 10560 1164
rect 10520 600 10548 1158
rect 10796 600 10824 1226
rect 11060 1216 11112 1222
rect 11060 1158 11112 1164
rect 11072 600 11100 1158
rect 11348 600 11376 1294
rect 11624 600 11652 1838
rect 12992 1352 13044 1358
rect 12992 1294 13044 1300
rect 11888 1284 11940 1290
rect 12808 1284 12860 1290
rect 11888 1226 11940 1232
rect 12728 1244 12808 1272
rect 11900 600 11928 1226
rect 12164 1216 12216 1222
rect 12164 1158 12216 1164
rect 12176 600 12204 1158
rect 12440 740 12492 746
rect 12440 682 12492 688
rect 12452 600 12480 682
rect 12728 600 12756 1244
rect 12808 1226 12860 1232
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12912 746 12940 1158
rect 12900 740 12952 746
rect 12900 682 12952 688
rect 13004 600 13032 1294
rect 13238 1114 13338 2150
rect 19238 2746 19338 3312
rect 19536 3194 19564 3454
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19628 2990 19656 3800
rect 19904 3058 19932 3800
rect 20180 3126 20208 3800
rect 20456 3194 20484 3800
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 20732 2990 20760 3800
rect 21008 3058 21036 3800
rect 21284 3126 21312 3800
rect 21560 3194 21588 3800
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21836 3074 21864 3800
rect 22112 3176 22140 3800
rect 22112 3148 22232 3176
rect 21836 3058 22140 3074
rect 20996 3052 21048 3058
rect 21836 3052 22152 3058
rect 21836 3046 22100 3052
rect 20996 2994 21048 3000
rect 22100 2994 22152 3000
rect 22204 2990 22232 3148
rect 22388 3126 22416 3800
rect 22664 3194 22692 3800
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22940 3058 22968 3800
rect 23216 3176 23244 3800
rect 23492 3210 23520 3800
rect 23492 3182 23612 3210
rect 23768 3194 23796 3800
rect 23216 3148 23428 3176
rect 23400 3108 23428 3148
rect 23480 3120 23532 3126
rect 23400 3080 23480 3108
rect 23480 3062 23532 3068
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23584 2990 23612 3182
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 24044 3058 24072 3800
rect 24320 3126 24348 3800
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24596 3074 24624 3800
rect 24872 3398 24900 3800
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 25148 3194 25176 3800
rect 25238 3290 25338 3312
rect 25238 3238 25262 3290
rect 25314 3238 25338 3290
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 24032 3052 24084 3058
rect 24596 3046 24900 3074
rect 24032 2994 24084 3000
rect 24872 2990 24900 3046
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 19238 2694 19262 2746
rect 19314 2694 19338 2746
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13238 1062 13262 1114
rect 13314 1062 13338 1114
rect 13238 1040 13338 1062
rect 13464 626 13492 1158
rect 13280 600 13492 626
rect 13556 600 13584 1838
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 15752 1352 15804 1358
rect 15752 1294 15804 1300
rect 13832 600 13860 1294
rect 14096 1284 14148 1290
rect 14740 1284 14792 1290
rect 14096 1226 14148 1232
rect 14660 1244 14740 1272
rect 14108 600 14136 1226
rect 14372 1216 14424 1222
rect 14372 1158 14424 1164
rect 14384 600 14412 1158
rect 14660 600 14688 1244
rect 15292 1284 15344 1290
rect 14740 1226 14792 1232
rect 15212 1244 15292 1272
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15028 626 15056 1158
rect 14936 600 15056 626
rect 15212 600 15240 1244
rect 15292 1226 15344 1232
rect 15476 740 15528 746
rect 15476 682 15528 688
rect 15488 600 15516 682
rect 15764 600 15792 1294
rect 16028 1216 16080 1222
rect 16028 1158 16080 1164
rect 16040 746 16068 1158
rect 16028 740 16080 746
rect 16028 682 16080 688
rect 16132 626 16160 1838
rect 19238 1658 19338 2694
rect 25238 2348 25338 3238
rect 25424 3040 25452 3800
rect 25504 3052 25556 3058
rect 25424 3012 25504 3040
rect 25504 2994 25556 3000
rect 25700 2938 25728 3800
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 25884 2990 25912 3334
rect 25976 3126 26004 3800
rect 26252 3210 26280 3800
rect 26252 3194 26372 3210
rect 26252 3188 26384 3194
rect 26252 3182 26332 3188
rect 26332 3130 26384 3136
rect 25964 3120 26016 3126
rect 25964 3062 26016 3068
rect 26528 3074 26556 3800
rect 26528 3058 26648 3074
rect 26528 3052 26660 3058
rect 26528 3046 26608 3052
rect 26608 2994 26660 3000
rect 25872 2984 25924 2990
rect 25700 2922 25820 2938
rect 26804 2972 26832 3800
rect 27080 3210 27108 3800
rect 27356 3210 27384 3800
rect 27632 3346 27660 3800
rect 27632 3318 27844 3346
rect 27080 3182 27292 3210
rect 27356 3194 27660 3210
rect 27356 3188 27672 3194
rect 27356 3182 27620 3188
rect 27264 3126 27292 3182
rect 27620 3130 27672 3136
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 27816 3058 27844 3318
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 26884 2984 26936 2990
rect 26804 2944 26884 2972
rect 25872 2926 25924 2932
rect 27908 2972 27936 3800
rect 28080 2984 28132 2990
rect 27908 2944 28080 2972
rect 26884 2926 26936 2932
rect 28080 2926 28132 2932
rect 28184 2922 28212 3800
rect 25700 2916 25832 2922
rect 25700 2910 25780 2916
rect 25780 2858 25832 2864
rect 28172 2916 28224 2922
rect 28172 2858 28224 2864
rect 28460 2514 28488 3800
rect 28736 3194 28764 3800
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 29012 3126 29040 3800
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 29288 3058 29316 3800
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 29564 2990 29592 3800
rect 29840 3194 29868 3800
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 30116 3126 30144 3800
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 30392 3058 30420 3800
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30668 2990 30696 3800
rect 30944 3194 30972 3800
rect 31220 3380 31248 3800
rect 31496 3482 31524 3800
rect 31772 3618 31800 3800
rect 32048 3754 32076 3800
rect 32048 3726 32168 3754
rect 31772 3590 32076 3618
rect 31496 3454 31892 3482
rect 31220 3352 31800 3380
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 31238 2746 31338 3312
rect 31772 3126 31800 3352
rect 31760 3120 31812 3126
rect 31760 3062 31812 3068
rect 31864 3058 31892 3454
rect 32048 3194 32076 3590
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 32140 2990 32168 3726
rect 32324 3108 32352 3800
rect 32404 3120 32456 3126
rect 32324 3080 32404 3108
rect 32404 3062 32456 3068
rect 32600 3074 32628 3800
rect 32876 3346 32904 3800
rect 33152 3482 33180 3800
rect 33152 3454 33272 3482
rect 32876 3318 33180 3346
rect 33152 3194 33180 3318
rect 33140 3188 33192 3194
rect 33140 3130 33192 3136
rect 32600 3058 32720 3074
rect 32600 3052 32732 3058
rect 32600 3046 32680 3052
rect 32680 2994 32732 3000
rect 33244 2990 33272 3454
rect 33428 3108 33456 3800
rect 33508 3120 33560 3126
rect 33428 3080 33508 3108
rect 33508 3062 33560 3068
rect 33704 3074 33732 3800
rect 33980 3210 34008 3800
rect 33980 3194 34100 3210
rect 33980 3188 34112 3194
rect 33980 3182 34060 3188
rect 34060 3130 34112 3136
rect 33704 3058 33824 3074
rect 33704 3052 33836 3058
rect 33704 3046 33784 3052
rect 33784 2994 33836 3000
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 33232 2984 33284 2990
rect 34256 2972 34284 3800
rect 34532 3074 34560 3800
rect 34808 3126 34836 3800
rect 34796 3120 34848 3126
rect 34532 3046 34652 3074
rect 34796 3062 34848 3068
rect 35084 3058 35112 3800
rect 35360 3194 35388 3800
rect 35348 3188 35400 3194
rect 35348 3130 35400 3136
rect 34520 2984 34572 2990
rect 34256 2944 34520 2972
rect 33232 2926 33284 2932
rect 34520 2926 34572 2932
rect 34624 2922 34652 3046
rect 35072 3052 35124 3058
rect 35072 2994 35124 3000
rect 35636 2972 35664 3800
rect 35912 3074 35940 3800
rect 35912 3046 36032 3074
rect 35900 2984 35952 2990
rect 35636 2944 35900 2972
rect 35900 2926 35952 2932
rect 36004 2922 36032 3046
rect 34612 2916 34664 2922
rect 34612 2858 34664 2864
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 31238 2694 31262 2746
rect 31314 2694 31338 2746
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 25238 2292 25260 2348
rect 25316 2292 25338 2348
rect 25238 2202 25338 2292
rect 25238 2150 25262 2202
rect 25314 2150 25338 2202
rect 19616 1896 19668 1902
rect 19616 1838 19668 1844
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 24308 1896 24360 1902
rect 24308 1838 24360 1844
rect 19238 1606 19262 1658
rect 19314 1606 19338 1658
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 17684 1352 17736 1358
rect 17684 1294 17736 1300
rect 16580 1284 16632 1290
rect 16580 1226 16632 1232
rect 16396 1216 16448 1222
rect 16396 1158 16448 1164
rect 16408 626 16436 1158
rect 16040 600 16160 626
rect 16316 600 16436 626
rect 16592 600 16620 1226
rect 16868 600 16896 1294
rect 17408 1284 17460 1290
rect 17408 1226 17460 1232
rect 17132 1216 17184 1222
rect 17132 1158 17184 1164
rect 17144 600 17172 1158
rect 17420 600 17448 1226
rect 17696 600 17724 1294
rect 17960 1284 18012 1290
rect 17960 1226 18012 1232
rect 19064 1284 19116 1290
rect 19064 1226 19116 1232
rect 19238 1268 19338 1606
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 17972 600 18000 1226
rect 18236 1216 18288 1222
rect 18972 1216 19024 1222
rect 18236 1158 18288 1164
rect 18524 1176 18972 1204
rect 18248 600 18276 1158
rect 18524 600 18552 1176
rect 18972 1158 19024 1164
rect 18788 740 18840 746
rect 18788 682 18840 688
rect 18800 600 18828 682
rect 19076 600 19104 1226
rect 19238 1212 19260 1268
rect 19316 1212 19338 1268
rect 19238 1040 19338 1212
rect 19444 626 19472 1294
rect 19352 600 19472 626
rect 19628 600 19656 1838
rect 20168 1352 20220 1358
rect 20168 1294 20220 1300
rect 20996 1352 21048 1358
rect 20996 1294 21048 1300
rect 19892 1284 19944 1290
rect 19892 1226 19944 1232
rect 19904 600 19932 1226
rect 20180 600 20208 1294
rect 20720 1284 20772 1290
rect 20720 1226 20772 1232
rect 20260 1216 20312 1222
rect 20628 1216 20680 1222
rect 20260 1158 20312 1164
rect 20456 1176 20628 1204
rect 20272 746 20300 1158
rect 20260 740 20312 746
rect 20260 682 20312 688
rect 20456 600 20484 1176
rect 20628 1158 20680 1164
rect 20732 600 20760 1226
rect 21008 600 21036 1294
rect 21272 1216 21324 1222
rect 21272 1158 21324 1164
rect 21284 600 21312 1158
rect 21560 600 21588 1838
rect 22376 1352 22428 1358
rect 22376 1294 22428 1300
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 21824 1284 21876 1290
rect 21824 1226 21876 1232
rect 21836 600 21864 1226
rect 22100 1216 22152 1222
rect 22100 1158 22152 1164
rect 22112 600 22140 1158
rect 22388 600 22416 1294
rect 22652 1284 22704 1290
rect 22652 1226 22704 1232
rect 22928 1284 22980 1290
rect 22928 1226 22980 1232
rect 22664 600 22692 1226
rect 22940 600 22968 1226
rect 23388 1216 23440 1222
rect 23216 1176 23388 1204
rect 23216 600 23244 1176
rect 23388 1158 23440 1164
rect 23492 600 23520 1294
rect 23756 1284 23808 1290
rect 23756 1226 23808 1232
rect 23768 600 23796 1226
rect 24032 1216 24084 1222
rect 24032 1158 24084 1164
rect 24044 600 24072 1158
rect 24320 600 24348 1838
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 24676 1284 24728 1290
rect 24676 1226 24728 1232
rect 24688 626 24716 1226
rect 24596 600 24716 626
rect 24872 600 24900 1294
rect 25136 1216 25188 1222
rect 25136 1158 25188 1164
rect 25148 600 25176 1158
rect 25238 1114 25338 2150
rect 28448 1896 28500 1902
rect 28448 1838 28500 1844
rect 30656 1896 30708 1902
rect 30656 1838 30708 1844
rect 26516 1420 26568 1426
rect 26516 1362 26568 1368
rect 27896 1420 27948 1426
rect 27896 1362 27948 1368
rect 25964 1352 26016 1358
rect 25964 1294 26016 1300
rect 25688 1284 25740 1290
rect 25688 1226 25740 1232
rect 25238 1062 25262 1114
rect 25314 1062 25338 1114
rect 25238 1040 25338 1062
rect 25412 740 25464 746
rect 25412 682 25464 688
rect 25424 600 25452 682
rect 25700 600 25728 1226
rect 25976 600 26004 1294
rect 26148 1216 26200 1222
rect 26148 1158 26200 1164
rect 26240 1216 26292 1222
rect 26240 1158 26292 1164
rect 26160 746 26188 1158
rect 26148 740 26200 746
rect 26148 682 26200 688
rect 26252 600 26280 1158
rect 26528 600 26556 1362
rect 27344 1352 27396 1358
rect 27344 1294 27396 1300
rect 26792 1284 26844 1290
rect 26792 1226 26844 1232
rect 26804 600 26832 1226
rect 27068 740 27120 746
rect 27068 682 27120 688
rect 27080 600 27108 682
rect 27356 600 27384 1294
rect 27620 1284 27672 1290
rect 27620 1226 27672 1232
rect 27632 600 27660 1226
rect 27908 600 27936 1362
rect 28172 1284 28224 1290
rect 28172 1226 28224 1232
rect 28184 600 28212 1226
rect 28460 600 28488 1838
rect 29552 1352 29604 1358
rect 29552 1294 29604 1300
rect 29000 1284 29052 1290
rect 29000 1226 29052 1232
rect 28632 1216 28684 1222
rect 28632 1158 28684 1164
rect 28724 1216 28776 1222
rect 28724 1158 28776 1164
rect 28644 746 28672 1158
rect 28632 740 28684 746
rect 28632 682 28684 688
rect 28736 600 28764 1158
rect 29012 600 29040 1226
rect 29276 808 29328 814
rect 29276 750 29328 756
rect 29288 600 29316 750
rect 29564 600 29592 1294
rect 29920 1284 29972 1290
rect 29840 1244 29920 1272
rect 29840 600 29868 1244
rect 29920 1226 29972 1232
rect 30380 1216 30432 1222
rect 30380 1158 30432 1164
rect 30104 740 30156 746
rect 30104 682 30156 688
rect 30116 600 30144 682
rect 30392 600 30420 1158
rect 30668 600 30696 1838
rect 31238 1658 31338 2694
rect 36188 2514 36216 3800
rect 36464 3126 36492 3800
rect 36740 3194 36768 3800
rect 36728 3188 36780 3194
rect 36728 3130 36780 3136
rect 36452 3120 36504 3126
rect 36452 3062 36504 3068
rect 37016 3058 37044 3800
rect 37292 3482 37320 3800
rect 37292 3454 37412 3482
rect 37238 3290 37338 3312
rect 37238 3238 37262 3290
rect 37314 3238 37338 3290
rect 37004 3052 37056 3058
rect 37004 2994 37056 3000
rect 36176 2508 36228 2514
rect 36176 2450 36228 2456
rect 37238 2348 37338 3238
rect 37384 2990 37412 3454
rect 37568 3126 37596 3800
rect 37844 3194 37872 3800
rect 37832 3188 37884 3194
rect 37832 3130 37884 3136
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 38120 3058 38148 3800
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 38396 2990 38424 3800
rect 38672 3126 38700 3800
rect 38948 3194 38976 3800
rect 38936 3188 38988 3194
rect 38936 3130 38988 3136
rect 38660 3120 38712 3126
rect 38660 3062 38712 3068
rect 39224 3058 39252 3800
rect 39212 3052 39264 3058
rect 39212 2994 39264 3000
rect 39500 2990 39528 3800
rect 39776 3126 39804 3800
rect 40052 3176 40080 3800
rect 40132 3188 40184 3194
rect 40052 3148 40132 3176
rect 40132 3130 40184 3136
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 40328 3074 40356 3800
rect 40328 3058 40448 3074
rect 40328 3052 40460 3058
rect 40328 3046 40408 3052
rect 40408 2994 40460 3000
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 38384 2984 38436 2990
rect 38384 2926 38436 2932
rect 39488 2984 39540 2990
rect 40604 2972 40632 3800
rect 40684 2984 40736 2990
rect 40604 2944 40684 2972
rect 39488 2926 39540 2932
rect 40684 2926 40736 2932
rect 40880 2922 40908 3800
rect 41156 3176 41184 3800
rect 41236 3188 41288 3194
rect 41156 3148 41236 3176
rect 41236 3130 41288 3136
rect 40868 2916 40920 2922
rect 40868 2858 40920 2864
rect 41432 2514 41460 3800
rect 41708 3194 41736 3800
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 41984 3126 42012 3800
rect 41972 3120 42024 3126
rect 41972 3062 42024 3068
rect 42260 3074 42288 3800
rect 42536 3176 42564 3800
rect 42812 3346 42840 3800
rect 42812 3318 42932 3346
rect 42800 3188 42852 3194
rect 42536 3148 42800 3176
rect 42800 3130 42852 3136
rect 42260 3058 42380 3074
rect 42260 3052 42392 3058
rect 42260 3046 42340 3052
rect 42340 2994 42392 3000
rect 42904 2990 42932 3318
rect 43088 3126 43116 3800
rect 43364 3482 43392 3800
rect 43364 3454 43576 3482
rect 43076 3120 43128 3126
rect 43076 3062 43128 3068
rect 42892 2984 42944 2990
rect 42892 2926 42944 2932
rect 43238 2746 43338 3312
rect 43548 3194 43576 3454
rect 43536 3188 43588 3194
rect 43536 3130 43588 3136
rect 43640 3058 43668 3800
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43916 2990 43944 3800
rect 43904 2984 43956 2990
rect 43904 2926 43956 2932
rect 43238 2694 43262 2746
rect 43314 2694 43338 2746
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 37238 2292 37260 2348
rect 37316 2292 37338 2348
rect 37238 2202 37338 2292
rect 37238 2150 37262 2202
rect 37314 2150 37338 2202
rect 31760 1896 31812 1902
rect 31760 1838 31812 1844
rect 31238 1606 31262 1658
rect 31314 1606 31338 1658
rect 30932 1352 30984 1358
rect 30932 1294 30984 1300
rect 30840 1216 30892 1222
rect 30840 1158 30892 1164
rect 30852 814 30880 1158
rect 30840 808 30892 814
rect 30840 750 30892 756
rect 30944 600 30972 1294
rect 31238 1268 31338 1606
rect 31024 1216 31076 1222
rect 31024 1158 31076 1164
rect 31238 1212 31260 1268
rect 31316 1212 31338 1268
rect 31036 746 31064 1158
rect 31238 1040 31338 1212
rect 31576 1216 31628 1222
rect 31404 1176 31576 1204
rect 31024 740 31076 746
rect 31024 682 31076 688
rect 31404 626 31432 1176
rect 31576 1158 31628 1164
rect 31484 740 31536 746
rect 31484 682 31536 688
rect 31220 600 31432 626
rect 31496 600 31524 682
rect 31772 600 31800 1838
rect 32312 1352 32364 1358
rect 33232 1352 33284 1358
rect 32312 1294 32364 1300
rect 33152 1312 33232 1340
rect 32036 1284 32088 1290
rect 32036 1226 32088 1232
rect 32048 600 32076 1226
rect 32324 600 32352 1294
rect 32956 1284 33008 1290
rect 32876 1244 32956 1272
rect 32404 1216 32456 1222
rect 32680 1216 32732 1222
rect 32404 1158 32456 1164
rect 32600 1176 32680 1204
rect 32416 746 32444 1158
rect 32404 740 32456 746
rect 32404 682 32456 688
rect 32600 600 32628 1176
rect 32680 1158 32732 1164
rect 32876 600 32904 1244
rect 32956 1226 33008 1232
rect 33152 600 33180 1312
rect 34060 1352 34112 1358
rect 33232 1294 33284 1300
rect 33980 1312 34060 1340
rect 33784 1284 33836 1290
rect 33704 1244 33784 1272
rect 33508 1216 33560 1222
rect 33428 1176 33508 1204
rect 33428 600 33456 1176
rect 33508 1158 33560 1164
rect 33704 600 33732 1244
rect 33784 1226 33836 1232
rect 33980 600 34008 1312
rect 34060 1294 34112 1300
rect 35624 1352 35676 1358
rect 36636 1352 36688 1358
rect 35624 1294 35676 1300
rect 36464 1312 36636 1340
rect 34612 1284 34664 1290
rect 34532 1244 34612 1272
rect 34336 1216 34388 1222
rect 34256 1176 34336 1204
rect 34256 600 34284 1176
rect 34336 1158 34388 1164
rect 34532 600 34560 1244
rect 34612 1226 34664 1232
rect 35348 1284 35400 1290
rect 35348 1226 35400 1232
rect 34796 808 34848 814
rect 34796 750 34848 756
rect 34808 600 34836 750
rect 35072 740 35124 746
rect 35072 682 35124 688
rect 35084 600 35112 682
rect 35360 600 35388 1226
rect 35636 600 35664 1294
rect 36360 1284 36412 1290
rect 36188 1244 36360 1272
rect 35716 1216 35768 1222
rect 35716 1158 35768 1164
rect 35808 1216 35860 1222
rect 36084 1216 36136 1222
rect 35808 1158 35860 1164
rect 35912 1176 36084 1204
rect 35728 814 35756 1158
rect 35716 808 35768 814
rect 35716 750 35768 756
rect 35820 746 35848 1158
rect 35808 740 35860 746
rect 35808 682 35860 688
rect 35912 600 35940 1176
rect 36084 1158 36136 1164
rect 36188 600 36216 1244
rect 36360 1226 36412 1232
rect 36464 600 36492 1312
rect 36636 1294 36688 1300
rect 36912 1216 36964 1222
rect 36740 1176 36912 1204
rect 36740 600 36768 1176
rect 36912 1158 36964 1164
rect 37238 1114 37338 2150
rect 43238 1658 43338 2694
rect 44192 2514 44220 3800
rect 44468 3194 44496 3800
rect 44456 3188 44508 3194
rect 44456 3130 44508 3136
rect 44744 3126 44772 3800
rect 44732 3120 44784 3126
rect 44732 3062 44784 3068
rect 45020 3058 45048 3800
rect 45008 3052 45060 3058
rect 45008 2994 45060 3000
rect 45296 2514 45324 3800
rect 45572 2514 45600 3800
rect 45848 2514 45876 3800
rect 46124 2514 46152 3800
rect 46400 2514 46428 3800
rect 46676 2514 46704 3800
rect 46952 2514 46980 3800
rect 47228 2514 47256 3800
rect 47504 3194 47532 3800
rect 47492 3188 47544 3194
rect 47492 3130 47544 3136
rect 47780 3058 47808 3800
rect 47768 3052 47820 3058
rect 47768 2994 47820 3000
rect 48056 2514 48084 3800
rect 48332 2514 48360 3800
rect 48608 3194 48636 3800
rect 48884 3194 48912 3800
rect 49160 3194 49188 3800
rect 49238 3290 49338 3312
rect 49238 3238 49262 3290
rect 49314 3238 49338 3290
rect 48596 3188 48648 3194
rect 48596 3130 48648 3136
rect 48872 3188 48924 3194
rect 48872 3130 48924 3136
rect 49148 3188 49200 3194
rect 49148 3130 49200 3136
rect 44180 2508 44232 2514
rect 44180 2450 44232 2456
rect 45284 2508 45336 2514
rect 45284 2450 45336 2456
rect 45560 2508 45612 2514
rect 45560 2450 45612 2456
rect 45836 2508 45888 2514
rect 45836 2450 45888 2456
rect 46112 2508 46164 2514
rect 46112 2450 46164 2456
rect 46388 2508 46440 2514
rect 46388 2450 46440 2456
rect 46664 2508 46716 2514
rect 46664 2450 46716 2456
rect 46940 2508 46992 2514
rect 46940 2450 46992 2456
rect 47216 2508 47268 2514
rect 47216 2450 47268 2456
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 48320 2508 48372 2514
rect 48320 2450 48372 2456
rect 49238 2348 49338 3238
rect 49436 3194 49464 3800
rect 49712 3194 49740 3800
rect 49988 3194 50016 3800
rect 49424 3188 49476 3194
rect 49424 3130 49476 3136
rect 49700 3188 49752 3194
rect 49700 3130 49752 3136
rect 49976 3188 50028 3194
rect 49976 3130 50028 3136
rect 50264 3126 50292 3800
rect 50540 3194 50568 3800
rect 50528 3188 50580 3194
rect 50816 3176 50844 3800
rect 51092 3346 51120 3800
rect 51092 3318 51212 3346
rect 51080 3188 51132 3194
rect 50816 3148 51080 3176
rect 50528 3130 50580 3136
rect 51080 3130 51132 3136
rect 50252 3120 50304 3126
rect 50252 3062 50304 3068
rect 51184 3058 51212 3318
rect 51368 3194 51396 3800
rect 51356 3188 51408 3194
rect 51356 3130 51408 3136
rect 51644 3126 51672 3800
rect 51920 3194 51948 3800
rect 51908 3188 51960 3194
rect 52196 3176 52224 3800
rect 52472 3346 52500 3800
rect 52472 3318 52592 3346
rect 52460 3188 52512 3194
rect 52196 3148 52460 3176
rect 51908 3130 51960 3136
rect 52460 3130 52512 3136
rect 51632 3120 51684 3126
rect 51632 3062 51684 3068
rect 52564 3058 52592 3318
rect 52748 3194 52776 3800
rect 52736 3188 52788 3194
rect 52736 3130 52788 3136
rect 53024 3126 53052 3800
rect 53300 3194 53328 3800
rect 53288 3188 53340 3194
rect 53576 3176 53604 3800
rect 53852 3346 53880 3800
rect 53852 3318 53972 3346
rect 53840 3188 53892 3194
rect 53576 3148 53840 3176
rect 53288 3130 53340 3136
rect 53840 3130 53892 3136
rect 53944 3126 53972 3318
rect 54128 3194 54156 3800
rect 54116 3188 54168 3194
rect 54116 3130 54168 3136
rect 54404 3126 54432 3800
rect 54680 3194 54708 3800
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54956 3126 54984 3800
rect 55232 3482 55260 3800
rect 55232 3454 55444 3482
rect 53012 3120 53064 3126
rect 53012 3062 53064 3068
rect 53932 3120 53984 3126
rect 53932 3062 53984 3068
rect 54392 3120 54444 3126
rect 54392 3062 54444 3068
rect 54944 3120 54996 3126
rect 54944 3062 54996 3068
rect 51172 3052 51224 3058
rect 51172 2994 51224 3000
rect 52552 3052 52604 3058
rect 52552 2994 52604 3000
rect 49238 2292 49260 2348
rect 49316 2292 49338 2348
rect 49238 2202 49338 2292
rect 49238 2150 49262 2202
rect 49314 2150 49338 2202
rect 45008 1964 45060 1970
rect 45008 1906 45060 1912
rect 43444 1896 43496 1902
rect 43444 1838 43496 1844
rect 44456 1896 44508 1902
rect 44456 1838 44508 1844
rect 43238 1606 43262 1658
rect 43314 1606 43338 1658
rect 38936 1420 38988 1426
rect 38936 1362 38988 1368
rect 41420 1420 41472 1426
rect 41420 1362 41472 1368
rect 37556 1352 37608 1358
rect 37476 1312 37556 1340
rect 37372 1284 37424 1290
rect 37372 1226 37424 1232
rect 37238 1062 37262 1114
rect 37314 1062 37338 1114
rect 37238 1040 37338 1062
rect 37384 762 37412 1226
rect 37016 734 37412 762
rect 37016 600 37044 734
rect 37476 626 37504 1312
rect 38384 1352 38436 1358
rect 37556 1294 37608 1300
rect 38212 1312 38384 1340
rect 38108 1284 38160 1290
rect 37936 1244 38108 1272
rect 37832 1216 37884 1222
rect 37292 600 37504 626
rect 37568 1176 37832 1204
rect 37568 600 37596 1176
rect 37832 1158 37884 1164
rect 37936 626 37964 1244
rect 38108 1226 38160 1232
rect 38212 626 38240 1312
rect 38384 1294 38436 1300
rect 38660 1216 38712 1222
rect 37844 600 37964 626
rect 38120 600 38240 626
rect 38396 1176 38660 1204
rect 38396 600 38424 1176
rect 38660 1158 38712 1164
rect 38660 740 38712 746
rect 38660 682 38712 688
rect 38672 600 38700 682
rect 38948 600 38976 1362
rect 39488 1352 39540 1358
rect 40776 1352 40828 1358
rect 39488 1294 39540 1300
rect 40604 1312 40776 1340
rect 39212 1284 39264 1290
rect 39212 1226 39264 1232
rect 39224 600 39252 1226
rect 39500 600 39528 1294
rect 39672 1216 39724 1222
rect 39672 1158 39724 1164
rect 39764 1216 39816 1222
rect 40500 1216 40552 1222
rect 39764 1158 39816 1164
rect 40328 1176 40500 1204
rect 39684 746 39712 1158
rect 39672 740 39724 746
rect 39672 682 39724 688
rect 39776 600 39804 1158
rect 40040 740 40092 746
rect 40040 682 40092 688
rect 40052 600 40080 682
rect 40328 600 40356 1176
rect 40500 1158 40552 1164
rect 40604 600 40632 1312
rect 40776 1294 40828 1300
rect 40880 1278 41368 1306
rect 40880 600 40908 1278
rect 41340 1222 41368 1278
rect 41236 1216 41288 1222
rect 41236 1158 41288 1164
rect 41328 1216 41380 1222
rect 41328 1158 41380 1164
rect 41144 808 41196 814
rect 41144 750 41196 756
rect 41156 600 41184 750
rect 41248 746 41276 1158
rect 41236 740 41288 746
rect 41236 682 41288 688
rect 41432 600 41460 1362
rect 43076 1352 43128 1358
rect 43076 1294 43128 1300
rect 42524 1284 42576 1290
rect 42524 1226 42576 1232
rect 42248 944 42300 950
rect 42248 886 42300 892
rect 41972 876 42024 882
rect 41972 818 42024 824
rect 41696 740 41748 746
rect 41696 682 41748 688
rect 41708 600 41736 682
rect 41984 600 42012 818
rect 42260 600 42288 886
rect 42536 600 42564 1226
rect 42616 1216 42668 1222
rect 42616 1158 42668 1164
rect 42800 1216 42852 1222
rect 42800 1158 42852 1164
rect 42628 814 42656 1158
rect 42616 808 42668 814
rect 42616 750 42668 756
rect 42812 746 42840 1158
rect 42800 740 42852 746
rect 42800 682 42852 688
rect 42892 672 42944 678
rect 42812 620 42892 626
rect 42812 614 42944 620
rect 42812 600 42932 614
rect 43088 600 43116 1294
rect 43238 1268 43338 1606
rect 43238 1212 43260 1268
rect 43316 1212 43338 1268
rect 43238 1040 43338 1212
rect 43456 898 43484 1838
rect 43628 1284 43680 1290
rect 43628 1226 43680 1232
rect 43364 870 43484 898
rect 43364 600 43392 870
rect 43640 600 43668 1226
rect 43812 1216 43864 1222
rect 43812 1158 43864 1164
rect 44088 1216 44140 1222
rect 44088 1158 44140 1164
rect 43824 882 43852 1158
rect 44100 950 44128 1158
rect 44088 944 44140 950
rect 44088 886 44140 892
rect 43812 876 43864 882
rect 43812 818 43864 824
rect 44180 808 44232 814
rect 44180 750 44232 756
rect 43904 740 43956 746
rect 43904 682 43956 688
rect 43916 600 43944 682
rect 44192 600 44220 750
rect 44468 600 44496 1838
rect 44732 1284 44784 1290
rect 44732 1226 44784 1232
rect 44640 1216 44692 1222
rect 44640 1158 44692 1164
rect 44652 678 44680 1158
rect 44640 672 44692 678
rect 44640 614 44692 620
rect 44744 600 44772 1226
rect 45020 600 45048 1906
rect 45836 1420 45888 1426
rect 45836 1362 45888 1368
rect 47400 1420 47452 1426
rect 47400 1362 47452 1368
rect 48872 1420 48924 1426
rect 48872 1362 48924 1368
rect 45284 1352 45336 1358
rect 45284 1294 45336 1300
rect 45296 600 45324 1294
rect 45468 1216 45520 1222
rect 45468 1158 45520 1164
rect 45560 1216 45612 1222
rect 45560 1158 45612 1164
rect 45480 746 45508 1158
rect 45468 740 45520 746
rect 45468 682 45520 688
rect 45572 600 45600 1158
rect 45848 600 45876 1362
rect 46480 1352 46532 1358
rect 46400 1312 46480 1340
rect 46112 1216 46164 1222
rect 46112 1158 46164 1164
rect 46204 1216 46256 1222
rect 46204 1158 46256 1164
rect 46124 814 46152 1158
rect 46112 808 46164 814
rect 46112 750 46164 756
rect 46216 626 46244 1158
rect 46124 600 46244 626
rect 46400 600 46428 1312
rect 46480 1294 46532 1300
rect 47308 1284 47360 1290
rect 47308 1226 47360 1232
rect 46940 1216 46992 1222
rect 46676 1176 46940 1204
rect 46676 600 46704 1176
rect 46940 1158 46992 1164
rect 47320 728 47348 1226
rect 46952 700 47348 728
rect 46952 600 46980 700
rect 47412 626 47440 1362
rect 48688 1352 48740 1358
rect 48516 1312 48688 1340
rect 48412 1284 48464 1290
rect 48412 1226 48464 1232
rect 48136 1216 48188 1222
rect 47228 600 47440 626
rect 47504 1176 48136 1204
rect 47504 600 47532 1176
rect 48136 1158 48188 1164
rect 47768 740 47820 746
rect 48424 728 48452 1226
rect 47768 682 47820 688
rect 48056 700 48452 728
rect 47780 600 47808 682
rect 48056 600 48084 700
rect 48516 626 48544 1312
rect 48688 1294 48740 1300
rect 48596 808 48648 814
rect 48596 750 48648 756
rect 48332 600 48544 626
rect 48608 600 48636 750
rect 48884 600 48912 1362
rect 49148 1216 49200 1222
rect 49148 1158 49200 1164
rect 49160 746 49188 1158
rect 49238 1114 49338 2150
rect 55238 2746 55338 3312
rect 55416 3194 55444 3454
rect 55404 3188 55456 3194
rect 55404 3130 55456 3136
rect 55508 2990 55536 3800
rect 55784 3058 55812 3800
rect 56060 3194 56088 3800
rect 56048 3188 56100 3194
rect 56048 3130 56100 3136
rect 56336 3074 56364 3800
rect 56612 3210 56640 3800
rect 56612 3194 56732 3210
rect 56612 3188 56744 3194
rect 56612 3182 56692 3188
rect 56692 3130 56744 3136
rect 56888 3108 56916 3800
rect 56968 3120 57020 3126
rect 56888 3080 56968 3108
rect 56336 3058 56640 3074
rect 56968 3062 57020 3068
rect 57164 3058 57192 3800
rect 57440 3210 57468 3800
rect 57716 3210 57744 3800
rect 57992 3346 58020 3800
rect 57992 3318 58112 3346
rect 57440 3194 57560 3210
rect 57440 3188 57572 3194
rect 57440 3182 57520 3188
rect 57716 3182 58020 3210
rect 57520 3130 57572 3136
rect 57992 3126 58020 3182
rect 57980 3120 58032 3126
rect 57980 3062 58032 3068
rect 58084 3058 58112 3318
rect 58268 3194 58296 3800
rect 58256 3188 58308 3194
rect 58256 3130 58308 3136
rect 58544 3126 58572 3800
rect 58532 3120 58584 3126
rect 58532 3062 58584 3068
rect 58820 3058 58848 3800
rect 59096 3194 59124 3800
rect 59084 3188 59136 3194
rect 59084 3130 59136 3136
rect 59372 3126 59400 3800
rect 59360 3120 59412 3126
rect 59360 3062 59412 3068
rect 59648 3058 59676 3800
rect 59924 3194 59952 3800
rect 59912 3188 59964 3194
rect 59912 3130 59964 3136
rect 60200 3126 60228 3800
rect 60476 3210 60504 3800
rect 60752 3346 60780 3800
rect 60752 3318 60872 3346
rect 60476 3194 60780 3210
rect 60476 3188 60792 3194
rect 60476 3182 60740 3188
rect 60740 3130 60792 3136
rect 60188 3120 60240 3126
rect 60188 3062 60240 3068
rect 60844 3058 60872 3318
rect 61028 3126 61056 3800
rect 61304 3482 61332 3800
rect 61304 3454 61424 3482
rect 61238 3290 61338 3312
rect 61238 3238 61262 3290
rect 61314 3238 61338 3290
rect 61016 3120 61068 3126
rect 61016 3062 61068 3068
rect 55772 3052 55824 3058
rect 56336 3052 56652 3058
rect 56336 3046 56600 3052
rect 55772 2994 55824 3000
rect 56600 2994 56652 3000
rect 57152 3052 57204 3058
rect 57152 2994 57204 3000
rect 58072 3052 58124 3058
rect 58072 2994 58124 3000
rect 58808 3052 58860 3058
rect 58808 2994 58860 3000
rect 59636 3052 59688 3058
rect 59636 2994 59688 3000
rect 60832 3052 60884 3058
rect 60832 2994 60884 3000
rect 55496 2984 55548 2990
rect 55496 2926 55548 2932
rect 55238 2694 55262 2746
rect 55314 2694 55338 2746
rect 51080 1896 51132 1902
rect 51080 1838 51132 1844
rect 49884 1420 49936 1426
rect 49884 1362 49936 1368
rect 50804 1420 50856 1426
rect 50804 1362 50856 1368
rect 49516 1284 49568 1290
rect 49516 1226 49568 1232
rect 49238 1062 49262 1114
rect 49314 1062 49338 1114
rect 49238 1040 49338 1062
rect 49148 740 49200 746
rect 49528 728 49556 1226
rect 49148 682 49200 688
rect 49252 700 49556 728
rect 49252 626 49280 700
rect 49896 626 49924 1362
rect 49976 1216 50028 1222
rect 49976 1158 50028 1164
rect 50068 1216 50120 1222
rect 50068 1158 50120 1164
rect 49988 814 50016 1158
rect 49976 808 50028 814
rect 49976 750 50028 756
rect 50080 626 50108 1158
rect 50528 808 50580 814
rect 50528 750 50580 756
rect 50252 740 50304 746
rect 50252 682 50304 688
rect 49160 600 49280 626
rect 49436 610 49556 626
rect 49436 604 49568 610
rect 49436 600 49516 604
rect 4066 575 4122 584
rect 4158 0 4214 600
rect 4434 598 4568 600
rect 4434 0 4490 598
rect 4710 0 4766 600
rect 4986 0 5042 600
rect 5262 0 5318 600
rect 5538 0 5594 600
rect 5814 0 5870 600
rect 6090 598 6224 600
rect 6090 0 6146 598
rect 6366 0 6422 600
rect 6642 0 6698 600
rect 6918 0 6974 600
rect 7194 598 7420 600
rect 7194 0 7250 598
rect 7470 0 7526 600
rect 7746 0 7802 600
rect 8022 0 8078 600
rect 8298 0 8354 600
rect 8574 0 8630 600
rect 8850 0 8906 600
rect 9126 598 9260 600
rect 9126 0 9182 598
rect 9402 0 9458 600
rect 9678 0 9734 600
rect 9954 0 10010 600
rect 10230 0 10286 600
rect 10506 0 10562 600
rect 10782 0 10838 600
rect 11058 0 11114 600
rect 11334 0 11390 600
rect 11610 0 11666 600
rect 11886 0 11942 600
rect 12162 0 12218 600
rect 12438 0 12494 600
rect 12714 0 12770 600
rect 12990 0 13046 600
rect 13266 598 13492 600
rect 13266 0 13322 598
rect 13542 0 13598 600
rect 13818 0 13874 600
rect 14094 0 14150 600
rect 14370 0 14426 600
rect 14646 0 14702 600
rect 14922 598 15056 600
rect 14922 0 14978 598
rect 15198 0 15254 600
rect 15474 0 15530 600
rect 15750 0 15806 600
rect 16026 598 16160 600
rect 16302 598 16436 600
rect 16026 0 16082 598
rect 16302 0 16358 598
rect 16578 0 16634 600
rect 16854 0 16910 600
rect 17130 0 17186 600
rect 17406 0 17462 600
rect 17682 0 17738 600
rect 17958 0 18014 600
rect 18234 0 18290 600
rect 18510 0 18566 600
rect 18786 0 18842 600
rect 19062 0 19118 600
rect 19338 598 19472 600
rect 19338 0 19394 598
rect 19614 0 19670 600
rect 19890 0 19946 600
rect 20166 0 20222 600
rect 20442 0 20498 600
rect 20718 0 20774 600
rect 20994 0 21050 600
rect 21270 0 21326 600
rect 21546 0 21602 600
rect 21822 0 21878 600
rect 22098 0 22154 600
rect 22374 0 22430 600
rect 22650 0 22706 600
rect 22926 0 22982 600
rect 23202 0 23258 600
rect 23478 0 23534 600
rect 23754 0 23810 600
rect 24030 0 24086 600
rect 24306 0 24362 600
rect 24582 598 24716 600
rect 24582 0 24638 598
rect 24858 0 24914 600
rect 25134 0 25190 600
rect 25410 0 25466 600
rect 25686 0 25742 600
rect 25962 0 26018 600
rect 26238 0 26294 600
rect 26514 0 26570 600
rect 26790 0 26846 600
rect 27066 0 27122 600
rect 27342 0 27398 600
rect 27618 0 27674 600
rect 27894 0 27950 600
rect 28170 0 28226 600
rect 28446 0 28502 600
rect 28722 0 28778 600
rect 28998 0 29054 600
rect 29274 0 29330 600
rect 29550 0 29606 600
rect 29826 0 29882 600
rect 30102 0 30158 600
rect 30378 0 30434 600
rect 30654 0 30710 600
rect 30930 0 30986 600
rect 31206 598 31432 600
rect 31206 0 31262 598
rect 31482 0 31538 600
rect 31758 0 31814 600
rect 32034 0 32090 600
rect 32310 0 32366 600
rect 32586 0 32642 600
rect 32862 0 32918 600
rect 33138 0 33194 600
rect 33414 0 33470 600
rect 33690 0 33746 600
rect 33966 0 34022 600
rect 34242 0 34298 600
rect 34518 0 34574 600
rect 34794 0 34850 600
rect 35070 0 35126 600
rect 35346 0 35402 600
rect 35622 0 35678 600
rect 35898 0 35954 600
rect 36174 0 36230 600
rect 36450 0 36506 600
rect 36726 0 36782 600
rect 37002 0 37058 600
rect 37278 598 37504 600
rect 37278 0 37334 598
rect 37554 0 37610 600
rect 37830 598 37964 600
rect 38106 598 38240 600
rect 37830 0 37886 598
rect 38106 0 38162 598
rect 38382 0 38438 600
rect 38658 0 38714 600
rect 38934 0 38990 600
rect 39210 0 39266 600
rect 39486 0 39542 600
rect 39762 0 39818 600
rect 40038 0 40094 600
rect 40314 0 40370 600
rect 40590 0 40646 600
rect 40866 0 40922 600
rect 41142 0 41198 600
rect 41418 0 41474 600
rect 41694 0 41750 600
rect 41970 0 42026 600
rect 42246 0 42302 600
rect 42522 0 42578 600
rect 42798 598 42932 600
rect 42798 0 42854 598
rect 43074 0 43130 600
rect 43350 0 43406 600
rect 43626 0 43682 600
rect 43902 0 43958 600
rect 44178 0 44234 600
rect 44454 0 44510 600
rect 44730 0 44786 600
rect 45006 0 45062 600
rect 45282 0 45338 600
rect 45558 0 45614 600
rect 45834 0 45890 600
rect 46110 598 46244 600
rect 46110 0 46166 598
rect 46386 0 46442 600
rect 46662 0 46718 600
rect 46938 0 46994 600
rect 47214 598 47440 600
rect 47214 0 47270 598
rect 47490 0 47546 600
rect 47766 0 47822 600
rect 48042 0 48098 600
rect 48318 598 48544 600
rect 48318 0 48374 598
rect 48594 0 48650 600
rect 48870 0 48926 600
rect 49146 598 49280 600
rect 49422 598 49516 600
rect 49146 0 49202 598
rect 49422 0 49478 598
rect 49712 600 49924 626
rect 49988 600 50108 626
rect 50264 600 50292 682
rect 50540 600 50568 750
rect 50816 600 50844 1362
rect 50896 1216 50948 1222
rect 50896 1158 50948 1164
rect 50908 610 50936 1158
rect 50896 604 50948 610
rect 49516 546 49568 552
rect 49698 598 49924 600
rect 49974 598 50108 600
rect 49698 0 49754 598
rect 49974 0 50030 598
rect 50250 0 50306 600
rect 50526 0 50582 600
rect 50802 0 50858 600
rect 51092 600 51120 1838
rect 55238 1658 55338 2694
rect 55238 1606 55262 1658
rect 55314 1606 55338 1658
rect 51632 1352 51684 1358
rect 53012 1352 53064 1358
rect 51632 1294 51684 1300
rect 52748 1312 53012 1340
rect 51356 1284 51408 1290
rect 51356 1226 51408 1232
rect 51368 600 51396 1226
rect 51644 600 51672 1294
rect 52644 1284 52696 1290
rect 52644 1226 52696 1232
rect 51724 1216 51776 1222
rect 51724 1158 51776 1164
rect 51816 1216 51868 1222
rect 52368 1216 52420 1222
rect 51816 1158 51868 1164
rect 51920 1176 52368 1204
rect 51736 746 51764 1158
rect 51828 814 51856 1158
rect 51816 808 51868 814
rect 51816 750 51868 756
rect 51724 740 51776 746
rect 51724 682 51776 688
rect 51920 600 51948 1176
rect 52368 1158 52420 1164
rect 52656 728 52684 1226
rect 52196 700 52684 728
rect 52196 600 52224 700
rect 52472 610 52592 626
rect 52472 604 52604 610
rect 52472 600 52552 604
rect 50896 546 50948 552
rect 51078 0 51134 600
rect 51354 0 51410 600
rect 51630 0 51686 600
rect 51906 0 51962 600
rect 52182 0 52238 600
rect 52458 598 52552 600
rect 52458 0 52514 598
rect 52748 600 52776 1312
rect 54668 1352 54720 1358
rect 53012 1294 53064 1300
rect 53576 1278 53880 1306
rect 54668 1294 54720 1300
rect 53288 1216 53340 1222
rect 53024 1176 53288 1204
rect 53024 600 53052 1176
rect 53288 1158 53340 1164
rect 53288 876 53340 882
rect 53288 818 53340 824
rect 53300 600 53328 818
rect 53576 600 53604 1278
rect 53852 1222 53880 1278
rect 53748 1216 53800 1222
rect 53748 1158 53800 1164
rect 53840 1216 53892 1222
rect 53840 1158 53892 1164
rect 54576 1216 54628 1222
rect 54576 1158 54628 1164
rect 53760 610 53788 1158
rect 53840 944 53892 950
rect 53840 886 53892 892
rect 53748 604 53800 610
rect 52552 546 52604 552
rect 52734 0 52790 600
rect 53010 0 53066 600
rect 53286 0 53342 600
rect 53562 0 53618 600
rect 53852 600 53880 886
rect 54588 882 54616 1158
rect 54576 876 54628 882
rect 54576 818 54628 824
rect 54392 808 54444 814
rect 54392 750 54444 756
rect 54116 740 54168 746
rect 54116 682 54168 688
rect 54128 600 54156 682
rect 54404 600 54432 750
rect 54680 600 54708 1294
rect 54944 1284 54996 1290
rect 54944 1226 54996 1232
rect 55238 1268 55338 1606
rect 54956 600 54984 1226
rect 55128 1216 55180 1222
rect 55128 1158 55180 1164
rect 55238 1212 55260 1268
rect 55316 1212 55338 1268
rect 61238 2348 61338 3238
rect 61396 3194 61424 3454
rect 61384 3188 61436 3194
rect 61384 3130 61436 3136
rect 61580 3058 61608 3800
rect 61856 3210 61884 3800
rect 62132 3346 62160 3800
rect 62132 3318 62252 3346
rect 61856 3194 62160 3210
rect 61856 3188 62172 3194
rect 61856 3182 62120 3188
rect 62120 3130 62172 3136
rect 62224 3126 62252 3318
rect 62212 3120 62264 3126
rect 62212 3062 62264 3068
rect 62408 3058 62436 3800
rect 62684 3194 62712 3800
rect 62672 3188 62724 3194
rect 62672 3130 62724 3136
rect 62960 3126 62988 3800
rect 63236 3210 63264 3800
rect 63512 3346 63540 3800
rect 63512 3318 63632 3346
rect 63236 3182 63540 3210
rect 62948 3120 63000 3126
rect 62948 3062 63000 3068
rect 61568 3052 61620 3058
rect 61568 2994 61620 3000
rect 62396 3052 62448 3058
rect 62396 2994 62448 3000
rect 63512 2990 63540 3182
rect 63604 3058 63632 3318
rect 63592 3052 63644 3058
rect 63592 2994 63644 3000
rect 63500 2984 63552 2990
rect 63500 2926 63552 2932
rect 63788 2922 63816 3800
rect 64064 3126 64092 3800
rect 64340 3194 64368 3800
rect 64328 3188 64380 3194
rect 64328 3130 64380 3136
rect 64052 3120 64104 3126
rect 64052 3062 64104 3068
rect 64616 3074 64644 3800
rect 64616 3058 64736 3074
rect 64616 3052 64748 3058
rect 64616 3046 64696 3052
rect 64696 2994 64748 3000
rect 63776 2916 63828 2922
rect 63776 2858 63828 2864
rect 64892 2514 64920 3800
rect 65168 3210 65196 3800
rect 65168 3182 65288 3210
rect 65260 3126 65288 3182
rect 65248 3120 65300 3126
rect 65248 3062 65300 3068
rect 65444 2514 65472 3800
rect 65720 3194 65748 3800
rect 65708 3188 65760 3194
rect 65708 3130 65760 3136
rect 65996 2514 66024 3800
rect 66272 2514 66300 3800
rect 66548 3194 66576 3800
rect 66536 3188 66588 3194
rect 66536 3130 66588 3136
rect 66824 2514 66852 3800
rect 67100 3194 67128 3800
rect 67376 3346 67404 3800
rect 67376 3318 67496 3346
rect 67088 3188 67140 3194
rect 67088 3130 67140 3136
rect 67238 2746 67338 3312
rect 67468 3194 67496 3318
rect 67652 3194 67680 3800
rect 67456 3188 67508 3194
rect 67456 3130 67508 3136
rect 67640 3188 67692 3194
rect 67640 3130 67692 3136
rect 67928 3058 67956 3800
rect 67916 3052 67968 3058
rect 67916 2994 67968 3000
rect 67238 2694 67262 2746
rect 67314 2694 67338 2746
rect 64880 2508 64932 2514
rect 64880 2450 64932 2456
rect 65432 2508 65484 2514
rect 65432 2450 65484 2456
rect 65984 2508 66036 2514
rect 65984 2450 66036 2456
rect 66260 2508 66312 2514
rect 66260 2450 66312 2456
rect 66812 2508 66864 2514
rect 66812 2450 66864 2456
rect 61238 2292 61260 2348
rect 61316 2292 61338 2348
rect 61238 2202 61338 2292
rect 61238 2150 61262 2202
rect 61314 2150 61338 2202
rect 55140 950 55168 1158
rect 55238 1040 55338 1212
rect 55496 1216 55548 1222
rect 55496 1158 55548 1164
rect 56324 1216 56376 1222
rect 56324 1158 56376 1164
rect 55128 944 55180 950
rect 55128 886 55180 892
rect 55508 746 55536 1158
rect 56336 814 56364 1158
rect 61238 1114 61338 2150
rect 61238 1062 61262 1114
rect 61314 1062 61338 1114
rect 61238 1040 61338 1062
rect 67238 1658 67338 2694
rect 67238 1606 67262 1658
rect 67314 1606 67338 1658
rect 67238 1268 67338 1606
rect 67238 1212 67260 1268
rect 67316 1212 67338 1268
rect 67238 1040 67338 1212
rect 56324 808 56376 814
rect 56324 750 56376 756
rect 55496 740 55548 746
rect 55496 682 55548 688
rect 53748 546 53800 552
rect 53838 0 53894 600
rect 54114 0 54170 600
rect 54390 0 54446 600
rect 54666 0 54722 600
rect 54942 0 54998 600
<< via2 >>
rect 2962 3712 3018 3768
rect 3698 3304 3754 3360
rect 3790 3032 3846 3088
rect 4066 3712 4122 3768
rect 3974 3576 4030 3632
rect 4066 2488 4122 2544
rect 4250 2760 4306 2816
rect 2778 1980 2780 2000
rect 2780 1980 2832 2000
rect 2832 1980 2834 2000
rect 2778 1944 2834 1980
rect 2870 1672 2926 1728
rect 2962 1400 3018 1456
rect 3606 2080 3662 2136
rect 3514 856 3570 912
rect 3422 584 3478 640
rect 3698 992 3754 1048
rect 3790 584 3846 640
rect 4066 584 4122 640
rect 13260 2292 13316 2348
rect 7260 1212 7316 1268
rect 25260 2292 25316 2348
rect 19260 1212 19316 1268
rect 37260 2292 37316 2348
rect 31260 1212 31316 1268
rect 49260 2292 49316 2348
rect 43260 1212 43316 1268
rect 55260 1212 55316 1268
rect 61260 2292 61316 2348
rect 67260 1212 67316 1268
<< metal3 >>
rect 0 4178 600 4208
rect 0 4118 3618 4178
rect 0 4088 600 4118
rect 0 3906 600 3936
rect 0 3846 2882 3906
rect 0 3816 600 3846
rect 2822 3770 2882 3846
rect 2957 3770 3023 3773
rect 2822 3768 3023 3770
rect 2822 3712 2962 3768
rect 3018 3712 3023 3768
rect 2822 3710 3023 3712
rect 3558 3770 3618 4118
rect 4061 3770 4127 3773
rect 3558 3768 4127 3770
rect 3558 3712 4066 3768
rect 4122 3712 4127 3768
rect 3558 3710 4127 3712
rect 2957 3707 3023 3710
rect 4061 3707 4127 3710
rect 0 3634 600 3664
rect 3969 3634 4035 3637
rect 0 3632 4035 3634
rect 0 3576 3974 3632
rect 4030 3576 4035 3632
rect 0 3574 4035 3576
rect 0 3544 600 3574
rect 3969 3571 4035 3574
rect 0 3362 600 3392
rect 3693 3362 3759 3365
rect 0 3360 3759 3362
rect 0 3304 3698 3360
rect 3754 3304 3759 3360
rect 0 3302 3759 3304
rect 0 3272 600 3302
rect 3693 3299 3759 3302
rect 0 3090 600 3120
rect 3785 3090 3851 3093
rect 0 3088 3851 3090
rect 0 3032 3790 3088
rect 3846 3032 3851 3088
rect 0 3030 3851 3032
rect 0 3000 600 3030
rect 3785 3027 3851 3030
rect 0 2818 600 2848
rect 4245 2818 4311 2821
rect 0 2816 4311 2818
rect 0 2760 4250 2816
rect 4306 2760 4311 2816
rect 0 2758 4311 2760
rect 0 2728 600 2758
rect 4245 2755 4311 2758
rect 0 2546 600 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 600 2486
rect 4061 2483 4127 2486
rect 1288 2348 68816 2370
rect 0 2274 600 2304
rect 1288 2292 13260 2348
rect 13316 2292 25260 2348
rect 25316 2292 37260 2348
rect 37316 2292 49260 2348
rect 49316 2292 61260 2348
rect 61316 2292 68816 2348
rect 0 2214 1226 2274
rect 1288 2270 68816 2292
rect 0 2184 600 2214
rect 1166 2138 1226 2214
rect 3601 2138 3667 2141
rect 1166 2136 3667 2138
rect 1166 2080 3606 2136
rect 3662 2080 3667 2136
rect 1166 2078 3667 2080
rect 3601 2075 3667 2078
rect 0 2002 600 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 600 1942
rect 2773 1939 2839 1942
rect 0 1730 600 1760
rect 2865 1730 2931 1733
rect 0 1728 2931 1730
rect 0 1672 2870 1728
rect 2926 1672 2931 1728
rect 0 1670 2931 1672
rect 0 1640 600 1670
rect 2865 1667 2931 1670
rect 0 1458 600 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 600 1398
rect 2957 1395 3023 1398
rect 1288 1268 68816 1290
rect 0 1186 600 1216
rect 1288 1212 7260 1268
rect 7316 1212 19260 1268
rect 19316 1212 31260 1268
rect 31316 1212 43260 1268
rect 43316 1212 55260 1268
rect 55316 1212 67260 1268
rect 67316 1212 68816 1268
rect 1288 1190 68816 1212
rect 0 1126 1226 1186
rect 0 1096 600 1126
rect 1166 1050 1226 1126
rect 3693 1050 3759 1053
rect 1166 1048 3759 1050
rect 1166 992 3698 1048
rect 3754 992 3759 1048
rect 1166 990 3759 992
rect 3693 987 3759 990
rect 0 914 600 944
rect 3509 914 3575 917
rect 0 912 3575 914
rect 0 856 3514 912
rect 3570 856 3575 912
rect 0 854 3575 856
rect 0 824 600 854
rect 3509 851 3575 854
rect 0 642 600 672
rect 3417 642 3483 645
rect 3785 642 3851 645
rect 4061 642 4127 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 0 552 600 582
rect 3417 579 3483 582
rect 3558 640 3851 642
rect 3558 584 3790 640
rect 3846 584 3851 640
rect 3558 582 3851 584
rect 0 370 600 400
rect 3558 370 3618 582
rect 3785 579 3851 582
rect 3926 640 4127 642
rect 3926 584 4066 640
rect 4122 584 4127 640
rect 3926 582 4127 584
rect 0 310 3618 370
rect 0 280 600 310
rect 0 98 600 128
rect 3926 98 3986 582
rect 4061 579 4127 582
rect 0 38 3986 98
rect 0 8 600 38
use sky130_fd_sc_hd__conb_1  insts\[327\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform -1 0 2208 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[321\]
timestamp 1637331468
transform 1 0 2208 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[2\]
timestamp 1637331468
transform -1 0 1932 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[297\]
timestamp 1637331468
transform -1 0 2208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[288\]
timestamp 1637331468
transform -1 0 2484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 1288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1637331468
transform 1 0 1288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 1564 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 1564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[28\]
timestamp 1637331468
transform -1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[284\]
timestamp 1637331468
transform 1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[260\]
timestamp 1637331468
transform 1 0 2484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[228\]
timestamp 1637331468
transform 1 0 2760 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[280\]
timestamp 1637331468
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[210\]
timestamp 1637331468
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[17\]
timestamp 1637331468
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[158\]
timestamp 1637331468
transform 1 0 3312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[156\]
timestamp 1637331468
transform 1 0 3588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[113\]
timestamp 1637331468
transform 1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[155\]
timestamp 1637331468
transform 1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[111\]
timestamp 1637331468
transform 1 0 4692 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[110\]
timestamp 1637331468
transform 1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[109\]
timestamp 1637331468
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[107\]
timestamp 1637331468
transform 1 0 4692 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[106\]
timestamp 1637331468
transform 1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[103\]
timestamp 1637331468
transform 1 0 4140 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 3956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[262\]
timestamp 1637331468
transform 1 0 5520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[222\]
timestamp 1637331468
transform 1 0 5796 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[209\]
timestamp 1637331468
transform 1 0 5796 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[206\]
timestamp 1637331468
transform 1 0 5520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[18\]
timestamp 1637331468
transform 1 0 5244 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[161\]
timestamp 1637331468
transform 1 0 5244 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[112\]
timestamp 1637331468
transform 1 0 4968 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[108\]
timestamp 1637331468
transform 1 0 4968 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1637331468
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1637331468
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[277\]
timestamp 1637331468
transform 1 0 6072 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[214\]
timestamp 1637331468
transform 1 0 6072 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1637331468
transform 1 0 6532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_9
timestamp 1637331468
transform 1 0 6440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1637331468
transform 1 0 6440 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[291\]
timestamp 1637331468
transform 1 0 6532 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[177\]
timestamp 1637331468
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[31\]
timestamp 1637331468
transform 1 0 6808 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[185\]
timestamp 1637331468
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1637331468
transform 1 0 7084 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[26\]
timestamp 1637331468
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[282\]
timestamp 1637331468
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[271\]
timestamp 1637331468
transform 1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[221\]
timestamp 1637331468
transform 1 0 7820 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[168\]
timestamp 1637331468
transform 1 0 8096 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 7544 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1637331468
transform 1 0 8372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1637331468
transform 1 0 7452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[329\]
timestamp 1637331468
transform 1 0 8464 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[195\]
timestamp 1637331468
transform 1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[179\]
timestamp 1637331468
transform 1 0 8740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[169\]
timestamp 1637331468
transform 1 0 9108 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10
timestamp 1637331468
transform 1 0 9016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1637331468
transform 1 0 8648 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[336\]
timestamp 1637331468
transform 1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[335\]
timestamp 1637331468
transform 1 0 10396 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[293\]
timestamp 1637331468
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[196\]
timestamp 1637331468
transform 1 0 9660 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[174\]
timestamp 1637331468
transform 1 0 10672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1637331468
transform 1 0 9936 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1637331468
transform 1 0 10120 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1637331468
transform 1 0 9752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[273\]
timestamp 1637331468
transform 1 0 10948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[171\]
timestamp 1637331468
transform 1 0 11224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[166\]
timestamp 1637331468
transform 1 0 11684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1637331468
transform 1 0 11592 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_11
timestamp 1637331468
transform 1 0 11592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1637331468
transform 1 0 11684 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1637331468
transform 1 0 11224 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1637331468
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[340\]
timestamp 1637331468
transform 1 0 12144 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[310\]
timestamp 1637331468
transform 1 0 12972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[241\]
timestamp 1637331468
transform 1 0 12696 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[193\]
timestamp 1637331468
transform 1 0 11960 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[163\]
timestamp 1637331468
transform 1 0 12420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_119
timestamp 1637331468
transform 1 0 12236 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_121
timestamp 1637331468
transform 1 0 12420 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1637331468
transform 1 0 12052 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[303\]
timestamp 1637331468
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[243\]
timestamp 1637331468
transform 1 0 13800 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[230\]
timestamp 1637331468
transform 1 0 13248 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[200\]
timestamp 1637331468
transform 1 0 13524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1637331468
transform 1 0 14168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_133 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 13524 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1637331468
transform 1 0 14260 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1637331468
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[264\]
timestamp 1637331468
transform 1 0 14904 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[255\]
timestamp 1637331468
transform 1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[247\]
timestamp 1637331468
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[188\]
timestamp 1637331468
transform 1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[182\]
timestamp 1637331468
transform 1 0 14628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1637331468
transform 1 0 15456 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_142
timestamp 1637331468
transform 1 0 14352 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[316\]
timestamp 1637331468
transform 1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[312\]
timestamp 1637331468
transform 1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[254\]
timestamp 1637331468
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1637331468
transform 1 0 16560 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1637331468
transform 1 0 16560 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[325\]
timestamp 1637331468
transform 1 0 16836 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[263\]
timestamp 1637331468
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[25\]
timestamp 1637331468
transform 1 0 17204 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[258\]
timestamp 1637331468
transform 1 0 16836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[190\]
timestamp 1637331468
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1637331468
transform 1 0 16744 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1637331468
transform 1 0 16744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1637331468
transform 1 0 17112 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_172
timestamp 1637331468
transform 1 0 17112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[339\]
timestamp 1637331468
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[270\]
timestamp 1637331468
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[267\]
timestamp 1637331468
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[165\]
timestamp 1637331468
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1637331468
transform 1 0 18216 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[278\]
timestamp 1637331468
transform 1 0 19964 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[217\]
timestamp 1637331468
transform 1 0 19412 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[176\]
timestamp 1637331468
transform 1 0 19688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1637331468
transform 1 0 19320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1637331468
transform 1 0 20056 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1637331468
transform 1 0 19136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_196 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1637331468
transform 1 0 19320 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[338\]
timestamp 1637331468
transform 1 0 20240 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[332\]
timestamp 1637331468
transform 1 0 20240 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[318\]
timestamp 1637331468
transform 1 0 20516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[285\]
timestamp 1637331468
transform 1 0 21068 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[236\]
timestamp 1637331468
transform 1 0 20792 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[192\]
timestamp 1637331468
transform 1 0 21344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_209
timestamp 1637331468
transform 1 0 20516 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1637331468
transform 1 0 21620 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1637331468
transform 1 0 21896 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1637331468
transform 1 0 21896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[244\]
timestamp 1637331468
transform 1 0 21620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1637331468
transform 1 0 21988 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_228
timestamp 1637331468
transform 1 0 22264 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[292\]
timestamp 1637331468
transform 1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[202\]
timestamp 1637331468
transform 1 0 22448 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[198\]
timestamp 1637331468
transform 1 0 21988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1637331468
transform 1 0 22448 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[29\]
timestamp 1637331468
transform 1 0 23276 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[252\]
timestamp 1637331468
transform 1 0 22724 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[213\]
timestamp 1637331468
transform 1 0 23552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[208\]
timestamp 1637331468
transform 1 0 23000 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_242
timestamp 1637331468
transform 1 0 23552 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[302\]
timestamp 1637331468
transform 1 0 23920 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[224\]
timestamp 1637331468
transform 1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[219\]
timestamp 1637331468
transform 1 0 24196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[181\]
timestamp 1637331468
transform 1 0 24564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1637331468
transform 1 0 24472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1637331468
transform 1 0 24656 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_245
timestamp 1637331468
transform 1 0 23828 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[274\]
timestamp 1637331468
transform 1 0 25024 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[235\]
timestamp 1637331468
transform 1 0 25852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[22\]
timestamp 1637331468
transform 1 0 25300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[205\]
timestamp 1637331468
transform 1 0 25576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_259
timestamp 1637331468
transform 1 0 25116 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1637331468
transform 1 0 25300 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[317\]
timestamp 1637331468
transform 1 0 26128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[240\]
timestamp 1637331468
transform 1 0 26404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1637331468
transform 1 0 26956 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1637331468
transform 1 0 26956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1637331468
transform 1 0 27048 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1637331468
transform 1 0 27048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[320\]
timestamp 1637331468
transform 1 0 26680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[246\]
timestamp 1637331468
transform 1 0 27140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1637331468
transform 1 0 27140 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1637331468
transform 1 0 26404 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[324\]
timestamp 1637331468
transform 1 0 27784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[305\]
timestamp 1637331468
transform 1 0 28336 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[257\]
timestamp 1637331468
transform 1 0 28060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[251\]
timestamp 1637331468
transform 1 0 27508 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_284
timestamp 1637331468
transform 1 0 27416 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1637331468
transform 1 0 28244 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[33\]
timestamp 1637331468
transform 1 0 29256 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[334\]
timestamp 1637331468
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[328\]
timestamp 1637331468
transform 1 0 28612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[266\]
timestamp 1637331468
transform 1 0 28888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1637331468
transform 1 0 29624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_301
timestamp 1637331468
transform 1 0 28980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1637331468
transform 1 0 29440 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_307
timestamp 1637331468
transform 1 0 29532 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[227\]
timestamp 1637331468
transform 1 0 30084 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[172\]
timestamp 1637331468
transform 1 0 30636 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[16\]
timestamp 1637331468
transform 1 0 30360 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[164\]
timestamp 1637331468
transform 1 0 29808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1637331468
transform 1 0 29716 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_319
timestamp 1637331468
transform 1 0 30636 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[296\]
timestamp 1637331468
transform 1 0 31464 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[289\]
timestamp 1637331468
transform 1 0 31464 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[279\]
timestamp 1637331468
transform 1 0 30912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[183\]
timestamp 1637331468
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[178\]
timestamp 1637331468
transform 1 0 31188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1637331468
transform 1 0 31740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_327
timestamp 1637331468
transform 1 0 31372 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1637331468
transform 1 0 32108 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1637331468
transform 1 0 32016 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1637331468
transform 1 0 32292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1637331468
transform 1 0 32200 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1637331468
transform 1 0 32200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[30\]
timestamp 1637331468
transform 1 0 32568 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[189\]
timestamp 1637331468
transform 1 0 32568 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[186\]
timestamp 1637331468
transform 1 0 32292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[286\]
timestamp 1637331468
transform 1 0 32844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[197\]
timestamp 1637331468
transform 1 0 33120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_343
timestamp 1637331468
transform 1 0 32844 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[24\]
timestamp 1637331468
transform 1 0 34224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[204\]
timestamp 1637331468
transform 1 0 33948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[201\]
timestamp 1637331468
transform 1 0 33672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[19\]
timestamp 1637331468
transform 1 0 33396 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_355
timestamp 1637331468
transform 1 0 33948 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[299\]
timestamp 1637331468
transform 1 0 34500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[218\]
timestamp 1637331468
transform 1 0 35420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[215\]
timestamp 1637331468
transform 1 0 35144 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[212\]
timestamp 1637331468
transform 1 0 34868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1637331468
transform 1 0 34776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1637331468
transform 1 0 35052 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[229\]
timestamp 1637331468
transform 1 0 36524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[226\]
timestamp 1637331468
transform 1 0 36248 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[223\]
timestamp 1637331468
transform 1 0 35972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[220\]
timestamp 1637331468
transform 1 0 35696 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1637331468
transform 1 0 36156 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[23\]
timestamp 1637331468
transform 1 0 37720 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[237\]
timestamp 1637331468
transform 1 0 37444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[234\]
timestamp 1637331468
transform 1 0 37076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[231\]
timestamp 1637331468
transform 1 0 36800 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1637331468
transform 1 0 37352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1637331468
transform 1 0 37352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1637331468
transform 1 0 37444 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1637331468
transform 1 0 37260 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[250\]
timestamp 1637331468
transform 1 0 38824 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[248\]
timestamp 1637331468
transform 1 0 38548 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[245\]
timestamp 1637331468
transform 1 0 38272 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[242\]
timestamp 1637331468
transform 1 0 37996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1637331468
transform 1 0 38548 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[259\]
timestamp 1637331468
transform 1 0 39652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[256\]
timestamp 1637331468
transform 1 0 39376 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[253\]
timestamp 1637331468
transform 1 0 39100 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[232\]
timestamp 1637331468
transform 1 0 40112 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1637331468
transform 1 0 39928 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1637331468
transform 1 0 39652 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1637331468
transform 1 0 40020 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[276\]
timestamp 1637331468
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[272\]
timestamp 1637331468
transform 1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[269\]
timestamp 1637331468
transform 1 0 40664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[261\]
timestamp 1637331468
transform 1 0 40388 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1637331468
transform 1 0 40756 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[283\]
timestamp 1637331468
transform 1 0 41768 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[27\]
timestamp 1637331468
transform 1 0 41492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1637331468
transform 1 0 42412 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1637331468
transform 1 0 42320 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1637331468
transform 1 0 42504 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1637331468
transform 1 0 42504 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[290\]
timestamp 1637331468
transform 1 0 42596 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[287\]
timestamp 1637331468
transform 1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1637331468
transform 1 0 42596 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1637331468
transform 1 0 41860 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[300\]
timestamp 1637331468
transform 1 0 43792 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[298\]
timestamp 1637331468
transform 1 0 43148 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[294\]
timestamp 1637331468
transform 1 0 42872 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[268\]
timestamp 1637331468
transform 1 0 43516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_461
timestamp 1637331468
transform 1 0 43700 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_458
timestamp 1637331468
transform 1 0 43424 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[319\]
timestamp 1637331468
transform 1 0 44344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[311\]
timestamp 1637331468
transform 1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[309\]
timestamp 1637331468
transform 1 0 44344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[304\]
timestamp 1637331468
transform 1 0 44068 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1637331468
transform 1 0 44896 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1637331468
transform 1 0 44252 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_471
timestamp 1637331468
transform 1 0 44620 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1637331468
transform 1 0 45080 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[313\]
timestamp 1637331468
transform 1 0 45172 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_479
timestamp 1637331468
transform 1 0 45356 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[333\]
timestamp 1637331468
transform 1 0 45540 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[326\]
timestamp 1637331468
transform 1 0 45448 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 1637331468
transform 1 0 45724 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_484
timestamp 1637331468
transform 1 0 45816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[315\]
timestamp 1637331468
transform 1 0 45816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[342\]
timestamp 1637331468
transform 1 0 46092 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[32\]
timestamp 1637331468
transform 1 0 46092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[322\]
timestamp 1637331468
transform 1 0 46920 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[180\]
timestamp 1637331468
transform 1 0 47196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[170\]
timestamp 1637331468
transform 1 0 46644 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[167\]
timestamp 1637331468
transform 1 0 46368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_490
timestamp 1637331468
transform 1 0 46368 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[199\]
timestamp 1637331468
transform 1 0 48300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[191\]
timestamp 1637331468
transform 1 0 48024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[187\]
timestamp 1637331468
transform 1 0 47748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1637331468
transform 1 0 47656 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1637331468
transform 1 0 47656 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1637331468
transform 1 0 47472 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1637331468
transform 1 0 47472 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1637331468
transform 1 0 47748 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[21\]
timestamp 1637331468
transform 1 0 49680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[216\]
timestamp 1637331468
transform 1 0 49404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[211\]
timestamp 1637331468
transform 1 0 49128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[207\]
timestamp 1637331468
transform 1 0 48852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[203\]
timestamp 1637331468
transform 1 0 48576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1637331468
transform 1 0 48852 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[281\]
timestamp 1637331468
transform 1 0 50876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[275\]
timestamp 1637331468
transform 1 0 50600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[265\]
timestamp 1637331468
transform 1 0 50324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[233\]
timestamp 1637331468
transform 1 0 49956 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1637331468
transform 1 0 50232 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1637331468
transform 1 0 49956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[314\]
timestamp 1637331468
transform 1 0 51980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[306\]
timestamp 1637331468
transform 1 0 51704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[301\]
timestamp 1637331468
transform 1 0 51428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[295\]
timestamp 1637331468
transform 1 0 51152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1637331468
transform 1 0 51060 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_553
timestamp 1637331468
transform 1 0 52164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1637331468
transform 1 0 52532 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[337\]
timestamp 1637331468
transform 1 0 52256 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[323\]
timestamp 1637331468
transform 1 0 52256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[173\]
timestamp 1637331468
transform 1 0 52532 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1637331468
transform 1 0 52808 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1637331468
transform 1 0 52808 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[194\]
timestamp 1637331468
transform 1 0 53176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[184\]
timestamp 1637331468
transform 1 0 52900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1637331468
transform 1 0 52900 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[249\]
timestamp 1637331468
transform 1 0 54280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[238\]
timestamp 1637331468
transform 1 0 54004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[225\]
timestamp 1637331468
transform 1 0 53728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[1\]
timestamp 1637331468
transform 1 0 53452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1637331468
transform 1 0 54004 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[341\]
timestamp 1637331468
transform 1 0 55108 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[331\]
timestamp 1637331468
transform 1 0 54832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[307\]
timestamp 1637331468
transform 1 0 54556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[20\]
timestamp 1637331468
transform 1 0 55476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1637331468
transform 1 0 55384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1637331468
transform 1 0 55108 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[308\]
timestamp 1637331468
transform 1 0 56304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[239\]
timestamp 1637331468
transform 1 0 56028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[175\]
timestamp 1637331468
transform 1 0 55752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1637331468
transform 1 0 56212 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_601
timestamp 1637331468
transform 1 0 56580 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1637331468
transform 1 0 57960 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1637331468
transform 1 0 57960 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1637331468
transform 1 0 57684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1637331468
transform 1 0 57316 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1637331468
transform 1 0 57868 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1637331468
transform 1 0 59156 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1637331468
transform 1 0 58052 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_629
timestamp 1637331468
transform 1 0 59156 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1637331468
transform 1 0 58052 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1637331468
transform 1 0 60260 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_641
timestamp 1637331468
transform 1 0 60260 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1637331468
transform 1 0 60536 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1637331468
transform 1 0 61364 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_645
timestamp 1637331468
transform 1 0 60628 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1637331468
transform 1 0 62468 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_657
timestamp 1637331468
transform 1 0 61732 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1637331468
transform 1 0 63112 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1637331468
transform 1 0 63112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1637331468
transform 1 0 62836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1637331468
transform 1 0 63204 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_673
timestamp 1637331468
transform 1 0 63204 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1637331468
transform 1 0 63020 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1637331468
transform 1 0 64308 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_685
timestamp 1637331468
transform 1 0 64308 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1637331468
transform 1 0 65688 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1637331468
transform 1 0 65412 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_697
timestamp 1637331468
transform 1 0 65412 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_701
timestamp 1637331468
transform 1 0 65780 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_709
timestamp 1637331468
transform 1 0 66516 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_713
timestamp 1637331468
transform 1 0 66884 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1637331468
transform 1 0 68264 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1637331468
transform 1 0 68264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1637331468
transform -1 0 68816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1637331468
transform -1 0 68816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1637331468
transform 1 0 67988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_729
timestamp 1637331468
transform 1 0 68356 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_729
timestamp 1637331468
transform 1 0 68356 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1637331468
transform 1 0 67620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1637331468
transform 1 0 68172 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1637331468
transform 1 0 1288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1637331468
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1637331468
transform 1 0 1564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[162\]
timestamp 1637331468
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[159\]
timestamp 1637331468
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[157\]
timestamp 1637331468
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[151\]
timestamp 1637331468
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[105\]
timestamp 1637331468
transform 1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[101\]
timestamp 1637331468
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[100\]
timestamp 1637331468
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[0\]
timestamp 1637331468
transform 1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1637331468
transform 1 0 3864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1637331468
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[154\]
timestamp 1637331468
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[150\]
timestamp 1637331468
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[14\]
timestamp 1637331468
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[102\]
timestamp 1637331468
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[330\]
timestamp 1637331468
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[145\]
timestamp 1637331468
transform 1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1637331468
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_60
timestamp 1637331468
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1637331468
transform 1 0 7912 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1637331468
transform 1 0 9016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1637331468
transform 1 0 9108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1637331468
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[125\]
timestamp 1637331468
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1637331468
transform 1 0 11316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_118
timestamp 1637331468
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1637331468
transform 1 0 14168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1637331468
transform 1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1637331468
transform 1 0 14260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1637331468
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1637331468
transform 1 0 15364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1637331468
transform 1 0 16468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1637331468
transform 1 0 17572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1637331468
transform 1 0 18676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1637331468
transform 1 0 19320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1637331468
transform 1 0 19412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1637331468
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1637331468
transform 1 0 20516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1637331468
transform 1 0 21620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1637331468
transform 1 0 22724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1637331468
transform 1 0 24472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1637331468
transform 1 0 23828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1637331468
transform 1 0 24564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1637331468
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1637331468
transform 1 0 25668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1637331468
transform 1 0 26772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1637331468
transform 1 0 27876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[389\]
timestamp 1637331468
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1637331468
transform 1 0 29624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1637331468
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1637331468
transform 1 0 29072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1637331468
transform 1 0 29716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1637331468
transform 1 0 31924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1637331468
transform 1 0 30820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1637331468
transform 1 0 33028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1637331468
transform 1 0 34132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1637331468
transform 1 0 34776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1637331468
transform 1 0 34868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1637331468
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[413\]
timestamp 1637331468
transform 1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1637331468
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_386
timestamp 1637331468
transform 1 0 36800 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1637331468
transform 1 0 37904 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1637331468
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1637331468
transform 1 0 39928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1637331468
transform 1 0 39744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1637331468
transform 1 0 40020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_433
timestamp 1637331468
transform 1 0 41124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[430\]
timestamp 1637331468
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_442
timestamp 1637331468
transform 1 0 41952 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_454
timestamp 1637331468
transform 1 0 43056 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[43\]
timestamp 1637331468
transform 1 0 44252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1637331468
transform 1 0 44528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_466
timestamp 1637331468
transform 1 0 44160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[446\]
timestamp 1637331468
transform 1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[445\]
timestamp 1637331468
transform 1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[444\]
timestamp 1637331468
transform 1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[443\]
timestamp 1637331468
transform 1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1637331468
transform 1 0 45080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_477
timestamp 1637331468
transform 1 0 45172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[44\]
timestamp 1637331468
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[449\]
timestamp 1637331468
transform 1 0 46920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[448\]
timestamp 1637331468
transform 1 0 46644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[447\]
timestamp 1637331468
transform 1 0 46368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[453\]
timestamp 1637331468
transform 1 0 48300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[452\]
timestamp 1637331468
transform 1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_502
timestamp 1637331468
transform 1 0 47472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_526
timestamp 1637331468
transform 1 0 49680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_514
timestamp 1637331468
transform 1 0 48576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1637331468
transform 1 0 50232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1637331468
transform 1 0 50324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1637331468
transform 1 0 51428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1637331468
transform 1 0 52532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1637331468
transform 1 0 53636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1637331468
transform 1 0 55384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1637331468
transform 1 0 54740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1637331468
transform 1 0 55476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1637331468
transform 1 0 55292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1637331468
transform 1 0 56580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1637331468
transform 1 0 57684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1637331468
transform 1 0 58788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1637331468
transform 1 0 59892 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1637331468
transform 1 0 60536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1637331468
transform 1 0 60628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1637331468
transform 1 0 60444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1637331468
transform 1 0 61732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1637331468
transform 1 0 62836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  insts\[90\]
timestamp 1637331468
transform 1 0 64952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_689
timestamp 1637331468
transform 1 0 64676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_681
timestamp 1637331468
transform 1 0 63940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[95\]
timestamp 1637331468
transform -1 0 66332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[94\]
timestamp 1637331468
transform -1 0 66056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[92\]
timestamp 1637331468
transform 1 0 65412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1637331468
transform 1 0 65688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_695
timestamp 1637331468
transform 1 0 65228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[97\]
timestamp 1637331468
transform -1 0 66608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_710
timestamp 1637331468
transform 1 0 66608 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1637331468
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_730
timestamp 1637331468
transform 1 0 68448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_722
timestamp 1637331468
transform 1 0 67712 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  insts\[160\]
timestamp 1637331468
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1637331468
transform 1 0 1288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1637331468
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1637331468
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[153\]
timestamp 1637331468
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[152\]
timestamp 1637331468
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[149\]
timestamp 1637331468
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[146\]
timestamp 1637331468
transform -1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[144\]
timestamp 1637331468
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[12\]
timestamp 1637331468
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[10\]
timestamp 1637331468
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[104\]
timestamp 1637331468
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1637331468
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1637331468
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[148\]
timestamp 1637331468
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[147\]
timestamp 1637331468
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[139\]
timestamp 1637331468
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[133\]
timestamp 1637331468
transform 1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_50
timestamp 1637331468
transform 1 0 5888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1637331468
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[143\]
timestamp 1637331468
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[142\]
timestamp 1637331468
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[122\]
timestamp 1637331468
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1637331468
transform 1 0 6440 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1637331468
transform 1 0 6256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[141\]
timestamp 1637331468
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[140\]
timestamp 1637331468
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[138\]
timestamp 1637331468
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[132\]
timestamp 1637331468
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[137\]
timestamp 1637331468
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[136\]
timestamp 1637331468
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[135\]
timestamp 1637331468
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[134\]
timestamp 1637331468
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1637331468
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[131\]
timestamp 1637331468
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[130\]
timestamp 1637331468
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[126\]
timestamp 1637331468
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[118\]
timestamp 1637331468
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[129\]
timestamp 1637331468
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[128\]
timestamp 1637331468
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[127\]
timestamp 1637331468
transform 1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[120\]
timestamp 1637331468
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1637331468
transform 1 0 11592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[124\]
timestamp 1637331468
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[123\]
timestamp 1637331468
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[121\]
timestamp 1637331468
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[11\]
timestamp 1637331468
transform 1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1637331468
transform 1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[119\]
timestamp 1637331468
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[117\]
timestamp 1637331468
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[115\]
timestamp 1637331468
transform 1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1637331468
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_141
timestamp 1637331468
transform 1 0 14260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_139
timestamp 1637331468
transform 1 0 14076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[344\]
timestamp 1637331468
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[15\]
timestamp 1637331468
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[13\]
timestamp 1637331468
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[116\]
timestamp 1637331468
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[114\]
timestamp 1637331468
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[347\]
timestamp 1637331468
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[346\]
timestamp 1637331468
transform 1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[345\]
timestamp 1637331468
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1637331468
transform 1 0 16560 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[350\]
timestamp 1637331468
transform 1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[34\]
timestamp 1637331468
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[349\]
timestamp 1637331468
transform 1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[348\]
timestamp 1637331468
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1637331468
transform 1 0 16744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[354\]
timestamp 1637331468
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[353\]
timestamp 1637331468
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[352\]
timestamp 1637331468
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[351\]
timestamp 1637331468
transform 1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[358\]
timestamp 1637331468
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[357\]
timestamp 1637331468
transform 1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[356\]
timestamp 1637331468
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[355\]
timestamp 1637331468
transform 1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1637331468
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[362\]
timestamp 1637331468
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[361\]
timestamp 1637331468
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[360\]
timestamp 1637331468
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[35\]
timestamp 1637331468
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[359\]
timestamp 1637331468
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[366\]
timestamp 1637331468
transform 1 0 22540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[365\]
timestamp 1637331468
transform 1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[364\]
timestamp 1637331468
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[363\]
timestamp 1637331468
transform 1 0 21620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1637331468
transform 1 0 21896 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[36\]
timestamp 1637331468
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[369\]
timestamp 1637331468
transform 1 0 23368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[368\]
timestamp 1637331468
transform 1 0 23092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[367\]
timestamp 1637331468
transform 1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[373\]
timestamp 1637331468
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[372\]
timestamp 1637331468
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[371\]
timestamp 1637331468
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[370\]
timestamp 1637331468
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1637331468
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[377\]
timestamp 1637331468
transform 1 0 25944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[376\]
timestamp 1637331468
transform 1 0 25668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[375\]
timestamp 1637331468
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[374\]
timestamp 1637331468
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[380\]
timestamp 1637331468
transform 1 0 27140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[37\]
timestamp 1637331468
transform 1 0 26772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[379\]
timestamp 1637331468
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[378\]
timestamp 1637331468
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1637331468
transform 1 0 27048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[384\]
timestamp 1637331468
transform 1 0 28244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[383\]
timestamp 1637331468
transform 1 0 27968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[382\]
timestamp 1637331468
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[381\]
timestamp 1637331468
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[388\]
timestamp 1637331468
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[387\]
timestamp 1637331468
transform 1 0 29072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[386\]
timestamp 1637331468
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[385\]
timestamp 1637331468
transform 1 0 28520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1637331468
transform 1 0 29624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[392\]
timestamp 1637331468
transform 1 0 30544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[391\]
timestamp 1637331468
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[390\]
timestamp 1637331468
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[38\]
timestamp 1637331468
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[397\]
timestamp 1637331468
transform 1 0 31924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[396\]
timestamp 1637331468
transform 1 0 31648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[395\]
timestamp 1637331468
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[394\]
timestamp 1637331468
transform 1 0 31096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[393\]
timestamp 1637331468
transform 1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[3\]
timestamp 1637331468
transform 1 0 33120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[39\]
timestamp 1637331468
transform 1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[399\]
timestamp 1637331468
transform 1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[398\]
timestamp 1637331468
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1637331468
transform 1 0 32200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[403\]
timestamp 1637331468
transform 1 0 34224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[402\]
timestamp 1637331468
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[401\]
timestamp 1637331468
transform 1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[400\]
timestamp 1637331468
transform 1 0 33396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[407\]
timestamp 1637331468
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[406\]
timestamp 1637331468
transform 1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[405\]
timestamp 1637331468
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[404\]
timestamp 1637331468
transform 1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1637331468
transform 1 0 34776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[410\]
timestamp 1637331468
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[40\]
timestamp 1637331468
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[409\]
timestamp 1637331468
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[408\]
timestamp 1637331468
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[415\]
timestamp 1637331468
transform 1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[414\]
timestamp 1637331468
transform 1 0 37444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[412\]
timestamp 1637331468
transform 1 0 37076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[411\]
timestamp 1637331468
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1637331468
transform 1 0 37352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[419\]
timestamp 1637331468
transform 1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[418\]
timestamp 1637331468
transform 1 0 38548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[417\]
timestamp 1637331468
transform 1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[416\]
timestamp 1637331468
transform 1 0 37996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[422\]
timestamp 1637331468
transform 1 0 40020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[421\]
timestamp 1637331468
transform 1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[420\]
timestamp 1637331468
transform 1 0 39376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[41\]
timestamp 1637331468
transform 1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1637331468
transform 1 0 39928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[427\]
timestamp 1637331468
transform 1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[426\]
timestamp 1637331468
transform 1 0 41124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[425\]
timestamp 1637331468
transform 1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[424\]
timestamp 1637331468
transform 1 0 40572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[423\]
timestamp 1637331468
transform 1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[431\]
timestamp 1637331468
transform 1 0 42596 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[42\]
timestamp 1637331468
transform 1 0 42228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[429\]
timestamp 1637331468
transform 1 0 41952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[428\]
timestamp 1637331468
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1637331468
transform 1 0 42504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[435\]
timestamp 1637331468
transform 1 0 43700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[434\]
timestamp 1637331468
transform 1 0 43424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[433\]
timestamp 1637331468
transform 1 0 43148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[432\]
timestamp 1637331468
transform 1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[439\]
timestamp 1637331468
transform 1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[438\]
timestamp 1637331468
transform 1 0 44528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[437\]
timestamp 1637331468
transform 1 0 44252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[436\]
timestamp 1637331468
transform 1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[442\]
timestamp 1637331468
transform 1 0 45724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[441\]
timestamp 1637331468
transform 1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[440\]
timestamp 1637331468
transform 1 0 45172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1637331468
transform 1 0 45080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_486
timestamp 1637331468
transform 1 0 46000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_498
timestamp 1637331468
transform 1 0 47104 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  insts\[451\]
timestamp 1637331468
transform 1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[450\]
timestamp 1637331468
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1637331468
transform 1 0 47656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_511
timestamp 1637331468
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  insts\[457\]
timestamp 1637331468
transform 1 0 49496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[456\]
timestamp 1637331468
transform 1 0 49220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[455\]
timestamp 1637331468
transform 1 0 48944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[454\]
timestamp 1637331468
transform 1 0 48668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[460\]
timestamp 1637331468
transform 1 0 50876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[45\]
timestamp 1637331468
transform 1 0 50600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[459\]
timestamp 1637331468
transform 1 0 50324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[458\]
timestamp 1637331468
transform 1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1637331468
transform 1 0 50232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_530
timestamp 1637331468
transform 1 0 50048 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  insts\[47\]
timestamp 1637331468
transform 1 0 51980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[46\]
timestamp 1637331468
transform 1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[462\]
timestamp 1637331468
transform 1 0 51428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[461\]
timestamp 1637331468
transform 1 0 51152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[50\]
timestamp 1637331468
transform 1 0 53176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[4\]
timestamp 1637331468
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[49\]
timestamp 1637331468
transform 1 0 52532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[48\]
timestamp 1637331468
transform 1 0 52256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1637331468
transform 1 0 52808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[54\]
timestamp 1637331468
transform 1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[53\]
timestamp 1637331468
transform 1 0 54004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[52\]
timestamp 1637331468
transform 1 0 53728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[51\]
timestamp 1637331468
transform 1 0 53452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[58\]
timestamp 1637331468
transform 1 0 55476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[57\]
timestamp 1637331468
transform 1 0 55108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[56\]
timestamp 1637331468
transform 1 0 54832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[55\]
timestamp 1637331468
transform 1 0 54556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1637331468
transform 1 0 55384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[61\]
timestamp 1637331468
transform 1 0 56580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[60\]
timestamp 1637331468
transform 1 0 56304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[5\]
timestamp 1637331468
transform 1 0 56028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[59\]
timestamp 1637331468
transform 1 0 55752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[65\]
timestamp 1637331468
transform 1 0 57684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[64\]
timestamp 1637331468
transform 1 0 57408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[63\]
timestamp 1637331468
transform 1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[62\]
timestamp 1637331468
transform 1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1637331468
transform 1 0 57960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[6\]
timestamp 1637331468
transform 1 0 59156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[69\]
timestamp 1637331468
transform 1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[68\]
timestamp 1637331468
transform 1 0 58604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[67\]
timestamp 1637331468
transform 1 0 58328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[66\]
timestamp 1637331468
transform 1 0 58052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[73\]
timestamp 1637331468
transform 1 0 60260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[72\]
timestamp 1637331468
transform 1 0 59984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[71\]
timestamp 1637331468
transform 1 0 59708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[70\]
timestamp 1637331468
transform 1 0 59432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[77\]
timestamp 1637331468
transform 1 0 61456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[76\]
timestamp 1637331468
transform 1 0 61180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[75\]
timestamp 1637331468
transform 1 0 60904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[74\]
timestamp 1637331468
transform 1 0 60628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1637331468
transform 1 0 60536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[80\]
timestamp 1637331468
transform 1 0 62560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[7\]
timestamp 1637331468
transform 1 0 62284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[79\]
timestamp 1637331468
transform 1 0 62008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[78\]
timestamp 1637331468
transform 1 0 61732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[84\]
timestamp 1637331468
transform 1 0 63756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[83\]
timestamp 1637331468
transform 1 0 63480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[82\]
timestamp 1637331468
transform 1 0 63204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[81\]
timestamp 1637331468
transform 1 0 62836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1637331468
transform 1 0 63112 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[88\]
timestamp 1637331468
transform 1 0 64860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[87\]
timestamp 1637331468
transform 1 0 64584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[86\]
timestamp 1637331468
transform 1 0 64308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[85\]
timestamp 1637331468
transform 1 0 64032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[91\]
timestamp 1637331468
transform 1 0 66056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[8\]
timestamp 1637331468
transform 1 0 65412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[89\]
timestamp 1637331468
transform 1 0 65136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[343\]
timestamp 1637331468
transform -1 0 66056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1637331468
transform 1 0 65688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  insts\[99\]
timestamp 1637331468
transform -1 0 67436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[98\]
timestamp 1637331468
transform -1 0 67160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[96\]
timestamp 1637331468
transform 1 0 66608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[93\]
timestamp 1637331468
transform 1 0 66332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  insts\[9\]
timestamp 1637331468
transform -1 0 67712 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1637331468
transform 1 0 68264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1637331468
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_729
timestamp 1637331468
transform 1 0 68356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_722
timestamp 1637331468
transform 1 0 67712 0 -1 3264
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 3816 600 3936 6 HI[0]
port 0 nsew signal tristate
rlabel metal3 s 0 3544 600 3664 6 HI[100]
port 1 nsew signal tristate
rlabel metal3 s 0 3272 600 3392 6 HI[101]
port 2 nsew signal tristate
rlabel metal3 s 0 3000 600 3120 6 HI[102]
port 3 nsew signal tristate
rlabel metal3 s 0 2728 600 2848 6 HI[103]
port 4 nsew signal tristate
rlabel metal3 s 0 2456 600 2576 6 HI[104]
port 5 nsew signal tristate
rlabel metal3 s 0 2184 600 2304 6 HI[105]
port 6 nsew signal tristate
rlabel metal3 s 0 1912 600 2032 6 HI[106]
port 7 nsew signal tristate
rlabel metal3 s 0 1640 600 1760 6 HI[107]
port 8 nsew signal tristate
rlabel metal3 s 0 1368 600 1488 6 HI[108]
port 9 nsew signal tristate
rlabel metal3 s 0 1096 600 1216 6 HI[109]
port 10 nsew signal tristate
rlabel metal3 s 0 4088 600 4208 6 HI[10]
port 11 nsew signal tristate
rlabel metal3 s 0 824 600 944 6 HI[110]
port 12 nsew signal tristate
rlabel metal3 s 0 280 600 400 6 HI[111]
port 13 nsew signal tristate
rlabel metal3 s 0 8 600 128 6 HI[112]
port 14 nsew signal tristate
rlabel metal3 s 0 552 600 672 6 HI[113]
port 15 nsew signal tristate
rlabel metal2 s 14094 3800 14150 4400 6 HI[114]
port 16 nsew signal tristate
rlabel metal2 s 12990 3800 13046 4400 6 HI[115]
port 17 nsew signal tristate
rlabel metal2 s 13818 3800 13874 4400 6 HI[116]
port 18 nsew signal tristate
rlabel metal2 s 13542 3800 13598 4400 6 HI[117]
port 19 nsew signal tristate
rlabel metal2 s 9402 3800 9458 4400 6 HI[118]
port 20 nsew signal tristate
rlabel metal2 s 13266 3800 13322 4400 6 HI[119]
port 21 nsew signal tristate
rlabel metal2 s 12438 3800 12494 4400 6 HI[11]
port 22 nsew signal tristate
rlabel metal2 s 11334 3800 11390 4400 6 HI[120]
port 23 nsew signal tristate
rlabel metal2 s 12714 3800 12770 4400 6 HI[121]
port 24 nsew signal tristate
rlabel metal2 s 6366 3800 6422 4400 6 HI[122]
port 25 nsew signal tristate
rlabel metal2 s 12162 3800 12218 4400 6 HI[123]
port 26 nsew signal tristate
rlabel metal2 s 11886 3800 11942 4400 6 HI[124]
port 27 nsew signal tristate
rlabel metal2 s 11610 3800 11666 4400 6 HI[125]
port 28 nsew signal tristate
rlabel metal2 s 9678 3800 9734 4400 6 HI[126]
port 29 nsew signal tristate
rlabel metal2 s 11058 3800 11114 4400 6 HI[127]
port 30 nsew signal tristate
rlabel metal2 s 10782 3800 10838 4400 6 HI[128]
port 31 nsew signal tristate
rlabel metal2 s 10506 3800 10562 4400 6 HI[129]
port 32 nsew signal tristate
rlabel metal2 s 570 3800 626 4400 6 HI[12]
port 33 nsew signal tristate
rlabel metal2 s 10230 3800 10286 4400 6 HI[130]
port 34 nsew signal tristate
rlabel metal2 s 9954 3800 10010 4400 6 HI[131]
port 35 nsew signal tristate
rlabel metal2 s 7746 3800 7802 4400 6 HI[132]
port 36 nsew signal tristate
rlabel metal2 s 4986 3800 5042 4400 6 HI[133]
port 37 nsew signal tristate
rlabel metal2 s 9126 3800 9182 4400 6 HI[134]
port 38 nsew signal tristate
rlabel metal2 s 8850 3800 8906 4400 6 HI[135]
port 39 nsew signal tristate
rlabel metal2 s 8574 3800 8630 4400 6 HI[136]
port 40 nsew signal tristate
rlabel metal2 s 8298 3800 8354 4400 6 HI[137]
port 41 nsew signal tristate
rlabel metal2 s 8022 3800 8078 4400 6 HI[138]
port 42 nsew signal tristate
rlabel metal2 s 5814 3800 5870 4400 6 HI[139]
port 43 nsew signal tristate
rlabel metal2 s 14370 3800 14426 4400 6 HI[13]
port 44 nsew signal tristate
rlabel metal2 s 7470 3800 7526 4400 6 HI[140]
port 45 nsew signal tristate
rlabel metal2 s 7194 3800 7250 4400 6 HI[141]
port 46 nsew signal tristate
rlabel metal2 s 6918 3800 6974 4400 6 HI[142]
port 47 nsew signal tristate
rlabel metal2 s 6642 3800 6698 4400 6 HI[143]
port 48 nsew signal tristate
rlabel metal2 s 18 3800 74 4400 6 HI[144]
port 49 nsew signal tristate
rlabel metal2 s 6090 3800 6146 4400 6 HI[145]
port 50 nsew signal tristate
rlabel metal2 s 3606 3800 3662 4400 6 HI[146]
port 51 nsew signal tristate
rlabel metal2 s 5538 3800 5594 4400 6 HI[147]
port 52 nsew signal tristate
rlabel metal2 s 5262 3800 5318 4400 6 HI[148]
port 53 nsew signal tristate
rlabel metal2 s 294 3800 350 4400 6 HI[149]
port 54 nsew signal tristate
rlabel metal2 s 4434 3800 4490 4400 6 HI[14]
port 55 nsew signal tristate
rlabel metal2 s 4710 3800 4766 4400 6 HI[150]
port 56 nsew signal tristate
rlabel metal2 s 3882 3800 3938 4400 6 HI[151]
port 57 nsew signal tristate
rlabel metal2 s 4158 3800 4214 4400 6 HI[152]
port 58 nsew signal tristate
rlabel metal2 s 3330 3800 3386 4400 6 HI[153]
port 59 nsew signal tristate
rlabel metal2 s 1122 3800 1178 4400 6 HI[154]
port 60 nsew signal tristate
rlabel metal2 s 3054 3800 3110 4400 6 HI[155]
port 61 nsew signal tristate
rlabel metal2 s 2778 3800 2834 4400 6 HI[156]
port 62 nsew signal tristate
rlabel metal2 s 2502 3800 2558 4400 6 HI[157]
port 63 nsew signal tristate
rlabel metal2 s 2226 3800 2282 4400 6 HI[158]
port 64 nsew signal tristate
rlabel metal2 s 1950 3800 2006 4400 6 HI[159]
port 65 nsew signal tristate
rlabel metal2 s 14646 3800 14702 4400 6 HI[15]
port 66 nsew signal tristate
rlabel metal2 s 1398 3800 1454 4400 6 HI[160]
port 67 nsew signal tristate
rlabel metal2 s 1674 3800 1730 4400 6 HI[161]
port 68 nsew signal tristate
rlabel metal2 s 846 3800 902 4400 6 HI[162]
port 69 nsew signal tristate
rlabel metal2 s 11886 0 11942 600 6 HI[163]
port 70 nsew signal tristate
rlabel metal2 s 28998 0 29054 600 6 HI[164]
port 71 nsew signal tristate
rlabel metal2 s 17958 0 18014 600 6 HI[165]
port 72 nsew signal tristate
rlabel metal2 s 11058 0 11114 600 6 HI[166]
port 73 nsew signal tristate
rlabel metal2 s 45282 0 45338 600 6 HI[167]
port 74 nsew signal tristate
rlabel metal2 s 7746 0 7802 600 6 HI[168]
port 75 nsew signal tristate
rlabel metal2 s 8574 0 8630 600 6 HI[169]
port 76 nsew signal tristate
rlabel metal2 s 29550 0 29606 600 6 HI[16]
port 77 nsew signal tristate
rlabel metal2 s 45558 0 45614 600 6 HI[170]
port 78 nsew signal tristate
rlabel metal2 s 10782 0 10838 600 6 HI[171]
port 79 nsew signal tristate
rlabel metal2 s 29826 0 29882 600 6 HI[172]
port 80 nsew signal tristate
rlabel metal2 s 51354 0 51410 600 6 HI[173]
port 81 nsew signal tristate
rlabel metal2 s 10230 0 10286 600 6 HI[174]
port 82 nsew signal tristate
rlabel metal2 s 54666 0 54722 600 6 HI[175]
port 83 nsew signal tristate
rlabel metal2 s 19062 0 19118 600 6 HI[176]
port 84 nsew signal tristate
rlabel metal2 s 6366 0 6422 600 6 HI[177]
port 85 nsew signal tristate
rlabel metal2 s 30378 0 30434 600 6 HI[178]
port 86 nsew signal tristate
rlabel metal2 s 8298 0 8354 600 6 HI[179]
port 87 nsew signal tristate
rlabel metal2 s 294 0 350 600 6 HI[17]
port 88 nsew signal tristate
rlabel metal2 s 46110 0 46166 600 6 HI[180]
port 89 nsew signal tristate
rlabel metal2 s 23754 0 23810 600 6 HI[181]
port 90 nsew signal tristate
rlabel metal2 s 14094 0 14150 600 6 HI[182]
port 91 nsew signal tristate
rlabel metal2 s 30930 0 30986 600 6 HI[183]
port 92 nsew signal tristate
rlabel metal2 s 51630 0 51686 600 6 HI[184]
port 93 nsew signal tristate
rlabel metal2 s 6090 0 6146 600 6 HI[185]
port 94 nsew signal tristate
rlabel metal2 s 31206 0 31262 600 6 HI[186]
port 95 nsew signal tristate
rlabel metal2 s 46386 0 46442 600 6 HI[187]
port 96 nsew signal tristate
rlabel metal2 s 13818 0 13874 600 6 HI[188]
port 97 nsew signal tristate
rlabel metal2 s 31482 0 31538 600 6 HI[189]
port 98 nsew signal tristate
rlabel metal2 s 2778 0 2834 600 6 HI[18]
port 99 nsew signal tristate
rlabel metal2 s 16854 0 16910 600 6 HI[190]
port 100 nsew signal tristate
rlabel metal2 s 46662 0 46718 600 6 HI[191]
port 101 nsew signal tristate
rlabel metal2 s 20718 0 20774 600 6 HI[192]
port 102 nsew signal tristate
rlabel metal2 s 11334 0 11390 600 6 HI[193]
port 103 nsew signal tristate
rlabel metal2 s 51906 0 51962 600 6 HI[194]
port 104 nsew signal tristate
rlabel metal2 s 8850 0 8906 600 6 HI[195]
port 105 nsew signal tristate
rlabel metal2 s 9126 0 9182 600 6 HI[196]
port 106 nsew signal tristate
rlabel metal2 s 32310 0 32366 600 6 HI[197]
port 107 nsew signal tristate
rlabel metal2 s 21270 0 21326 600 6 HI[198]
port 108 nsew signal tristate
rlabel metal2 s 46938 0 46994 600 6 HI[199]
port 109 nsew signal tristate
rlabel metal2 s 32586 0 32642 600 6 HI[19]
port 110 nsew signal tristate
rlabel metal2 s 52182 0 52238 600 6 HI[1]
port 111 nsew signal tristate
rlabel metal2 s 12990 0 13046 600 6 HI[200]
port 112 nsew signal tristate
rlabel metal2 s 32862 0 32918 600 6 HI[201]
port 113 nsew signal tristate
rlabel metal2 s 21822 0 21878 600 6 HI[202]
port 114 nsew signal tristate
rlabel metal2 s 47214 0 47270 600 6 HI[203]
port 115 nsew signal tristate
rlabel metal2 s 33138 0 33194 600 6 HI[204]
port 116 nsew signal tristate
rlabel metal2 s 24858 0 24914 600 6 HI[205]
port 117 nsew signal tristate
rlabel metal2 s 4986 0 5042 600 6 HI[206]
port 118 nsew signal tristate
rlabel metal2 s 47490 0 47546 600 6 HI[207]
port 119 nsew signal tristate
rlabel metal2 s 22374 0 22430 600 6 HI[208]
port 120 nsew signal tristate
rlabel metal2 s 846 0 902 600 6 HI[209]
port 121 nsew signal tristate
rlabel metal2 s 54114 0 54170 600 6 HI[20]
port 122 nsew signal tristate
rlabel metal2 s 2226 0 2282 600 6 HI[210]
port 123 nsew signal tristate
rlabel metal2 s 47766 0 47822 600 6 HI[211]
port 124 nsew signal tristate
rlabel metal2 s 33966 0 34022 600 6 HI[212]
port 125 nsew signal tristate
rlabel metal2 s 22926 0 22982 600 6 HI[213]
port 126 nsew signal tristate
rlabel metal2 s 4434 0 4490 600 6 HI[214]
port 127 nsew signal tristate
rlabel metal2 s 34242 0 34298 600 6 HI[215]
port 128 nsew signal tristate
rlabel metal2 s 48042 0 48098 600 6 HI[216]
port 129 nsew signal tristate
rlabel metal2 s 18510 0 18566 600 6 HI[217]
port 130 nsew signal tristate
rlabel metal2 s 34518 0 34574 600 6 HI[218]
port 131 nsew signal tristate
rlabel metal2 s 23478 0 23534 600 6 HI[219]
port 132 nsew signal tristate
rlabel metal2 s 48318 0 48374 600 6 HI[21]
port 133 nsew signal tristate
rlabel metal2 s 34794 0 34850 600 6 HI[220]
port 134 nsew signal tristate
rlabel metal2 s 7470 0 7526 600 6 HI[221]
port 135 nsew signal tristate
rlabel metal2 s 5538 0 5594 600 6 HI[222]
port 136 nsew signal tristate
rlabel metal2 s 35070 0 35126 600 6 HI[223]
port 137 nsew signal tristate
rlabel metal2 s 24030 0 24086 600 6 HI[224]
port 138 nsew signal tristate
rlabel metal2 s 52458 0 52514 600 6 HI[225]
port 139 nsew signal tristate
rlabel metal2 s 35346 0 35402 600 6 HI[226]
port 140 nsew signal tristate
rlabel metal2 s 28722 0 28778 600 6 HI[227]
port 141 nsew signal tristate
rlabel metal2 s 18 0 74 600 6 HI[228]
port 142 nsew signal tristate
rlabel metal2 s 35622 0 35678 600 6 HI[229]
port 143 nsew signal tristate
rlabel metal2 s 24582 0 24638 600 6 HI[22]
port 144 nsew signal tristate
rlabel metal2 s 12714 0 12770 600 6 HI[230]
port 145 nsew signal tristate
rlabel metal2 s 35898 0 35954 600 6 HI[231]
port 146 nsew signal tristate
rlabel metal2 s 39210 0 39266 600 6 HI[232]
port 147 nsew signal tristate
rlabel metal2 s 48594 0 48650 600 6 HI[233]
port 148 nsew signal tristate
rlabel metal2 s 36174 0 36230 600 6 HI[234]
port 149 nsew signal tristate
rlabel metal2 s 25134 0 25190 600 6 HI[235]
port 150 nsew signal tristate
rlabel metal2 s 20166 0 20222 600 6 HI[236]
port 151 nsew signal tristate
rlabel metal2 s 36450 0 36506 600 6 HI[237]
port 152 nsew signal tristate
rlabel metal2 s 52734 0 52790 600 6 HI[238]
port 153 nsew signal tristate
rlabel metal2 s 54942 0 54998 600 6 HI[239]
port 154 nsew signal tristate
rlabel metal2 s 36726 0 36782 600 6 HI[23]
port 155 nsew signal tristate
rlabel metal2 s 25686 0 25742 600 6 HI[240]
port 156 nsew signal tristate
rlabel metal2 s 12162 0 12218 600 6 HI[241]
port 157 nsew signal tristate
rlabel metal2 s 37002 0 37058 600 6 HI[242]
port 158 nsew signal tristate
rlabel metal2 s 13266 0 13322 600 6 HI[243]
port 159 nsew signal tristate
rlabel metal2 s 20994 0 21050 600 6 HI[244]
port 160 nsew signal tristate
rlabel metal2 s 37278 0 37334 600 6 HI[245]
port 161 nsew signal tristate
rlabel metal2 s 26238 0 26294 600 6 HI[246]
port 162 nsew signal tristate
rlabel metal2 s 14646 0 14702 600 6 HI[247]
port 163 nsew signal tristate
rlabel metal2 s 37554 0 37610 600 6 HI[248]
port 164 nsew signal tristate
rlabel metal2 s 53010 0 53066 600 6 HI[249]
port 165 nsew signal tristate
rlabel metal2 s 33414 0 33470 600 6 HI[24]
port 166 nsew signal tristate
rlabel metal2 s 37830 0 37886 600 6 HI[250]
port 167 nsew signal tristate
rlabel metal2 s 26790 0 26846 600 6 HI[251]
port 168 nsew signal tristate
rlabel metal2 s 22098 0 22154 600 6 HI[252]
port 169 nsew signal tristate
rlabel metal2 s 38106 0 38162 600 6 HI[253]
port 170 nsew signal tristate
rlabel metal2 s 15750 0 15806 600 6 HI[254]
port 171 nsew signal tristate
rlabel metal2 s 14922 0 14978 600 6 HI[255]
port 172 nsew signal tristate
rlabel metal2 s 38382 0 38438 600 6 HI[256]
port 173 nsew signal tristate
rlabel metal2 s 27342 0 27398 600 6 HI[257]
port 174 nsew signal tristate
rlabel metal2 s 16302 0 16358 600 6 HI[258]
port 175 nsew signal tristate
rlabel metal2 s 38658 0 38714 600 6 HI[259]
port 176 nsew signal tristate
rlabel metal2 s 16578 0 16634 600 6 HI[25]
port 177 nsew signal tristate
rlabel metal2 s 1950 0 2006 600 6 HI[260]
port 178 nsew signal tristate
rlabel metal2 s 38934 0 38990 600 6 HI[261]
port 179 nsew signal tristate
rlabel metal2 s 1674 0 1730 600 6 HI[262]
port 180 nsew signal tristate
rlabel metal2 s 17130 0 17186 600 6 HI[263]
port 181 nsew signal tristate
rlabel metal2 s 14370 0 14426 600 6 HI[264]
port 182 nsew signal tristate
rlabel metal2 s 48870 0 48926 600 6 HI[265]
port 183 nsew signal tristate
rlabel metal2 s 28170 0 28226 600 6 HI[266]
port 184 nsew signal tristate
rlabel metal2 s 17682 0 17738 600 6 HI[267]
port 185 nsew signal tristate
rlabel metal2 s 42522 0 42578 600 6 HI[268]
port 186 nsew signal tristate
rlabel metal2 s 39486 0 39542 600 6 HI[269]
port 187 nsew signal tristate
rlabel metal2 s 6642 0 6698 600 6 HI[26]
port 188 nsew signal tristate
rlabel metal2 s 18234 0 18290 600 6 HI[270]
port 189 nsew signal tristate
rlabel metal2 s 7194 0 7250 600 6 HI[271]
port 190 nsew signal tristate
rlabel metal2 s 39762 0 39818 600 6 HI[272]
port 191 nsew signal tristate
rlabel metal2 s 10506 0 10562 600 6 HI[273]
port 192 nsew signal tristate
rlabel metal2 s 24306 0 24362 600 6 HI[274]
port 193 nsew signal tristate
rlabel metal2 s 49146 0 49202 600 6 HI[275]
port 194 nsew signal tristate
rlabel metal2 s 40038 0 40094 600 6 HI[276]
port 195 nsew signal tristate
rlabel metal2 s 5262 0 5318 600 6 HI[277]
port 196 nsew signal tristate
rlabel metal2 s 19338 0 19394 600 6 HI[278]
port 197 nsew signal tristate
rlabel metal2 s 29274 0 29330 600 6 HI[279]
port 198 nsew signal tristate
rlabel metal2 s 40314 0 40370 600 6 HI[27]
port 199 nsew signal tristate
rlabel metal2 s 3054 0 3110 600 6 HI[280]
port 200 nsew signal tristate
rlabel metal2 s 49422 0 49478 600 6 HI[281]
port 201 nsew signal tristate
rlabel metal2 s 6918 0 6974 600 6 HI[282]
port 202 nsew signal tristate
rlabel metal2 s 40590 0 40646 600 6 HI[283]
port 203 nsew signal tristate
rlabel metal2 s 1398 0 1454 600 6 HI[284]
port 204 nsew signal tristate
rlabel metal2 s 20442 0 20498 600 6 HI[285]
port 205 nsew signal tristate
rlabel metal2 s 32034 0 32090 600 6 HI[286]
port 206 nsew signal tristate
rlabel metal2 s 40866 0 40922 600 6 HI[287]
port 207 nsew signal tristate
rlabel metal2 s 3330 0 3386 600 6 HI[288]
port 208 nsew signal tristate
rlabel metal2 s 30102 0 30158 600 6 HI[289]
port 209 nsew signal tristate
rlabel metal2 s 3882 0 3938 600 6 HI[28]
port 210 nsew signal tristate
rlabel metal2 s 41142 0 41198 600 6 HI[290]
port 211 nsew signal tristate
rlabel metal2 s 4710 0 4766 600 6 HI[291]
port 212 nsew signal tristate
rlabel metal2 s 21546 0 21602 600 6 HI[292]
port 213 nsew signal tristate
rlabel metal2 s 9678 0 9734 600 6 HI[293]
port 214 nsew signal tristate
rlabel metal2 s 41418 0 41474 600 6 HI[294]
port 215 nsew signal tristate
rlabel metal2 s 49698 0 49754 600 6 HI[295]
port 216 nsew signal tristate
rlabel metal2 s 30654 0 30710 600 6 HI[296]
port 217 nsew signal tristate
rlabel metal2 s 2502 0 2558 600 6 HI[297]
port 218 nsew signal tristate
rlabel metal2 s 41694 0 41750 600 6 HI[298]
port 219 nsew signal tristate
rlabel metal2 s 33690 0 33746 600 6 HI[299]
port 220 nsew signal tristate
rlabel metal2 s 22650 0 22706 600 6 HI[29]
port 221 nsew signal tristate
rlabel metal2 s 4158 0 4214 600 6 HI[2]
port 222 nsew signal tristate
rlabel metal2 s 41970 0 42026 600 6 HI[300]
port 223 nsew signal tristate
rlabel metal2 s 49974 0 50030 600 6 HI[301]
port 224 nsew signal tristate
rlabel metal2 s 23202 0 23258 600 6 HI[302]
port 225 nsew signal tristate
rlabel metal2 s 13542 0 13598 600 6 HI[303]
port 226 nsew signal tristate
rlabel metal2 s 42246 0 42302 600 6 HI[304]
port 227 nsew signal tristate
rlabel metal2 s 27618 0 27674 600 6 HI[305]
port 228 nsew signal tristate
rlabel metal2 s 50250 0 50306 600 6 HI[306]
port 229 nsew signal tristate
rlabel metal2 s 53286 0 53342 600 6 HI[307]
port 230 nsew signal tristate
rlabel metal2 s 54390 0 54446 600 6 HI[308]
port 231 nsew signal tristate
rlabel metal2 s 43074 0 43130 600 6 HI[309]
port 232 nsew signal tristate
rlabel metal2 s 31758 0 31814 600 6 HI[30]
port 233 nsew signal tristate
rlabel metal2 s 12438 0 12494 600 6 HI[310]
port 234 nsew signal tristate
rlabel metal2 s 42798 0 42854 600 6 HI[311]
port 235 nsew signal tristate
rlabel metal2 s 15198 0 15254 600 6 HI[312]
port 236 nsew signal tristate
rlabel metal2 s 43626 0 43682 600 6 HI[313]
port 237 nsew signal tristate
rlabel metal2 s 50526 0 50582 600 6 HI[314]
port 238 nsew signal tristate
rlabel metal2 s 44730 0 44786 600 6 HI[315]
port 239 nsew signal tristate
rlabel metal2 s 15474 0 15530 600 6 HI[316]
port 240 nsew signal tristate
rlabel metal2 s 25410 0 25466 600 6 HI[317]
port 241 nsew signal tristate
rlabel metal2 s 19890 0 19946 600 6 HI[318]
port 242 nsew signal tristate
rlabel metal2 s 43350 0 43406 600 6 HI[319]
port 243 nsew signal tristate
rlabel metal2 s 570 0 626 600 6 HI[31]
port 244 nsew signal tristate
rlabel metal2 s 25962 0 26018 600 6 HI[320]
port 245 nsew signal tristate
rlabel metal2 s 1122 0 1178 600 6 HI[321]
port 246 nsew signal tristate
rlabel metal2 s 45834 0 45890 600 6 HI[322]
port 247 nsew signal tristate
rlabel metal2 s 50802 0 50858 600 6 HI[323]
port 248 nsew signal tristate
rlabel metal2 s 26514 0 26570 600 6 HI[324]
port 249 nsew signal tristate
rlabel metal2 s 16026 0 16082 600 6 HI[325]
port 250 nsew signal tristate
rlabel metal2 s 43902 0 43958 600 6 HI[326]
port 251 nsew signal tristate
rlabel metal2 s 3606 0 3662 600 6 HI[327]
port 252 nsew signal tristate
rlabel metal2 s 27066 0 27122 600 6 HI[328]
port 253 nsew signal tristate
rlabel metal2 s 8022 0 8078 600 6 HI[329]
port 254 nsew signal tristate
rlabel metal2 s 44178 0 44234 600 6 HI[32]
port 255 nsew signal tristate
rlabel metal2 s 5814 0 5870 600 6 HI[330]
port 256 nsew signal tristate
rlabel metal2 s 53562 0 53618 600 6 HI[331]
port 257 nsew signal tristate
rlabel metal2 s 18786 0 18842 600 6 HI[332]
port 258 nsew signal tristate
rlabel metal2 s 44454 0 44510 600 6 HI[333]
port 259 nsew signal tristate
rlabel metal2 s 27894 0 27950 600 6 HI[334]
port 260 nsew signal tristate
rlabel metal2 s 9954 0 10010 600 6 HI[335]
port 261 nsew signal tristate
rlabel metal2 s 9402 0 9458 600 6 HI[336]
port 262 nsew signal tristate
rlabel metal2 s 51078 0 51134 600 6 HI[337]
port 263 nsew signal tristate
rlabel metal2 s 19614 0 19670 600 6 HI[338]
port 264 nsew signal tristate
rlabel metal2 s 17406 0 17462 600 6 HI[339]
port 265 nsew signal tristate
rlabel metal2 s 28446 0 28502 600 6 HI[33]
port 266 nsew signal tristate
rlabel metal2 s 11610 0 11666 600 6 HI[340]
port 267 nsew signal tristate
rlabel metal2 s 53838 0 53894 600 6 HI[341]
port 268 nsew signal tristate
rlabel metal2 s 45006 0 45062 600 6 HI[342]
port 269 nsew signal tristate
rlabel metal2 s 67914 3800 67970 4400 6 HI[343]
port 270 nsew signal tristate
rlabel metal2 s 14922 3800 14978 4400 6 HI[344]
port 271 nsew signal tristate
rlabel metal2 s 15198 3800 15254 4400 6 HI[345]
port 272 nsew signal tristate
rlabel metal2 s 15474 3800 15530 4400 6 HI[346]
port 273 nsew signal tristate
rlabel metal2 s 15750 3800 15806 4400 6 HI[347]
port 274 nsew signal tristate
rlabel metal2 s 16026 3800 16082 4400 6 HI[348]
port 275 nsew signal tristate
rlabel metal2 s 16302 3800 16358 4400 6 HI[349]
port 276 nsew signal tristate
rlabel metal2 s 16578 3800 16634 4400 6 HI[34]
port 277 nsew signal tristate
rlabel metal2 s 16854 3800 16910 4400 6 HI[350]
port 278 nsew signal tristate
rlabel metal2 s 17130 3800 17186 4400 6 HI[351]
port 279 nsew signal tristate
rlabel metal2 s 17406 3800 17462 4400 6 HI[352]
port 280 nsew signal tristate
rlabel metal2 s 17682 3800 17738 4400 6 HI[353]
port 281 nsew signal tristate
rlabel metal2 s 17958 3800 18014 4400 6 HI[354]
port 282 nsew signal tristate
rlabel metal2 s 18234 3800 18290 4400 6 HI[355]
port 283 nsew signal tristate
rlabel metal2 s 18510 3800 18566 4400 6 HI[356]
port 284 nsew signal tristate
rlabel metal2 s 18786 3800 18842 4400 6 HI[357]
port 285 nsew signal tristate
rlabel metal2 s 19062 3800 19118 4400 6 HI[358]
port 286 nsew signal tristate
rlabel metal2 s 19338 3800 19394 4400 6 HI[359]
port 287 nsew signal tristate
rlabel metal2 s 19614 3800 19670 4400 6 HI[35]
port 288 nsew signal tristate
rlabel metal2 s 19890 3800 19946 4400 6 HI[360]
port 289 nsew signal tristate
rlabel metal2 s 20166 3800 20222 4400 6 HI[361]
port 290 nsew signal tristate
rlabel metal2 s 20442 3800 20498 4400 6 HI[362]
port 291 nsew signal tristate
rlabel metal2 s 20718 3800 20774 4400 6 HI[363]
port 292 nsew signal tristate
rlabel metal2 s 20994 3800 21050 4400 6 HI[364]
port 293 nsew signal tristate
rlabel metal2 s 21270 3800 21326 4400 6 HI[365]
port 294 nsew signal tristate
rlabel metal2 s 21546 3800 21602 4400 6 HI[366]
port 295 nsew signal tristate
rlabel metal2 s 21822 3800 21878 4400 6 HI[367]
port 296 nsew signal tristate
rlabel metal2 s 22098 3800 22154 4400 6 HI[368]
port 297 nsew signal tristate
rlabel metal2 s 22374 3800 22430 4400 6 HI[369]
port 298 nsew signal tristate
rlabel metal2 s 22650 3800 22706 4400 6 HI[36]
port 299 nsew signal tristate
rlabel metal2 s 22926 3800 22982 4400 6 HI[370]
port 300 nsew signal tristate
rlabel metal2 s 23202 3800 23258 4400 6 HI[371]
port 301 nsew signal tristate
rlabel metal2 s 23478 3800 23534 4400 6 HI[372]
port 302 nsew signal tristate
rlabel metal2 s 23754 3800 23810 4400 6 HI[373]
port 303 nsew signal tristate
rlabel metal2 s 24030 3800 24086 4400 6 HI[374]
port 304 nsew signal tristate
rlabel metal2 s 24306 3800 24362 4400 6 HI[375]
port 305 nsew signal tristate
rlabel metal2 s 24582 3800 24638 4400 6 HI[376]
port 306 nsew signal tristate
rlabel metal2 s 24858 3800 24914 4400 6 HI[377]
port 307 nsew signal tristate
rlabel metal2 s 25134 3800 25190 4400 6 HI[378]
port 308 nsew signal tristate
rlabel metal2 s 25410 3800 25466 4400 6 HI[379]
port 309 nsew signal tristate
rlabel metal2 s 25686 3800 25742 4400 6 HI[37]
port 310 nsew signal tristate
rlabel metal2 s 25962 3800 26018 4400 6 HI[380]
port 311 nsew signal tristate
rlabel metal2 s 26238 3800 26294 4400 6 HI[381]
port 312 nsew signal tristate
rlabel metal2 s 26514 3800 26570 4400 6 HI[382]
port 313 nsew signal tristate
rlabel metal2 s 26790 3800 26846 4400 6 HI[383]
port 314 nsew signal tristate
rlabel metal2 s 27066 3800 27122 4400 6 HI[384]
port 315 nsew signal tristate
rlabel metal2 s 27342 3800 27398 4400 6 HI[385]
port 316 nsew signal tristate
rlabel metal2 s 27618 3800 27674 4400 6 HI[386]
port 317 nsew signal tristate
rlabel metal2 s 27894 3800 27950 4400 6 HI[387]
port 318 nsew signal tristate
rlabel metal2 s 28170 3800 28226 4400 6 HI[388]
port 319 nsew signal tristate
rlabel metal2 s 28446 3800 28502 4400 6 HI[389]
port 320 nsew signal tristate
rlabel metal2 s 28722 3800 28778 4400 6 HI[38]
port 321 nsew signal tristate
rlabel metal2 s 28998 3800 29054 4400 6 HI[390]
port 322 nsew signal tristate
rlabel metal2 s 29274 3800 29330 4400 6 HI[391]
port 323 nsew signal tristate
rlabel metal2 s 29550 3800 29606 4400 6 HI[392]
port 324 nsew signal tristate
rlabel metal2 s 29826 3800 29882 4400 6 HI[393]
port 325 nsew signal tristate
rlabel metal2 s 30102 3800 30158 4400 6 HI[394]
port 326 nsew signal tristate
rlabel metal2 s 30378 3800 30434 4400 6 HI[395]
port 327 nsew signal tristate
rlabel metal2 s 30654 3800 30710 4400 6 HI[396]
port 328 nsew signal tristate
rlabel metal2 s 30930 3800 30986 4400 6 HI[397]
port 329 nsew signal tristate
rlabel metal2 s 31206 3800 31262 4400 6 HI[398]
port 330 nsew signal tristate
rlabel metal2 s 31482 3800 31538 4400 6 HI[399]
port 331 nsew signal tristate
rlabel metal2 s 31758 3800 31814 4400 6 HI[39]
port 332 nsew signal tristate
rlabel metal2 s 32034 3800 32090 4400 6 HI[3]
port 333 nsew signal tristate
rlabel metal2 s 32310 3800 32366 4400 6 HI[400]
port 334 nsew signal tristate
rlabel metal2 s 32586 3800 32642 4400 6 HI[401]
port 335 nsew signal tristate
rlabel metal2 s 32862 3800 32918 4400 6 HI[402]
port 336 nsew signal tristate
rlabel metal2 s 33138 3800 33194 4400 6 HI[403]
port 337 nsew signal tristate
rlabel metal2 s 33414 3800 33470 4400 6 HI[404]
port 338 nsew signal tristate
rlabel metal2 s 33690 3800 33746 4400 6 HI[405]
port 339 nsew signal tristate
rlabel metal2 s 33966 3800 34022 4400 6 HI[406]
port 340 nsew signal tristate
rlabel metal2 s 34242 3800 34298 4400 6 HI[407]
port 341 nsew signal tristate
rlabel metal2 s 34518 3800 34574 4400 6 HI[408]
port 342 nsew signal tristate
rlabel metal2 s 34794 3800 34850 4400 6 HI[409]
port 343 nsew signal tristate
rlabel metal2 s 35070 3800 35126 4400 6 HI[40]
port 344 nsew signal tristate
rlabel metal2 s 35346 3800 35402 4400 6 HI[410]
port 345 nsew signal tristate
rlabel metal2 s 35622 3800 35678 4400 6 HI[411]
port 346 nsew signal tristate
rlabel metal2 s 35898 3800 35954 4400 6 HI[412]
port 347 nsew signal tristate
rlabel metal2 s 36174 3800 36230 4400 6 HI[413]
port 348 nsew signal tristate
rlabel metal2 s 36450 3800 36506 4400 6 HI[414]
port 349 nsew signal tristate
rlabel metal2 s 36726 3800 36782 4400 6 HI[415]
port 350 nsew signal tristate
rlabel metal2 s 37002 3800 37058 4400 6 HI[416]
port 351 nsew signal tristate
rlabel metal2 s 37278 3800 37334 4400 6 HI[417]
port 352 nsew signal tristate
rlabel metal2 s 37554 3800 37610 4400 6 HI[418]
port 353 nsew signal tristate
rlabel metal2 s 37830 3800 37886 4400 6 HI[419]
port 354 nsew signal tristate
rlabel metal2 s 38106 3800 38162 4400 6 HI[41]
port 355 nsew signal tristate
rlabel metal2 s 38382 3800 38438 4400 6 HI[420]
port 356 nsew signal tristate
rlabel metal2 s 38658 3800 38714 4400 6 HI[421]
port 357 nsew signal tristate
rlabel metal2 s 38934 3800 38990 4400 6 HI[422]
port 358 nsew signal tristate
rlabel metal2 s 39210 3800 39266 4400 6 HI[423]
port 359 nsew signal tristate
rlabel metal2 s 39486 3800 39542 4400 6 HI[424]
port 360 nsew signal tristate
rlabel metal2 s 39762 3800 39818 4400 6 HI[425]
port 361 nsew signal tristate
rlabel metal2 s 40038 3800 40094 4400 6 HI[426]
port 362 nsew signal tristate
rlabel metal2 s 40314 3800 40370 4400 6 HI[427]
port 363 nsew signal tristate
rlabel metal2 s 40590 3800 40646 4400 6 HI[428]
port 364 nsew signal tristate
rlabel metal2 s 40866 3800 40922 4400 6 HI[429]
port 365 nsew signal tristate
rlabel metal2 s 41142 3800 41198 4400 6 HI[42]
port 366 nsew signal tristate
rlabel metal2 s 41418 3800 41474 4400 6 HI[430]
port 367 nsew signal tristate
rlabel metal2 s 41694 3800 41750 4400 6 HI[431]
port 368 nsew signal tristate
rlabel metal2 s 41970 3800 42026 4400 6 HI[432]
port 369 nsew signal tristate
rlabel metal2 s 42246 3800 42302 4400 6 HI[433]
port 370 nsew signal tristate
rlabel metal2 s 42522 3800 42578 4400 6 HI[434]
port 371 nsew signal tristate
rlabel metal2 s 42798 3800 42854 4400 6 HI[435]
port 372 nsew signal tristate
rlabel metal2 s 43074 3800 43130 4400 6 HI[436]
port 373 nsew signal tristate
rlabel metal2 s 43350 3800 43406 4400 6 HI[437]
port 374 nsew signal tristate
rlabel metal2 s 43626 3800 43682 4400 6 HI[438]
port 375 nsew signal tristate
rlabel metal2 s 43902 3800 43958 4400 6 HI[439]
port 376 nsew signal tristate
rlabel metal2 s 44178 3800 44234 4400 6 HI[43]
port 377 nsew signal tristate
rlabel metal2 s 44454 3800 44510 4400 6 HI[440]
port 378 nsew signal tristate
rlabel metal2 s 44730 3800 44786 4400 6 HI[441]
port 379 nsew signal tristate
rlabel metal2 s 45006 3800 45062 4400 6 HI[442]
port 380 nsew signal tristate
rlabel metal2 s 45282 3800 45338 4400 6 HI[443]
port 381 nsew signal tristate
rlabel metal2 s 45558 3800 45614 4400 6 HI[444]
port 382 nsew signal tristate
rlabel metal2 s 45834 3800 45890 4400 6 HI[445]
port 383 nsew signal tristate
rlabel metal2 s 46110 3800 46166 4400 6 HI[446]
port 384 nsew signal tristate
rlabel metal2 s 46386 3800 46442 4400 6 HI[447]
port 385 nsew signal tristate
rlabel metal2 s 46662 3800 46718 4400 6 HI[448]
port 386 nsew signal tristate
rlabel metal2 s 46938 3800 46994 4400 6 HI[449]
port 387 nsew signal tristate
rlabel metal2 s 47214 3800 47270 4400 6 HI[44]
port 388 nsew signal tristate
rlabel metal2 s 47490 3800 47546 4400 6 HI[450]
port 389 nsew signal tristate
rlabel metal2 s 47766 3800 47822 4400 6 HI[451]
port 390 nsew signal tristate
rlabel metal2 s 48042 3800 48098 4400 6 HI[452]
port 391 nsew signal tristate
rlabel metal2 s 48318 3800 48374 4400 6 HI[453]
port 392 nsew signal tristate
rlabel metal2 s 48594 3800 48650 4400 6 HI[454]
port 393 nsew signal tristate
rlabel metal2 s 48870 3800 48926 4400 6 HI[455]
port 394 nsew signal tristate
rlabel metal2 s 49146 3800 49202 4400 6 HI[456]
port 395 nsew signal tristate
rlabel metal2 s 49422 3800 49478 4400 6 HI[457]
port 396 nsew signal tristate
rlabel metal2 s 49698 3800 49754 4400 6 HI[458]
port 397 nsew signal tristate
rlabel metal2 s 49974 3800 50030 4400 6 HI[459]
port 398 nsew signal tristate
rlabel metal2 s 50250 3800 50306 4400 6 HI[45]
port 399 nsew signal tristate
rlabel metal2 s 50526 3800 50582 4400 6 HI[460]
port 400 nsew signal tristate
rlabel metal2 s 50802 3800 50858 4400 6 HI[461]
port 401 nsew signal tristate
rlabel metal2 s 51078 3800 51134 4400 6 HI[462]
port 402 nsew signal tristate
rlabel metal2 s 51354 3800 51410 4400 6 HI[46]
port 403 nsew signal tristate
rlabel metal2 s 51630 3800 51686 4400 6 HI[47]
port 404 nsew signal tristate
rlabel metal2 s 51906 3800 51962 4400 6 HI[48]
port 405 nsew signal tristate
rlabel metal2 s 52182 3800 52238 4400 6 HI[49]
port 406 nsew signal tristate
rlabel metal2 s 52458 3800 52514 4400 6 HI[4]
port 407 nsew signal tristate
rlabel metal2 s 52734 3800 52790 4400 6 HI[50]
port 408 nsew signal tristate
rlabel metal2 s 53010 3800 53066 4400 6 HI[51]
port 409 nsew signal tristate
rlabel metal2 s 53286 3800 53342 4400 6 HI[52]
port 410 nsew signal tristate
rlabel metal2 s 53562 3800 53618 4400 6 HI[53]
port 411 nsew signal tristate
rlabel metal2 s 53838 3800 53894 4400 6 HI[54]
port 412 nsew signal tristate
rlabel metal2 s 54114 3800 54170 4400 6 HI[55]
port 413 nsew signal tristate
rlabel metal2 s 54390 3800 54446 4400 6 HI[56]
port 414 nsew signal tristate
rlabel metal2 s 54666 3800 54722 4400 6 HI[57]
port 415 nsew signal tristate
rlabel metal2 s 54942 3800 54998 4400 6 HI[58]
port 416 nsew signal tristate
rlabel metal2 s 55218 3800 55274 4400 6 HI[59]
port 417 nsew signal tristate
rlabel metal2 s 55494 3800 55550 4400 6 HI[5]
port 418 nsew signal tristate
rlabel metal2 s 55770 3800 55826 4400 6 HI[60]
port 419 nsew signal tristate
rlabel metal2 s 56046 3800 56102 4400 6 HI[61]
port 420 nsew signal tristate
rlabel metal2 s 56322 3800 56378 4400 6 HI[62]
port 421 nsew signal tristate
rlabel metal2 s 56598 3800 56654 4400 6 HI[63]
port 422 nsew signal tristate
rlabel metal2 s 56874 3800 56930 4400 6 HI[64]
port 423 nsew signal tristate
rlabel metal2 s 57150 3800 57206 4400 6 HI[65]
port 424 nsew signal tristate
rlabel metal2 s 57426 3800 57482 4400 6 HI[66]
port 425 nsew signal tristate
rlabel metal2 s 57702 3800 57758 4400 6 HI[67]
port 426 nsew signal tristate
rlabel metal2 s 57978 3800 58034 4400 6 HI[68]
port 427 nsew signal tristate
rlabel metal2 s 58254 3800 58310 4400 6 HI[69]
port 428 nsew signal tristate
rlabel metal2 s 58530 3800 58586 4400 6 HI[6]
port 429 nsew signal tristate
rlabel metal2 s 58806 3800 58862 4400 6 HI[70]
port 430 nsew signal tristate
rlabel metal2 s 59082 3800 59138 4400 6 HI[71]
port 431 nsew signal tristate
rlabel metal2 s 59358 3800 59414 4400 6 HI[72]
port 432 nsew signal tristate
rlabel metal2 s 59634 3800 59690 4400 6 HI[73]
port 433 nsew signal tristate
rlabel metal2 s 59910 3800 59966 4400 6 HI[74]
port 434 nsew signal tristate
rlabel metal2 s 60186 3800 60242 4400 6 HI[75]
port 435 nsew signal tristate
rlabel metal2 s 60462 3800 60518 4400 6 HI[76]
port 436 nsew signal tristate
rlabel metal2 s 60738 3800 60794 4400 6 HI[77]
port 437 nsew signal tristate
rlabel metal2 s 61014 3800 61070 4400 6 HI[78]
port 438 nsew signal tristate
rlabel metal2 s 61290 3800 61346 4400 6 HI[79]
port 439 nsew signal tristate
rlabel metal2 s 61566 3800 61622 4400 6 HI[7]
port 440 nsew signal tristate
rlabel metal2 s 61842 3800 61898 4400 6 HI[80]
port 441 nsew signal tristate
rlabel metal2 s 62118 3800 62174 4400 6 HI[81]
port 442 nsew signal tristate
rlabel metal2 s 62394 3800 62450 4400 6 HI[82]
port 443 nsew signal tristate
rlabel metal2 s 62670 3800 62726 4400 6 HI[83]
port 444 nsew signal tristate
rlabel metal2 s 62946 3800 63002 4400 6 HI[84]
port 445 nsew signal tristate
rlabel metal2 s 63222 3800 63278 4400 6 HI[85]
port 446 nsew signal tristate
rlabel metal2 s 63498 3800 63554 4400 6 HI[86]
port 447 nsew signal tristate
rlabel metal2 s 63774 3800 63830 4400 6 HI[87]
port 448 nsew signal tristate
rlabel metal2 s 64050 3800 64106 4400 6 HI[88]
port 449 nsew signal tristate
rlabel metal2 s 64326 3800 64382 4400 6 HI[89]
port 450 nsew signal tristate
rlabel metal2 s 64602 3800 64658 4400 6 HI[8]
port 451 nsew signal tristate
rlabel metal2 s 64878 3800 64934 4400 6 HI[90]
port 452 nsew signal tristate
rlabel metal2 s 65154 3800 65210 4400 6 HI[91]
port 453 nsew signal tristate
rlabel metal2 s 65430 3800 65486 4400 6 HI[92]
port 454 nsew signal tristate
rlabel metal2 s 65706 3800 65762 4400 6 HI[93]
port 455 nsew signal tristate
rlabel metal2 s 65982 3800 66038 4400 6 HI[94]
port 456 nsew signal tristate
rlabel metal2 s 66258 3800 66314 4400 6 HI[95]
port 457 nsew signal tristate
rlabel metal2 s 66534 3800 66590 4400 6 HI[96]
port 458 nsew signal tristate
rlabel metal2 s 66810 3800 66866 4400 6 HI[97]
port 459 nsew signal tristate
rlabel metal2 s 67086 3800 67142 4400 6 HI[98]
port 460 nsew signal tristate
rlabel metal2 s 67362 3800 67418 4400 6 HI[99]
port 461 nsew signal tristate
rlabel metal2 s 67638 3800 67694 4400 6 HI[9]
port 462 nsew signal tristate
rlabel metal3 s 1288 1190 68816 1290 6 vccd1
port 463 nsew power input
rlabel metal2 s 7238 1040 7338 3312 6 vccd1
port 463 nsew power input
rlabel metal2 s 19238 1040 19338 3312 6 vccd1
port 463 nsew power input
rlabel metal2 s 31238 1040 31338 3312 6 vccd1
port 463 nsew power input
rlabel metal2 s 43238 1040 43338 3312 6 vccd1
port 463 nsew power input
rlabel metal2 s 55238 1040 55338 3312 6 vccd1
port 463 nsew power input
rlabel metal2 s 67238 1040 67338 3312 6 vccd1
port 463 nsew power input
rlabel metal3 s 1288 2270 68816 2370 6 vssd1
port 464 nsew ground input
rlabel metal2 s 13238 1040 13338 3312 6 vssd1
port 464 nsew ground input
rlabel metal2 s 25238 1040 25338 3312 6 vssd1
port 464 nsew ground input
rlabel metal2 s 37238 1040 37338 3312 6 vssd1
port 464 nsew ground input
rlabel metal2 s 49238 1040 49338 3312 6 vssd1
port 464 nsew ground input
rlabel metal2 s 61238 1040 61338 3312 6 vssd1
port 464 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 70000 4400
<< end >>
