magic
tech sky130A
magscale 1 2
timestamp 1666119982
<< checkpaint >>
rect -1260 -1260 35260 14274
<< isosubstrate >>
rect 1090 4514 2656 4518
rect 1090 1592 2678 4514
rect 1090 1552 2656 1592
<< viali >>
rect 3985 11849 4019 11883
rect 1317 11713 1351 11747
rect 5457 11713 5491 11747
rect 6561 11713 6595 11747
rect 8585 11713 8619 11747
rect 9321 11713 9355 11747
rect 1409 11645 1443 11679
rect 3433 11645 3467 11679
rect 3617 11645 3651 11679
rect 3801 11645 3835 11679
rect 4077 11645 4111 11679
rect 6469 11645 6503 11679
rect 9873 11645 9907 11679
rect 10057 11645 10091 11679
rect 6837 11577 6871 11611
rect 9505 11577 9539 11611
rect 9597 11577 9631 11611
rect 2513 11509 2547 11543
rect 6285 11509 6319 11543
rect 8769 11509 8803 11543
rect 1317 11305 1351 11339
rect 1685 11305 1719 11339
rect 7205 11237 7239 11271
rect 1501 11169 1535 11203
rect 3433 11169 3467 11203
rect 3893 11169 3927 11203
rect 5365 11169 5399 11203
rect 7021 11169 7055 11203
rect 9413 11169 9447 11203
rect 3525 11101 3559 11135
rect 6193 11101 6227 11135
rect 7297 11101 7331 11135
rect 7573 11101 7607 11135
rect 7941 11101 7975 11135
rect 5925 11033 5959 11067
rect 9973 11033 10007 11067
rect 3175 10965 3209 10999
rect 6837 10965 6871 10999
rect 1317 10761 1351 10795
rect 3709 10693 3743 10727
rect 8769 10693 8803 10727
rect 1685 10625 1719 10659
rect 3985 10625 4019 10659
rect 6009 10625 6043 10659
rect 6101 10625 6135 10659
rect 9321 10625 9355 10659
rect 1409 10557 1443 10591
rect 3893 10557 3927 10591
rect 6469 10557 6503 10591
rect 7941 10557 7975 10591
rect 9597 10557 9631 10591
rect 10057 10557 10091 10591
rect 3433 10489 3467 10523
rect 4261 10489 4295 10523
rect 8505 10489 8539 10523
rect 9781 10489 9815 10523
rect 6929 10217 6963 10251
rect 1685 10149 1719 10183
rect 3433 10149 3467 10183
rect 9965 10149 9999 10183
rect 5365 10081 5399 10115
rect 7389 10081 7423 10115
rect 8861 10081 8895 10115
rect 9597 10081 9631 10115
rect 1409 10013 1443 10047
rect 3525 10013 3559 10047
rect 3893 10013 3927 10047
rect 6285 10013 6319 10047
rect 7021 10013 7055 10047
rect 9781 10013 9815 10047
rect 1317 9877 1351 9911
rect 5929 9877 5963 9911
rect 9421 9877 9455 9911
rect 6757 9673 6791 9707
rect 1685 9537 1719 9571
rect 3433 9537 3467 9571
rect 4353 9537 4387 9571
rect 4721 9537 4755 9571
rect 7481 9537 7515 9571
rect 8217 9537 8251 9571
rect 1409 9469 1443 9503
rect 4169 9469 4203 9503
rect 6193 9469 6227 9503
rect 8401 9469 8435 9503
rect 8769 9469 8803 9503
rect 9597 9469 9631 9503
rect 9965 9469 9999 9503
rect 1317 9401 1351 9435
rect 9781 9401 9815 9435
rect 3617 9333 3651 9367
rect 6929 9333 6963 9367
rect 7665 9333 7699 9367
rect 8493 9333 8527 9367
rect 9413 9333 9447 9367
rect 6009 9061 6043 9095
rect 3893 8993 3927 9027
rect 8217 8993 8251 9027
rect 1317 8925 1351 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6837 8925 6871 8959
rect 9689 8925 9723 8959
rect 10057 8925 10091 8959
rect 2789 8857 2823 8891
rect 7652 8857 7686 8891
rect 1869 8789 1903 8823
rect 6285 8789 6319 8823
rect 7389 8789 7423 8823
rect 1593 8585 1627 8619
rect 9689 8585 9723 8619
rect 2145 8517 2179 8551
rect 6009 8517 6043 8551
rect 8493 8517 8527 8551
rect 1225 8449 1259 8483
rect 3617 8449 3651 8483
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 8401 8449 8435 8483
rect 1409 8381 1443 8415
rect 3433 8381 3467 8415
rect 5641 8381 5675 8415
rect 5917 8381 5951 8415
rect 6193 8381 6227 8415
rect 9321 8381 9355 8415
rect 9597 8381 9631 8415
rect 9965 8381 9999 8415
rect 8769 8245 8803 8279
rect 1317 8041 1351 8075
rect 9689 7973 9723 8007
rect 1409 7905 1443 7939
rect 3157 7905 3191 7939
rect 3893 7905 3927 7939
rect 5365 7905 5399 7939
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 6837 7905 6871 7939
rect 7205 7905 7239 7939
rect 8677 7905 8711 7939
rect 9505 7905 9539 7939
rect 2605 7837 2639 7871
rect 3525 7837 3559 7871
rect 9781 7837 9815 7871
rect 5929 7701 5963 7735
rect 6377 7701 6411 7735
rect 9237 7701 9271 7735
rect 8861 7497 8895 7531
rect 1409 7361 1443 7395
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 4445 7361 4479 7395
rect 4721 7361 4755 7395
rect 6469 7361 6503 7395
rect 8585 7361 8619 7395
rect 9781 7361 9815 7395
rect 3709 7293 3743 7327
rect 6561 7293 6595 7327
rect 8769 7293 8803 7327
rect 9689 7293 9723 7327
rect 6837 7225 6871 7259
rect 9045 7225 9079 7259
rect 9551 7225 9585 7259
rect 1317 7157 1351 7191
rect 4353 7157 4387 7191
rect 10057 6953 10091 6987
rect 3433 6885 3467 6919
rect 6929 6885 6963 6919
rect 1225 6817 1259 6851
rect 3525 6817 3559 6851
rect 5365 6817 5399 6851
rect 6193 6817 6227 6851
rect 8953 6817 8987 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3893 6749 3927 6783
rect 6745 6749 6779 6783
rect 7113 6749 7147 6783
rect 7481 6749 7515 6783
rect 9873 6749 9907 6783
rect 9689 6681 9723 6715
rect 5929 6613 5963 6647
rect 9137 6613 9171 6647
rect 9513 6613 9547 6647
rect 8401 6409 8435 6443
rect 1593 6341 1627 6375
rect 8769 6341 8803 6375
rect 1225 6273 1259 6307
rect 5365 6273 5399 6307
rect 5825 6273 5859 6307
rect 8217 6273 8251 6307
rect 1409 6205 1443 6239
rect 3433 6205 3467 6239
rect 5457 6205 5491 6239
rect 7297 6205 7331 6239
rect 8493 6205 8527 6239
rect 9137 6205 9171 6239
rect 9505 6205 9539 6239
rect 9781 6205 9815 6239
rect 3617 6137 3651 6171
rect 10057 6137 10091 6171
rect 2145 6069 2179 6103
rect 7861 6069 7895 6103
rect 2145 5865 2179 5899
rect 9965 5865 9999 5899
rect 1225 5797 1259 5831
rect 3433 5797 3467 5831
rect 4261 5797 4295 5831
rect 6009 5797 6043 5831
rect 6561 5797 6595 5831
rect 9137 5797 9171 5831
rect 9459 5797 9493 5831
rect 9873 5797 9907 5831
rect 1409 5729 1443 5763
rect 3617 5729 3651 5763
rect 6193 5729 6227 5763
rect 8585 5729 8619 5763
rect 9229 5729 9263 5763
rect 1593 5661 1627 5695
rect 3985 5661 4019 5695
rect 6377 5661 6411 5695
rect 7941 5661 7975 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 3801 5525 3835 5559
rect 9505 5525 9539 5559
rect 5825 5321 5859 5355
rect 3341 5185 3375 5219
rect 5457 5185 5491 5219
rect 6745 5185 6779 5219
rect 9413 5185 9447 5219
rect 3525 5117 3559 5151
rect 3801 5117 3835 5151
rect 6009 5117 6043 5151
rect 8033 5117 8067 5151
rect 10057 5117 10091 5151
rect 3709 5049 3743 5083
rect 3433 4777 3467 4811
rect 7573 4777 7607 4811
rect 8401 4777 8435 4811
rect 9597 4777 9631 4811
rect 3985 4709 4019 4743
rect 8125 4709 8159 4743
rect 9137 4709 9171 4743
rect 3617 4641 3651 4675
rect 3801 4641 3835 4675
rect 4721 4641 4755 4675
rect 6193 4641 6227 4675
rect 7021 4641 7055 4675
rect 8677 4641 8711 4675
rect 8953 4641 8987 4675
rect 10057 4641 10091 4675
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 7757 4573 7791 4607
rect 7941 4573 7975 4607
rect 8585 4573 8619 4607
rect 9413 4505 9447 4539
rect 6753 4437 6787 4471
rect 9873 4437 9907 4471
rect 5549 4165 5583 4199
rect 5089 4097 5123 4131
rect 3341 4029 3375 4063
rect 5181 4029 5215 4063
rect 5365 4029 5399 4063
rect 6009 4029 6043 4063
rect 6193 4029 6227 4063
rect 8125 4029 8159 4063
rect 10057 4029 10091 4063
rect 8033 3961 8067 3995
rect 5825 3893 5859 3927
rect 3341 3689 3375 3723
rect 8769 3621 8803 3655
rect 9689 3621 9723 3655
rect 3617 3553 3651 3587
rect 5733 3553 5767 3587
rect 6193 3553 6227 3587
rect 8861 3553 8895 3587
rect 9045 3553 9079 3587
rect 9873 3553 9907 3587
rect 3893 3485 3927 3519
rect 3985 3485 4019 3519
rect 5365 3485 5399 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9597 3485 9631 3519
rect 8125 3417 8159 3451
rect 9229 3349 9263 3383
rect 5273 3145 5307 3179
rect 5825 3145 5859 3179
rect 6101 3145 6135 3179
rect 6377 3145 6411 3179
rect 7021 3145 7055 3179
rect 7297 3145 7331 3179
rect 6653 3077 6687 3111
rect 5089 3009 5123 3043
rect 5365 2941 5399 2975
rect 5917 2941 5951 2975
rect 6193 2941 6227 2975
rect 7113 2941 7147 2975
rect 7205 2941 7239 2975
rect 3341 2873 3375 2907
rect 5457 2805 5491 2839
rect 6745 2805 6779 2839
rect 8953 2601 8987 2635
rect 9597 2533 9631 2567
rect 3617 2465 3651 2499
rect 6101 2465 6135 2499
rect 8125 2465 8159 2499
rect 8677 2465 8711 2499
rect 8769 2465 8803 2499
rect 9505 2465 9539 2499
rect 9781 2465 9815 2499
rect 3893 2397 3927 2431
rect 3985 2397 4019 2431
rect 5457 2397 5491 2431
rect 6745 2397 6779 2431
rect 9965 2397 9999 2431
rect 9321 2329 9355 2363
rect 3433 2261 3467 2295
rect 8493 2261 8527 2295
rect 3525 2057 3559 2091
rect 3801 2057 3835 2091
rect 4077 2057 4111 2091
rect 4353 2057 4387 2091
rect 4905 2057 4939 2091
rect 5825 2057 5859 2091
rect 6009 2057 6043 2091
rect 4537 1989 4571 2023
rect 5549 1989 5583 2023
rect 4721 1921 4755 1955
rect 5089 1921 5123 1955
rect 9413 1921 9447 1955
rect 3341 1853 3375 1887
rect 3893 1853 3927 1887
rect 4169 1853 4203 1887
rect 4261 1853 4295 1887
rect 6469 1853 6503 1887
rect 9873 1853 9907 1887
rect 8033 1785 8067 1819
rect 5273 1717 5307 1751
rect 3433 1513 3467 1547
rect 3709 1513 3743 1547
rect 7021 1513 7055 1547
rect 9229 1513 9263 1547
rect 9965 1513 9999 1547
rect 3341 1377 3375 1411
rect 3801 1377 3835 1411
rect 6101 1377 6135 1411
rect 8033 1377 8067 1411
rect 9045 1377 9079 1411
rect 9413 1377 9447 1411
rect 9781 1377 9815 1411
rect 3985 1309 4019 1343
rect 5457 1309 5491 1343
rect 8401 1309 8435 1343
rect 8493 1309 8527 1343
rect 8861 1309 8895 1343
rect 9597 1241 9631 1275
rect 8677 1173 8711 1207
rect 1685 969 1719 1003
rect 5089 969 5123 1003
rect 9229 969 9263 1003
rect 9873 969 9907 1003
rect 3065 901 3099 935
rect 3341 901 3375 935
rect 6561 901 6595 935
rect 8585 901 8619 935
rect 3985 833 4019 867
rect 2973 765 3007 799
rect 6009 765 6043 799
rect 6653 765 6687 799
rect 9413 765 9447 799
rect 10057 765 10091 799
rect 3709 697 3743 731
rect 9597 697 9631 731
rect 6285 629 6319 663
rect 8861 629 8895 663
rect 9137 629 9171 663
<< metal1 >>
rect 1302 12044 1308 12096
rect 1360 12084 1366 12096
rect 3786 12084 3792 12096
rect 1360 12056 3792 12084
rect 1360 12044 1366 12056
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 5718 12084 5724 12096
rect 3844 12056 5724 12084
rect 3844 12044 3850 12056
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 920 11994 10396 12016
rect 920 11942 2566 11994
rect 2618 11942 2630 11994
rect 2682 11942 2694 11994
rect 2746 11942 2758 11994
rect 2810 11942 2822 11994
rect 2874 11942 7566 11994
rect 7618 11942 7630 11994
rect 7682 11942 7694 11994
rect 7746 11942 7758 11994
rect 7810 11942 7822 11994
rect 7874 11942 10396 11994
rect 920 11920 10396 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3510 11880 3516 11892
rect 3016 11852 3516 11880
rect 3016 11840 3022 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 8018 11880 8024 11892
rect 4019 11852 8024 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 4798 11812 4804 11824
rect 3436 11784 4804 11812
rect 1305 11747 1363 11753
rect 1305 11713 1317 11747
rect 1351 11744 1363 11747
rect 1351 11716 3372 11744
rect 1351 11713 1363 11716
rect 1305 11707 1363 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2958 11676 2964 11688
rect 1443 11648 2964 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 3344 11608 3372 11716
rect 3436 11685 3464 11784
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 4338 11744 4344 11756
rect 3528 11716 4344 11744
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3528 11608 3556 11716
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5684 11716 6561 11744
rect 5684 11704 5690 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 7524 11716 8585 11744
rect 7524 11704 7530 11716
rect 8573 11713 8585 11716
rect 8619 11744 8631 11747
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8619 11716 9321 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11645 3663 11679
rect 3786 11676 3792 11688
rect 3747 11648 3792 11676
rect 3605 11639 3663 11645
rect 3344 11580 3556 11608
rect 3620 11608 3648 11639
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 4065 11679 4123 11685
rect 4065 11676 4077 11679
rect 3936 11648 4077 11676
rect 3936 11636 3942 11648
rect 4065 11645 4077 11648
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 4982 11676 4988 11688
rect 4488 11648 4988 11676
rect 4488 11636 4494 11648
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 6270 11636 6276 11688
rect 6328 11676 6334 11688
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 6328 11648 6469 11676
rect 6328 11636 6334 11648
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 9088 11648 9873 11676
rect 9088 11636 9094 11648
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11676 10103 11679
rect 10226 11676 10232 11688
rect 10091 11648 10232 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 4706 11608 4712 11620
rect 3620 11580 4712 11608
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 6288 11608 6316 11636
rect 5644 11580 6316 11608
rect 6825 11611 6883 11617
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 5644 11540 5672 11580
rect 6825 11577 6837 11611
rect 6871 11608 6883 11611
rect 6914 11608 6920 11620
rect 6871 11580 6920 11608
rect 6871 11577 6883 11580
rect 6825 11571 6883 11577
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 8202 11608 8208 11620
rect 8050 11580 8208 11608
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 9490 11608 9496 11620
rect 9451 11580 9496 11608
rect 9490 11568 9496 11580
rect 9548 11568 9554 11620
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 9640 11580 9685 11608
rect 9640 11568 9646 11580
rect 3660 11512 5672 11540
rect 6273 11543 6331 11549
rect 3660 11500 3666 11512
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6638 11540 6644 11552
rect 6319 11512 6644 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8168 11512 8769 11540
rect 8168 11500 8174 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 920 11450 10396 11472
rect 920 11398 5066 11450
rect 5118 11398 5130 11450
rect 5182 11398 5194 11450
rect 5246 11398 5258 11450
rect 5310 11398 5322 11450
rect 5374 11398 10396 11450
rect 920 11376 10396 11398
rect 1302 11336 1308 11348
rect 1263 11308 1308 11336
rect 1302 11296 1308 11308
rect 1360 11296 1366 11348
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 3878 11336 3884 11348
rect 1719 11308 3884 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6546 11336 6552 11348
rect 6052 11308 6552 11336
rect 6052 11296 6058 11308
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 2406 11228 2412 11280
rect 2464 11228 2470 11280
rect 7193 11271 7251 11277
rect 7193 11268 7205 11271
rect 5014 11240 7205 11268
rect 7193 11237 7205 11240
rect 7239 11237 7251 11271
rect 10318 11268 10324 11280
rect 9062 11240 10324 11268
rect 7193 11231 7251 11237
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 1489 11163 1547 11169
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 3694 11200 3700 11212
rect 3467 11172 3700 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 1504 11132 1532 11163
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 5353 11203 5411 11209
rect 3936 11172 3981 11200
rect 3936 11160 3942 11172
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 6086 11200 6092 11212
rect 5399 11172 6092 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7098 11200 7104 11212
rect 7055 11172 7104 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 9398 11200 9404 11212
rect 9359 11172 9404 11200
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 2130 11132 2136 11144
rect 1504 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3786 11132 3792 11144
rect 3559 11104 3792 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6052 11104 6193 11132
rect 6052 11092 6058 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 6181 11095 6239 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7432 11104 7573 11132
rect 7432 11092 7438 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8110 11132 8116 11144
rect 7975 11104 8116 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 5913 11067 5971 11073
rect 5913 11064 5925 11067
rect 5868 11036 5925 11064
rect 5868 11024 5874 11036
rect 5913 11033 5925 11036
rect 5959 11033 5971 11067
rect 7466 11064 7472 11076
rect 5913 11027 5971 11033
rect 6380 11036 7472 11064
rect 3163 10999 3221 11005
rect 3163 10965 3175 10999
rect 3209 10996 3221 10999
rect 6380 10996 6408 11036
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 9961 11067 10019 11073
rect 9961 11064 9973 11067
rect 9916 11036 9973 11064
rect 9916 11024 9922 11036
rect 9961 11033 9973 11036
rect 10007 11033 10019 11067
rect 9961 11027 10019 11033
rect 3209 10968 6408 10996
rect 3209 10965 3221 10968
rect 3163 10959 3221 10965
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6825 10999 6883 11005
rect 6825 10996 6837 10999
rect 6512 10968 6837 10996
rect 6512 10956 6518 10968
rect 6825 10965 6837 10968
rect 6871 10965 6883 10999
rect 6825 10959 6883 10965
rect 920 10906 10396 10928
rect 920 10854 2566 10906
rect 2618 10854 2630 10906
rect 2682 10854 2694 10906
rect 2746 10854 2758 10906
rect 2810 10854 2822 10906
rect 2874 10854 7566 10906
rect 7618 10854 7630 10906
rect 7682 10854 7694 10906
rect 7746 10854 7758 10906
rect 7810 10854 7822 10906
rect 7874 10854 10396 10906
rect 920 10832 10396 10854
rect 1305 10795 1363 10801
rect 1305 10761 1317 10795
rect 1351 10792 1363 10795
rect 1486 10792 1492 10804
rect 1351 10764 1492 10792
rect 1351 10761 1363 10764
rect 1305 10755 1363 10761
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 2746 10764 5764 10792
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2746 10656 2774 10764
rect 3234 10684 3240 10736
rect 3292 10724 3298 10736
rect 3697 10727 3755 10733
rect 3697 10724 3709 10727
rect 3292 10696 3709 10724
rect 3292 10684 3298 10696
rect 3697 10693 3709 10696
rect 3743 10724 3755 10727
rect 3786 10724 3792 10736
rect 3743 10696 3792 10724
rect 3743 10693 3755 10696
rect 3697 10687 3755 10693
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 1719 10628 2774 10656
rect 3973 10659 4031 10665
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 5626 10656 5632 10668
rect 4019 10628 5632 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 3881 10591 3939 10597
rect 3881 10588 3893 10591
rect 3660 10560 3893 10588
rect 3660 10548 3666 10560
rect 3881 10557 3893 10560
rect 3927 10557 3939 10591
rect 3881 10551 3939 10557
rect 5350 10548 5356 10600
rect 5408 10592 5414 10600
rect 5408 10564 5580 10592
rect 5408 10548 5414 10564
rect 3142 10520 3148 10532
rect 2898 10492 3148 10520
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 3421 10523 3479 10529
rect 3421 10489 3433 10523
rect 3467 10489 3479 10523
rect 3421 10483 3479 10489
rect 4249 10523 4307 10529
rect 4249 10489 4261 10523
rect 4295 10520 4307 10523
rect 4522 10520 4528 10532
rect 4295 10492 4528 10520
rect 4295 10489 4307 10492
rect 4249 10483 4307 10489
rect 3436 10452 3464 10483
rect 4522 10480 4528 10492
rect 4580 10480 4586 10532
rect 5552 10520 5580 10564
rect 5736 10588 5764 10764
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 5960 10764 9352 10792
rect 5960 10752 5966 10764
rect 8754 10724 8760 10736
rect 8715 10696 8760 10724
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 5994 10656 6000 10668
rect 5955 10628 6000 10656
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 7006 10656 7012 10668
rect 6135 10628 7012 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 9324 10665 9352 10764
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 6454 10588 6460 10600
rect 5736 10560 6460 10588
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 9214 10588 9220 10600
rect 7975 10560 9220 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9548 10560 9597 10588
rect 9548 10548 9554 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 10042 10588 10048 10600
rect 10003 10560 10048 10588
rect 9585 10551 9643 10557
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 5994 10520 6000 10532
rect 5552 10492 6000 10520
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 7466 10480 7472 10532
rect 7524 10480 7530 10532
rect 8493 10523 8551 10529
rect 8493 10489 8505 10523
rect 8539 10520 8551 10523
rect 9508 10520 9536 10548
rect 9766 10520 9772 10532
rect 8539 10492 9536 10520
rect 9727 10492 9772 10520
rect 8539 10489 8551 10492
rect 8493 10483 8551 10489
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 8386 10452 8392 10464
rect 3436 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 920 10362 10396 10384
rect 920 10310 5066 10362
rect 5118 10310 5130 10362
rect 5182 10310 5194 10362
rect 5246 10310 5258 10362
rect 5310 10310 5322 10362
rect 5374 10310 10396 10362
rect 920 10288 10396 10310
rect 6730 10248 6736 10260
rect 3436 10220 6736 10248
rect 1670 10180 1676 10192
rect 1631 10152 1676 10180
rect 1670 10140 1676 10152
rect 1728 10140 1734 10192
rect 3142 10180 3148 10192
rect 2898 10152 3148 10180
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 3436 10189 3464 10220
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 10042 10248 10048 10260
rect 7248 10220 10048 10248
rect 7248 10208 7254 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10149 3479 10183
rect 3421 10143 3479 10149
rect 4246 10140 4252 10192
rect 4304 10140 4310 10192
rect 5074 10140 5080 10192
rect 5132 10180 5138 10192
rect 5902 10180 5908 10192
rect 5132 10152 5908 10180
rect 5132 10140 5138 10152
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 6454 10180 6460 10192
rect 6328 10152 6460 10180
rect 6328 10140 6334 10152
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 4948 10084 5365 10112
rect 4948 10072 4954 10084
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 6932 10112 6960 10208
rect 8294 10140 8300 10192
rect 8352 10140 8358 10192
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 8628 10152 8984 10180
rect 8628 10140 8634 10152
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 6932 10084 7389 10112
rect 5353 10075 5411 10081
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 8846 10112 8852 10124
rect 8807 10084 8852 10112
rect 7377 10075 7435 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 8956 10112 8984 10152
rect 9214 10140 9220 10192
rect 9272 10180 9278 10192
rect 9953 10183 10011 10189
rect 9953 10180 9965 10183
rect 9272 10152 9965 10180
rect 9272 10140 9278 10152
rect 9953 10149 9965 10152
rect 9999 10149 10011 10183
rect 9953 10143 10011 10149
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 8956 10084 9597 10112
rect 9585 10081 9597 10084
rect 9631 10081 9643 10115
rect 9585 10075 9643 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10044 3571 10047
rect 3786 10044 3792 10056
rect 3559 10016 3792 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 4154 10044 4160 10056
rect 3927 10016 4160 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 6270 10044 6276 10056
rect 6231 10016 6276 10044
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 7009 10007 7067 10013
rect 8864 10016 9781 10044
rect 7024 9976 7052 10007
rect 4816 9948 7052 9976
rect 1305 9911 1363 9917
rect 1305 9877 1317 9911
rect 1351 9908 1363 9911
rect 3878 9908 3884 9920
rect 1351 9880 3884 9908
rect 1351 9877 1363 9880
rect 1305 9871 1363 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4816 9908 4844 9948
rect 4580 9880 4844 9908
rect 5917 9911 5975 9917
rect 4580 9868 4586 9880
rect 5917 9877 5929 9911
rect 5963 9908 5975 9911
rect 7926 9908 7932 9920
rect 5963 9880 7932 9908
rect 5963 9877 5975 9880
rect 5917 9871 5975 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 8864 9908 8892 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 8168 9880 8892 9908
rect 8168 9868 8174 9880
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9409 9911 9467 9917
rect 9409 9908 9421 9911
rect 9180 9880 9421 9908
rect 9180 9868 9186 9880
rect 9409 9877 9421 9880
rect 9455 9877 9467 9911
rect 9409 9871 9467 9877
rect 920 9818 10396 9840
rect 920 9766 2566 9818
rect 2618 9766 2630 9818
rect 2682 9766 2694 9818
rect 2746 9766 2758 9818
rect 2810 9766 2822 9818
rect 2874 9766 7566 9818
rect 7618 9766 7630 9818
rect 7682 9766 7694 9818
rect 7746 9766 7758 9818
rect 7810 9766 7822 9818
rect 7874 9766 10396 9818
rect 920 9744 10396 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 5074 9704 5080 9716
rect 3476 9676 5080 9704
rect 3476 9664 3482 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 5408 9676 5672 9704
rect 5408 9664 5414 9676
rect 5644 9636 5672 9676
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6745 9707 6803 9713
rect 6052 9676 6500 9704
rect 6052 9664 6058 9676
rect 5902 9636 5908 9648
rect 3252 9608 4476 9636
rect 5644 9608 5908 9636
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 3252 9568 3280 9608
rect 3418 9568 3424 9580
rect 1719 9540 3280 9568
rect 3379 9540 3424 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4338 9568 4344 9580
rect 4299 9540 4344 9568
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4448 9568 4476 9608
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4448 9540 4721 9568
rect 4709 9537 4721 9540
rect 4755 9568 4767 9571
rect 5350 9568 5356 9580
rect 4755 9540 5356 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3660 9472 4169 9500
rect 3660 9460 3666 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 5994 9500 6000 9512
rect 5776 9472 6000 9500
rect 5776 9460 5782 9472
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6178 9500 6184 9512
rect 6139 9472 6184 9500
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6472 9500 6500 9676
rect 6745 9673 6757 9707
rect 6791 9704 6803 9707
rect 6791 9676 8524 9704
rect 6791 9673 6803 9676
rect 6745 9667 6803 9673
rect 8386 9636 8392 9648
rect 8220 9608 8392 9636
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 8220 9577 8248 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 8496 9636 8524 9676
rect 9950 9636 9956 9648
rect 8496 9608 9956 9636
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 6788 9540 7481 9568
rect 6788 9528 6794 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8312 9540 9628 9568
rect 8312 9500 8340 9540
rect 6472 9472 8340 9500
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9600 9509 9628 9540
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9732 9472 9965 9500
rect 9732 9460 9738 9472
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 1302 9432 1308 9444
rect 1263 9404 1308 9432
rect 1302 9392 1308 9404
rect 1360 9392 1366 9444
rect 3142 9432 3148 9444
rect 2898 9404 3148 9432
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 9769 9435 9827 9441
rect 9769 9432 9781 9435
rect 5842 9404 9781 9432
rect 9769 9401 9781 9404
rect 9815 9401 9827 9435
rect 9769 9395 9827 9401
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 3568 9336 3617 9364
rect 3568 9324 3574 9336
rect 3605 9333 3617 9336
rect 3651 9333 3663 9367
rect 3605 9327 3663 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 4212 9336 6929 9364
rect 4212 9324 4218 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 6917 9327 6975 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9272 9336 9413 9364
rect 9272 9324 9278 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 920 9274 10396 9296
rect 920 9222 5066 9274
rect 5118 9222 5130 9274
rect 5182 9222 5194 9274
rect 5246 9222 5258 9274
rect 5310 9222 5322 9274
rect 5374 9222 10396 9274
rect 920 9200 10396 9222
rect 5718 9160 5724 9172
rect 3988 9132 5724 9160
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 3988 9024 4016 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 8662 9160 8668 9172
rect 6604 9132 8668 9160
rect 6604 9120 6610 9132
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 9674 9160 9680 9172
rect 9416 9132 9680 9160
rect 5997 9095 6055 9101
rect 5997 9061 6009 9095
rect 6043 9092 6055 9095
rect 6270 9092 6276 9104
rect 6043 9064 6276 9092
rect 6043 9061 6055 9064
rect 5997 9055 6055 9061
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 7098 9092 7104 9104
rect 6380 9064 7104 9092
rect 5902 9024 5908 9036
rect 3927 8996 4016 9024
rect 5382 8996 5908 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 1302 8956 1308 8968
rect 1263 8928 1308 8956
rect 1302 8916 1308 8928
rect 1360 8916 1366 8968
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 3142 8956 3148 8968
rect 1452 8928 3148 8956
rect 1452 8916 1458 8928
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3200 8928 3985 8956
rect 3200 8916 3206 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 5534 8956 5540 8968
rect 4295 8928 5540 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 6380 8956 6408 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 9416 9092 9444 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9338 9064 9444 9092
rect 8202 9024 8208 9036
rect 8163 8996 8208 9024
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 6380 8928 6469 8956
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6604 8928 6653 8956
rect 6604 8916 6610 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6822 8956 6828 8968
rect 6783 8928 6828 8956
rect 6641 8919 6699 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9272 8928 9689 8956
rect 9272 8916 9278 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 9677 8919 9735 8925
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 2777 8891 2835 8897
rect 2777 8888 2789 8891
rect 2740 8860 2789 8888
rect 2740 8848 2746 8860
rect 2777 8857 2789 8860
rect 2823 8857 2835 8891
rect 2777 8851 2835 8857
rect 5258 8848 5264 8900
rect 5316 8888 5322 8900
rect 7640 8891 7698 8897
rect 7640 8888 7652 8891
rect 5316 8860 6408 8888
rect 5316 8848 5322 8860
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1728 8792 1869 8820
rect 1728 8780 1734 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 6273 8823 6331 8829
rect 6273 8820 6285 8823
rect 6144 8792 6285 8820
rect 6144 8780 6150 8792
rect 6273 8789 6285 8792
rect 6319 8789 6331 8823
rect 6380 8820 6408 8860
rect 6840 8860 7652 8888
rect 6840 8820 6868 8860
rect 7640 8857 7652 8860
rect 7686 8857 7698 8891
rect 7640 8851 7698 8857
rect 6380 8792 6868 8820
rect 6273 8783 6331 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 7156 8792 7389 8820
rect 7156 8780 7162 8792
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 920 8730 10396 8752
rect 920 8678 2566 8730
rect 2618 8678 2630 8730
rect 2682 8678 2694 8730
rect 2746 8678 2758 8730
rect 2810 8678 2822 8730
rect 2874 8678 7566 8730
rect 7618 8678 7630 8730
rect 7682 8678 7694 8730
rect 7746 8678 7758 8730
rect 7810 8678 7822 8730
rect 7874 8678 10396 8730
rect 920 8656 10396 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 6178 8616 6184 8628
rect 1627 8588 6184 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 6788 8588 9689 8616
rect 6788 8576 6794 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 2133 8551 2191 8557
rect 2133 8517 2145 8551
rect 2179 8548 2191 8551
rect 3418 8548 3424 8560
rect 2179 8520 3424 8548
rect 2179 8517 2191 8520
rect 2133 8511 2191 8517
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 5997 8551 6055 8557
rect 5997 8517 6009 8551
rect 6043 8548 6055 8551
rect 6270 8548 6276 8560
rect 6043 8520 6276 8548
rect 6043 8517 6055 8520
rect 5997 8511 6055 8517
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 7742 8508 7748 8560
rect 7800 8548 7806 8560
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 7800 8520 8493 8548
rect 7800 8508 7806 8520
rect 8481 8517 8493 8520
rect 8527 8517 8539 8551
rect 8481 8511 8539 8517
rect 1213 8483 1271 8489
rect 1213 8449 1225 8483
rect 1259 8480 1271 8483
rect 1486 8480 1492 8492
rect 1259 8452 1492 8480
rect 1259 8449 1271 8452
rect 1213 8443 1271 8449
rect 1486 8440 1492 8452
rect 1544 8480 1550 8492
rect 2774 8480 2780 8492
rect 1544 8452 2780 8480
rect 1544 8440 1550 8452
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3602 8480 3608 8492
rect 3563 8452 3608 8480
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 4212 8452 5365 8480
rect 4212 8440 4218 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5353 8443 5411 8449
rect 5644 8452 6377 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2038 8412 2044 8424
rect 1443 8384 2044 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2038 8372 2044 8384
rect 2096 8412 2102 8424
rect 3252 8412 3280 8440
rect 5644 8424 5672 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7098 8480 7104 8492
rect 6687 8452 7104 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 7098 8440 7104 8452
rect 7156 8480 7162 8492
rect 7650 8480 7656 8492
rect 7156 8452 7656 8480
rect 7156 8440 7162 8452
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8754 8480 8760 8492
rect 8435 8452 8760 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 8996 8452 9996 8480
rect 8996 8440 9002 8452
rect 2096 8384 3280 8412
rect 3421 8415 3479 8421
rect 2096 8372 2102 8384
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 3878 8412 3884 8424
rect 3467 8384 3884 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 5905 8415 5963 8421
rect 5684 8384 5729 8412
rect 5684 8372 5690 8384
rect 5905 8381 5917 8415
rect 5951 8412 5963 8415
rect 6086 8412 6092 8424
rect 5951 8384 6092 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 9306 8412 9312 8424
rect 6236 8384 6281 8412
rect 9267 8384 9312 8412
rect 6236 8372 6242 8384
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9968 8421 9996 8452
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 5994 8344 6000 8356
rect 4922 8316 6000 8344
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 6196 8344 6224 8372
rect 7098 8344 7104 8356
rect 6196 8316 7104 8344
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 9600 8344 9628 8375
rect 8996 8316 9628 8344
rect 8996 8304 9002 8316
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 5258 8276 5264 8288
rect 3384 8248 5264 8276
rect 3384 8236 3390 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 7558 8276 7564 8288
rect 6328 8248 7564 8276
rect 6328 8236 6334 8248
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8754 8276 8760 8288
rect 8715 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 19334 8276 19340 8288
rect 18012 8248 19340 8276
rect 18012 8236 18018 8248
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 920 8186 10396 8208
rect 920 8134 5066 8186
rect 5118 8134 5130 8186
rect 5182 8134 5194 8186
rect 5246 8134 5258 8186
rect 5310 8134 5322 8186
rect 5374 8134 10396 8186
rect 920 8112 10396 8134
rect 1305 8075 1363 8081
rect 1305 8041 1317 8075
rect 1351 8072 1363 8075
rect 1351 8044 6868 8072
rect 1351 8041 1363 8044
rect 1305 8035 1363 8041
rect 1578 7964 1584 8016
rect 1636 8004 1642 8016
rect 3050 8004 3056 8016
rect 1636 7976 3056 8004
rect 1636 7964 1642 7976
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 3326 8004 3332 8016
rect 3160 7976 3332 8004
rect 3160 7945 3188 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 3510 7964 3516 8016
rect 3568 7964 3574 8016
rect 6730 8004 6736 8016
rect 5014 7976 6736 8004
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 3145 7939 3203 7945
rect 1443 7908 2774 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2590 7868 2596 7880
rect 2551 7840 2596 7868
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2746 7732 2774 7908
rect 3145 7905 3157 7939
rect 3191 7905 3203 7939
rect 3528 7936 3556 7964
rect 3881 7939 3939 7945
rect 3881 7936 3893 7939
rect 3145 7899 3203 7905
rect 3252 7908 3893 7936
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 3252 7800 3280 7908
rect 3881 7905 3893 7908
rect 3927 7905 3939 7939
rect 3881 7899 3939 7905
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 4856 7908 5365 7936
rect 4856 7896 4862 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 6052 7908 6285 7936
rect 6052 7896 6058 7908
rect 6273 7905 6285 7908
rect 6319 7936 6331 7939
rect 6546 7936 6552 7948
rect 6319 7908 6408 7936
rect 6507 7908 6552 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 3510 7868 3516 7880
rect 3471 7840 3516 7868
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 6380 7868 6408 7908
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6840 7945 6868 8044
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7282 8072 7288 8084
rect 7156 8044 7288 8072
rect 7156 8032 7162 8044
rect 7282 8032 7288 8044
rect 7340 8072 7346 8084
rect 7340 8044 9536 8072
rect 7340 8032 7346 8044
rect 7558 7964 7564 8016
rect 7616 7964 7622 8016
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 6638 7868 6644 7880
rect 6380 7840 6644 7868
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7208 7868 7236 7899
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 9508 7945 9536 8044
rect 9674 8004 9680 8016
rect 9635 7976 9680 8004
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 8168 7908 8677 7936
rect 8168 7896 8174 7908
rect 8665 7905 8677 7908
rect 8711 7905 8723 7939
rect 8665 7899 8723 7905
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 7650 7868 7656 7880
rect 7208 7840 7656 7868
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 3200 7772 3280 7800
rect 3200 7760 3206 7772
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 6086 7800 6092 7812
rect 5040 7772 6092 7800
rect 5040 7760 5046 7772
rect 6086 7760 6092 7772
rect 6144 7760 6150 7812
rect 9784 7800 9812 7831
rect 8128 7772 9812 7800
rect 5442 7732 5448 7744
rect 2746 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 5917 7735 5975 7741
rect 5917 7701 5929 7735
rect 5963 7732 5975 7735
rect 6178 7732 6184 7744
rect 5963 7704 6184 7732
rect 5963 7701 5975 7704
rect 5917 7695 5975 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6362 7732 6368 7744
rect 6323 7704 6368 7732
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 8128 7732 8156 7772
rect 6696 7704 8156 7732
rect 6696 7692 6702 7704
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9225 7735 9283 7741
rect 9225 7732 9237 7735
rect 8812 7704 9237 7732
rect 8812 7692 8818 7704
rect 9225 7701 9237 7704
rect 9271 7701 9283 7735
rect 9225 7695 9283 7701
rect 920 7642 10396 7664
rect 920 7590 2566 7642
rect 2618 7590 2630 7642
rect 2682 7590 2694 7642
rect 2746 7590 2758 7642
rect 2810 7590 2822 7642
rect 2874 7590 7566 7642
rect 7618 7590 7630 7642
rect 7682 7590 7694 7642
rect 7746 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 10396 7642
rect 920 7568 10396 7590
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 8849 7531 8907 7537
rect 3016 7500 8248 7528
rect 3016 7488 3022 7500
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1360 7364 1409 7392
rect 1360 7352 1366 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 1397 7355 1455 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3878 7392 3884 7404
rect 3467 7364 3884 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3878 7352 3884 7364
rect 3936 7392 3942 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3936 7364 4445 7392
rect 3936 7352 3942 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 6086 7392 6092 7404
rect 4755 7364 6092 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7392 6515 7395
rect 6822 7392 6828 7404
rect 6503 7364 6828 7392
rect 6503 7361 6515 7364
rect 6457 7355 6515 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7293 3755 7327
rect 3697 7287 3755 7293
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 8220 7324 8248 7500
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 10042 7528 10048 7540
rect 8895 7500 10048 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 9646 7432 9812 7460
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 9306 7392 9312 7404
rect 8619 7364 9312 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9646 7392 9674 7432
rect 9784 7401 9812 7432
rect 9416 7364 9674 7392
rect 9769 7395 9827 7401
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8220 7296 8769 7324
rect 6549 7287 6607 7293
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 9416 7324 9444 7364
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9815 7364 12434 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 9674 7324 9680 7336
rect 8757 7287 8815 7293
rect 9324 7296 9444 7324
rect 9635 7296 9680 7324
rect 3142 7256 3148 7268
rect 2714 7228 3148 7256
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3712 7256 3740 7287
rect 4706 7256 4712 7268
rect 3292 7228 3740 7256
rect 4172 7228 4712 7256
rect 3292 7216 3298 7228
rect 4172 7200 4200 7228
rect 4706 7216 4712 7228
rect 4764 7256 4770 7268
rect 4982 7256 4988 7268
rect 4764 7228 4988 7256
rect 4764 7216 4770 7228
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 5994 7256 6000 7268
rect 5934 7228 6000 7256
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 1305 7191 1363 7197
rect 1305 7157 1317 7191
rect 1351 7188 1363 7191
rect 4154 7188 4160 7200
rect 1351 7160 4160 7188
rect 1351 7157 1363 7160
rect 1305 7151 1363 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4338 7188 4344 7200
rect 4299 7160 4344 7188
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6564 7188 6592 7287
rect 9324 7268 9352 7296
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 12406 7324 12434 7364
rect 20714 7324 20720 7336
rect 12406 7296 20720 7324
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 6825 7259 6883 7265
rect 6825 7225 6837 7259
rect 6871 7225 6883 7259
rect 6825 7219 6883 7225
rect 5592 7160 6592 7188
rect 6840 7188 6868 7219
rect 7282 7216 7288 7268
rect 7340 7216 7346 7268
rect 8662 7216 8668 7268
rect 8720 7256 8726 7268
rect 9033 7259 9091 7265
rect 9033 7256 9045 7259
rect 8720 7228 9045 7256
rect 8720 7216 8726 7228
rect 9033 7225 9045 7228
rect 9079 7225 9091 7259
rect 9033 7219 9091 7225
rect 9306 7216 9312 7268
rect 9364 7216 9370 7268
rect 9490 7216 9496 7268
rect 9548 7265 9554 7268
rect 9548 7259 9597 7265
rect 9548 7225 9551 7259
rect 9585 7225 9597 7259
rect 9548 7219 9597 7225
rect 9548 7216 9554 7219
rect 9214 7188 9220 7200
rect 6840 7160 9220 7188
rect 5592 7148 5598 7160
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 920 7098 10396 7120
rect 920 7046 5066 7098
rect 5118 7046 5130 7098
rect 5182 7046 5194 7098
rect 5246 7046 5258 7098
rect 5310 7046 5322 7098
rect 5374 7046 10396 7098
rect 920 7024 10396 7046
rect 5442 6944 5448 6996
rect 5500 6984 5506 6996
rect 8386 6984 8392 6996
rect 5500 6956 8392 6984
rect 5500 6944 5506 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 9732 6956 10057 6984
rect 9732 6944 9738 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 8576 6928 8628 6934
rect 2406 6876 2412 6928
rect 2464 6876 2470 6928
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 3421 6919 3479 6925
rect 3421 6916 3433 6919
rect 3384 6888 3433 6916
rect 3384 6876 3390 6888
rect 3421 6885 3433 6888
rect 3467 6885 3479 6919
rect 3421 6879 3479 6885
rect 4798 6876 4804 6928
rect 4856 6876 4862 6928
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 6917 6919 6975 6925
rect 6917 6916 6929 6919
rect 6604 6888 6929 6916
rect 6604 6876 6610 6888
rect 6917 6885 6929 6888
rect 6963 6885 6975 6919
rect 6917 6879 6975 6885
rect 8576 6870 8628 6876
rect 1210 6848 1216 6860
rect 1171 6820 1216 6848
rect 1210 6808 1216 6820
rect 1268 6808 1274 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 5353 6851 5411 6857
rect 3559 6820 4016 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1397 6743 1455 6749
rect 1412 6644 1440 6743
rect 1670 6740 1676 6752
rect 1728 6780 1734 6792
rect 2222 6780 2228 6792
rect 1728 6752 2228 6780
rect 1728 6740 1734 6752
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3528 6752 3893 6780
rect 2682 6672 2688 6724
rect 2740 6712 2746 6724
rect 3528 6712 3556 6752
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 3988 6780 4016 6820
rect 5353 6817 5365 6851
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 4430 6780 4436 6792
rect 3988 6752 4436 6780
rect 3881 6743 3939 6749
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 2740 6684 3556 6712
rect 2740 6672 2746 6684
rect 4982 6672 4988 6724
rect 5040 6712 5046 6724
rect 5368 6712 5396 6811
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 6144 6820 6193 6848
rect 6144 6808 6150 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 8938 6848 8944 6860
rect 8899 6820 8944 6848
rect 6181 6811 6239 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9490 6848 9496 6860
rect 9180 6820 9496 6848
rect 9180 6808 9186 6820
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6733 6783 6791 6789
rect 6733 6780 6745 6783
rect 6052 6752 6745 6780
rect 6052 6740 6058 6752
rect 6733 6749 6745 6752
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 8018 6780 8024 6792
rect 7515 6752 8024 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 5040 6684 5396 6712
rect 5040 6672 5046 6684
rect 3878 6644 3884 6656
rect 1412 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 5917 6647 5975 6653
rect 5917 6613 5929 6647
rect 5963 6644 5975 6647
rect 6638 6644 6644 6656
rect 5963 6616 6644 6644
rect 5963 6613 5975 6616
rect 5917 6607 5975 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 7116 6644 7144 6743
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9364 6752 9873 6780
rect 9364 6740 9370 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 9950 6712 9956 6724
rect 9723 6684 9956 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 8478 6644 8484 6656
rect 7116 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9501 6647 9559 6653
rect 9501 6644 9513 6647
rect 9272 6616 9513 6644
rect 9272 6604 9278 6616
rect 9501 6613 9513 6616
rect 9547 6613 9559 6647
rect 9501 6607 9559 6613
rect 920 6554 10396 6576
rect 920 6502 2566 6554
rect 2618 6502 2630 6554
rect 2682 6502 2694 6554
rect 2746 6502 2758 6554
rect 2810 6502 2822 6554
rect 2874 6502 7566 6554
rect 7618 6502 7630 6554
rect 7682 6502 7694 6554
rect 7746 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 10396 6554
rect 920 6480 10396 6502
rect 7282 6400 7288 6452
rect 7340 6440 7346 6452
rect 8018 6440 8024 6452
rect 7340 6412 8024 6440
rect 7340 6400 7346 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8570 6440 8576 6452
rect 8435 6412 8576 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 1581 6375 1639 6381
rect 1581 6341 1593 6375
rect 1627 6372 1639 6375
rect 4706 6372 4712 6384
rect 1627 6344 4712 6372
rect 1627 6341 1639 6344
rect 1581 6335 1639 6341
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 6880 6344 8769 6372
rect 6880 6332 6886 6344
rect 1118 6264 1124 6316
rect 1176 6304 1182 6316
rect 1213 6307 1271 6313
rect 1213 6304 1225 6307
rect 1176 6276 1225 6304
rect 1176 6264 1182 6276
rect 1213 6273 1225 6276
rect 1259 6273 1271 6307
rect 1213 6267 1271 6273
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5534 6304 5540 6316
rect 5399 6276 5540 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6086 6304 6092 6316
rect 5859 6276 6092 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 8220 6313 8248 6344
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 9214 6372 9220 6384
rect 8757 6335 8815 6341
rect 8864 6344 9220 6372
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8386 6304 8392 6316
rect 8251 6276 8392 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 1394 6236 1400 6248
rect 1307 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 2406 6236 2412 6248
rect 1452 6208 2412 6236
rect 1452 6196 1458 6208
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3384 6208 3433 6236
rect 3384 6196 3390 6208
rect 3421 6205 3433 6208
rect 3467 6236 3479 6239
rect 3970 6236 3976 6248
rect 3467 6208 3976 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5718 6236 5724 6248
rect 5491 6208 5724 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8018 6236 8024 6248
rect 7892 6208 8024 6236
rect 7892 6196 7898 6208
rect 8018 6196 8024 6208
rect 8076 6236 8082 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8076 6208 8493 6236
rect 8076 6196 8082 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 3602 6168 3608 6180
rect 3563 6140 3608 6168
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 6362 6128 6368 6180
rect 6420 6128 6426 6180
rect 8864 6168 8892 6344
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9214 6236 9220 6248
rect 9171 6208 9220 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 9582 6236 9588 6248
rect 9539 6208 9588 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9766 6236 9772 6248
rect 9727 6208 9772 6236
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 10042 6168 10048 6180
rect 7024 6140 8892 6168
rect 10003 6140 10048 6168
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 3620 6100 3648 6128
rect 2179 6072 3648 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 7024 6100 7052 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 6880 6072 7052 6100
rect 7849 6103 7907 6109
rect 6880 6060 6886 6072
rect 7849 6069 7861 6103
rect 7895 6100 7907 6103
rect 8018 6100 8024 6112
rect 7895 6072 8024 6100
rect 7895 6069 7907 6072
rect 7849 6063 7907 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 920 6010 10396 6032
rect 920 5958 5066 6010
rect 5118 5958 5130 6010
rect 5182 5958 5194 6010
rect 5246 5958 5258 6010
rect 5310 5958 5322 6010
rect 5374 5958 10396 6010
rect 920 5936 10396 5958
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2958 5896 2964 5908
rect 2179 5868 2964 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 4982 5896 4988 5908
rect 3252 5868 4988 5896
rect 1213 5831 1271 5837
rect 1213 5797 1225 5831
rect 1259 5828 1271 5831
rect 3252 5828 3280 5868
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 7156 5868 7420 5896
rect 7156 5856 7162 5868
rect 3418 5828 3424 5840
rect 1259 5800 3280 5828
rect 3379 5800 3424 5828
rect 1259 5797 1271 5800
rect 1213 5791 1271 5797
rect 3418 5788 3424 5800
rect 3476 5788 3482 5840
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 4338 5828 4344 5840
rect 4295 5800 4344 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5258 5788 5264 5840
rect 5316 5788 5322 5840
rect 5994 5828 6000 5840
rect 5955 5800 6000 5828
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 7282 5828 7288 5840
rect 6595 5800 7288 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 3605 5763 3663 5769
rect 3605 5729 3617 5763
rect 3651 5729 3663 5763
rect 3605 5723 3663 5729
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 6454 5760 6460 5772
rect 6227 5732 6460 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 3620 5624 3648 5723
rect 6454 5720 6460 5732
rect 6512 5760 6518 5772
rect 7098 5760 7104 5772
rect 6512 5732 7104 5760
rect 6512 5720 6518 5732
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7392 5760 7420 5868
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 8444 5868 9965 5896
rect 8444 5856 8450 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 9953 5859 10011 5865
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 9125 5831 9183 5837
rect 9125 5828 9137 5831
rect 8996 5800 9137 5828
rect 8996 5788 9002 5800
rect 9125 5797 9137 5800
rect 9171 5797 9183 5831
rect 9125 5791 9183 5797
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9447 5831 9505 5837
rect 9447 5828 9459 5831
rect 9364 5800 9459 5828
rect 9364 5788 9370 5800
rect 9447 5797 9459 5800
rect 9493 5797 9505 5831
rect 9858 5828 9864 5840
rect 9819 5800 9864 5828
rect 9447 5791 9505 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 17954 5828 17960 5840
rect 11112 5800 17960 5828
rect 11112 5788 11118 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 8570 5760 8576 5772
rect 7300 5732 7420 5760
rect 8531 5732 8576 5760
rect 7300 5704 7328 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 8720 5732 8984 5760
rect 8720 5720 8726 5732
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 5902 5692 5908 5704
rect 3973 5655 4031 5661
rect 4080 5664 5908 5692
rect 4080 5624 4108 5664
rect 5902 5652 5908 5664
rect 5960 5692 5966 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 5960 5664 6377 5692
rect 5960 5652 5966 5664
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 3200 5596 4108 5624
rect 7944 5624 7972 5655
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8956 5701 8984 5732
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 9088 5732 9229 5760
rect 9088 5720 9094 5732
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8444 5664 8769 5692
rect 8444 5652 8450 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 19334 5624 19340 5636
rect 7944 5596 19340 5624
rect 3200 5584 3206 5596
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 2464 5528 3801 5556
rect 2464 5516 2470 5528
rect 3789 5525 3801 5528
rect 3835 5556 3847 5559
rect 5258 5556 5264 5568
rect 3835 5528 5264 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9490 5556 9496 5568
rect 8628 5528 9496 5556
rect 8628 5516 8634 5528
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 920 5466 10396 5488
rect 920 5414 2566 5466
rect 2618 5414 2630 5466
rect 2682 5414 2694 5466
rect 2746 5414 2758 5466
rect 2810 5414 2822 5466
rect 2874 5414 7566 5466
rect 7618 5414 7630 5466
rect 7682 5414 7694 5466
rect 7746 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 10396 5466
rect 920 5392 10396 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 3108 5256 6040 5284
rect 3108 5244 3114 5256
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3292 5188 3341 5216
rect 3292 5176 3298 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 5442 5216 5448 5228
rect 3476 5188 3832 5216
rect 5403 5188 5448 5216
rect 3476 5176 3482 5188
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3804 5157 3832 5188
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 6012 5157 6040 5256
rect 6730 5216 6736 5228
rect 6691 5188 6736 5216
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 12434 5216 12440 5228
rect 9447 5188 12440 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3200 5120 3525 5148
rect 3200 5108 3206 5120
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 5997 5151 6055 5157
rect 5997 5117 6009 5151
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8110 5148 8116 5160
rect 8067 5120 8116 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 3697 5083 3755 5089
rect 3697 5049 3709 5083
rect 3743 5080 3755 5083
rect 5902 5080 5908 5092
rect 3743 5052 5908 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 6012 5080 6040 5111
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 10042 5148 10048 5160
rect 10003 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 9766 5080 9772 5092
rect 6012 5052 9772 5080
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 7742 5012 7748 5024
rect 6144 4984 7748 5012
rect 6144 4972 6150 4984
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 3036 4922 10396 4944
rect 3036 4870 5066 4922
rect 5118 4870 5130 4922
rect 5182 4870 5194 4922
rect 5246 4870 5258 4922
rect 5310 4870 5322 4922
rect 5374 4870 10396 4922
rect 3036 4848 10396 4870
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4672 4780 6960 4808
rect 4672 4768 4678 4780
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 3142 4740 3148 4752
rect 1636 4712 3148 4740
rect 1636 4700 1642 4712
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3436 4740 3464 4768
rect 3973 4743 4031 4749
rect 3436 4712 3832 4740
rect 2038 4632 2044 4684
rect 2096 4672 2102 4684
rect 3804 4681 3832 4712
rect 3973 4709 3985 4743
rect 4019 4740 4031 4743
rect 4246 4740 4252 4752
rect 4019 4712 4252 4740
rect 4019 4709 4031 4712
rect 3973 4703 4031 4709
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 4338 4700 4344 4752
rect 4396 4700 4402 4752
rect 4982 4700 4988 4752
rect 5040 4740 5046 4752
rect 5040 4712 5106 4740
rect 5040 4700 5046 4712
rect 3605 4675 3663 4681
rect 3605 4672 3617 4675
rect 2096 4644 3617 4672
rect 2096 4632 2102 4644
rect 3605 4641 3617 4644
rect 3651 4641 3663 4675
rect 3605 4635 3663 4641
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4641 3847 4675
rect 4356 4672 4384 4700
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 4356 4644 4721 4672
rect 3789 4635 3847 4641
rect 4709 4641 4721 4644
rect 4755 4641 4767 4675
rect 4709 4635 4767 4641
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5960 4644 6193 4672
rect 5960 4632 5966 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 4065 4607 4123 4613
rect 2004 4576 2774 4604
rect 2004 4564 2010 4576
rect 2746 4468 2774 4576
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4080 4468 4108 4567
rect 4246 4468 4252 4480
rect 2746 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4356 4468 4384 4567
rect 6086 4468 6092 4480
rect 4356 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6741 4471 6799 4477
rect 6741 4468 6753 4471
rect 6512 4440 6753 4468
rect 6512 4428 6518 4440
rect 6741 4437 6753 4440
rect 6787 4437 6799 4471
rect 6932 4468 6960 4780
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7156 4780 7573 4808
rect 7156 4768 7162 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7561 4771 7619 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 9272 4780 9597 4808
rect 9272 4768 9278 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 8202 4740 8208 4752
rect 8159 4712 8208 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 9122 4740 9128 4752
rect 8312 4712 8984 4740
rect 9083 4712 9128 4740
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7098 4672 7104 4684
rect 7055 4644 7104 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7098 4632 7104 4644
rect 7156 4672 7162 4684
rect 7208 4672 7328 4674
rect 8312 4672 8340 4712
rect 7156 4646 8340 4672
rect 7156 4644 7236 4646
rect 7300 4644 8340 4646
rect 7156 4632 7162 4644
rect 8220 4616 8248 4644
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 8444 4644 8677 4672
rect 8444 4632 8450 4644
rect 8665 4641 8677 4644
rect 8711 4672 8723 4675
rect 8754 4672 8760 4684
rect 8711 4644 8760 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 8956 4681 8984 4712
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 10008 4644 10057 4672
rect 10008 4632 10014 4644
rect 10045 4641 10057 4644
rect 10091 4672 10103 4675
rect 10134 4672 10140 4684
rect 10091 4644 10140 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7466 4604 7472 4616
rect 7423 4576 7472 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7300 4536 7328 4567
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7892 4576 7941 4604
rect 7892 4564 7898 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8202 4564 8208 4616
rect 8260 4564 8266 4616
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8352 4576 8585 4604
rect 8352 4564 8358 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 8478 4536 8484 4548
rect 7300 4508 8484 4536
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 9030 4496 9036 4548
rect 9088 4536 9094 4548
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 9088 4508 9413 4536
rect 9088 4496 9094 4508
rect 9401 4505 9413 4508
rect 9447 4505 9459 4539
rect 9401 4499 9459 4505
rect 9861 4471 9919 4477
rect 9861 4468 9873 4471
rect 6932 4440 9873 4468
rect 6741 4431 6799 4437
rect 9861 4437 9873 4440
rect 9907 4437 9919 4471
rect 9861 4431 9919 4437
rect 3036 4378 10396 4400
rect 3036 4326 7566 4378
rect 7618 4326 7630 4378
rect 7682 4326 7694 4378
rect 7746 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 10396 4378
rect 3036 4304 10396 4326
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4614 4264 4620 4276
rect 4212 4236 4620 4264
rect 4212 4224 4218 4236
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8478 4264 8484 4276
rect 8352 4236 8484 4264
rect 8352 4224 8358 4236
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 5537 4199 5595 4205
rect 5537 4196 5549 4199
rect 5000 4168 5549 4196
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5000 4128 5028 4168
rect 5537 4165 5549 4168
rect 5583 4165 5595 4199
rect 5537 4159 5595 4165
rect 4948 4100 5028 4128
rect 5077 4131 5135 4137
rect 4948 4088 4954 4100
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 11054 4128 11060 4140
rect 5123 4100 11060 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 16574 4128 16580 4140
rect 16546 4088 16580 4128
rect 16632 4088 16638 4140
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 3016 4032 3341 4060
rect 3016 4020 3022 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 4304 4032 5181 4060
rect 4304 4020 4310 4032
rect 4908 4004 4936 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 6178 4060 6184 4072
rect 6139 4032 6184 4060
rect 5997 4023 6055 4029
rect 4890 3952 4896 4004
rect 4948 3952 4954 4004
rect 3418 3884 3424 3936
rect 3476 3924 3482 3936
rect 5368 3924 5396 4023
rect 6012 3992 6040 4023
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7984 4032 8125 4060
rect 7984 4020 7990 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10686 4060 10692 4072
rect 10091 4032 10692 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 6362 3992 6368 4004
rect 6012 3964 6368 3992
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 16546 3992 16574 4088
rect 8067 3964 16574 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 3476 3896 5396 3924
rect 5813 3927 5871 3933
rect 3476 3884 3482 3896
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 7926 3924 7932 3936
rect 5859 3896 7932 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 3036 3834 10396 3856
rect 3036 3782 5066 3834
rect 5118 3782 5130 3834
rect 5182 3782 5194 3834
rect 5246 3782 5258 3834
rect 5310 3782 5322 3834
rect 5374 3782 10396 3834
rect 3036 3760 10396 3782
rect 3326 3720 3332 3732
rect 3287 3692 3332 3720
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 8846 3720 8852 3732
rect 5644 3692 8708 3720
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 3326 3584 3332 3596
rect 2740 3556 3332 3584
rect 2740 3544 2746 3556
rect 3326 3544 3332 3556
rect 3384 3584 3390 3596
rect 3605 3587 3663 3593
rect 3605 3584 3617 3587
rect 3384 3556 3617 3584
rect 3384 3544 3390 3556
rect 3605 3553 3617 3556
rect 3651 3553 3663 3587
rect 3605 3547 3663 3553
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3418 3516 3424 3528
rect 3292 3488 3424 3516
rect 3292 3476 3298 3488
rect 3418 3476 3424 3488
rect 3476 3516 3482 3528
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3476 3488 3893 3516
rect 3476 3476 3482 3488
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4982 3516 4988 3528
rect 4019 3488 4988 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5350 3516 5356 3528
rect 5311 3488 5356 3516
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 5644 3448 5672 3692
rect 6822 3652 6828 3664
rect 5736 3624 6828 3652
rect 5736 3593 5764 3624
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 5868 3556 6193 3584
rect 5868 3544 5874 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 8680 3584 8708 3692
rect 8772 3692 8852 3720
rect 8772 3661 8800 3692
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3621 8815 3655
rect 8757 3615 8815 3621
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 10318 3652 10324 3664
rect 9723 3624 10324 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 16666 3652 16672 3664
rect 16546 3624 16672 3652
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8260 3556 8616 3584
rect 8680 3556 8861 3584
rect 8260 3544 8266 3556
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8588 3525 8616 3556
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 9030 3584 9036 3596
rect 8991 3556 9036 3584
rect 8849 3547 8907 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9824 3556 9873 3584
rect 9824 3544 9830 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 9582 3516 9588 3528
rect 9543 3488 9588 3516
rect 8573 3479 8631 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 2740 3420 5672 3448
rect 8113 3451 8171 3457
rect 2740 3408 2746 3420
rect 8113 3417 8125 3451
rect 8159 3448 8171 3451
rect 16546 3448 16574 3624
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 8159 3420 16574 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 4764 3352 9229 3380
rect 4764 3340 4770 3352
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 9217 3343 9275 3349
rect 3036 3290 10396 3312
rect 3036 3238 7566 3290
rect 7618 3238 7630 3290
rect 7682 3238 7694 3290
rect 7746 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 10396 3290
rect 3036 3216 10396 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4488 3148 5273 3176
rect 4488 3136 4494 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 5813 3179 5871 3185
rect 5813 3176 5825 3179
rect 5776 3148 5825 3176
rect 5776 3136 5782 3148
rect 5813 3145 5825 3148
rect 5859 3145 5871 3179
rect 6086 3176 6092 3188
rect 6047 3148 6092 3176
rect 5813 3139 5871 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7374 3176 7380 3188
rect 7331 3148 7380 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 6641 3111 6699 3117
rect 6641 3077 6653 3111
rect 6687 3108 6699 3111
rect 7190 3108 7196 3120
rect 6687 3080 7196 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 6914 3040 6920 3052
rect 5123 3012 6920 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5040 2944 5365 2972
rect 5040 2932 5046 2944
rect 5353 2941 5365 2944
rect 5399 2972 5411 2975
rect 5442 2972 5448 2984
rect 5399 2944 5448 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5442 2932 5448 2944
rect 5500 2972 5506 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 5500 2944 5917 2972
rect 5500 2932 5506 2944
rect 5905 2941 5917 2944
rect 5951 2972 5963 2975
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 5951 2944 6193 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6181 2941 6193 2944
rect 6227 2941 6239 2975
rect 6181 2935 6239 2941
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 7064 2944 7113 2972
rect 7064 2932 7070 2944
rect 7101 2941 7113 2944
rect 7147 2972 7159 2975
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 7147 2944 7205 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 5534 2904 5540 2916
rect 3375 2876 5540 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5994 2864 6000 2916
rect 6052 2864 6058 2916
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4890 2836 4896 2848
rect 4304 2808 4896 2836
rect 4304 2796 4310 2808
rect 4890 2796 4896 2808
rect 4948 2836 4954 2848
rect 5445 2839 5503 2845
rect 5445 2836 5457 2839
rect 4948 2808 5457 2836
rect 4948 2796 4954 2808
rect 5445 2805 5457 2808
rect 5491 2805 5503 2839
rect 6012 2836 6040 2864
rect 6733 2839 6791 2845
rect 6733 2836 6745 2839
rect 6012 2808 6745 2836
rect 5445 2799 5503 2805
rect 6733 2805 6745 2808
rect 6779 2805 6791 2839
rect 6733 2799 6791 2805
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 9490 2836 9496 2848
rect 8260 2808 9496 2836
rect 8260 2796 8266 2808
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 3036 2746 10396 2768
rect 3036 2694 5066 2746
rect 5118 2694 5130 2746
rect 5182 2694 5194 2746
rect 5246 2694 5258 2746
rect 5310 2694 5322 2746
rect 5374 2694 10396 2746
rect 3036 2672 10396 2694
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 6972 2604 8953 2632
rect 6972 2592 6978 2604
rect 8941 2601 8953 2604
rect 8987 2632 8999 2635
rect 9214 2632 9220 2644
rect 8987 2604 9220 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9490 2592 9496 2644
rect 9548 2632 9554 2644
rect 9548 2604 9812 2632
rect 9548 2592 9554 2604
rect 7098 2564 7104 2576
rect 4816 2536 7104 2564
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 3605 2499 3663 2505
rect 3605 2496 3617 2499
rect 3384 2468 3617 2496
rect 3384 2456 3390 2468
rect 3605 2465 3617 2468
rect 3651 2465 3663 2499
rect 4338 2496 4344 2508
rect 3605 2459 3663 2465
rect 3896 2468 4344 2496
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3896 2437 3924 2468
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 3200 2400 3893 2428
rect 3200 2388 3206 2400
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4706 2428 4712 2440
rect 4019 2400 4712 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 4816 2360 4844 2536
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7926 2524 7932 2576
rect 7984 2564 7990 2576
rect 7984 2536 8800 2564
rect 7984 2524 7990 2536
rect 6089 2499 6147 2505
rect 6089 2465 6101 2499
rect 6135 2496 6147 2499
rect 8113 2499 8171 2505
rect 6135 2468 8064 2496
rect 6135 2465 6147 2468
rect 6089 2459 6147 2465
rect 5442 2428 5448 2440
rect 5403 2400 5448 2428
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 8036 2428 8064 2468
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8570 2496 8576 2508
rect 8159 2468 8576 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8772 2505 8800 2536
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 9456 2536 9597 2564
rect 9456 2524 9462 2536
rect 9585 2533 9597 2536
rect 9631 2533 9643 2567
rect 9585 2527 9643 2533
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2465 8723 2499
rect 8665 2459 8723 2465
rect 8757 2499 8815 2505
rect 8757 2465 8769 2499
rect 8803 2465 8815 2499
rect 9490 2496 9496 2508
rect 9451 2468 9496 2496
rect 8757 2459 8815 2465
rect 8294 2428 8300 2440
rect 8036 2400 8300 2428
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8680 2428 8708 2459
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9784 2505 9812 2604
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 9030 2428 9036 2440
rect 8680 2400 9036 2428
rect 9030 2388 9036 2400
rect 9088 2428 9094 2440
rect 9088 2400 9352 2428
rect 9088 2388 9094 2400
rect 2976 2332 4844 2360
rect 2976 2088 3004 2332
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 8846 2360 8852 2372
rect 5868 2332 8852 2360
rect 5868 2320 5874 2332
rect 8846 2320 8852 2332
rect 8904 2360 8910 2372
rect 9324 2369 9352 2400
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9640 2400 9965 2428
rect 9640 2388 9646 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 9309 2363 9367 2369
rect 8904 2332 9260 2360
rect 8904 2320 8910 2332
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 6086 2252 6092 2304
rect 6144 2292 6150 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 6144 2264 8493 2292
rect 6144 2252 6150 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 9232 2292 9260 2332
rect 9309 2329 9321 2363
rect 9355 2329 9367 2363
rect 9309 2323 9367 2329
rect 9490 2320 9496 2372
rect 9548 2360 9554 2372
rect 16942 2360 16948 2372
rect 9548 2332 16948 2360
rect 9548 2320 9554 2332
rect 16942 2320 16948 2332
rect 17000 2320 17006 2372
rect 9582 2292 9588 2304
rect 9232 2264 9588 2292
rect 8481 2255 8539 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 3036 2202 10396 2224
rect 3036 2150 7566 2202
rect 7618 2150 7630 2202
rect 7682 2150 7694 2202
rect 7746 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 10396 2202
rect 3036 2128 10396 2150
rect 3513 2091 3571 2097
rect 3513 2088 3525 2091
rect 2976 2060 3525 2088
rect 3513 2057 3525 2060
rect 3559 2057 3571 2091
rect 3786 2088 3792 2100
rect 3747 2060 3792 2088
rect 3513 2051 3571 2057
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 4062 2088 4068 2100
rect 4023 2060 4068 2088
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 4341 2091 4399 2097
rect 4341 2057 4353 2091
rect 4387 2088 4399 2091
rect 4430 2088 4436 2100
rect 4387 2060 4436 2088
rect 4387 2057 4399 2060
rect 4341 2051 4399 2057
rect 4430 2048 4436 2060
rect 4488 2048 4494 2100
rect 4614 2048 4620 2100
rect 4672 2088 4678 2100
rect 4893 2091 4951 2097
rect 4893 2088 4905 2091
rect 4672 2060 4905 2088
rect 4672 2048 4678 2060
rect 4893 2057 4905 2060
rect 4939 2057 4951 2091
rect 5810 2088 5816 2100
rect 5771 2060 5816 2088
rect 4893 2051 4951 2057
rect 5810 2048 5816 2060
rect 5868 2048 5874 2100
rect 5997 2091 6055 2097
rect 5997 2057 6009 2091
rect 6043 2088 6055 2091
rect 7282 2088 7288 2100
rect 6043 2060 7288 2088
rect 6043 2057 6055 2060
rect 5997 2051 6055 2057
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 4525 2023 4583 2029
rect 4525 2020 4537 2023
rect 3476 1992 4537 2020
rect 3476 1980 3482 1992
rect 4525 1989 4537 1992
rect 4571 1989 4583 2023
rect 4525 1983 4583 1989
rect 5537 2023 5595 2029
rect 5537 1989 5549 2023
rect 5583 2020 5595 2023
rect 9490 2020 9496 2032
rect 5583 1992 9496 2020
rect 5583 1989 5595 1992
rect 5537 1983 5595 1989
rect 9490 1980 9496 1992
rect 9548 1980 9554 2032
rect 2958 1912 2964 1964
rect 3016 1952 3022 1964
rect 3016 1924 3924 1952
rect 3016 1912 3022 1924
rect 2682 1844 2688 1896
rect 2740 1884 2746 1896
rect 3896 1893 3924 1924
rect 4338 1912 4344 1964
rect 4396 1952 4402 1964
rect 4709 1955 4767 1961
rect 4709 1952 4721 1955
rect 4396 1924 4721 1952
rect 4396 1912 4402 1924
rect 4709 1921 4721 1924
rect 4755 1952 4767 1955
rect 5077 1955 5135 1961
rect 5077 1952 5089 1955
rect 4755 1924 5089 1952
rect 4755 1921 4767 1924
rect 4709 1915 4767 1921
rect 5077 1921 5089 1924
rect 5123 1921 5135 1955
rect 7006 1952 7012 1964
rect 5077 1915 5135 1921
rect 6288 1924 7012 1952
rect 3329 1887 3387 1893
rect 3329 1884 3341 1887
rect 2740 1856 3341 1884
rect 2740 1844 2746 1856
rect 3329 1853 3341 1856
rect 3375 1853 3387 1887
rect 3329 1847 3387 1853
rect 3881 1887 3939 1893
rect 3881 1853 3893 1887
rect 3927 1884 3939 1887
rect 4157 1887 4215 1893
rect 4157 1884 4169 1887
rect 3927 1856 4169 1884
rect 3927 1853 3939 1856
rect 3881 1847 3939 1853
rect 4157 1853 4169 1856
rect 4203 1884 4215 1887
rect 4249 1887 4307 1893
rect 4249 1884 4261 1887
rect 4203 1856 4261 1884
rect 4203 1853 4215 1856
rect 4157 1847 4215 1853
rect 4249 1853 4261 1856
rect 4295 1884 4307 1887
rect 6288 1884 6316 1924
rect 7006 1912 7012 1924
rect 7064 1912 7070 1964
rect 9401 1955 9459 1961
rect 9401 1921 9413 1955
rect 9447 1952 9459 1955
rect 9447 1924 16574 1952
rect 9447 1921 9459 1924
rect 9401 1915 9459 1921
rect 6454 1884 6460 1896
rect 4295 1856 6316 1884
rect 6415 1856 6460 1884
rect 4295 1853 4307 1856
rect 4249 1847 4307 1853
rect 3344 1748 3372 1847
rect 6454 1844 6460 1856
rect 6512 1844 6518 1896
rect 9858 1884 9864 1896
rect 9819 1856 9864 1884
rect 9858 1844 9864 1856
rect 9916 1844 9922 1896
rect 8021 1819 8079 1825
rect 8021 1785 8033 1819
rect 8067 1816 8079 1819
rect 16546 1816 16574 1924
rect 16850 1816 16856 1828
rect 8067 1788 12664 1816
rect 16546 1788 16856 1816
rect 8067 1785 8079 1788
rect 8021 1779 8079 1785
rect 4154 1748 4160 1760
rect 3344 1720 4160 1748
rect 4154 1708 4160 1720
rect 4212 1748 4218 1760
rect 5261 1751 5319 1757
rect 5261 1748 5273 1751
rect 4212 1720 5273 1748
rect 4212 1708 4218 1720
rect 5261 1717 5273 1720
rect 5307 1717 5319 1751
rect 12636 1748 12664 1788
rect 16850 1776 16856 1788
rect 16908 1776 16914 1828
rect 16666 1748 16672 1760
rect 12636 1720 16672 1748
rect 5261 1711 5319 1717
rect 16666 1708 16672 1720
rect 16724 1708 16730 1760
rect 3036 1658 10396 1680
rect 3036 1606 5066 1658
rect 5118 1606 5130 1658
rect 5182 1606 5194 1658
rect 5246 1606 5258 1658
rect 5310 1606 5322 1658
rect 5374 1606 10396 1658
rect 3036 1584 10396 1606
rect 3421 1547 3479 1553
rect 3421 1513 3433 1547
rect 3467 1544 3479 1547
rect 3510 1544 3516 1556
rect 3467 1516 3516 1544
rect 3467 1513 3479 1516
rect 3421 1507 3479 1513
rect 3510 1504 3516 1516
rect 3568 1504 3574 1556
rect 3694 1544 3700 1556
rect 3655 1516 3700 1544
rect 3694 1504 3700 1516
rect 3752 1504 3758 1556
rect 6822 1504 6828 1556
rect 6880 1544 6886 1556
rect 7009 1547 7067 1553
rect 7009 1544 7021 1547
rect 6880 1516 7021 1544
rect 6880 1504 6886 1516
rect 7009 1513 7021 1516
rect 7055 1513 7067 1547
rect 7009 1507 7067 1513
rect 9217 1547 9275 1553
rect 9217 1513 9229 1547
rect 9263 1544 9275 1547
rect 9306 1544 9312 1556
rect 9263 1516 9312 1544
rect 9263 1513 9275 1516
rect 9217 1507 9275 1513
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 9766 1504 9772 1556
rect 9824 1544 9830 1556
rect 9953 1547 10011 1553
rect 9953 1544 9965 1547
rect 9824 1516 9965 1544
rect 9824 1504 9830 1516
rect 9953 1513 9965 1516
rect 9999 1513 10011 1547
rect 9953 1507 10011 1513
rect 4982 1476 4988 1488
rect 3344 1448 4988 1476
rect 3344 1417 3372 1448
rect 4982 1436 4988 1448
rect 5040 1436 5046 1488
rect 3329 1411 3387 1417
rect 3329 1377 3341 1411
rect 3375 1377 3387 1411
rect 3329 1371 3387 1377
rect 3789 1411 3847 1417
rect 3789 1377 3801 1411
rect 3835 1408 3847 1411
rect 3878 1408 3884 1420
rect 3835 1380 3884 1408
rect 3835 1377 3847 1380
rect 3789 1371 3847 1377
rect 3878 1368 3884 1380
rect 3936 1368 3942 1420
rect 6086 1408 6092 1420
rect 6047 1380 6092 1408
rect 6086 1368 6092 1380
rect 6144 1368 6150 1420
rect 8018 1408 8024 1420
rect 7979 1380 8024 1408
rect 8018 1368 8024 1380
rect 8076 1368 8082 1420
rect 8570 1368 8576 1420
rect 8628 1408 8634 1420
rect 9030 1408 9036 1420
rect 8628 1380 9036 1408
rect 8628 1368 8634 1380
rect 9030 1368 9036 1380
rect 9088 1368 9094 1420
rect 9214 1368 9220 1420
rect 9272 1408 9278 1420
rect 9401 1411 9459 1417
rect 9401 1408 9413 1411
rect 9272 1380 9413 1408
rect 9272 1368 9278 1380
rect 9401 1377 9413 1380
rect 9447 1377 9459 1411
rect 9769 1411 9827 1417
rect 9769 1408 9781 1411
rect 9401 1371 9459 1377
rect 9600 1380 9781 1408
rect 3973 1343 4031 1349
rect 3973 1309 3985 1343
rect 4019 1340 4031 1343
rect 4246 1340 4252 1352
rect 4019 1312 4252 1340
rect 4019 1309 4031 1312
rect 3973 1303 4031 1309
rect 4246 1300 4252 1312
rect 4304 1300 4310 1352
rect 5442 1340 5448 1352
rect 5403 1312 5448 1340
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 8389 1343 8447 1349
rect 8389 1309 8401 1343
rect 8435 1340 8447 1343
rect 8478 1340 8484 1352
rect 8435 1312 8484 1340
rect 8435 1309 8447 1312
rect 8389 1303 8447 1309
rect 8478 1300 8484 1312
rect 8536 1300 8542 1352
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 8849 1343 8907 1349
rect 8849 1340 8861 1343
rect 8720 1312 8861 1340
rect 8720 1300 8726 1312
rect 8849 1309 8861 1312
rect 8895 1340 8907 1343
rect 9600 1340 9628 1380
rect 9769 1377 9781 1380
rect 9815 1377 9827 1411
rect 9769 1371 9827 1377
rect 8895 1312 9628 1340
rect 8895 1309 8907 1312
rect 8849 1303 8907 1309
rect 8938 1272 8944 1284
rect 8680 1244 8944 1272
rect 5258 1164 5264 1216
rect 5316 1204 5322 1216
rect 8680 1213 8708 1244
rect 8938 1232 8944 1244
rect 8996 1232 9002 1284
rect 9600 1281 9628 1312
rect 9585 1275 9643 1281
rect 9585 1241 9597 1275
rect 9631 1241 9643 1275
rect 9585 1235 9643 1241
rect 8665 1207 8723 1213
rect 8665 1204 8677 1207
rect 5316 1176 8677 1204
rect 5316 1164 5322 1176
rect 8665 1173 8677 1176
rect 8711 1173 8723 1207
rect 8665 1167 8723 1173
rect 920 1114 10396 1136
rect 920 1062 2566 1114
rect 2618 1062 2630 1114
rect 2682 1062 2694 1114
rect 2746 1062 2758 1114
rect 2810 1062 2822 1114
rect 2874 1062 7566 1114
rect 7618 1062 7630 1114
rect 7682 1062 7694 1114
rect 7746 1062 7758 1114
rect 7810 1062 7822 1114
rect 7874 1062 10396 1114
rect 920 1040 10396 1062
rect 1673 1003 1731 1009
rect 1673 969 1685 1003
rect 1719 1000 1731 1003
rect 3878 1000 3884 1012
rect 1719 972 3884 1000
rect 1719 969 1731 972
rect 1673 963 1731 969
rect 3878 960 3884 972
rect 3936 960 3942 1012
rect 5074 1000 5080 1012
rect 5035 972 5080 1000
rect 5074 960 5080 972
rect 5132 960 5138 1012
rect 8386 960 8392 1012
rect 8444 1000 8450 1012
rect 9217 1003 9275 1009
rect 9217 1000 9229 1003
rect 8444 972 9229 1000
rect 8444 960 8450 972
rect 9217 969 9229 972
rect 9263 969 9275 1003
rect 9217 963 9275 969
rect 9861 1003 9919 1009
rect 9861 969 9873 1003
rect 9907 1000 9919 1003
rect 10226 1000 10232 1012
rect 9907 972 10232 1000
rect 9907 969 9919 972
rect 9861 963 9919 969
rect 10226 960 10232 972
rect 10284 960 10290 1012
rect 1118 892 1124 944
rect 1176 932 1182 944
rect 3053 935 3111 941
rect 3053 932 3065 935
rect 1176 904 3065 932
rect 1176 892 1182 904
rect 3053 901 3065 904
rect 3099 901 3111 935
rect 3053 895 3111 901
rect 3329 935 3387 941
rect 3329 901 3341 935
rect 3375 932 3387 935
rect 5258 932 5264 944
rect 3375 904 5264 932
rect 3375 901 3387 904
rect 3329 895 3387 901
rect 5258 892 5264 904
rect 5316 892 5322 944
rect 6549 935 6607 941
rect 6549 901 6561 935
rect 6595 932 6607 935
rect 8478 932 8484 944
rect 6595 904 8484 932
rect 6595 901 6607 904
rect 6549 895 6607 901
rect 8478 892 8484 904
rect 8536 892 8542 944
rect 8573 935 8631 941
rect 8573 901 8585 935
rect 8619 932 8631 935
rect 8619 904 16574 932
rect 8619 901 8631 904
rect 8573 895 8631 901
rect 3973 867 4031 873
rect 3973 833 3985 867
rect 4019 864 4031 867
rect 16546 864 16574 904
rect 16758 864 16764 876
rect 4019 836 10088 864
rect 16546 836 16764 864
rect 4019 833 4031 836
rect 3973 827 4031 833
rect 2961 799 3019 805
rect 2961 765 2973 799
rect 3007 796 3019 799
rect 3602 796 3608 808
rect 3007 768 3608 796
rect 3007 765 3019 768
rect 2961 759 3019 765
rect 3602 756 3608 768
rect 3660 756 3666 808
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 6638 796 6644 808
rect 6599 768 6644 796
rect 5997 759 6055 765
rect 3697 731 3755 737
rect 3697 697 3709 731
rect 3743 728 3755 731
rect 4154 728 4160 740
rect 3743 700 4160 728
rect 3743 697 3755 700
rect 3697 691 3755 697
rect 4154 688 4160 700
rect 4212 688 4218 740
rect 6012 728 6040 759
rect 6638 756 6644 768
rect 6696 756 6702 808
rect 8294 756 8300 808
rect 8352 796 8358 808
rect 10060 805 10088 836
rect 16758 824 16764 836
rect 16816 824 16822 876
rect 9401 799 9459 805
rect 9401 796 9413 799
rect 8352 768 9413 796
rect 8352 756 8358 768
rect 9401 765 9413 768
rect 9447 765 9459 799
rect 9401 759 9459 765
rect 10045 799 10103 805
rect 10045 765 10057 799
rect 10091 796 10103 799
rect 16574 796 16580 808
rect 10091 768 16580 796
rect 10091 765 10103 768
rect 10045 759 10103 765
rect 16574 756 16580 768
rect 16632 756 16638 808
rect 9585 731 9643 737
rect 9585 728 9597 731
rect 6012 700 9597 728
rect 9585 697 9597 700
rect 9631 697 9643 731
rect 9585 691 9643 697
rect 4172 660 4200 688
rect 6273 663 6331 669
rect 6273 660 6285 663
rect 4172 632 6285 660
rect 6273 629 6285 632
rect 6319 660 6331 663
rect 8662 660 8668 672
rect 6319 632 8668 660
rect 6319 629 6331 632
rect 6273 623 6331 629
rect 8662 620 8668 632
rect 8720 620 8726 672
rect 8846 660 8852 672
rect 8807 632 8852 660
rect 8846 620 8852 632
rect 8904 620 8910 672
rect 9125 663 9183 669
rect 9125 629 9137 663
rect 9171 660 9183 663
rect 9950 660 9956 672
rect 9171 632 9956 660
rect 9171 629 9183 632
rect 9125 623 9183 629
rect 9950 620 9956 632
rect 10008 620 10014 672
rect 920 570 10396 592
rect 920 518 5066 570
rect 5118 518 5130 570
rect 5182 518 5194 570
rect 5246 518 5258 570
rect 5310 518 5322 570
rect 5374 518 10396 570
rect 920 496 10396 518
<< via1 >>
rect 1308 12044 1360 12096
rect 3792 12044 3844 12096
rect 5724 12044 5776 12096
rect 2566 11942 2618 11994
rect 2630 11942 2682 11994
rect 2694 11942 2746 11994
rect 2758 11942 2810 11994
rect 2822 11942 2874 11994
rect 7566 11942 7618 11994
rect 7630 11942 7682 11994
rect 7694 11942 7746 11994
rect 7758 11942 7810 11994
rect 7822 11942 7874 11994
rect 2964 11840 3016 11892
rect 3516 11840 3568 11892
rect 8024 11840 8076 11892
rect 2964 11636 3016 11688
rect 4804 11772 4856 11824
rect 4344 11704 4396 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 5632 11704 5684 11756
rect 7472 11704 7524 11756
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 3884 11636 3936 11688
rect 4436 11636 4488 11688
rect 4988 11636 5040 11688
rect 6276 11636 6328 11688
rect 9036 11636 9088 11688
rect 10232 11636 10284 11688
rect 4712 11568 4764 11620
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 3608 11500 3660 11552
rect 6920 11568 6972 11620
rect 8208 11568 8260 11620
rect 9496 11611 9548 11620
rect 9496 11577 9505 11611
rect 9505 11577 9539 11611
rect 9539 11577 9548 11611
rect 9496 11568 9548 11577
rect 9588 11611 9640 11620
rect 9588 11577 9597 11611
rect 9597 11577 9631 11611
rect 9631 11577 9640 11611
rect 9588 11568 9640 11577
rect 6644 11500 6696 11552
rect 8116 11500 8168 11552
rect 5066 11398 5118 11450
rect 5130 11398 5182 11450
rect 5194 11398 5246 11450
rect 5258 11398 5310 11450
rect 5322 11398 5374 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 3884 11296 3936 11348
rect 6000 11296 6052 11348
rect 6552 11296 6604 11348
rect 2412 11228 2464 11280
rect 10324 11228 10376 11280
rect 3700 11160 3752 11212
rect 3884 11203 3936 11212
rect 3884 11169 3893 11203
rect 3893 11169 3927 11203
rect 3927 11169 3936 11203
rect 3884 11160 3936 11169
rect 6092 11160 6144 11212
rect 7104 11160 7156 11212
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 2136 11092 2188 11144
rect 3792 11092 3844 11144
rect 6000 11092 6052 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7380 11092 7432 11144
rect 8116 11092 8168 11144
rect 5816 11024 5868 11076
rect 7472 11024 7524 11076
rect 9864 11024 9916 11076
rect 6460 10956 6512 11008
rect 2566 10854 2618 10906
rect 2630 10854 2682 10906
rect 2694 10854 2746 10906
rect 2758 10854 2810 10906
rect 2822 10854 2874 10906
rect 7566 10854 7618 10906
rect 7630 10854 7682 10906
rect 7694 10854 7746 10906
rect 7758 10854 7810 10906
rect 7822 10854 7874 10906
rect 1492 10752 1544 10804
rect 3240 10684 3292 10736
rect 3792 10684 3844 10736
rect 5632 10616 5684 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 3608 10548 3660 10600
rect 5356 10548 5408 10600
rect 3148 10480 3200 10532
rect 4528 10480 4580 10532
rect 5908 10752 5960 10804
rect 8760 10727 8812 10736
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 7012 10616 7064 10668
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 9220 10548 9272 10600
rect 9496 10548 9548 10600
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 6000 10480 6052 10532
rect 7472 10480 7524 10532
rect 9772 10523 9824 10532
rect 9772 10489 9781 10523
rect 9781 10489 9815 10523
rect 9815 10489 9824 10523
rect 9772 10480 9824 10489
rect 8392 10412 8444 10464
rect 5066 10310 5118 10362
rect 5130 10310 5182 10362
rect 5194 10310 5246 10362
rect 5258 10310 5310 10362
rect 5322 10310 5374 10362
rect 1676 10183 1728 10192
rect 1676 10149 1685 10183
rect 1685 10149 1719 10183
rect 1719 10149 1728 10183
rect 1676 10140 1728 10149
rect 3148 10140 3200 10192
rect 6736 10208 6788 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7196 10208 7248 10260
rect 10048 10208 10100 10260
rect 4252 10140 4304 10192
rect 5080 10140 5132 10192
rect 5908 10140 5960 10192
rect 6276 10140 6328 10192
rect 6460 10140 6512 10192
rect 4896 10072 4948 10124
rect 8300 10140 8352 10192
rect 8576 10140 8628 10192
rect 8852 10115 8904 10124
rect 8852 10081 8861 10115
rect 8861 10081 8895 10115
rect 8895 10081 8904 10115
rect 8852 10072 8904 10081
rect 9220 10140 9272 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3792 10004 3844 10056
rect 4160 10004 4212 10056
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 3884 9868 3936 9920
rect 4528 9868 4580 9920
rect 7932 9868 7984 9920
rect 8116 9868 8168 9920
rect 9128 9868 9180 9920
rect 2566 9766 2618 9818
rect 2630 9766 2682 9818
rect 2694 9766 2746 9818
rect 2758 9766 2810 9818
rect 2822 9766 2874 9818
rect 7566 9766 7618 9818
rect 7630 9766 7682 9818
rect 7694 9766 7746 9818
rect 7758 9766 7810 9818
rect 7822 9766 7874 9818
rect 3424 9664 3476 9716
rect 5080 9664 5132 9716
rect 5356 9664 5408 9716
rect 6000 9664 6052 9716
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 5908 9596 5960 9648
rect 5356 9528 5408 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 3608 9460 3660 9512
rect 5724 9460 5776 9512
rect 6000 9460 6052 9512
rect 6184 9503 6236 9512
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 6736 9528 6788 9580
rect 8392 9596 8444 9648
rect 9956 9596 10008 9648
rect 8484 9460 8536 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9680 9460 9732 9512
rect 1308 9435 1360 9444
rect 1308 9401 1317 9435
rect 1317 9401 1351 9435
rect 1351 9401 1360 9435
rect 1308 9392 1360 9401
rect 3148 9392 3200 9444
rect 3516 9324 3568 9376
rect 4160 9324 4212 9376
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9220 9324 9272 9376
rect 5066 9222 5118 9274
rect 5130 9222 5182 9274
rect 5194 9222 5246 9274
rect 5258 9222 5310 9274
rect 5322 9222 5374 9274
rect 5724 9120 5776 9172
rect 6552 9120 6604 9172
rect 8668 9120 8720 9172
rect 6276 9052 6328 9104
rect 5908 8984 5960 9036
rect 1308 8959 1360 8968
rect 1308 8925 1317 8959
rect 1317 8925 1351 8959
rect 1351 8925 1360 8959
rect 1308 8916 1360 8925
rect 1400 8916 1452 8968
rect 3148 8916 3200 8968
rect 5540 8916 5592 8968
rect 7104 9052 7156 9104
rect 9680 9120 9732 9172
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 6552 8916 6604 8968
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 9220 8916 9272 8968
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 2688 8848 2740 8900
rect 5264 8848 5316 8900
rect 1676 8780 1728 8832
rect 6092 8780 6144 8832
rect 7104 8780 7156 8832
rect 2566 8678 2618 8730
rect 2630 8678 2682 8730
rect 2694 8678 2746 8730
rect 2758 8678 2810 8730
rect 2822 8678 2874 8730
rect 7566 8678 7618 8730
rect 7630 8678 7682 8730
rect 7694 8678 7746 8730
rect 7758 8678 7810 8730
rect 7822 8678 7874 8730
rect 6184 8576 6236 8628
rect 6736 8576 6788 8628
rect 3424 8508 3476 8560
rect 6276 8508 6328 8560
rect 7748 8508 7800 8560
rect 1492 8440 1544 8492
rect 2780 8440 2832 8492
rect 3240 8440 3292 8492
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 4160 8440 4212 8492
rect 2044 8372 2096 8424
rect 7104 8440 7156 8492
rect 7656 8440 7708 8492
rect 8760 8440 8812 8492
rect 8944 8440 8996 8492
rect 3884 8372 3936 8424
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 6092 8372 6144 8424
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 9312 8415 9364 8424
rect 6184 8372 6236 8381
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 6000 8304 6052 8356
rect 7104 8304 7156 8356
rect 8944 8304 8996 8356
rect 3332 8236 3384 8288
rect 5264 8236 5316 8288
rect 6276 8236 6328 8288
rect 7564 8236 7616 8288
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 17960 8236 18012 8288
rect 19340 8236 19392 8288
rect 5066 8134 5118 8186
rect 5130 8134 5182 8186
rect 5194 8134 5246 8186
rect 5258 8134 5310 8186
rect 5322 8134 5374 8186
rect 1584 7964 1636 8016
rect 3056 7964 3108 8016
rect 3332 7964 3384 8016
rect 3516 7964 3568 8016
rect 6736 7964 6788 8016
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 3148 7760 3200 7812
rect 4804 7896 4856 7948
rect 6000 7896 6052 7948
rect 6552 7939 6604 7948
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 7104 8032 7156 8084
rect 7288 8032 7340 8084
rect 7564 7964 7616 8016
rect 6644 7828 6696 7880
rect 8116 7896 8168 7948
rect 9680 8007 9732 8016
rect 9680 7973 9689 8007
rect 9689 7973 9723 8007
rect 9723 7973 9732 8007
rect 9680 7964 9732 7973
rect 7656 7828 7708 7880
rect 4988 7760 5040 7812
rect 6092 7760 6144 7812
rect 5448 7692 5500 7744
rect 6184 7692 6236 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 6644 7692 6696 7744
rect 8760 7692 8812 7744
rect 2566 7590 2618 7642
rect 2630 7590 2682 7642
rect 2694 7590 2746 7642
rect 2758 7590 2810 7642
rect 2822 7590 2874 7642
rect 7566 7590 7618 7642
rect 7630 7590 7682 7642
rect 7694 7590 7746 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 2964 7488 3016 7540
rect 1308 7352 1360 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3884 7352 3936 7404
rect 6092 7352 6144 7404
rect 6828 7352 6880 7404
rect 10048 7488 10100 7540
rect 9312 7352 9364 7404
rect 9680 7327 9732 7336
rect 3148 7216 3200 7268
rect 3240 7216 3292 7268
rect 4712 7216 4764 7268
rect 4988 7216 5040 7268
rect 6000 7216 6052 7268
rect 4160 7148 4212 7200
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 5540 7148 5592 7200
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 20720 7284 20772 7336
rect 7288 7216 7340 7268
rect 8668 7216 8720 7268
rect 9312 7216 9364 7268
rect 9496 7216 9548 7268
rect 9220 7148 9272 7200
rect 5066 7046 5118 7098
rect 5130 7046 5182 7098
rect 5194 7046 5246 7098
rect 5258 7046 5310 7098
rect 5322 7046 5374 7098
rect 5448 6944 5500 6996
rect 8392 6944 8444 6996
rect 9680 6944 9732 6996
rect 2412 6876 2464 6928
rect 3332 6876 3384 6928
rect 4804 6876 4856 6928
rect 6552 6876 6604 6928
rect 8576 6876 8628 6928
rect 1216 6851 1268 6860
rect 1216 6817 1225 6851
rect 1225 6817 1259 6851
rect 1259 6817 1268 6851
rect 1216 6808 1268 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2228 6740 2280 6792
rect 2688 6672 2740 6724
rect 4436 6740 4488 6792
rect 4988 6672 5040 6724
rect 6092 6808 6144 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9128 6808 9180 6860
rect 9496 6808 9548 6860
rect 6000 6740 6052 6792
rect 3884 6604 3936 6656
rect 6644 6604 6696 6656
rect 8024 6740 8076 6792
rect 9312 6740 9364 6792
rect 9956 6672 10008 6724
rect 8484 6604 8536 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9220 6604 9272 6656
rect 2566 6502 2618 6554
rect 2630 6502 2682 6554
rect 2694 6502 2746 6554
rect 2758 6502 2810 6554
rect 2822 6502 2874 6554
rect 7566 6502 7618 6554
rect 7630 6502 7682 6554
rect 7694 6502 7746 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 7288 6400 7340 6452
rect 8024 6400 8076 6452
rect 8576 6400 8628 6452
rect 4712 6332 4764 6384
rect 6828 6332 6880 6384
rect 1124 6264 1176 6316
rect 5540 6264 5592 6316
rect 6092 6264 6144 6316
rect 8392 6264 8444 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2412 6196 2464 6248
rect 3332 6196 3384 6248
rect 3976 6196 4028 6248
rect 5724 6196 5776 6248
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 7840 6196 7892 6248
rect 8024 6196 8076 6248
rect 3608 6171 3660 6180
rect 3608 6137 3617 6171
rect 3617 6137 3651 6171
rect 3651 6137 3660 6171
rect 3608 6128 3660 6137
rect 6368 6128 6420 6180
rect 9220 6332 9272 6384
rect 9220 6196 9272 6248
rect 9588 6196 9640 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10048 6171 10100 6180
rect 6828 6060 6880 6112
rect 10048 6137 10057 6171
rect 10057 6137 10091 6171
rect 10091 6137 10100 6171
rect 10048 6128 10100 6137
rect 8024 6060 8076 6112
rect 5066 5958 5118 6010
rect 5130 5958 5182 6010
rect 5194 5958 5246 6010
rect 5258 5958 5310 6010
rect 5322 5958 5374 6010
rect 2964 5856 3016 5908
rect 4988 5856 5040 5908
rect 7104 5856 7156 5908
rect 3424 5831 3476 5840
rect 3424 5797 3433 5831
rect 3433 5797 3467 5831
rect 3467 5797 3476 5831
rect 3424 5788 3476 5797
rect 4344 5788 4396 5840
rect 5264 5788 5316 5840
rect 6000 5831 6052 5840
rect 6000 5797 6009 5831
rect 6009 5797 6043 5831
rect 6043 5797 6052 5831
rect 6000 5788 6052 5797
rect 7288 5788 7340 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 3148 5584 3200 5636
rect 6460 5720 6512 5772
rect 7104 5720 7156 5772
rect 8392 5856 8444 5908
rect 8944 5788 8996 5840
rect 9312 5788 9364 5840
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 11060 5788 11112 5840
rect 17960 5788 18012 5840
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 8668 5720 8720 5772
rect 3884 5652 3936 5704
rect 5908 5652 5960 5704
rect 7288 5652 7340 5704
rect 8392 5652 8444 5704
rect 9036 5720 9088 5772
rect 19340 5584 19392 5636
rect 2412 5516 2464 5568
rect 5264 5516 5316 5568
rect 8576 5516 8628 5568
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 2566 5414 2618 5466
rect 2630 5414 2682 5466
rect 2694 5414 2746 5466
rect 2758 5414 2810 5466
rect 2822 5414 2874 5466
rect 7566 5414 7618 5466
rect 7630 5414 7682 5466
rect 7694 5414 7746 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 5632 5312 5684 5364
rect 3056 5244 3108 5296
rect 3240 5176 3292 5228
rect 3424 5176 3476 5228
rect 5448 5219 5500 5228
rect 3148 5108 3200 5160
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 12440 5176 12492 5228
rect 5908 5040 5960 5092
rect 8116 5108 8168 5160
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 9772 5040 9824 5092
rect 6092 4972 6144 5024
rect 7748 4972 7800 5024
rect 5066 4870 5118 4922
rect 5130 4870 5182 4922
rect 5194 4870 5246 4922
rect 5258 4870 5310 4922
rect 5322 4870 5374 4922
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 4620 4768 4672 4820
rect 1584 4700 1636 4752
rect 3148 4700 3200 4752
rect 2044 4632 2096 4684
rect 4252 4700 4304 4752
rect 4344 4700 4396 4752
rect 4988 4700 5040 4752
rect 5908 4632 5960 4684
rect 1952 4564 2004 4616
rect 4252 4428 4304 4480
rect 6092 4428 6144 4480
rect 6460 4428 6512 4480
rect 7104 4768 7156 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9220 4768 9272 4820
rect 8208 4700 8260 4752
rect 9128 4743 9180 4752
rect 7104 4632 7156 4684
rect 8392 4632 8444 4684
rect 8760 4632 8812 4684
rect 9128 4709 9137 4743
rect 9137 4709 9171 4743
rect 9171 4709 9180 4743
rect 9128 4700 9180 4709
rect 9956 4632 10008 4684
rect 10140 4632 10192 4684
rect 7472 4564 7524 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 7840 4564 7892 4616
rect 8208 4564 8260 4616
rect 8300 4564 8352 4616
rect 8484 4496 8536 4548
rect 9036 4496 9088 4548
rect 7566 4326 7618 4378
rect 7630 4326 7682 4378
rect 7694 4326 7746 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 4160 4224 4212 4276
rect 4620 4224 4672 4276
rect 8300 4224 8352 4276
rect 8484 4224 8536 4276
rect 4896 4088 4948 4140
rect 11060 4088 11112 4140
rect 16580 4088 16632 4140
rect 2964 4020 3016 4072
rect 4252 4020 4304 4072
rect 6184 4063 6236 4072
rect 4896 3952 4948 4004
rect 3424 3884 3476 3936
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 7932 4020 7984 4072
rect 10692 4020 10744 4072
rect 6368 3952 6420 4004
rect 7932 3884 7984 3936
rect 5066 3782 5118 3834
rect 5130 3782 5182 3834
rect 5194 3782 5246 3834
rect 5258 3782 5310 3834
rect 5322 3782 5374 3834
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 2688 3544 2740 3596
rect 3332 3544 3384 3596
rect 3240 3476 3292 3528
rect 3424 3476 3476 3528
rect 4988 3476 5040 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 2688 3408 2740 3460
rect 6828 3612 6880 3664
rect 5816 3544 5868 3596
rect 8208 3544 8260 3596
rect 8852 3680 8904 3732
rect 10324 3612 10376 3664
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9036 3587 9088 3596
rect 9036 3553 9045 3587
rect 9045 3553 9079 3587
rect 9079 3553 9088 3587
rect 9036 3544 9088 3553
rect 9772 3544 9824 3596
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 16672 3612 16724 3664
rect 4712 3340 4764 3392
rect 7566 3238 7618 3290
rect 7630 3238 7682 3290
rect 7694 3238 7746 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 4436 3136 4488 3188
rect 5724 3136 5776 3188
rect 6092 3179 6144 3188
rect 6092 3145 6101 3179
rect 6101 3145 6135 3179
rect 6135 3145 6144 3179
rect 6092 3136 6144 3145
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7380 3136 7432 3188
rect 7196 3068 7248 3120
rect 6920 3000 6972 3052
rect 4988 2932 5040 2984
rect 5448 2932 5500 2984
rect 7012 2932 7064 2984
rect 5540 2864 5592 2916
rect 6000 2864 6052 2916
rect 4252 2796 4304 2848
rect 4896 2796 4948 2848
rect 8208 2796 8260 2848
rect 9496 2796 9548 2848
rect 5066 2694 5118 2746
rect 5130 2694 5182 2746
rect 5194 2694 5246 2746
rect 5258 2694 5310 2746
rect 5322 2694 5374 2746
rect 6920 2592 6972 2644
rect 9220 2592 9272 2644
rect 9496 2592 9548 2644
rect 3332 2456 3384 2508
rect 3148 2388 3200 2440
rect 4344 2456 4396 2508
rect 4712 2388 4764 2440
rect 7104 2524 7156 2576
rect 7932 2524 7984 2576
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 8576 2456 8628 2508
rect 9404 2524 9456 2576
rect 9496 2499 9548 2508
rect 8300 2388 8352 2440
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 9036 2388 9088 2440
rect 5816 2320 5868 2372
rect 8852 2320 8904 2372
rect 9588 2388 9640 2440
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 6092 2252 6144 2304
rect 9496 2320 9548 2372
rect 16948 2320 17000 2372
rect 9588 2252 9640 2304
rect 7566 2150 7618 2202
rect 7630 2150 7682 2202
rect 7694 2150 7746 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 3792 2091 3844 2100
rect 3792 2057 3801 2091
rect 3801 2057 3835 2091
rect 3835 2057 3844 2091
rect 3792 2048 3844 2057
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 4436 2048 4488 2100
rect 4620 2048 4672 2100
rect 5816 2091 5868 2100
rect 5816 2057 5825 2091
rect 5825 2057 5859 2091
rect 5859 2057 5868 2091
rect 5816 2048 5868 2057
rect 7288 2048 7340 2100
rect 3424 1980 3476 2032
rect 9496 1980 9548 2032
rect 2964 1912 3016 1964
rect 2688 1844 2740 1896
rect 4344 1912 4396 1964
rect 7012 1912 7064 1964
rect 6460 1887 6512 1896
rect 6460 1853 6469 1887
rect 6469 1853 6503 1887
rect 6503 1853 6512 1887
rect 6460 1844 6512 1853
rect 9864 1887 9916 1896
rect 9864 1853 9873 1887
rect 9873 1853 9907 1887
rect 9907 1853 9916 1887
rect 9864 1844 9916 1853
rect 4160 1708 4212 1760
rect 16856 1776 16908 1828
rect 16672 1708 16724 1760
rect 5066 1606 5118 1658
rect 5130 1606 5182 1658
rect 5194 1606 5246 1658
rect 5258 1606 5310 1658
rect 5322 1606 5374 1658
rect 3516 1504 3568 1556
rect 3700 1547 3752 1556
rect 3700 1513 3709 1547
rect 3709 1513 3743 1547
rect 3743 1513 3752 1547
rect 3700 1504 3752 1513
rect 6828 1504 6880 1556
rect 9312 1504 9364 1556
rect 9772 1504 9824 1556
rect 4988 1436 5040 1488
rect 3884 1368 3936 1420
rect 6092 1411 6144 1420
rect 6092 1377 6101 1411
rect 6101 1377 6135 1411
rect 6135 1377 6144 1411
rect 6092 1368 6144 1377
rect 8024 1411 8076 1420
rect 8024 1377 8033 1411
rect 8033 1377 8067 1411
rect 8067 1377 8076 1411
rect 8024 1368 8076 1377
rect 8576 1368 8628 1420
rect 9036 1411 9088 1420
rect 9036 1377 9045 1411
rect 9045 1377 9079 1411
rect 9079 1377 9088 1411
rect 9036 1368 9088 1377
rect 9220 1368 9272 1420
rect 4252 1300 4304 1352
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 8484 1343 8536 1352
rect 8484 1309 8493 1343
rect 8493 1309 8527 1343
rect 8527 1309 8536 1343
rect 8484 1300 8536 1309
rect 8668 1300 8720 1352
rect 5264 1164 5316 1216
rect 8944 1232 8996 1284
rect 2566 1062 2618 1114
rect 2630 1062 2682 1114
rect 2694 1062 2746 1114
rect 2758 1062 2810 1114
rect 2822 1062 2874 1114
rect 7566 1062 7618 1114
rect 7630 1062 7682 1114
rect 7694 1062 7746 1114
rect 7758 1062 7810 1114
rect 7822 1062 7874 1114
rect 3884 960 3936 1012
rect 5080 1003 5132 1012
rect 5080 969 5089 1003
rect 5089 969 5123 1003
rect 5123 969 5132 1003
rect 5080 960 5132 969
rect 8392 960 8444 1012
rect 10232 960 10284 1012
rect 1124 892 1176 944
rect 5264 892 5316 944
rect 8484 892 8536 944
rect 3608 756 3660 808
rect 6644 799 6696 808
rect 4160 688 4212 740
rect 6644 765 6653 799
rect 6653 765 6687 799
rect 6687 765 6696 799
rect 6644 756 6696 765
rect 8300 756 8352 808
rect 16764 824 16816 876
rect 16580 756 16632 808
rect 8668 620 8720 672
rect 8852 663 8904 672
rect 8852 629 8861 663
rect 8861 629 8895 663
rect 8895 629 8904 663
rect 8852 620 8904 629
rect 9956 620 10008 672
rect 5066 518 5118 570
rect 5130 518 5182 570
rect 5194 518 5246 570
rect 5258 518 5310 570
rect 5322 518 5374 570
<< metal2 >>
rect 938 12322 994 13000
rect 938 12294 1256 12322
rect 938 12200 994 12294
rect 1228 10713 1256 12294
rect 1398 12200 1454 13000
rect 1858 12322 1914 13000
rect 2318 12322 2374 13000
rect 1504 12294 1914 12322
rect 1308 12096 1360 12102
rect 1308 12038 1360 12044
rect 1320 11354 1348 12038
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1214 10704 1270 10713
rect 1412 10690 1440 12200
rect 1504 10826 1532 12294
rect 1858 12200 1914 12294
rect 1964 12294 2374 12322
rect 1674 11112 1730 11121
rect 1674 11047 1730 11056
rect 1504 10810 1624 10826
rect 1492 10804 1624 10810
rect 1544 10798 1624 10804
rect 1492 10746 1544 10752
rect 1412 10662 1532 10690
rect 1214 10639 1270 10648
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 10062 1440 10542
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1400 9512 1452 9518
rect 1306 9480 1362 9489
rect 1400 9454 1452 9460
rect 1136 9424 1306 9432
rect 1136 9404 1308 9424
rect 1136 6322 1164 9404
rect 1360 9415 1362 9424
rect 1308 9386 1360 9392
rect 1412 8974 1440 9454
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1214 7984 1270 7993
rect 1214 7919 1270 7928
rect 1228 6866 1256 7919
rect 1320 7410 1348 8910
rect 1504 8498 1532 10662
rect 1596 8537 1624 10798
rect 1688 10198 1716 11047
rect 1676 10192 1728 10198
rect 1676 10134 1728 10140
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1582 8528 1638 8537
rect 1492 8492 1544 8498
rect 1582 8463 1638 8472
rect 1492 8434 1544 8440
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1124 6316 1176 6322
rect 1124 6258 1176 6264
rect 1136 950 1164 6258
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5778 1440 6190
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1596 5710 1624 7958
rect 1688 6798 1716 8774
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 4758 1624 5646
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 1964 4622 1992 12294
rect 2318 12200 2374 12294
rect 2778 12322 2834 13000
rect 3238 12322 3294 13000
rect 3698 12322 3754 13000
rect 2778 12294 3004 12322
rect 2778 12200 2834 12294
rect 2566 11996 2874 12005
rect 2566 11994 2572 11996
rect 2628 11994 2652 11996
rect 2708 11994 2732 11996
rect 2788 11994 2812 11996
rect 2868 11994 2874 11996
rect 2628 11942 2630 11994
rect 2810 11942 2812 11994
rect 2566 11940 2572 11942
rect 2628 11940 2652 11942
rect 2708 11940 2732 11942
rect 2788 11940 2812 11942
rect 2868 11940 2874 11942
rect 2566 11931 2874 11940
rect 2976 11898 3004 12294
rect 3068 12294 3294 12322
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2964 11688 3016 11694
rect 2502 11656 2558 11665
rect 2964 11630 3016 11636
rect 2502 11591 2558 11600
rect 2516 11558 2544 11591
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2056 4690 2084 8366
rect 2148 5386 2176 11086
rect 2424 7177 2452 11222
rect 2566 10908 2874 10917
rect 2566 10906 2572 10908
rect 2628 10906 2652 10908
rect 2708 10906 2732 10908
rect 2788 10906 2812 10908
rect 2868 10906 2874 10908
rect 2628 10854 2630 10906
rect 2810 10854 2812 10906
rect 2566 10852 2572 10854
rect 2628 10852 2652 10854
rect 2708 10852 2732 10854
rect 2788 10852 2812 10854
rect 2868 10852 2874 10854
rect 2566 10843 2874 10852
rect 2566 9820 2874 9829
rect 2566 9818 2572 9820
rect 2628 9818 2652 9820
rect 2708 9818 2732 9820
rect 2788 9818 2812 9820
rect 2868 9818 2874 9820
rect 2628 9766 2630 9818
rect 2810 9766 2812 9818
rect 2566 9764 2572 9766
rect 2628 9764 2652 9766
rect 2708 9764 2732 9766
rect 2788 9764 2812 9766
rect 2868 9764 2874 9766
rect 2566 9755 2874 9764
rect 2686 8936 2742 8945
rect 2686 8871 2688 8880
rect 2740 8871 2742 8880
rect 2688 8842 2740 8848
rect 2566 8732 2874 8741
rect 2566 8730 2572 8732
rect 2628 8730 2652 8732
rect 2708 8730 2732 8732
rect 2788 8730 2812 8732
rect 2868 8730 2874 8732
rect 2628 8678 2630 8730
rect 2810 8678 2812 8730
rect 2566 8676 2572 8678
rect 2628 8676 2652 8678
rect 2708 8676 2732 8678
rect 2788 8676 2812 8678
rect 2868 8676 2874 8678
rect 2566 8667 2874 8676
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2792 7970 2820 8434
rect 2870 7984 2926 7993
rect 2792 7942 2870 7970
rect 2870 7919 2926 7928
rect 2596 7880 2648 7886
rect 2594 7848 2596 7857
rect 2648 7848 2650 7857
rect 2594 7783 2650 7792
rect 2566 7644 2874 7653
rect 2566 7642 2572 7644
rect 2628 7642 2652 7644
rect 2708 7642 2732 7644
rect 2788 7642 2812 7644
rect 2868 7642 2874 7644
rect 2628 7590 2630 7642
rect 2810 7590 2812 7642
rect 2566 7588 2572 7590
rect 2628 7588 2652 7590
rect 2708 7588 2732 7590
rect 2788 7588 2812 7590
rect 2868 7588 2874 7590
rect 2566 7579 2874 7588
rect 2976 7546 3004 11630
rect 3068 8022 3096 12294
rect 3238 12200 3294 12294
rect 3344 12294 3754 12322
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 10198 3188 10474
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3160 9625 3188 10134
rect 3146 9616 3202 9625
rect 3146 9551 3202 9560
rect 3160 9450 3188 9551
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3160 8129 3188 8910
rect 3252 8498 3280 10678
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 8378 3372 12294
rect 3698 12200 3754 12294
rect 4158 12322 4214 13000
rect 4618 12322 4674 13000
rect 5078 12322 5134 13000
rect 4158 12294 4476 12322
rect 4158 12200 4214 12294
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3436 9586 3464 9658
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3528 9489 3556 11834
rect 3804 11694 3832 12038
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 10606 3648 11494
rect 3896 11354 3924 11630
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3608 9512 3660 9518
rect 3514 9480 3570 9489
rect 3608 9454 3660 9460
rect 3514 9415 3570 9424
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3252 8350 3372 8378
rect 3146 8120 3202 8129
rect 3146 8055 3202 8064
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2410 7168 2466 7177
rect 2410 7103 2466 7112
rect 2240 6990 2636 7018
rect 2240 6798 2268 6990
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2424 6254 2452 6870
rect 2608 6746 2636 6990
rect 2608 6730 2728 6746
rect 2608 6724 2740 6730
rect 2608 6718 2688 6724
rect 2688 6666 2740 6672
rect 2566 6556 2874 6565
rect 2566 6554 2572 6556
rect 2628 6554 2652 6556
rect 2708 6554 2732 6556
rect 2788 6554 2812 6556
rect 2868 6554 2874 6556
rect 2628 6502 2630 6554
rect 2810 6502 2812 6554
rect 2566 6500 2572 6502
rect 2628 6500 2652 6502
rect 2708 6500 2732 6502
rect 2788 6500 2812 6502
rect 2868 6500 2874 6502
rect 2566 6491 2874 6500
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5574 2452 6190
rect 2976 5914 3004 7482
rect 3160 7410 3188 7754
rect 3252 7449 3280 8350
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 8022 3372 8230
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3238 7440 3294 7449
rect 3148 7404 3200 7410
rect 3238 7375 3294 7384
rect 3148 7346 3200 7352
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3054 7168 3110 7177
rect 3054 7103 3110 7112
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2148 5358 2360 5386
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 2332 1986 2360 5358
rect 2424 3584 2452 5510
rect 2566 5468 2874 5477
rect 2566 5466 2572 5468
rect 2628 5466 2652 5468
rect 2708 5466 2732 5468
rect 2788 5466 2812 5468
rect 2868 5466 2874 5468
rect 2628 5414 2630 5466
rect 2810 5414 2812 5466
rect 2566 5412 2572 5414
rect 2628 5412 2652 5414
rect 2708 5412 2732 5414
rect 2788 5412 2812 5414
rect 2868 5412 2874 5414
rect 2566 5403 2874 5412
rect 2976 4078 3004 5850
rect 3068 5302 3096 7103
rect 3160 5642 3188 7210
rect 3252 7154 3280 7210
rect 3252 7126 3372 7154
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3160 5166 3188 5578
rect 3252 5234 3280 6967
rect 3344 6934 3372 7126
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2688 3596 2740 3602
rect 2424 3556 2688 3584
rect 2688 3538 2740 3544
rect 2688 3460 2740 3466
rect 2686 3428 2688 3437
rect 2740 3428 2742 3437
rect 2686 3363 2742 3372
rect 2332 1958 2728 1986
rect 2976 1970 3004 4014
rect 3160 2446 3188 4694
rect 3252 3534 3280 5170
rect 3344 3738 3372 6190
rect 3436 5846 3464 8502
rect 3528 8022 3556 9318
rect 3620 8498 3648 9454
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3436 5234 3464 5782
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3422 4856 3478 4865
rect 3422 4791 3424 4800
rect 3476 4791 3478 4800
rect 3424 4762 3476 4768
rect 3436 3942 3464 4762
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3344 2514 3372 3538
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3436 2310 3464 3470
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2038 3464 2246
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 2700 1902 2728 1958
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 3528 1562 3556 7822
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 2566 1116 2874 1125
rect 2566 1114 2572 1116
rect 2628 1114 2652 1116
rect 2708 1114 2732 1116
rect 2788 1114 2812 1116
rect 2868 1114 2874 1116
rect 2628 1062 2630 1114
rect 2810 1062 2812 1114
rect 2566 1060 2572 1062
rect 2628 1060 2652 1062
rect 2708 1060 2732 1062
rect 2788 1060 2812 1062
rect 2868 1060 2874 1062
rect 2566 1051 2874 1060
rect 1124 944 1176 950
rect 1124 886 1176 892
rect 3620 814 3648 6122
rect 3712 1562 3740 11154
rect 3792 11144 3844 11150
rect 3896 11121 3924 11154
rect 3792 11086 3844 11092
rect 3882 11112 3938 11121
rect 3804 10962 3832 11086
rect 3882 11047 3938 11056
rect 3804 10934 4108 10962
rect 3790 10840 3846 10849
rect 3790 10775 3846 10784
rect 3804 10742 3832 10775
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3882 10704 3938 10713
rect 3882 10639 3938 10648
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 2106 3832 9998
rect 3896 9926 3924 10639
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 8430 3924 9862
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3882 8120 3938 8129
rect 3882 8055 3938 8064
rect 3896 7410 3924 8055
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3896 6662 3924 7346
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 5710 3924 6598
rect 3988 6254 4016 9007
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3700 1556 3752 1562
rect 3700 1498 3752 1504
rect 3896 1426 3924 5646
rect 4080 2106 4108 10934
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9382 4200 9998
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 8498 4200 9318
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 4282 4200 7142
rect 4264 4758 4292 10134
rect 4356 9586 4384 11698
rect 4448 11694 4476 12294
rect 4618 12294 4752 12322
rect 4618 12200 4674 12294
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4724 11626 4752 12294
rect 4908 12294 5134 12322
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4540 10010 4568 10474
rect 4540 9982 4660 10010
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4342 9480 4398 9489
rect 4342 9415 4398 9424
rect 4356 8537 4384 9415
rect 4342 8528 4398 8537
rect 4342 8463 4398 8472
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 5846 4384 7142
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4356 4758 4384 5782
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4264 4078 4292 4422
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4448 3194 4476 6734
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 3884 1420 3936 1426
rect 3884 1362 3936 1368
rect 3896 1018 3924 1362
rect 3884 1012 3936 1018
rect 3884 954 3936 960
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 4172 746 4200 1702
rect 4264 1358 4292 2790
rect 4540 2774 4568 9862
rect 4632 4826 4660 9982
rect 4724 7274 4752 11562
rect 4816 9625 4844 11766
rect 4908 10441 4936 12294
rect 5078 12200 5134 12294
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4894 10432 4950 10441
rect 4894 10367 4950 10376
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4816 7018 4844 7890
rect 4724 6990 4844 7018
rect 4724 6390 4752 6990
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4710 6216 4766 6225
rect 4710 6151 4766 6160
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4448 2746 4568 2774
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4356 1970 4384 2450
rect 4448 2106 4476 2746
rect 4632 2106 4660 4218
rect 4724 3398 4752 6151
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4816 2774 4844 6870
rect 4908 4146 4936 10066
rect 5000 8673 5028 11630
rect 5066 11452 5374 11461
rect 5066 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5312 11452
rect 5368 11450 5374 11452
rect 5128 11398 5130 11450
rect 5310 11398 5312 11450
rect 5066 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5312 11398
rect 5368 11396 5374 11398
rect 5066 11387 5374 11396
rect 5354 10840 5410 10849
rect 5354 10775 5410 10784
rect 5368 10606 5396 10775
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5066 10364 5374 10373
rect 5066 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5312 10364
rect 5368 10362 5374 10364
rect 5128 10310 5130 10362
rect 5310 10310 5312 10362
rect 5066 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5312 10310
rect 5368 10308 5374 10310
rect 5066 10299 5374 10308
rect 5460 10305 5488 11698
rect 5446 10296 5502 10305
rect 5446 10231 5502 10240
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5092 9722 5120 10134
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5356 9716 5408 9722
rect 5552 9674 5580 12200
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 10674 5672 11698
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5356 9658 5408 9664
rect 5368 9586 5396 9658
rect 5460 9646 5580 9674
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5066 9276 5374 9285
rect 5066 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5312 9276
rect 5368 9274 5374 9276
rect 5128 9222 5130 9274
rect 5310 9222 5312 9274
rect 5066 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5312 9222
rect 5368 9220 5374 9222
rect 5066 9211 5374 9220
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4986 8664 5042 8673
rect 4986 8599 5042 8608
rect 5276 8294 5304 8842
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5066 8188 5374 8197
rect 5066 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5312 8188
rect 5368 8186 5374 8188
rect 5128 8134 5130 8186
rect 5310 8134 5312 8186
rect 5066 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5312 8134
rect 5368 8132 5374 8134
rect 5066 8123 5374 8132
rect 5460 7834 5488 9646
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8129 5580 8910
rect 5644 8430 5672 10610
rect 5736 9518 5764 12038
rect 6012 11354 6040 12200
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5538 8120 5594 8129
rect 5538 8055 5594 8064
rect 5644 7970 5672 8366
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5368 7806 5488 7834
rect 5552 7942 5672 7970
rect 5000 7274 5028 7754
rect 5368 7313 5396 7806
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5354 7304 5410 7313
rect 4988 7268 5040 7274
rect 5354 7239 5410 7248
rect 4988 7210 5040 7216
rect 5066 7100 5374 7109
rect 5066 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5312 7100
rect 5368 7098 5374 7100
rect 5128 7046 5130 7098
rect 5310 7046 5312 7098
rect 5066 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5312 7046
rect 5368 7044 5374 7046
rect 5066 7035 5374 7044
rect 5460 7002 5488 7686
rect 5552 7206 5580 7942
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 5000 5914 5028 6666
rect 5066 6012 5374 6021
rect 5066 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5312 6012
rect 5368 6010 5374 6012
rect 5128 5958 5130 6010
rect 5310 5958 5312 6010
rect 5066 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5312 5958
rect 5368 5956 5374 5958
rect 5066 5947 5374 5956
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 5264 5840 5316 5846
rect 5262 5808 5264 5817
rect 5316 5808 5318 5817
rect 5262 5743 5318 5752
rect 5276 5574 5304 5743
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5460 5234 5488 6938
rect 5552 6322 5580 7142
rect 5736 6474 5764 9114
rect 5644 6446 5764 6474
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5066 4924 5374 4933
rect 5066 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5312 4924
rect 5368 4922 5374 4924
rect 5128 4870 5130 4922
rect 5310 4870 5312 4922
rect 5066 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5312 4870
rect 5368 4868 5374 4870
rect 5066 4859 5374 4868
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4908 2854 4936 3946
rect 5000 3534 5028 4694
rect 5066 3836 5374 3845
rect 5066 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5312 3836
rect 5368 3834 5374 3836
rect 5128 3782 5130 3834
rect 5310 3782 5312 3834
rect 5066 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5312 3782
rect 5368 3780 5374 3782
rect 5066 3771 5374 3780
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5368 3534 5396 3567
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5460 2990 5488 5170
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4724 2746 4844 2774
rect 4724 2446 4752 2746
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 5000 1494 5028 2926
rect 5552 2922 5580 6258
rect 5644 5370 5672 6446
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5736 3194 5764 6190
rect 5828 3602 5856 11018
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5920 10198 5948 10746
rect 6012 10674 6040 11086
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 6012 9722 6040 10474
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5920 9353 5948 9590
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5906 9344 5962 9353
rect 5906 9279 5962 9288
rect 5906 9208 5962 9217
rect 5906 9143 5962 9152
rect 5920 9042 5948 9143
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6012 8514 6040 9454
rect 6104 8838 6132 11154
rect 6288 10198 6316 11630
rect 6472 11098 6500 12200
rect 7566 11996 7874 12005
rect 7566 11994 7572 11996
rect 7628 11994 7652 11996
rect 7708 11994 7732 11996
rect 7788 11994 7812 11996
rect 7868 11994 7874 11996
rect 7628 11942 7630 11994
rect 7810 11942 7812 11994
rect 7566 11940 7572 11942
rect 7628 11940 7652 11942
rect 7708 11940 7732 11942
rect 7788 11940 7812 11942
rect 7868 11940 7874 11942
rect 7566 11931 7874 11940
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6380 11070 6500 11098
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6196 8634 6224 9454
rect 6288 9110 6316 9998
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6276 8560 6328 8566
rect 6012 8486 6224 8514
rect 6276 8502 6328 8508
rect 6196 8430 6224 8486
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6012 7954 6040 8298
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7274 6040 7890
rect 6104 7818 6132 8366
rect 6288 8294 6316 8502
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6380 7834 6408 11070
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10606 6500 10950
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6472 8401 6500 10134
rect 6564 9178 6592 11290
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8809 6592 8910
rect 6550 8800 6606 8809
rect 6550 8735 6606 8744
rect 6550 8664 6606 8673
rect 6550 8599 6606 8608
rect 6458 8392 6514 8401
rect 6458 8327 6514 8336
rect 6458 8256 6514 8265
rect 6458 8191 6514 8200
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6288 7806 6408 7834
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6000 7268 6052 7274
rect 5920 7228 6000 7256
rect 5920 5710 5948 7228
rect 6000 7210 6052 7216
rect 6104 6866 6132 7346
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 5846 6040 6734
rect 6104 6322 6132 6802
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6090 6216 6146 6225
rect 6090 6151 6146 6160
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5920 4690 5948 5034
rect 6104 5030 6132 6151
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6104 4570 6132 4966
rect 6012 4542 6132 4570
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 6012 2922 6040 4542
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 3194 6132 4422
rect 6196 4078 6224 7686
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6288 2774 6316 7806
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 6186 6408 7686
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6472 5930 6500 8191
rect 6564 7954 6592 8599
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6564 6934 6592 7890
rect 6656 7886 6684 11494
rect 6932 10266 6960 11562
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6748 9586 6776 10202
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8022 6776 8570
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6644 7744 6696 7750
rect 6642 7712 6644 7721
rect 6696 7712 6698 7721
rect 6642 7647 6698 7656
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6380 5902 6500 5930
rect 6380 4010 6408 5902
rect 6460 5772 6512 5778
rect 6564 5760 6592 6870
rect 6656 6769 6684 7647
rect 6734 7440 6790 7449
rect 6840 7410 6868 8910
rect 6734 7375 6790 7384
rect 6828 7404 6880 7410
rect 6642 6760 6698 6769
rect 6642 6695 6698 6704
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6512 5732 6592 5760
rect 6460 5714 6512 5720
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6380 3194 6408 3946
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5066 2748 5374 2757
rect 5066 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5312 2748
rect 5368 2746 5374 2748
rect 5128 2694 5130 2746
rect 5310 2694 5312 2746
rect 5066 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5312 2694
rect 5368 2692 5374 2694
rect 5066 2683 5374 2692
rect 5828 2746 6316 2774
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5066 1660 5374 1669
rect 5066 1658 5072 1660
rect 5128 1658 5152 1660
rect 5208 1658 5232 1660
rect 5288 1658 5312 1660
rect 5368 1658 5374 1660
rect 5128 1606 5130 1658
rect 5310 1606 5312 1658
rect 5066 1604 5072 1606
rect 5128 1604 5152 1606
rect 5208 1604 5232 1606
rect 5288 1604 5312 1606
rect 5368 1604 5374 1606
rect 5066 1595 5374 1604
rect 4988 1488 5040 1494
rect 5460 1442 5488 2382
rect 5828 2378 5856 2746
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5828 2106 5856 2314
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 4988 1430 5040 1436
rect 5368 1414 5488 1442
rect 6104 1426 6132 2246
rect 6472 1902 6500 4422
rect 6564 2825 6592 5607
rect 6550 2816 6606 2825
rect 6550 2751 6606 2760
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6092 1420 6144 1426
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 5078 1320 5134 1329
rect 5078 1255 5134 1264
rect 5092 1018 5120 1255
rect 5264 1216 5316 1222
rect 5264 1158 5316 1164
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5276 950 5304 1158
rect 5264 944 5316 950
rect 5264 886 5316 892
rect 5368 762 5396 1414
rect 6092 1362 6144 1368
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5460 921 5488 1294
rect 5446 912 5502 921
rect 5446 847 5502 856
rect 6656 814 6684 6598
rect 6748 5234 6776 7375
rect 6828 7346 6880 7352
rect 6826 7304 6882 7313
rect 6826 7239 6882 7248
rect 6840 6390 6868 7239
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6734 4176 6790 4185
rect 6734 4111 6790 4120
rect 6748 2446 6776 4111
rect 6840 3670 6868 6054
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6932 3058 6960 9415
rect 7024 3194 7052 10610
rect 7116 9625 7144 11154
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7102 9616 7158 9625
rect 7102 9551 7158 9560
rect 7116 9110 7144 9551
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8498 7144 8774
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7116 8090 7144 8298
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7208 7868 7236 10202
rect 7300 8809 7328 11086
rect 7286 8800 7342 8809
rect 7286 8735 7342 8744
rect 7300 8401 7328 8735
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7116 7840 7236 7868
rect 7116 5914 7144 7840
rect 7194 7304 7250 7313
rect 7300 7274 7328 8026
rect 7194 7239 7250 7248
rect 7288 7268 7340 7274
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7116 4826 7144 5714
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7102 4720 7158 4729
rect 7102 4655 7104 4664
rect 7156 4655 7158 4664
rect 7104 4626 7156 4632
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7012 2984 7064 2990
rect 6826 2952 6882 2961
rect 7012 2926 7064 2932
rect 6826 2887 6882 2896
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6840 1562 6868 2887
rect 6918 2816 6974 2825
rect 6918 2751 6974 2760
rect 6932 2650 6960 2751
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7024 1970 7052 2926
rect 7116 2582 7144 4626
rect 7208 3126 7236 7239
rect 7288 7210 7340 7216
rect 7300 6458 7328 7210
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5846 7328 6190
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7300 2106 7328 5646
rect 7392 3194 7420 11086
rect 7484 11082 7512 11698
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7566 10908 7874 10917
rect 7566 10906 7572 10908
rect 7628 10906 7652 10908
rect 7708 10906 7732 10908
rect 7788 10906 7812 10908
rect 7868 10906 7874 10908
rect 7628 10854 7630 10906
rect 7810 10854 7812 10906
rect 7566 10852 7572 10854
rect 7628 10852 7652 10854
rect 7708 10852 7732 10854
rect 7788 10852 7812 10854
rect 7868 10852 7874 10854
rect 7566 10843 7874 10852
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 4622 7512 10474
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7566 9820 7874 9829
rect 7566 9818 7572 9820
rect 7628 9818 7652 9820
rect 7708 9818 7732 9820
rect 7788 9818 7812 9820
rect 7868 9818 7874 9820
rect 7628 9766 7630 9818
rect 7810 9766 7812 9818
rect 7566 9764 7572 9766
rect 7628 9764 7652 9766
rect 7708 9764 7732 9766
rect 7788 9764 7812 9766
rect 7868 9764 7874 9766
rect 7566 9755 7874 9764
rect 7656 9376 7708 9382
rect 7654 9344 7656 9353
rect 7708 9344 7710 9353
rect 7654 9279 7710 9288
rect 7566 8732 7874 8741
rect 7566 8730 7572 8732
rect 7628 8730 7652 8732
rect 7708 8730 7732 8732
rect 7788 8730 7812 8732
rect 7868 8730 7874 8732
rect 7628 8678 7630 8730
rect 7810 8678 7812 8730
rect 7566 8676 7572 8678
rect 7628 8676 7652 8678
rect 7708 8676 7732 8678
rect 7788 8676 7812 8678
rect 7868 8676 7874 8678
rect 7566 8667 7874 8676
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 8022 7604 8230
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7668 7886 7696 8434
rect 7760 8401 7788 8502
rect 7746 8392 7802 8401
rect 7746 8327 7802 8336
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7566 7644 7874 7653
rect 7566 7642 7572 7644
rect 7628 7642 7652 7644
rect 7708 7642 7732 7644
rect 7788 7642 7812 7644
rect 7868 7642 7874 7644
rect 7628 7590 7630 7642
rect 7810 7590 7812 7642
rect 7566 7588 7572 7590
rect 7628 7588 7652 7590
rect 7708 7588 7732 7590
rect 7788 7588 7812 7590
rect 7868 7588 7874 7590
rect 7566 7579 7874 7588
rect 7566 6556 7874 6565
rect 7566 6554 7572 6556
rect 7628 6554 7652 6556
rect 7708 6554 7732 6556
rect 7788 6554 7812 6556
rect 7868 6554 7874 6556
rect 7628 6502 7630 6554
rect 7810 6502 7812 6554
rect 7566 6500 7572 6502
rect 7628 6500 7652 6502
rect 7708 6500 7732 6502
rect 7788 6500 7812 6502
rect 7868 6500 7874 6502
rect 7566 6491 7874 6500
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5556 7880 6190
rect 7944 5681 7972 9862
rect 8036 9194 8064 11834
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11150 8156 11494
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8116 9920 8168 9926
rect 8220 9874 8248 11562
rect 8758 11112 8814 11121
rect 8758 11047 8814 11056
rect 8772 10742 8800 11047
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8168 9868 8248 9874
rect 8116 9862 8248 9868
rect 8128 9846 8248 9862
rect 8220 9217 8248 9846
rect 8206 9208 8262 9217
rect 8036 9166 8156 9194
rect 8022 8120 8078 8129
rect 8022 8055 8078 8064
rect 8036 6798 8064 8055
rect 8128 7954 8156 9166
rect 8206 9143 8262 9152
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8036 6254 8064 6394
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7930 5672 7986 5681
rect 7930 5607 7986 5616
rect 7852 5528 7972 5556
rect 7566 5468 7874 5477
rect 7566 5466 7572 5468
rect 7628 5466 7652 5468
rect 7708 5466 7732 5468
rect 7788 5466 7812 5468
rect 7868 5466 7874 5468
rect 7628 5414 7630 5466
rect 7810 5414 7812 5466
rect 7566 5412 7572 5414
rect 7628 5412 7652 5414
rect 7708 5412 7732 5414
rect 7788 5412 7812 5414
rect 7868 5412 7874 5414
rect 7566 5403 7874 5412
rect 7944 5352 7972 5528
rect 7852 5324 7972 5352
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4622 7788 4966
rect 7852 4622 7880 5324
rect 7930 5264 7986 5273
rect 7930 5199 7986 5208
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7566 4380 7874 4389
rect 7566 4378 7572 4380
rect 7628 4378 7652 4380
rect 7708 4378 7732 4380
rect 7788 4378 7812 4380
rect 7868 4378 7874 4380
rect 7628 4326 7630 4378
rect 7810 4326 7812 4378
rect 7566 4324 7572 4326
rect 7628 4324 7652 4326
rect 7708 4324 7732 4326
rect 7788 4324 7812 4326
rect 7868 4324 7874 4326
rect 7566 4315 7874 4324
rect 7944 4078 7972 5199
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7566 3292 7874 3301
rect 7566 3290 7572 3292
rect 7628 3290 7652 3292
rect 7708 3290 7732 3292
rect 7788 3290 7812 3292
rect 7868 3290 7874 3292
rect 7628 3238 7630 3290
rect 7810 3238 7812 3290
rect 7566 3236 7572 3238
rect 7628 3236 7652 3238
rect 7708 3236 7732 3238
rect 7788 3236 7812 3238
rect 7868 3236 7874 3238
rect 7566 3227 7874 3236
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7944 2582 7972 3878
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 7566 2204 7874 2213
rect 7566 2202 7572 2204
rect 7628 2202 7652 2204
rect 7708 2202 7732 2204
rect 7788 2202 7812 2204
rect 7868 2202 7874 2204
rect 7628 2150 7630 2202
rect 7810 2150 7812 2202
rect 7566 2148 7572 2150
rect 7628 2148 7652 2150
rect 7708 2148 7732 2150
rect 7788 2148 7812 2150
rect 7868 2148 7874 2150
rect 7566 2139 7874 2148
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 8036 1426 8064 6054
rect 8128 5166 8156 7511
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8220 4758 8248 8978
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8312 4622 8340 10134
rect 8404 9654 8432 10406
rect 8576 10192 8628 10198
rect 8574 10160 8576 10169
rect 8628 10160 8630 10169
rect 8574 10095 8630 10104
rect 8852 10124 8904 10130
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8484 9512 8536 9518
rect 8404 9460 8484 9466
rect 8404 9454 8536 9460
rect 8404 9438 8524 9454
rect 8404 7002 8432 9438
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6662 8524 9318
rect 8588 7041 8616 10095
rect 8852 10066 8904 10072
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8680 7426 8708 9114
rect 8772 8498 8800 9454
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 8129 8800 8230
rect 8758 8120 8814 8129
rect 8758 8055 8814 8064
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7585 8800 7686
rect 8758 7576 8814 7585
rect 8758 7511 8814 7520
rect 8680 7398 8800 7426
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8574 7032 8630 7041
rect 8574 6967 8630 6976
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8588 6458 8616 6870
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8680 6338 8708 7210
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8588 6310 8708 6338
rect 8404 5914 8432 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8404 5710 8432 5850
rect 8588 5778 8616 6310
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8576 5568 8628 5574
rect 8390 5536 8446 5545
rect 8576 5510 8628 5516
rect 8390 5471 8446 5480
rect 8404 4842 8432 5471
rect 8404 4826 8524 4842
rect 8392 4820 8524 4826
rect 8444 4814 8524 4820
rect 8392 4762 8444 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8220 3602 8248 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 2854 8248 3538
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8312 2774 8340 4218
rect 8404 3534 8432 4626
rect 8496 4554 8524 4814
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 4282 8524 4490
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 3528 8444 3534
rect 8444 3476 8524 3482
rect 8392 3470 8524 3476
rect 8404 3454 8524 3470
rect 8312 2746 8432 2774
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8024 1420 8076 1426
rect 8024 1362 8076 1368
rect 7566 1116 7874 1125
rect 7566 1114 7572 1116
rect 7628 1114 7652 1116
rect 7708 1114 7732 1116
rect 7788 1114 7812 1116
rect 7868 1114 7874 1116
rect 7628 1062 7630 1114
rect 7810 1062 7812 1114
rect 7566 1060 7572 1062
rect 7628 1060 7652 1062
rect 7708 1060 7732 1062
rect 7788 1060 7812 1062
rect 7868 1060 7874 1062
rect 7566 1051 7874 1060
rect 8312 814 8340 2382
rect 8404 1018 8432 2746
rect 8496 1358 8524 3454
rect 8588 2514 8616 5510
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8576 1420 8628 1426
rect 8576 1362 8628 1368
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 8588 1034 8616 1362
rect 8680 1358 8708 5714
rect 8772 4690 8800 7398
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8864 3738 8892 10066
rect 8942 8528 8998 8537
rect 8942 8463 8944 8472
rect 8996 8463 8998 8472
rect 8944 8434 8996 8440
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8956 7177 8984 8298
rect 8942 7168 8998 7177
rect 8942 7103 8998 7112
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8956 5846 8984 6802
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9048 5778 9076 11630
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9232 10198 9260 10542
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 6866 9168 9862
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8974 9260 9318
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9232 7206 9260 8910
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 7410 9352 8366
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9310 7304 9366 7313
rect 9310 7239 9312 7248
rect 9364 7239 9366 7248
rect 9312 7210 9364 7216
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9048 4554 9076 5714
rect 9140 4758 9168 6598
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 4826 9260 6190
rect 9324 5846 9352 6734
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8942 2544 8998 2553
rect 8942 2479 8998 2488
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8392 1012 8444 1018
rect 8392 954 8444 960
rect 8496 1006 8616 1034
rect 8496 950 8524 1006
rect 8484 944 8536 950
rect 8484 886 8536 892
rect 6644 808 6696 814
rect 4160 740 4212 746
rect 5368 734 5488 762
rect 6644 750 6696 756
rect 8300 808 8352 814
rect 8300 750 8352 756
rect 4160 682 4212 688
rect 5066 572 5374 581
rect 5066 570 5072 572
rect 5128 570 5152 572
rect 5208 570 5232 572
rect 5288 570 5312 572
rect 5368 570 5374 572
rect 5128 518 5130 570
rect 5310 518 5312 570
rect 5066 516 5072 518
rect 5128 516 5152 518
rect 5208 516 5232 518
rect 5288 516 5312 518
rect 5368 516 5374 518
rect 5066 507 5374 516
rect 5460 513 5488 734
rect 8680 678 8708 1294
rect 8864 678 8892 2314
rect 8956 1290 8984 2479
rect 9048 2446 9076 3538
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9034 1728 9090 1737
rect 9034 1663 9090 1672
rect 9048 1426 9076 1663
rect 9232 1426 9260 2586
rect 9324 1562 9352 5782
rect 9416 2582 9444 11154
rect 9508 10606 9536 11562
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 7274 9536 10542
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 5574 9536 6802
rect 9600 6254 9628 11562
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9353 9720 9454
rect 9678 9344 9734 9353
rect 9678 9279 9734 9288
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9692 8022 9720 9114
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 7002 9720 7278
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6254 9812 10474
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9876 5846 9904 11018
rect 10060 10606 10088 12271
rect 20718 11928 20774 11937
rect 20718 11863 20774 11872
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10060 10266 10088 10542
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10138 9888 10194 9897
rect 10138 9823 10194 9832
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9968 6730 9996 9590
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 7546 10088 8910
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 3602 9812 5034
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9508 2650 9536 2790
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9508 2378 9536 2450
rect 9600 2446 9628 3470
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9508 2038 9536 2314
rect 9600 2310 9628 2382
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 9784 1562 9812 3538
rect 9876 1902 9904 5782
rect 10060 5166 10088 6122
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10152 4690 10180 9823
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9036 1420 9088 1426
rect 9036 1362 9088 1368
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 8944 1284 8996 1290
rect 8944 1226 8996 1232
rect 9968 678 9996 4626
rect 10244 1018 10272 11630
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10336 3670 10364 11222
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19352 8294 19380 11047
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 12438 6624 12494 6633
rect 12438 6559 12494 6568
rect 10690 6216 10746 6225
rect 10690 6151 10746 6160
rect 10704 4078 10732 6151
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 4146 11100 5782
rect 12452 5234 12480 6559
rect 17972 5846 18000 8230
rect 20732 7342 20760 11863
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 17960 5840 18012 5846
rect 16946 5808 17002 5817
rect 17960 5782 18012 5788
rect 16946 5743 17002 5752
rect 16578 5400 16634 5409
rect 16578 5335 16634 5344
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 16592 4146 16620 5335
rect 16670 4992 16726 5001
rect 16670 4927 16726 4936
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 16684 3670 16712 4927
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16670 3360 16726 3369
rect 16670 3295 16726 3304
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 10232 1012 10284 1018
rect 10232 954 10284 960
rect 16592 814 16620 2071
rect 16684 1766 16712 3295
rect 16762 2544 16818 2553
rect 16762 2479 16818 2488
rect 16672 1760 16724 1766
rect 16672 1702 16724 1708
rect 16776 882 16804 2479
rect 16868 1834 16896 4519
rect 16960 2378 16988 5743
rect 19352 5642 19380 6967
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 16764 876 16816 882
rect 16764 818 16816 824
rect 16580 808 16632 814
rect 16580 750 16632 756
rect 8668 672 8720 678
rect 8668 614 8720 620
rect 8852 672 8904 678
rect 8852 614 8904 620
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 5446 504 5502 513
rect 5446 439 5502 448
<< via2 >>
rect 1214 10648 1270 10704
rect 1674 11056 1730 11112
rect 1306 9444 1362 9480
rect 1306 9424 1308 9444
rect 1308 9424 1360 9444
rect 1360 9424 1362 9444
rect 1214 7928 1270 7984
rect 1582 8472 1638 8528
rect 2572 11994 2628 11996
rect 2652 11994 2708 11996
rect 2732 11994 2788 11996
rect 2812 11994 2868 11996
rect 2572 11942 2618 11994
rect 2618 11942 2628 11994
rect 2652 11942 2682 11994
rect 2682 11942 2694 11994
rect 2694 11942 2708 11994
rect 2732 11942 2746 11994
rect 2746 11942 2758 11994
rect 2758 11942 2788 11994
rect 2812 11942 2822 11994
rect 2822 11942 2868 11994
rect 2572 11940 2628 11942
rect 2652 11940 2708 11942
rect 2732 11940 2788 11942
rect 2812 11940 2868 11942
rect 2502 11600 2558 11656
rect 2572 10906 2628 10908
rect 2652 10906 2708 10908
rect 2732 10906 2788 10908
rect 2812 10906 2868 10908
rect 2572 10854 2618 10906
rect 2618 10854 2628 10906
rect 2652 10854 2682 10906
rect 2682 10854 2694 10906
rect 2694 10854 2708 10906
rect 2732 10854 2746 10906
rect 2746 10854 2758 10906
rect 2758 10854 2788 10906
rect 2812 10854 2822 10906
rect 2822 10854 2868 10906
rect 2572 10852 2628 10854
rect 2652 10852 2708 10854
rect 2732 10852 2788 10854
rect 2812 10852 2868 10854
rect 2572 9818 2628 9820
rect 2652 9818 2708 9820
rect 2732 9818 2788 9820
rect 2812 9818 2868 9820
rect 2572 9766 2618 9818
rect 2618 9766 2628 9818
rect 2652 9766 2682 9818
rect 2682 9766 2694 9818
rect 2694 9766 2708 9818
rect 2732 9766 2746 9818
rect 2746 9766 2758 9818
rect 2758 9766 2788 9818
rect 2812 9766 2822 9818
rect 2822 9766 2868 9818
rect 2572 9764 2628 9766
rect 2652 9764 2708 9766
rect 2732 9764 2788 9766
rect 2812 9764 2868 9766
rect 2686 8900 2742 8936
rect 2686 8880 2688 8900
rect 2688 8880 2740 8900
rect 2740 8880 2742 8900
rect 2572 8730 2628 8732
rect 2652 8730 2708 8732
rect 2732 8730 2788 8732
rect 2812 8730 2868 8732
rect 2572 8678 2618 8730
rect 2618 8678 2628 8730
rect 2652 8678 2682 8730
rect 2682 8678 2694 8730
rect 2694 8678 2708 8730
rect 2732 8678 2746 8730
rect 2746 8678 2758 8730
rect 2758 8678 2788 8730
rect 2812 8678 2822 8730
rect 2822 8678 2868 8730
rect 2572 8676 2628 8678
rect 2652 8676 2708 8678
rect 2732 8676 2788 8678
rect 2812 8676 2868 8678
rect 2870 7928 2926 7984
rect 2594 7828 2596 7848
rect 2596 7828 2648 7848
rect 2648 7828 2650 7848
rect 2594 7792 2650 7828
rect 2572 7642 2628 7644
rect 2652 7642 2708 7644
rect 2732 7642 2788 7644
rect 2812 7642 2868 7644
rect 2572 7590 2618 7642
rect 2618 7590 2628 7642
rect 2652 7590 2682 7642
rect 2682 7590 2694 7642
rect 2694 7590 2708 7642
rect 2732 7590 2746 7642
rect 2746 7590 2758 7642
rect 2758 7590 2788 7642
rect 2812 7590 2822 7642
rect 2822 7590 2868 7642
rect 2572 7588 2628 7590
rect 2652 7588 2708 7590
rect 2732 7588 2788 7590
rect 2812 7588 2868 7590
rect 3146 9560 3202 9616
rect 3514 9424 3570 9480
rect 3146 8064 3202 8120
rect 2410 7112 2466 7168
rect 2572 6554 2628 6556
rect 2652 6554 2708 6556
rect 2732 6554 2788 6556
rect 2812 6554 2868 6556
rect 2572 6502 2618 6554
rect 2618 6502 2628 6554
rect 2652 6502 2682 6554
rect 2682 6502 2694 6554
rect 2694 6502 2708 6554
rect 2732 6502 2746 6554
rect 2746 6502 2758 6554
rect 2758 6502 2788 6554
rect 2812 6502 2822 6554
rect 2822 6502 2868 6554
rect 2572 6500 2628 6502
rect 2652 6500 2708 6502
rect 2732 6500 2788 6502
rect 2812 6500 2868 6502
rect 3238 7384 3294 7440
rect 3054 7112 3110 7168
rect 2572 5466 2628 5468
rect 2652 5466 2708 5468
rect 2732 5466 2788 5468
rect 2812 5466 2868 5468
rect 2572 5414 2618 5466
rect 2618 5414 2628 5466
rect 2652 5414 2682 5466
rect 2682 5414 2694 5466
rect 2694 5414 2708 5466
rect 2732 5414 2746 5466
rect 2746 5414 2758 5466
rect 2758 5414 2788 5466
rect 2812 5414 2822 5466
rect 2822 5414 2868 5466
rect 2572 5412 2628 5414
rect 2652 5412 2708 5414
rect 2732 5412 2788 5414
rect 2812 5412 2868 5414
rect 3238 6976 3294 7032
rect 2686 3408 2688 3428
rect 2688 3408 2740 3428
rect 2740 3408 2742 3428
rect 2686 3372 2742 3408
rect 3422 4820 3478 4856
rect 3422 4800 3424 4820
rect 3424 4800 3476 4820
rect 3476 4800 3478 4820
rect 2572 1114 2628 1116
rect 2652 1114 2708 1116
rect 2732 1114 2788 1116
rect 2812 1114 2868 1116
rect 2572 1062 2618 1114
rect 2618 1062 2628 1114
rect 2652 1062 2682 1114
rect 2682 1062 2694 1114
rect 2694 1062 2708 1114
rect 2732 1062 2746 1114
rect 2746 1062 2758 1114
rect 2758 1062 2788 1114
rect 2812 1062 2822 1114
rect 2822 1062 2868 1114
rect 2572 1060 2628 1062
rect 2652 1060 2708 1062
rect 2732 1060 2788 1062
rect 2812 1060 2868 1062
rect 3882 11056 3938 11112
rect 3790 10784 3846 10840
rect 3882 10648 3938 10704
rect 3974 9016 4030 9072
rect 3882 8064 3938 8120
rect 4342 9424 4398 9480
rect 4342 8472 4398 8528
rect 10046 12280 10102 12336
rect 4894 10376 4950 10432
rect 4802 9560 4858 9616
rect 4710 6160 4766 6216
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 5312 11450 5368 11452
rect 5072 11398 5118 11450
rect 5118 11398 5128 11450
rect 5152 11398 5182 11450
rect 5182 11398 5194 11450
rect 5194 11398 5208 11450
rect 5232 11398 5246 11450
rect 5246 11398 5258 11450
rect 5258 11398 5288 11450
rect 5312 11398 5322 11450
rect 5322 11398 5368 11450
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 5312 11396 5368 11398
rect 5354 10784 5410 10840
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 5312 10362 5368 10364
rect 5072 10310 5118 10362
rect 5118 10310 5128 10362
rect 5152 10310 5182 10362
rect 5182 10310 5194 10362
rect 5194 10310 5208 10362
rect 5232 10310 5246 10362
rect 5246 10310 5258 10362
rect 5258 10310 5288 10362
rect 5312 10310 5322 10362
rect 5322 10310 5368 10362
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 5312 10308 5368 10310
rect 5446 10240 5502 10296
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 5312 9274 5368 9276
rect 5072 9222 5118 9274
rect 5118 9222 5128 9274
rect 5152 9222 5182 9274
rect 5182 9222 5194 9274
rect 5194 9222 5208 9274
rect 5232 9222 5246 9274
rect 5246 9222 5258 9274
rect 5258 9222 5288 9274
rect 5312 9222 5322 9274
rect 5322 9222 5368 9274
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 5312 9220 5368 9222
rect 4986 8608 5042 8664
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 5312 8186 5368 8188
rect 5072 8134 5118 8186
rect 5118 8134 5128 8186
rect 5152 8134 5182 8186
rect 5182 8134 5194 8186
rect 5194 8134 5208 8186
rect 5232 8134 5246 8186
rect 5246 8134 5258 8186
rect 5258 8134 5288 8186
rect 5312 8134 5322 8186
rect 5322 8134 5368 8186
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 5312 8132 5368 8134
rect 5538 8064 5594 8120
rect 5354 7248 5410 7304
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 5312 7098 5368 7100
rect 5072 7046 5118 7098
rect 5118 7046 5128 7098
rect 5152 7046 5182 7098
rect 5182 7046 5194 7098
rect 5194 7046 5208 7098
rect 5232 7046 5246 7098
rect 5246 7046 5258 7098
rect 5258 7046 5288 7098
rect 5312 7046 5322 7098
rect 5322 7046 5368 7098
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 5312 7044 5368 7046
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 5312 6010 5368 6012
rect 5072 5958 5118 6010
rect 5118 5958 5128 6010
rect 5152 5958 5182 6010
rect 5182 5958 5194 6010
rect 5194 5958 5208 6010
rect 5232 5958 5246 6010
rect 5246 5958 5258 6010
rect 5258 5958 5288 6010
rect 5312 5958 5322 6010
rect 5322 5958 5368 6010
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 5312 5956 5368 5958
rect 5262 5788 5264 5808
rect 5264 5788 5316 5808
rect 5316 5788 5318 5808
rect 5262 5752 5318 5788
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 5312 4922 5368 4924
rect 5072 4870 5118 4922
rect 5118 4870 5128 4922
rect 5152 4870 5182 4922
rect 5182 4870 5194 4922
rect 5194 4870 5208 4922
rect 5232 4870 5246 4922
rect 5246 4870 5258 4922
rect 5258 4870 5288 4922
rect 5312 4870 5322 4922
rect 5322 4870 5368 4922
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 5312 4868 5368 4870
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 5312 3834 5368 3836
rect 5072 3782 5118 3834
rect 5118 3782 5128 3834
rect 5152 3782 5182 3834
rect 5182 3782 5194 3834
rect 5194 3782 5208 3834
rect 5232 3782 5246 3834
rect 5246 3782 5258 3834
rect 5258 3782 5288 3834
rect 5312 3782 5322 3834
rect 5322 3782 5368 3834
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5312 3780 5368 3782
rect 5354 3576 5410 3632
rect 5906 9288 5962 9344
rect 5906 9152 5962 9208
rect 7572 11994 7628 11996
rect 7652 11994 7708 11996
rect 7732 11994 7788 11996
rect 7812 11994 7868 11996
rect 7572 11942 7618 11994
rect 7618 11942 7628 11994
rect 7652 11942 7682 11994
rect 7682 11942 7694 11994
rect 7694 11942 7708 11994
rect 7732 11942 7746 11994
rect 7746 11942 7758 11994
rect 7758 11942 7788 11994
rect 7812 11942 7822 11994
rect 7822 11942 7868 11994
rect 7572 11940 7628 11942
rect 7652 11940 7708 11942
rect 7732 11940 7788 11942
rect 7812 11940 7868 11942
rect 6550 8744 6606 8800
rect 6550 8608 6606 8664
rect 6458 8336 6514 8392
rect 6458 8200 6514 8256
rect 6090 6160 6146 6216
rect 6918 9424 6974 9480
rect 6642 7692 6644 7712
rect 6644 7692 6696 7712
rect 6696 7692 6698 7712
rect 6642 7656 6698 7692
rect 6734 7384 6790 7440
rect 6642 6704 6698 6760
rect 6550 5616 6606 5672
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 5312 2746 5368 2748
rect 5072 2694 5118 2746
rect 5118 2694 5128 2746
rect 5152 2694 5182 2746
rect 5182 2694 5194 2746
rect 5194 2694 5208 2746
rect 5232 2694 5246 2746
rect 5246 2694 5258 2746
rect 5258 2694 5288 2746
rect 5312 2694 5322 2746
rect 5322 2694 5368 2746
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 5312 2692 5368 2694
rect 5072 1658 5128 1660
rect 5152 1658 5208 1660
rect 5232 1658 5288 1660
rect 5312 1658 5368 1660
rect 5072 1606 5118 1658
rect 5118 1606 5128 1658
rect 5152 1606 5182 1658
rect 5182 1606 5194 1658
rect 5194 1606 5208 1658
rect 5232 1606 5246 1658
rect 5246 1606 5258 1658
rect 5258 1606 5288 1658
rect 5312 1606 5322 1658
rect 5322 1606 5368 1658
rect 5072 1604 5128 1606
rect 5152 1604 5208 1606
rect 5232 1604 5288 1606
rect 5312 1604 5368 1606
rect 6550 2760 6606 2816
rect 5078 1264 5134 1320
rect 5446 856 5502 912
rect 6826 7248 6882 7304
rect 6734 4120 6790 4176
rect 7102 9560 7158 9616
rect 7286 8744 7342 8800
rect 7286 8336 7342 8392
rect 7194 7248 7250 7304
rect 7102 4684 7158 4720
rect 7102 4664 7104 4684
rect 7104 4664 7156 4684
rect 7156 4664 7158 4684
rect 6826 2896 6882 2952
rect 6918 2760 6974 2816
rect 7572 10906 7628 10908
rect 7652 10906 7708 10908
rect 7732 10906 7788 10908
rect 7812 10906 7868 10908
rect 7572 10854 7618 10906
rect 7618 10854 7628 10906
rect 7652 10854 7682 10906
rect 7682 10854 7694 10906
rect 7694 10854 7708 10906
rect 7732 10854 7746 10906
rect 7746 10854 7758 10906
rect 7758 10854 7788 10906
rect 7812 10854 7822 10906
rect 7822 10854 7868 10906
rect 7572 10852 7628 10854
rect 7652 10852 7708 10854
rect 7732 10852 7788 10854
rect 7812 10852 7868 10854
rect 7572 9818 7628 9820
rect 7652 9818 7708 9820
rect 7732 9818 7788 9820
rect 7812 9818 7868 9820
rect 7572 9766 7618 9818
rect 7618 9766 7628 9818
rect 7652 9766 7682 9818
rect 7682 9766 7694 9818
rect 7694 9766 7708 9818
rect 7732 9766 7746 9818
rect 7746 9766 7758 9818
rect 7758 9766 7788 9818
rect 7812 9766 7822 9818
rect 7822 9766 7868 9818
rect 7572 9764 7628 9766
rect 7652 9764 7708 9766
rect 7732 9764 7788 9766
rect 7812 9764 7868 9766
rect 7654 9324 7656 9344
rect 7656 9324 7708 9344
rect 7708 9324 7710 9344
rect 7654 9288 7710 9324
rect 7572 8730 7628 8732
rect 7652 8730 7708 8732
rect 7732 8730 7788 8732
rect 7812 8730 7868 8732
rect 7572 8678 7618 8730
rect 7618 8678 7628 8730
rect 7652 8678 7682 8730
rect 7682 8678 7694 8730
rect 7694 8678 7708 8730
rect 7732 8678 7746 8730
rect 7746 8678 7758 8730
rect 7758 8678 7788 8730
rect 7812 8678 7822 8730
rect 7822 8678 7868 8730
rect 7572 8676 7628 8678
rect 7652 8676 7708 8678
rect 7732 8676 7788 8678
rect 7812 8676 7868 8678
rect 7746 8336 7802 8392
rect 7572 7642 7628 7644
rect 7652 7642 7708 7644
rect 7732 7642 7788 7644
rect 7812 7642 7868 7644
rect 7572 7590 7618 7642
rect 7618 7590 7628 7642
rect 7652 7590 7682 7642
rect 7682 7590 7694 7642
rect 7694 7590 7708 7642
rect 7732 7590 7746 7642
rect 7746 7590 7758 7642
rect 7758 7590 7788 7642
rect 7812 7590 7822 7642
rect 7822 7590 7868 7642
rect 7572 7588 7628 7590
rect 7652 7588 7708 7590
rect 7732 7588 7788 7590
rect 7812 7588 7868 7590
rect 7572 6554 7628 6556
rect 7652 6554 7708 6556
rect 7732 6554 7788 6556
rect 7812 6554 7868 6556
rect 7572 6502 7618 6554
rect 7618 6502 7628 6554
rect 7652 6502 7682 6554
rect 7682 6502 7694 6554
rect 7694 6502 7708 6554
rect 7732 6502 7746 6554
rect 7746 6502 7758 6554
rect 7758 6502 7788 6554
rect 7812 6502 7822 6554
rect 7822 6502 7868 6554
rect 7572 6500 7628 6502
rect 7652 6500 7708 6502
rect 7732 6500 7788 6502
rect 7812 6500 7868 6502
rect 8758 11056 8814 11112
rect 8022 8064 8078 8120
rect 8206 9152 8262 9208
rect 8114 7520 8170 7576
rect 7930 5616 7986 5672
rect 7572 5466 7628 5468
rect 7652 5466 7708 5468
rect 7732 5466 7788 5468
rect 7812 5466 7868 5468
rect 7572 5414 7618 5466
rect 7618 5414 7628 5466
rect 7652 5414 7682 5466
rect 7682 5414 7694 5466
rect 7694 5414 7708 5466
rect 7732 5414 7746 5466
rect 7746 5414 7758 5466
rect 7758 5414 7788 5466
rect 7812 5414 7822 5466
rect 7822 5414 7868 5466
rect 7572 5412 7628 5414
rect 7652 5412 7708 5414
rect 7732 5412 7788 5414
rect 7812 5412 7868 5414
rect 7930 5208 7986 5264
rect 7572 4378 7628 4380
rect 7652 4378 7708 4380
rect 7732 4378 7788 4380
rect 7812 4378 7868 4380
rect 7572 4326 7618 4378
rect 7618 4326 7628 4378
rect 7652 4326 7682 4378
rect 7682 4326 7694 4378
rect 7694 4326 7708 4378
rect 7732 4326 7746 4378
rect 7746 4326 7758 4378
rect 7758 4326 7788 4378
rect 7812 4326 7822 4378
rect 7822 4326 7868 4378
rect 7572 4324 7628 4326
rect 7652 4324 7708 4326
rect 7732 4324 7788 4326
rect 7812 4324 7868 4326
rect 7572 3290 7628 3292
rect 7652 3290 7708 3292
rect 7732 3290 7788 3292
rect 7812 3290 7868 3292
rect 7572 3238 7618 3290
rect 7618 3238 7628 3290
rect 7652 3238 7682 3290
rect 7682 3238 7694 3290
rect 7694 3238 7708 3290
rect 7732 3238 7746 3290
rect 7746 3238 7758 3290
rect 7758 3238 7788 3290
rect 7812 3238 7822 3290
rect 7822 3238 7868 3290
rect 7572 3236 7628 3238
rect 7652 3236 7708 3238
rect 7732 3236 7788 3238
rect 7812 3236 7868 3238
rect 7572 2202 7628 2204
rect 7652 2202 7708 2204
rect 7732 2202 7788 2204
rect 7812 2202 7868 2204
rect 7572 2150 7618 2202
rect 7618 2150 7628 2202
rect 7652 2150 7682 2202
rect 7682 2150 7694 2202
rect 7694 2150 7708 2202
rect 7732 2150 7746 2202
rect 7746 2150 7758 2202
rect 7758 2150 7788 2202
rect 7812 2150 7822 2202
rect 7822 2150 7868 2202
rect 7572 2148 7628 2150
rect 7652 2148 7708 2150
rect 7732 2148 7788 2150
rect 7812 2148 7868 2150
rect 8574 10140 8576 10160
rect 8576 10140 8628 10160
rect 8628 10140 8630 10160
rect 8574 10104 8630 10140
rect 8758 8064 8814 8120
rect 8758 7520 8814 7576
rect 8574 6976 8630 7032
rect 8390 5480 8446 5536
rect 7572 1114 7628 1116
rect 7652 1114 7708 1116
rect 7732 1114 7788 1116
rect 7812 1114 7868 1116
rect 7572 1062 7618 1114
rect 7618 1062 7628 1114
rect 7652 1062 7682 1114
rect 7682 1062 7694 1114
rect 7694 1062 7708 1114
rect 7732 1062 7746 1114
rect 7746 1062 7758 1114
rect 7758 1062 7788 1114
rect 7812 1062 7822 1114
rect 7822 1062 7868 1114
rect 7572 1060 7628 1062
rect 7652 1060 7708 1062
rect 7732 1060 7788 1062
rect 7812 1060 7868 1062
rect 8942 8492 8998 8528
rect 8942 8472 8944 8492
rect 8944 8472 8996 8492
rect 8996 8472 8998 8492
rect 8942 7112 8998 7168
rect 9310 7268 9366 7304
rect 9310 7248 9312 7268
rect 9312 7248 9364 7268
rect 9364 7248 9366 7268
rect 8942 2488 8998 2544
rect 5072 570 5128 572
rect 5152 570 5208 572
rect 5232 570 5288 572
rect 5312 570 5368 572
rect 5072 518 5118 570
rect 5118 518 5128 570
rect 5152 518 5182 570
rect 5182 518 5194 570
rect 5194 518 5208 570
rect 5232 518 5246 570
rect 5246 518 5258 570
rect 5258 518 5288 570
rect 5312 518 5322 570
rect 5322 518 5368 570
rect 5072 516 5128 518
rect 5152 516 5208 518
rect 5232 516 5288 518
rect 5312 516 5368 518
rect 9034 1672 9090 1728
rect 9678 9288 9734 9344
rect 20718 11872 20774 11928
rect 10138 9832 10194 9888
rect 19338 11056 19394 11112
rect 12438 6568 12494 6624
rect 10690 6160 10746 6216
rect 19338 6976 19394 7032
rect 16946 5752 17002 5808
rect 16578 5344 16634 5400
rect 16670 4936 16726 4992
rect 16854 4528 16910 4584
rect 16670 3304 16726 3360
rect 16578 2080 16634 2136
rect 16762 2488 16818 2544
rect 5446 448 5502 504
<< metal3 >>
rect 10041 12338 10107 12341
rect 14000 12338 34000 12368
rect 10041 12336 34000 12338
rect 10041 12280 10046 12336
rect 10102 12280 34000 12336
rect 10041 12278 34000 12280
rect 10041 12275 10107 12278
rect 14000 12248 34000 12278
rect 2562 12000 2878 12001
rect 2562 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2878 12000
rect 2562 11935 2878 11936
rect 7562 12000 7878 12001
rect 7562 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7878 12000
rect 7562 11935 7878 11936
rect 14000 11928 34000 11960
rect 14000 11872 20718 11928
rect 20774 11872 34000 11928
rect 14000 11840 34000 11872
rect 2497 11658 2563 11661
rect 2497 11656 12450 11658
rect 2497 11600 2502 11656
rect 2558 11600 12450 11656
rect 2497 11598 12450 11600
rect 2497 11595 2563 11598
rect 12390 11522 12450 11598
rect 14000 11522 34000 11552
rect 12390 11462 34000 11522
rect 5062 11456 5378 11457
rect 5062 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5378 11456
rect 14000 11432 34000 11462
rect 5062 11391 5378 11392
rect 1669 11114 1735 11117
rect 3877 11114 3943 11117
rect 8753 11114 8819 11117
rect 1669 11112 8819 11114
rect 1669 11056 1674 11112
rect 1730 11056 3882 11112
rect 3938 11056 8758 11112
rect 8814 11056 8819 11112
rect 1669 11054 8819 11056
rect 1669 11051 1735 11054
rect 3877 11051 3943 11054
rect 8753 11051 8819 11054
rect 14000 11112 34000 11144
rect 14000 11056 19338 11112
rect 19394 11056 34000 11112
rect 14000 11024 34000 11056
rect 2562 10912 2878 10913
rect 2562 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2878 10912
rect 2562 10847 2878 10848
rect 7562 10912 7878 10913
rect 7562 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7878 10912
rect 7562 10847 7878 10848
rect 3785 10842 3851 10845
rect 5349 10842 5415 10845
rect 3785 10840 5415 10842
rect 3785 10784 3790 10840
rect 3846 10784 5354 10840
rect 5410 10784 5415 10840
rect 3785 10782 5415 10784
rect 3785 10779 3851 10782
rect 5349 10779 5415 10782
rect 1209 10706 1275 10709
rect 3877 10706 3943 10709
rect 14000 10706 34000 10736
rect 1209 10704 2790 10706
rect 1209 10648 1214 10704
rect 1270 10648 2790 10704
rect 1209 10646 2790 10648
rect 1209 10643 1275 10646
rect 2730 10162 2790 10646
rect 3877 10704 34000 10706
rect 3877 10648 3882 10704
rect 3938 10648 34000 10704
rect 3877 10646 34000 10648
rect 3877 10643 3943 10646
rect 14000 10616 34000 10646
rect 2998 10372 3004 10436
rect 3068 10434 3074 10436
rect 4889 10434 4955 10437
rect 3068 10432 4955 10434
rect 3068 10376 4894 10432
rect 4950 10376 4955 10432
rect 3068 10374 4955 10376
rect 3068 10372 3074 10374
rect 4889 10371 4955 10374
rect 5062 10368 5378 10369
rect 5062 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5378 10368
rect 5062 10303 5378 10304
rect 5441 10298 5507 10301
rect 14000 10298 34000 10328
rect 5441 10296 34000 10298
rect 5441 10240 5446 10296
rect 5502 10240 34000 10296
rect 5441 10238 34000 10240
rect 5441 10235 5507 10238
rect 14000 10208 34000 10238
rect 8569 10162 8635 10165
rect 2730 10160 8635 10162
rect 2730 10104 8574 10160
rect 8630 10104 8635 10160
rect 2730 10102 8635 10104
rect 8569 10099 8635 10102
rect 10133 9890 10199 9893
rect 14000 9890 34000 9920
rect 10133 9888 34000 9890
rect 10133 9832 10138 9888
rect 10194 9832 34000 9888
rect 10133 9830 34000 9832
rect 10133 9827 10199 9830
rect 2562 9824 2878 9825
rect 2562 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2878 9824
rect 2562 9759 2878 9760
rect 7562 9824 7878 9825
rect 7562 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7878 9824
rect 14000 9800 34000 9830
rect 7562 9759 7878 9760
rect 3141 9618 3207 9621
rect 3366 9618 3372 9620
rect 3141 9616 3372 9618
rect 3141 9560 3146 9616
rect 3202 9560 3372 9616
rect 3141 9558 3372 9560
rect 3141 9555 3207 9558
rect 3366 9556 3372 9558
rect 3436 9618 3442 9620
rect 3436 9558 4538 9618
rect 3436 9556 3442 9558
rect 1301 9482 1367 9485
rect 3509 9482 3575 9485
rect 4337 9482 4403 9485
rect 1301 9480 4403 9482
rect 1301 9424 1306 9480
rect 1362 9424 3514 9480
rect 3570 9424 4342 9480
rect 4398 9424 4403 9480
rect 1301 9422 4403 9424
rect 4478 9482 4538 9558
rect 4654 9556 4660 9620
rect 4724 9618 4730 9620
rect 4797 9618 4863 9621
rect 7097 9618 7163 9621
rect 4724 9616 4863 9618
rect 4724 9560 4802 9616
rect 4858 9560 4863 9616
rect 4724 9558 4863 9560
rect 4724 9556 4730 9558
rect 4797 9555 4863 9558
rect 5030 9616 7163 9618
rect 5030 9560 7102 9616
rect 7158 9560 7163 9616
rect 5030 9558 7163 9560
rect 5030 9482 5090 9558
rect 7097 9555 7163 9558
rect 4478 9422 5090 9482
rect 6913 9482 6979 9485
rect 14000 9482 34000 9512
rect 6913 9480 34000 9482
rect 6913 9424 6918 9480
rect 6974 9424 34000 9480
rect 6913 9422 34000 9424
rect 1301 9419 1367 9422
rect 3509 9419 3575 9422
rect 4337 9419 4403 9422
rect 6913 9419 6979 9422
rect 14000 9392 34000 9422
rect 5901 9346 5967 9349
rect 7649 9346 7715 9349
rect 5901 9344 7715 9346
rect 5901 9288 5906 9344
rect 5962 9288 7654 9344
rect 7710 9288 7715 9344
rect 5901 9286 7715 9288
rect 5901 9283 5967 9286
rect 7649 9283 7715 9286
rect 9070 9284 9076 9348
rect 9140 9346 9146 9348
rect 9673 9346 9739 9349
rect 9140 9344 9739 9346
rect 9140 9288 9678 9344
rect 9734 9288 9739 9344
rect 9140 9286 9739 9288
rect 9140 9284 9146 9286
rect 9673 9283 9739 9286
rect 5062 9280 5378 9281
rect 5062 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5378 9280
rect 5062 9215 5378 9216
rect 5901 9210 5967 9213
rect 7046 9210 7052 9212
rect 5901 9208 7052 9210
rect 5901 9152 5906 9208
rect 5962 9152 7052 9208
rect 5901 9150 7052 9152
rect 5901 9147 5967 9150
rect 7046 9148 7052 9150
rect 7116 9210 7122 9212
rect 8201 9210 8267 9213
rect 7116 9208 8267 9210
rect 7116 9152 8206 9208
rect 8262 9152 8267 9208
rect 7116 9150 8267 9152
rect 7116 9148 7122 9150
rect 8201 9147 8267 9150
rect 3969 9074 4035 9077
rect 14000 9074 34000 9104
rect 3969 9072 34000 9074
rect 3969 9016 3974 9072
rect 4030 9016 34000 9072
rect 3969 9014 34000 9016
rect 3969 9011 4035 9014
rect 14000 8984 34000 9014
rect 2681 8938 2747 8941
rect 2681 8936 12450 8938
rect 2681 8880 2686 8936
rect 2742 8880 12450 8936
rect 2681 8878 12450 8880
rect 2681 8875 2747 8878
rect 6545 8802 6611 8805
rect 7281 8802 7347 8805
rect 3236 8800 7347 8802
rect 3236 8744 6550 8800
rect 6606 8744 7286 8800
rect 7342 8744 7347 8800
rect 3236 8742 7347 8744
rect 2562 8736 2878 8737
rect 2562 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2878 8736
rect 2562 8671 2878 8672
rect 1577 8530 1643 8533
rect 3236 8530 3296 8742
rect 6545 8739 6611 8742
rect 7281 8739 7347 8742
rect 7562 8736 7878 8737
rect 7562 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7878 8736
rect 7562 8671 7878 8672
rect 4981 8666 5047 8669
rect 6545 8666 6611 8669
rect 4981 8664 6611 8666
rect 4981 8608 4986 8664
rect 5042 8608 6550 8664
rect 6606 8608 6611 8664
rect 4981 8606 6611 8608
rect 12390 8666 12450 8878
rect 14000 8666 34000 8696
rect 12390 8606 34000 8666
rect 4981 8603 5047 8606
rect 6545 8603 6611 8606
rect 14000 8576 34000 8606
rect 1577 8528 3296 8530
rect 1577 8472 1582 8528
rect 1638 8472 3296 8528
rect 1577 8470 3296 8472
rect 4337 8530 4403 8533
rect 8937 8530 9003 8533
rect 4337 8528 9003 8530
rect 4337 8472 4342 8528
rect 4398 8472 8942 8528
rect 8998 8472 9003 8528
rect 4337 8470 9003 8472
rect 1577 8467 1643 8470
rect 4337 8467 4403 8470
rect 8937 8467 9003 8470
rect 6453 8396 6519 8397
rect 6453 8394 6500 8396
rect 6408 8392 6500 8394
rect 6408 8336 6458 8392
rect 6408 8334 6500 8336
rect 6453 8332 6500 8334
rect 6564 8332 6570 8396
rect 7281 8394 7347 8397
rect 7741 8394 7807 8397
rect 7281 8392 7807 8394
rect 7281 8336 7286 8392
rect 7342 8336 7746 8392
rect 7802 8336 7807 8392
rect 7281 8334 7807 8336
rect 6453 8331 6519 8332
rect 7281 8331 7347 8334
rect 7741 8331 7807 8334
rect 6453 8258 6519 8261
rect 14000 8258 34000 8288
rect 6453 8256 34000 8258
rect 6453 8200 6458 8256
rect 6514 8200 34000 8256
rect 6453 8198 34000 8200
rect 6453 8195 6519 8198
rect 5062 8192 5378 8193
rect 5062 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5378 8192
rect 14000 8168 34000 8198
rect 5062 8127 5378 8128
rect 2998 8122 3004 8124
rect 2730 8062 3004 8122
rect 1209 7986 1275 7989
rect 2730 7986 2790 8062
rect 2998 8060 3004 8062
rect 3068 8060 3074 8124
rect 3141 8122 3207 8125
rect 3877 8122 3943 8125
rect 3141 8120 3943 8122
rect 3141 8064 3146 8120
rect 3202 8064 3882 8120
rect 3938 8064 3943 8120
rect 3141 8062 3943 8064
rect 3141 8059 3207 8062
rect 3877 8059 3943 8062
rect 5533 8122 5599 8125
rect 8017 8122 8083 8125
rect 8753 8122 8819 8125
rect 5533 8120 8819 8122
rect 5533 8064 5538 8120
rect 5594 8064 8022 8120
rect 8078 8064 8758 8120
rect 8814 8064 8819 8120
rect 5533 8062 8819 8064
rect 5533 8059 5599 8062
rect 8017 8059 8083 8062
rect 8753 8059 8819 8062
rect 1209 7984 2790 7986
rect 1209 7928 1214 7984
rect 1270 7928 2790 7984
rect 1209 7926 2790 7928
rect 2865 7986 2931 7989
rect 9070 7986 9076 7988
rect 2865 7984 9076 7986
rect 2865 7928 2870 7984
rect 2926 7928 9076 7984
rect 2865 7926 9076 7928
rect 1209 7923 1275 7926
rect 2865 7923 2931 7926
rect 9070 7924 9076 7926
rect 9140 7924 9146 7988
rect 2589 7850 2655 7853
rect 14000 7850 34000 7880
rect 2589 7848 34000 7850
rect 2589 7792 2594 7848
rect 2650 7792 34000 7848
rect 2589 7790 34000 7792
rect 2589 7787 2655 7790
rect 14000 7760 34000 7790
rect 2998 7652 3004 7716
rect 3068 7714 3074 7716
rect 6637 7714 6703 7717
rect 3068 7712 6703 7714
rect 3068 7656 6642 7712
rect 6698 7656 6703 7712
rect 3068 7654 6703 7656
rect 3068 7652 3074 7654
rect 6637 7651 6703 7654
rect 2562 7648 2878 7649
rect 2562 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2878 7648
rect 2562 7583 2878 7584
rect 7562 7648 7878 7649
rect 7562 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7878 7648
rect 7562 7583 7878 7584
rect 8109 7578 8175 7581
rect 8753 7578 8819 7581
rect 8109 7576 8819 7578
rect 8109 7520 8114 7576
rect 8170 7520 8758 7576
rect 8814 7520 8819 7576
rect 8109 7518 8819 7520
rect 8109 7515 8175 7518
rect 8753 7515 8819 7518
rect 3233 7442 3299 7445
rect 3190 7440 3299 7442
rect 3190 7384 3238 7440
rect 3294 7384 3299 7440
rect 3190 7379 3299 7384
rect 6729 7442 6795 7445
rect 14000 7442 34000 7472
rect 6729 7440 34000 7442
rect 6729 7384 6734 7440
rect 6790 7384 34000 7440
rect 6729 7382 34000 7384
rect 6729 7379 6795 7382
rect 2405 7170 2471 7173
rect 3049 7170 3115 7173
rect 2405 7168 3115 7170
rect 2405 7112 2410 7168
rect 2466 7112 3054 7168
rect 3110 7112 3115 7168
rect 2405 7110 3115 7112
rect 2405 7107 2471 7110
rect 3049 7107 3115 7110
rect 3190 7037 3250 7379
rect 14000 7352 34000 7382
rect 5349 7306 5415 7309
rect 6821 7306 6887 7309
rect 5349 7304 6887 7306
rect 5349 7248 5354 7304
rect 5410 7248 6826 7304
rect 6882 7248 6887 7304
rect 5349 7246 6887 7248
rect 5349 7243 5415 7246
rect 6821 7243 6887 7246
rect 7189 7306 7255 7309
rect 9305 7306 9371 7309
rect 7189 7304 9371 7306
rect 7189 7248 7194 7304
rect 7250 7248 9310 7304
rect 9366 7248 9371 7304
rect 7189 7246 9371 7248
rect 7189 7243 7255 7246
rect 9305 7243 9371 7246
rect 5574 7108 5580 7172
rect 5644 7170 5650 7172
rect 8937 7170 9003 7173
rect 5644 7168 9003 7170
rect 5644 7112 8942 7168
rect 8998 7112 9003 7168
rect 5644 7110 9003 7112
rect 5644 7108 5650 7110
rect 8937 7107 9003 7110
rect 5062 7104 5378 7105
rect 5062 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5378 7104
rect 5062 7039 5378 7040
rect 3190 7032 3299 7037
rect 8569 7034 8635 7037
rect 3190 6976 3238 7032
rect 3294 6976 3299 7032
rect 3190 6974 3299 6976
rect 3233 6971 3299 6974
rect 8526 7032 8635 7034
rect 8526 6976 8574 7032
rect 8630 6976 8635 7032
rect 8526 6971 8635 6976
rect 14000 7032 34000 7064
rect 14000 6976 19338 7032
rect 19394 6976 34000 7032
rect 6637 6762 6703 6765
rect 6318 6760 6703 6762
rect 6318 6704 6642 6760
rect 6698 6704 6703 6760
rect 6318 6702 6703 6704
rect 2562 6560 2878 6561
rect 2562 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2878 6560
rect 2562 6495 2878 6496
rect 4705 6220 4771 6221
rect 4654 6156 4660 6220
rect 4724 6218 4771 6220
rect 6085 6218 6151 6221
rect 6318 6218 6378 6702
rect 6637 6699 6703 6702
rect 7562 6560 7878 6561
rect 7562 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7878 6560
rect 7562 6495 7878 6496
rect 4724 6216 4816 6218
rect 4766 6160 4816 6216
rect 4724 6158 4816 6160
rect 6085 6216 6378 6218
rect 6085 6160 6090 6216
rect 6146 6160 6378 6216
rect 6085 6158 6378 6160
rect 4724 6156 4771 6158
rect 4705 6155 4771 6156
rect 6085 6155 6151 6158
rect 5062 6016 5378 6017
rect 5062 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5378 6016
rect 5062 5951 5378 5952
rect 5257 5810 5323 5813
rect 5574 5810 5580 5812
rect 5257 5808 5580 5810
rect 5257 5752 5262 5808
rect 5318 5752 5580 5808
rect 5257 5750 5580 5752
rect 5257 5747 5323 5750
rect 5574 5748 5580 5750
rect 5644 5748 5650 5812
rect 6545 5676 6611 5677
rect 6494 5674 6500 5676
rect 6454 5614 6500 5674
rect 6564 5672 6611 5676
rect 6606 5616 6611 5672
rect 6494 5612 6500 5614
rect 6564 5612 6611 5616
rect 6545 5611 6611 5612
rect 7925 5674 7991 5677
rect 7925 5672 8034 5674
rect 7925 5616 7930 5672
rect 7986 5616 8034 5672
rect 7925 5611 8034 5616
rect 2562 5472 2878 5473
rect 2562 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2878 5472
rect 2562 5407 2878 5408
rect 7562 5472 7878 5473
rect 7562 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7878 5472
rect 7562 5407 7878 5408
rect 7974 5269 8034 5611
rect 8385 5538 8451 5541
rect 8526 5538 8586 6971
rect 14000 6944 34000 6976
rect 12433 6626 12499 6629
rect 14000 6626 34000 6656
rect 12433 6624 34000 6626
rect 12433 6568 12438 6624
rect 12494 6568 34000 6624
rect 12433 6566 34000 6568
rect 12433 6563 12499 6566
rect 14000 6536 34000 6566
rect 10685 6218 10751 6221
rect 14000 6218 34000 6248
rect 10685 6216 34000 6218
rect 10685 6160 10690 6216
rect 10746 6160 34000 6216
rect 10685 6158 34000 6160
rect 10685 6155 10751 6158
rect 14000 6128 34000 6158
rect 14000 5808 34000 5840
rect 14000 5752 16946 5808
rect 17002 5752 34000 5808
rect 14000 5720 34000 5752
rect 8385 5536 8586 5538
rect 8385 5480 8390 5536
rect 8446 5480 8586 5536
rect 8385 5478 8586 5480
rect 8385 5475 8451 5478
rect 14000 5400 34000 5432
rect 14000 5344 16578 5400
rect 16634 5344 34000 5400
rect 14000 5312 34000 5344
rect 7925 5264 8034 5269
rect 7925 5208 7930 5264
rect 7986 5208 8034 5264
rect 7925 5206 8034 5208
rect 7925 5203 7991 5206
rect 14000 4992 34000 5024
rect 14000 4936 16670 4992
rect 16726 4936 34000 4992
rect 5062 4928 5378 4929
rect 5062 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5378 4928
rect 14000 4904 34000 4936
rect 5062 4863 5378 4864
rect 3417 4860 3483 4861
rect 3366 4796 3372 4860
rect 3436 4858 3483 4860
rect 3436 4856 3528 4858
rect 3478 4800 3528 4856
rect 3436 4798 3528 4800
rect 3436 4796 3483 4798
rect 3417 4795 3483 4796
rect 7097 4724 7163 4725
rect 7046 4660 7052 4724
rect 7116 4722 7163 4724
rect 7116 4720 7208 4722
rect 7158 4664 7208 4720
rect 7116 4662 7208 4664
rect 7116 4660 7163 4662
rect 7097 4659 7163 4660
rect 14000 4584 34000 4616
rect 14000 4528 16854 4584
rect 16910 4528 34000 4584
rect 14000 4496 34000 4528
rect 7562 4384 7878 4385
rect 7562 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7878 4384
rect 7562 4319 7878 4320
rect 6729 4178 6795 4181
rect 14000 4178 34000 4208
rect 6729 4176 34000 4178
rect 6729 4120 6734 4176
rect 6790 4120 34000 4176
rect 6729 4118 34000 4120
rect 6729 4115 6795 4118
rect 14000 4088 34000 4118
rect 5062 3840 5378 3841
rect 5062 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5378 3840
rect 5062 3775 5378 3776
rect 14000 3770 34000 3800
rect 12390 3710 34000 3770
rect 5349 3634 5415 3637
rect 12390 3634 12450 3710
rect 14000 3680 34000 3710
rect 5349 3632 12450 3634
rect 5349 3576 5354 3632
rect 5410 3576 12450 3632
rect 5349 3574 12450 3576
rect 5349 3571 5415 3574
rect 2681 3430 2747 3433
rect 2484 3428 2747 3430
rect 2484 3372 2686 3428
rect 2742 3372 2747 3428
rect 2484 3370 2747 3372
rect 2681 3367 2747 3370
rect 14000 3360 34000 3392
rect 14000 3304 16670 3360
rect 16726 3304 34000 3360
rect 7562 3296 7878 3297
rect 7562 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7878 3296
rect 14000 3272 34000 3304
rect 7562 3231 7878 3232
rect 6821 2954 6887 2957
rect 14000 2954 34000 2984
rect 6821 2952 34000 2954
rect 6821 2896 6826 2952
rect 6882 2896 34000 2952
rect 6821 2894 34000 2896
rect 6821 2891 6887 2894
rect 14000 2864 34000 2894
rect 6545 2818 6611 2821
rect 6913 2818 6979 2821
rect 6545 2816 6979 2818
rect 6545 2760 6550 2816
rect 6606 2760 6918 2816
rect 6974 2760 6979 2816
rect 6545 2758 6979 2760
rect 6545 2755 6611 2758
rect 6913 2755 6979 2758
rect 5062 2752 5378 2753
rect 5062 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5378 2752
rect 5062 2687 5378 2688
rect 8937 2546 9003 2549
rect 9070 2546 9076 2548
rect 8937 2544 9076 2546
rect 8937 2488 8942 2544
rect 8998 2488 9076 2544
rect 8937 2486 9076 2488
rect 8937 2483 9003 2486
rect 9070 2484 9076 2486
rect 9140 2484 9146 2548
rect 14000 2544 34000 2576
rect 14000 2488 16762 2544
rect 16818 2488 34000 2544
rect 14000 2456 34000 2488
rect 7562 2208 7878 2209
rect 7562 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7878 2208
rect 7562 2143 7878 2144
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 9029 1730 9095 1733
rect 14000 1730 34000 1760
rect 9029 1728 34000 1730
rect 9029 1672 9034 1728
rect 9090 1672 34000 1728
rect 9029 1670 34000 1672
rect 9029 1667 9095 1670
rect 5062 1664 5378 1665
rect 5062 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5378 1664
rect 14000 1640 34000 1670
rect 5062 1599 5378 1600
rect 5073 1322 5139 1325
rect 14000 1322 34000 1352
rect 5073 1320 34000 1322
rect 5073 1264 5078 1320
rect 5134 1264 34000 1320
rect 5073 1262 34000 1264
rect 5073 1259 5139 1262
rect 14000 1232 34000 1262
rect 2562 1120 2878 1121
rect 2562 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2878 1120
rect 2562 1055 2878 1056
rect 7562 1120 7878 1121
rect 7562 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7878 1120
rect 7562 1055 7878 1056
rect 5441 914 5507 917
rect 14000 914 34000 944
rect 5441 912 34000 914
rect 5441 856 5446 912
rect 5502 856 34000 912
rect 5441 854 34000 856
rect 5441 851 5507 854
rect 14000 824 34000 854
rect 5062 576 5378 577
rect 5062 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5378 576
rect 5062 511 5378 512
rect 5441 506 5507 509
rect 14000 506 34000 536
rect 5441 504 34000 506
rect 5441 448 5446 504
rect 5502 448 34000 504
rect 5441 446 34000 448
rect 5441 443 5507 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11996 2632 12000
rect 2568 11940 2572 11996
rect 2572 11940 2628 11996
rect 2628 11940 2632 11996
rect 2568 11936 2632 11940
rect 2648 11996 2712 12000
rect 2648 11940 2652 11996
rect 2652 11940 2708 11996
rect 2708 11940 2712 11996
rect 2648 11936 2712 11940
rect 2728 11996 2792 12000
rect 2728 11940 2732 11996
rect 2732 11940 2788 11996
rect 2788 11940 2792 11996
rect 2728 11936 2792 11940
rect 2808 11996 2872 12000
rect 2808 11940 2812 11996
rect 2812 11940 2868 11996
rect 2868 11940 2872 11996
rect 2808 11936 2872 11940
rect 7568 11996 7632 12000
rect 7568 11940 7572 11996
rect 7572 11940 7628 11996
rect 7628 11940 7632 11996
rect 7568 11936 7632 11940
rect 7648 11996 7712 12000
rect 7648 11940 7652 11996
rect 7652 11940 7708 11996
rect 7708 11940 7712 11996
rect 7648 11936 7712 11940
rect 7728 11996 7792 12000
rect 7728 11940 7732 11996
rect 7732 11940 7788 11996
rect 7788 11940 7792 11996
rect 7728 11936 7792 11940
rect 7808 11996 7872 12000
rect 7808 11940 7812 11996
rect 7812 11940 7868 11996
rect 7868 11940 7872 11996
rect 7808 11936 7872 11940
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 5308 11452 5372 11456
rect 5308 11396 5312 11452
rect 5312 11396 5368 11452
rect 5368 11396 5372 11452
rect 5308 11392 5372 11396
rect 2568 10908 2632 10912
rect 2568 10852 2572 10908
rect 2572 10852 2628 10908
rect 2628 10852 2632 10908
rect 2568 10848 2632 10852
rect 2648 10908 2712 10912
rect 2648 10852 2652 10908
rect 2652 10852 2708 10908
rect 2708 10852 2712 10908
rect 2648 10848 2712 10852
rect 2728 10908 2792 10912
rect 2728 10852 2732 10908
rect 2732 10852 2788 10908
rect 2788 10852 2792 10908
rect 2728 10848 2792 10852
rect 2808 10908 2872 10912
rect 2808 10852 2812 10908
rect 2812 10852 2868 10908
rect 2868 10852 2872 10908
rect 2808 10848 2872 10852
rect 7568 10908 7632 10912
rect 7568 10852 7572 10908
rect 7572 10852 7628 10908
rect 7628 10852 7632 10908
rect 7568 10848 7632 10852
rect 7648 10908 7712 10912
rect 7648 10852 7652 10908
rect 7652 10852 7708 10908
rect 7708 10852 7712 10908
rect 7648 10848 7712 10852
rect 7728 10908 7792 10912
rect 7728 10852 7732 10908
rect 7732 10852 7788 10908
rect 7788 10852 7792 10908
rect 7728 10848 7792 10852
rect 7808 10908 7872 10912
rect 7808 10852 7812 10908
rect 7812 10852 7868 10908
rect 7868 10852 7872 10908
rect 7808 10848 7872 10852
rect 3004 10372 3068 10436
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 5308 10364 5372 10368
rect 5308 10308 5312 10364
rect 5312 10308 5368 10364
rect 5368 10308 5372 10364
rect 5308 10304 5372 10308
rect 2568 9820 2632 9824
rect 2568 9764 2572 9820
rect 2572 9764 2628 9820
rect 2628 9764 2632 9820
rect 2568 9760 2632 9764
rect 2648 9820 2712 9824
rect 2648 9764 2652 9820
rect 2652 9764 2708 9820
rect 2708 9764 2712 9820
rect 2648 9760 2712 9764
rect 2728 9820 2792 9824
rect 2728 9764 2732 9820
rect 2732 9764 2788 9820
rect 2788 9764 2792 9820
rect 2728 9760 2792 9764
rect 2808 9820 2872 9824
rect 2808 9764 2812 9820
rect 2812 9764 2868 9820
rect 2868 9764 2872 9820
rect 2808 9760 2872 9764
rect 7568 9820 7632 9824
rect 7568 9764 7572 9820
rect 7572 9764 7628 9820
rect 7628 9764 7632 9820
rect 7568 9760 7632 9764
rect 7648 9820 7712 9824
rect 7648 9764 7652 9820
rect 7652 9764 7708 9820
rect 7708 9764 7712 9820
rect 7648 9760 7712 9764
rect 7728 9820 7792 9824
rect 7728 9764 7732 9820
rect 7732 9764 7788 9820
rect 7788 9764 7792 9820
rect 7728 9760 7792 9764
rect 7808 9820 7872 9824
rect 7808 9764 7812 9820
rect 7812 9764 7868 9820
rect 7868 9764 7872 9820
rect 7808 9760 7872 9764
rect 3372 9556 3436 9620
rect 4660 9556 4724 9620
rect 9076 9284 9140 9348
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 5308 9276 5372 9280
rect 5308 9220 5312 9276
rect 5312 9220 5368 9276
rect 5368 9220 5372 9276
rect 5308 9216 5372 9220
rect 7052 9148 7116 9212
rect 2568 8732 2632 8736
rect 2568 8676 2572 8732
rect 2572 8676 2628 8732
rect 2628 8676 2632 8732
rect 2568 8672 2632 8676
rect 2648 8732 2712 8736
rect 2648 8676 2652 8732
rect 2652 8676 2708 8732
rect 2708 8676 2712 8732
rect 2648 8672 2712 8676
rect 2728 8732 2792 8736
rect 2728 8676 2732 8732
rect 2732 8676 2788 8732
rect 2788 8676 2792 8732
rect 2728 8672 2792 8676
rect 2808 8732 2872 8736
rect 2808 8676 2812 8732
rect 2812 8676 2868 8732
rect 2868 8676 2872 8732
rect 2808 8672 2872 8676
rect 7568 8732 7632 8736
rect 7568 8676 7572 8732
rect 7572 8676 7628 8732
rect 7628 8676 7632 8732
rect 7568 8672 7632 8676
rect 7648 8732 7712 8736
rect 7648 8676 7652 8732
rect 7652 8676 7708 8732
rect 7708 8676 7712 8732
rect 7648 8672 7712 8676
rect 7728 8732 7792 8736
rect 7728 8676 7732 8732
rect 7732 8676 7788 8732
rect 7788 8676 7792 8732
rect 7728 8672 7792 8676
rect 7808 8732 7872 8736
rect 7808 8676 7812 8732
rect 7812 8676 7868 8732
rect 7868 8676 7872 8732
rect 7808 8672 7872 8676
rect 6500 8392 6564 8396
rect 6500 8336 6514 8392
rect 6514 8336 6564 8392
rect 6500 8332 6564 8336
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 5308 8188 5372 8192
rect 5308 8132 5312 8188
rect 5312 8132 5368 8188
rect 5368 8132 5372 8188
rect 5308 8128 5372 8132
rect 3004 8060 3068 8124
rect 9076 7924 9140 7988
rect 3004 7652 3068 7716
rect 2568 7644 2632 7648
rect 2568 7588 2572 7644
rect 2572 7588 2628 7644
rect 2628 7588 2632 7644
rect 2568 7584 2632 7588
rect 2648 7644 2712 7648
rect 2648 7588 2652 7644
rect 2652 7588 2708 7644
rect 2708 7588 2712 7644
rect 2648 7584 2712 7588
rect 2728 7644 2792 7648
rect 2728 7588 2732 7644
rect 2732 7588 2788 7644
rect 2788 7588 2792 7644
rect 2728 7584 2792 7588
rect 2808 7644 2872 7648
rect 2808 7588 2812 7644
rect 2812 7588 2868 7644
rect 2868 7588 2872 7644
rect 2808 7584 2872 7588
rect 7568 7644 7632 7648
rect 7568 7588 7572 7644
rect 7572 7588 7628 7644
rect 7628 7588 7632 7644
rect 7568 7584 7632 7588
rect 7648 7644 7712 7648
rect 7648 7588 7652 7644
rect 7652 7588 7708 7644
rect 7708 7588 7712 7644
rect 7648 7584 7712 7588
rect 7728 7644 7792 7648
rect 7728 7588 7732 7644
rect 7732 7588 7788 7644
rect 7788 7588 7792 7644
rect 7728 7584 7792 7588
rect 7808 7644 7872 7648
rect 7808 7588 7812 7644
rect 7812 7588 7868 7644
rect 7868 7588 7872 7644
rect 7808 7584 7872 7588
rect 5580 7108 5644 7172
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 5308 7100 5372 7104
rect 5308 7044 5312 7100
rect 5312 7044 5368 7100
rect 5368 7044 5372 7100
rect 5308 7040 5372 7044
rect 2568 6556 2632 6560
rect 2568 6500 2572 6556
rect 2572 6500 2628 6556
rect 2628 6500 2632 6556
rect 2568 6496 2632 6500
rect 2648 6556 2712 6560
rect 2648 6500 2652 6556
rect 2652 6500 2708 6556
rect 2708 6500 2712 6556
rect 2648 6496 2712 6500
rect 2728 6556 2792 6560
rect 2728 6500 2732 6556
rect 2732 6500 2788 6556
rect 2788 6500 2792 6556
rect 2728 6496 2792 6500
rect 2808 6556 2872 6560
rect 2808 6500 2812 6556
rect 2812 6500 2868 6556
rect 2868 6500 2872 6556
rect 2808 6496 2872 6500
rect 4660 6216 4724 6220
rect 7568 6556 7632 6560
rect 7568 6500 7572 6556
rect 7572 6500 7628 6556
rect 7628 6500 7632 6556
rect 7568 6496 7632 6500
rect 7648 6556 7712 6560
rect 7648 6500 7652 6556
rect 7652 6500 7708 6556
rect 7708 6500 7712 6556
rect 7648 6496 7712 6500
rect 7728 6556 7792 6560
rect 7728 6500 7732 6556
rect 7732 6500 7788 6556
rect 7788 6500 7792 6556
rect 7728 6496 7792 6500
rect 7808 6556 7872 6560
rect 7808 6500 7812 6556
rect 7812 6500 7868 6556
rect 7868 6500 7872 6556
rect 7808 6496 7872 6500
rect 4660 6160 4710 6216
rect 4710 6160 4724 6216
rect 4660 6156 4724 6160
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 5308 6012 5372 6016
rect 5308 5956 5312 6012
rect 5312 5956 5368 6012
rect 5368 5956 5372 6012
rect 5308 5952 5372 5956
rect 5580 5748 5644 5812
rect 6500 5672 6564 5676
rect 6500 5616 6550 5672
rect 6550 5616 6564 5672
rect 6500 5612 6564 5616
rect 2568 5468 2632 5472
rect 2568 5412 2572 5468
rect 2572 5412 2628 5468
rect 2628 5412 2632 5468
rect 2568 5408 2632 5412
rect 2648 5468 2712 5472
rect 2648 5412 2652 5468
rect 2652 5412 2708 5468
rect 2708 5412 2712 5468
rect 2648 5408 2712 5412
rect 2728 5468 2792 5472
rect 2728 5412 2732 5468
rect 2732 5412 2788 5468
rect 2788 5412 2792 5468
rect 2728 5408 2792 5412
rect 2808 5468 2872 5472
rect 2808 5412 2812 5468
rect 2812 5412 2868 5468
rect 2868 5412 2872 5468
rect 2808 5408 2872 5412
rect 7568 5468 7632 5472
rect 7568 5412 7572 5468
rect 7572 5412 7628 5468
rect 7628 5412 7632 5468
rect 7568 5408 7632 5412
rect 7648 5468 7712 5472
rect 7648 5412 7652 5468
rect 7652 5412 7708 5468
rect 7708 5412 7712 5468
rect 7648 5408 7712 5412
rect 7728 5468 7792 5472
rect 7728 5412 7732 5468
rect 7732 5412 7788 5468
rect 7788 5412 7792 5468
rect 7728 5408 7792 5412
rect 7808 5468 7872 5472
rect 7808 5412 7812 5468
rect 7812 5412 7868 5468
rect 7868 5412 7872 5468
rect 7808 5408 7872 5412
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 5308 4924 5372 4928
rect 5308 4868 5312 4924
rect 5312 4868 5368 4924
rect 5368 4868 5372 4924
rect 5308 4864 5372 4868
rect 3372 4856 3436 4860
rect 3372 4800 3422 4856
rect 3422 4800 3436 4856
rect 3372 4796 3436 4800
rect 7052 4720 7116 4724
rect 7052 4664 7102 4720
rect 7102 4664 7116 4720
rect 7052 4660 7116 4664
rect 7568 4380 7632 4384
rect 7568 4324 7572 4380
rect 7572 4324 7628 4380
rect 7628 4324 7632 4380
rect 7568 4320 7632 4324
rect 7648 4380 7712 4384
rect 7648 4324 7652 4380
rect 7652 4324 7708 4380
rect 7708 4324 7712 4380
rect 7648 4320 7712 4324
rect 7728 4380 7792 4384
rect 7728 4324 7732 4380
rect 7732 4324 7788 4380
rect 7788 4324 7792 4380
rect 7728 4320 7792 4324
rect 7808 4380 7872 4384
rect 7808 4324 7812 4380
rect 7812 4324 7868 4380
rect 7868 4324 7872 4380
rect 7808 4320 7872 4324
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 5308 3836 5372 3840
rect 5308 3780 5312 3836
rect 5312 3780 5368 3836
rect 5368 3780 5372 3836
rect 5308 3776 5372 3780
rect 7568 3292 7632 3296
rect 7568 3236 7572 3292
rect 7572 3236 7628 3292
rect 7628 3236 7632 3292
rect 7568 3232 7632 3236
rect 7648 3292 7712 3296
rect 7648 3236 7652 3292
rect 7652 3236 7708 3292
rect 7708 3236 7712 3292
rect 7648 3232 7712 3236
rect 7728 3292 7792 3296
rect 7728 3236 7732 3292
rect 7732 3236 7788 3292
rect 7788 3236 7792 3292
rect 7728 3232 7792 3236
rect 7808 3292 7872 3296
rect 7808 3236 7812 3292
rect 7812 3236 7868 3292
rect 7868 3236 7872 3292
rect 7808 3232 7872 3236
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 5308 2748 5372 2752
rect 5308 2692 5312 2748
rect 5312 2692 5368 2748
rect 5368 2692 5372 2748
rect 5308 2688 5372 2692
rect 9076 2484 9140 2548
rect 7568 2204 7632 2208
rect 7568 2148 7572 2204
rect 7572 2148 7628 2204
rect 7628 2148 7632 2204
rect 7568 2144 7632 2148
rect 7648 2204 7712 2208
rect 7648 2148 7652 2204
rect 7652 2148 7708 2204
rect 7708 2148 7712 2204
rect 7648 2144 7712 2148
rect 7728 2204 7792 2208
rect 7728 2148 7732 2204
rect 7732 2148 7788 2204
rect 7788 2148 7792 2204
rect 7728 2144 7792 2148
rect 7808 2204 7872 2208
rect 7808 2148 7812 2204
rect 7812 2148 7868 2204
rect 7868 2148 7872 2204
rect 7808 2144 7872 2148
rect 5068 1660 5132 1664
rect 5068 1604 5072 1660
rect 5072 1604 5128 1660
rect 5128 1604 5132 1660
rect 5068 1600 5132 1604
rect 5148 1660 5212 1664
rect 5148 1604 5152 1660
rect 5152 1604 5208 1660
rect 5208 1604 5212 1660
rect 5148 1600 5212 1604
rect 5228 1660 5292 1664
rect 5228 1604 5232 1660
rect 5232 1604 5288 1660
rect 5288 1604 5292 1660
rect 5228 1600 5292 1604
rect 5308 1660 5372 1664
rect 5308 1604 5312 1660
rect 5312 1604 5368 1660
rect 5368 1604 5372 1660
rect 5308 1600 5372 1604
rect 2568 1116 2632 1120
rect 2568 1060 2572 1116
rect 2572 1060 2628 1116
rect 2628 1060 2632 1116
rect 2568 1056 2632 1060
rect 2648 1116 2712 1120
rect 2648 1060 2652 1116
rect 2652 1060 2708 1116
rect 2708 1060 2712 1116
rect 2648 1056 2712 1060
rect 2728 1116 2792 1120
rect 2728 1060 2732 1116
rect 2732 1060 2788 1116
rect 2788 1060 2792 1116
rect 2728 1056 2792 1060
rect 2808 1116 2872 1120
rect 2808 1060 2812 1116
rect 2812 1060 2868 1116
rect 2868 1060 2872 1116
rect 2808 1056 2872 1060
rect 7568 1116 7632 1120
rect 7568 1060 7572 1116
rect 7572 1060 7628 1116
rect 7628 1060 7632 1116
rect 7568 1056 7632 1060
rect 7648 1116 7712 1120
rect 7648 1060 7652 1116
rect 7652 1060 7708 1116
rect 7708 1060 7712 1116
rect 7648 1056 7712 1060
rect 7728 1116 7792 1120
rect 7728 1060 7732 1116
rect 7732 1060 7788 1116
rect 7788 1060 7792 1116
rect 7728 1056 7792 1060
rect 7808 1116 7872 1120
rect 7808 1060 7812 1116
rect 7812 1060 7868 1116
rect 7868 1060 7872 1116
rect 7808 1056 7872 1060
rect 5068 572 5132 576
rect 5068 516 5072 572
rect 5072 516 5128 572
rect 5128 516 5132 572
rect 5068 512 5132 516
rect 5148 572 5212 576
rect 5148 516 5152 572
rect 5152 516 5208 572
rect 5208 516 5212 572
rect 5148 512 5212 516
rect 5228 572 5292 576
rect 5228 516 5232 572
rect 5232 516 5288 572
rect 5288 516 5292 572
rect 5228 512 5292 516
rect 5308 572 5372 576
rect 5308 516 5312 572
rect 5312 516 5368 572
rect 5368 516 5372 572
rect 5308 512 5372 516
<< metal4 >>
rect 2560 12000 2880 12016
rect 2560 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2880 12000
rect 2560 11598 2880 11936
rect 2560 11362 2602 11598
rect 2838 11362 2880 11598
rect 2560 10912 2880 11362
rect 2560 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2880 10912
rect 2560 9824 2880 10848
rect 3003 10436 3069 10437
rect 3003 10372 3004 10436
rect 3068 10372 3069 10436
rect 3003 10371 3069 10372
rect 2560 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2880 9824
rect 2560 8736 2880 9760
rect 2560 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2880 8736
rect 2560 8218 2880 8672
rect 2560 7982 2602 8218
rect 2838 7982 2880 8218
rect 3006 8125 3066 10371
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 3003 8124 3069 8125
rect 3003 8060 3004 8124
rect 3068 8060 3069 8124
rect 3003 8059 3069 8060
rect 2560 7648 2880 7982
rect 3006 7717 3066 8059
rect 3003 7716 3069 7717
rect 3003 7652 3004 7716
rect 3068 7652 3069 7716
rect 3003 7651 3069 7652
rect 2560 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2880 7648
rect 2560 6560 2880 7584
rect 2560 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2880 6560
rect 2560 5472 2880 6496
rect 2560 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2880 5472
rect 2560 4838 2880 5408
rect 3374 4861 3434 9555
rect 3560 9266 3880 12016
rect 5060 11456 5380 12016
rect 5060 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5380 11456
rect 5060 10368 5380 11392
rect 5060 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5380 10368
rect 5060 9908 5380 10304
rect 5060 9672 5102 9908
rect 5338 9672 5380 9908
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 4662 6221 4722 9555
rect 5060 9280 5380 9672
rect 5060 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5380 9280
rect 5060 8192 5380 9216
rect 5060 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5380 8192
rect 5060 7104 5380 8128
rect 6060 10956 6380 12016
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 7560 12000 7880 12016
rect 7560 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7880 12000
rect 7560 11598 7880 11936
rect 7560 11362 7602 11598
rect 7838 11362 7880 11598
rect 7560 10912 7880 11362
rect 7560 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7880 10912
rect 7560 9824 7880 10848
rect 7560 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7880 9824
rect 7051 9212 7117 9213
rect 7051 9148 7052 9212
rect 7116 9148 7117 9212
rect 7051 9147 7117 9148
rect 6499 8396 6565 8397
rect 6499 8332 6500 8396
rect 6564 8332 6565 8396
rect 6499 8331 6565 8332
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 5579 7172 5645 7173
rect 5579 7108 5580 7172
rect 5644 7108 5645 7172
rect 5579 7107 5645 7108
rect 5060 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5380 7104
rect 5060 6528 5380 7040
rect 5060 6292 5102 6528
rect 5338 6292 5380 6528
rect 4659 6220 4725 6221
rect 4659 6156 4660 6220
rect 4724 6156 4725 6220
rect 4659 6155 4725 6156
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 3371 4860 3437 4861
rect 3371 4796 3372 4860
rect 3436 4796 3437 4860
rect 3371 4795 3437 4796
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1120 2880 1222
rect 2560 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2880 1120
rect 2560 496 2880 1056
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 496 3880 2270
rect 5060 6016 5380 6292
rect 5060 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5380 6016
rect 5060 4928 5380 5952
rect 5582 5813 5642 7107
rect 5579 5812 5645 5813
rect 5579 5748 5580 5812
rect 5644 5748 5645 5812
rect 5579 5747 5645 5748
rect 5060 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5380 4928
rect 5060 3840 5380 4864
rect 5060 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5380 3840
rect 5060 3148 5380 3776
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2752 5380 2912
rect 5060 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5380 2752
rect 5060 1664 5380 2688
rect 5060 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5380 1664
rect 5060 576 5380 1600
rect 5060 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5380 576
rect 5060 496 5380 512
rect 6060 4196 6380 7340
rect 6502 5677 6562 8331
rect 6499 5676 6565 5677
rect 6499 5612 6500 5676
rect 6564 5612 6565 5676
rect 6499 5611 6565 5612
rect 7054 4725 7114 9147
rect 7560 8736 7880 9760
rect 7560 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7880 8736
rect 7560 8218 7880 8672
rect 7560 7982 7602 8218
rect 7838 7982 7880 8218
rect 7560 7648 7880 7982
rect 7560 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7880 7648
rect 7560 6560 7880 7584
rect 7560 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7880 6560
rect 7560 5472 7880 6496
rect 7560 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7880 5472
rect 7560 4838 7880 5408
rect 7051 4724 7117 4725
rect 7051 4660 7052 4724
rect 7116 4660 7117 4724
rect 7051 4659 7117 4660
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 496 6380 3960
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 4384 7880 4602
rect 7560 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7880 4384
rect 7560 3296 7880 4320
rect 7560 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7880 3296
rect 7560 2208 7880 3232
rect 7560 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7880 2208
rect 7560 1458 7880 2144
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 7560 1120 7880 1222
rect 7560 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7880 1120
rect 7560 496 7880 1056
rect 8560 9266 8880 12016
rect 9075 9348 9141 9349
rect 9075 9284 9076 9348
rect 9140 9284 9141 9348
rect 9075 9283 9141 9284
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 9078 7989 9138 9283
rect 9075 7988 9141 7989
rect 9075 7924 9076 7988
rect 9140 7924 9141 7988
rect 9075 7923 9141 7924
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 9078 2549 9138 7923
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 9075 2548 9141 2549
rect 9075 2484 9076 2548
rect 9140 2484 9141 2548
rect 9075 2483 9141 2484
rect 8560 496 8880 2270
<< via4 >>
rect 2602 11362 2838 11598
rect 2602 7982 2838 8218
rect 5102 9672 5338 9908
rect 3602 9030 3838 9266
rect 6102 10720 6338 10956
rect 7602 11362 7838 11598
rect 6102 7340 6338 7576
rect 5102 6292 5338 6528
rect 3602 5650 3838 5886
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 2270 3838 2506
rect 5102 2912 5338 3148
rect 7602 7982 7838 8218
rect 6102 3960 6338 4196
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 872 11598 10000 11640
rect 872 11362 2602 11598
rect 2838 11362 7602 11598
rect 7838 11362 10000 11598
rect 872 11320 10000 11362
rect 872 10956 10000 10998
rect 872 10720 6102 10956
rect 6338 10720 10000 10956
rect 872 10678 10000 10720
rect 872 9908 10000 9950
rect 872 9672 5102 9908
rect 5338 9672 10000 9908
rect 872 9630 10000 9672
rect 872 9266 10000 9308
rect 872 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 10000 9266
rect 872 8988 10000 9030
rect 872 8218 10000 8260
rect 872 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 10000 8218
rect 872 7940 10000 7982
rect 872 7576 10000 7618
rect 872 7340 6102 7576
rect 6338 7340 10000 7576
rect 872 7298 10000 7340
rect 872 6528 10000 6570
rect 872 6292 5102 6528
rect 5338 6292 10000 6528
rect 872 6250 10000 6292
rect 872 5886 10000 5928
rect 872 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 10000 5886
rect 872 5608 10000 5650
rect 872 4838 10000 4880
rect 872 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 10000 4838
rect 872 4560 10000 4602
rect 872 4196 10000 4238
rect 872 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 10000 4196
rect 872 3918 10000 3960
rect 872 3148 10000 3190
rect 872 2912 5102 3148
rect 5338 2912 10000 3148
rect 872 2870 10000 2912
rect 872 2506 10000 2548
rect 872 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 10000 2506
rect 872 2228 10000 2270
rect 872 1458 10000 1500
rect 872 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 10000 1458
rect 872 1180 10000 1222
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 6716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__B
timestamp 1663859327
transform -1 0 6072 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 1663859327
transform -1 0 9384 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 1663859327
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B
timestamp 1663859327
transform -1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 1663859327
transform -1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 1663859327
transform -1 0 5060 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 1663859327
transform -1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 1663859327
transform -1 0 6900 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 1663859327
transform -1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 1663859327
transform -1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 1663859327
transform -1 0 4048 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 1663859327
transform -1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 1663859327
transform 1 0 1196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1663859327
transform -1 0 3404 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 1663859327
transform 1 0 8648 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1663859327
transform 1 0 8832 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1663859327
transform -1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1663859327
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 1663859327
transform -1 0 8648 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 1663859327
transform -1 0 8464 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1663859327
transform -1 0 5888 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1663859327
transform -1 0 9016 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1663859327
transform -1 0 4876 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 1663859327
transform -1 0 5244 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 1663859327
transform 1 0 3312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1663859327
transform -1 0 4692 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1663859327
transform -1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B
timestamp 1663859327
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1663859327
transform -1 0 3496 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1663859327
transform -1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1663859327
transform -1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout28_A
timestamp 1663859327
transform 1 0 5244 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout29_A
timestamp 1663859327
transform -1 0 6440 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1663859327
transform -1 0 6624 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1663859327
transform -1 0 4048 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1663859327
transform -1 0 5612 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1663859327
transform -1 0 6440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1663859327
transform -1 0 9200 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 3404 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31
timestamp 1663859327
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1663859327
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1663859327
transform 1 0 8740 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95
timestamp 1663859327
transform 1 0 9660 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34
timestamp 1663859327
transform 1 0 4048 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1663859327
transform 1 0 8280 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_89
timestamp 1663859327
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1663859327
transform 1 0 10028 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1663859327
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1663859327
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1663859327
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1663859327
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_99
timestamp 1663859327
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1663859327
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_71
timestamp 1663859327
transform 1 0 7452 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1663859327
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1663859327
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1663859327
transform -1 0 10396 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1663859327
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1663859327
transform -1 0 10396 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1663859327
transform 1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1663859327
transform -1 0 10396 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1663859327
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1663859327
transform -1 0 10396 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1663859327
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1663859327
transform -1 0 10396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1663859327
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1663859327
transform -1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1663859327
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1663859327
transform -1 0 10396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1663859327
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1663859327
transform -1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1663859327
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1663859327
transform -1 0 10396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1663859327
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1663859327
transform -1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1663859327
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1663859327
transform -1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1663859327
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1663859327
transform -1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1663859327
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1663859327
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1663859327
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1663859327
transform -1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1663859327
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1663859327
transform -1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1663859327
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1663859327
transform -1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1663859327
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1663859327
transform -1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1663859327
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1663859327
transform -1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1663859327
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1663859327
transform -1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1663859327
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1663859327
transform -1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1663859327
transform 1 0 920 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1663859327
transform -1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 3496 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1663859327
transform 1 0 6072 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1663859327
transform 1 0 8648 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1663859327
transform 1 0 8188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1663859327
transform 1 0 5612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1663859327
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1663859327
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1663859327
transform 1 0 8188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1663859327
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1663859327
transform 1 0 8188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1663859327
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1663859327
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1663859327
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1663859327
transform 1 0 8648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1663859327
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1663859327
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1663859327
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1663859327
transform 1 0 3496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1663859327
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1663859327
transform 1 0 6072 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1663859327
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1663859327
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1663859327
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1663859327
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1663859327
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1663859327
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1663859327
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1663859327
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1663859327
transform 1 0 6072 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1663859327
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1663859327
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1663859327
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _058__1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059__14
timestamp 1663859327
transform -1 0 3864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 9660 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_2  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 9476 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 9936 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 9108 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 10120 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 8924 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 8832 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or2_0  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 9568 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _069_
timestamp 1663859327
transform 1 0 6900 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _070_
timestamp 1663859327
transform -1 0 6716 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _071_
timestamp 1663859327
transform 1 0 6900 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _072_
timestamp 1663859327
transform 1 0 3588 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _073_
timestamp 1663859327
transform -1 0 6348 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _074_
timestamp 1663859327
transform 1 0 7728 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _075_
timestamp 1663859327
transform 1 0 9384 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _076_
timestamp 1663859327
transform 1 0 5152 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _077_
timestamp 1663859327
transform 1 0 3680 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _078_
timestamp 1663859327
transform 1 0 1196 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _079_
timestamp 1663859327
transform 1 0 9476 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _080_
timestamp 1663859327
transform 1 0 1196 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _081_
timestamp 1663859327
transform 1 0 9476 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _082_
timestamp 1663859327
transform 1 0 8740 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _083_
timestamp 1663859327
transform -1 0 8648 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _084_
timestamp 1663859327
transform 1 0 8372 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _085_
timestamp 1663859327
transform -1 0 9108 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _086_
timestamp 1663859327
transform -1 0 10028 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _087_
timestamp 1663859327
transform -1 0 10028 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _088_
timestamp 1663859327
transform -1 0 1656 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _089_
timestamp 1663859327
transform 1 0 3496 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _090_
timestamp 1663859327
transform 1 0 3312 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _091_
timestamp 1663859327
transform 1 0 3496 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _092_
timestamp 1663859327
transform 1 0 6164 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _093_
timestamp 1663859327
transform 1 0 6164 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _094__2
timestamp 1663859327
transform -1 0 4232 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095__3
timestamp 1663859327
transform -1 0 1472 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096__4
timestamp 1663859327
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097__5
timestamp 1663859327
transform -1 0 3956 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__6
timestamp 1663859327
transform 1 0 3312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__7
timestamp 1663859327
transform -1 0 1472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__8
timestamp 1663859327
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__9
timestamp 1663859327
transform 1 0 4232 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__10
timestamp 1663859327
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__11
timestamp 1663859327
transform -1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__12
timestamp 1663859327
transform -1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105__13
timestamp 1663859327
transform -1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 6072 0 1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 1663859327
transform 1 0 3496 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 1663859327
transform 1 0 6808 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 1663859327
transform -1 0 10120 0 -1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1663859327
transform 1 0 3496 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1663859327
transform 1 0 3496 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1663859327
transform 1 0 4324 0 1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1663859327
transform 1 0 7084 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1663859327
transform 1 0 6992 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1663859327
transform 1 0 7544 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1663859327
transform 1 0 3496 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1663859327
transform 1 0 4324 0 -1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _118_
timestamp 1663859327
transform 1 0 5428 0 1 5984
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_4  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 3956 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _120_
timestamp 1663859327
transform 1 0 1380 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _121_
timestamp 1663859327
transform 1 0 1380 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _122_
timestamp 1663859327
transform 1 0 1380 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _123_
timestamp 1663859327
transform -1 0 5704 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _124_
timestamp 1663859327
transform -1 0 3496 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _125_
timestamp 1663859327
transform 1 0 1380 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _126_
timestamp 1663859327
transform 1 0 3956 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _127_
timestamp 1663859327
transform 1 0 4416 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _128_
timestamp 1663859327
transform 1 0 6348 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _129_
timestamp 1663859327
transform 1 0 6532 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _130_
timestamp 1663859327
transform 1 0 3956 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _131_
timestamp 1663859327
transform 1 0 6532 0 1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 3496 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1663859327
transform -1 0 6072 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 3496 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1663859327
transform -1 0 3496 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1663859327
transform -1 0 3036 0 1 544
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1663859327
transform 1 0 3772 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1663859327
transform 1 0 3588 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1663859327
transform -1 0 3496 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 9660 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1663859327
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1663859327
transform -1 0 6532 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1663859327
transform -1 0 3680 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1663859327
transform -1 0 3956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1663859327
transform -1 0 1564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1663859327
transform 1 0 3312 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1663859327
transform 1 0 9752 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1663859327
transform 1 0 9384 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1663859327
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use gpio_logic_high  gpio_logic_high
timestamp 1638030917
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1663859327
transform 1 0 8740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1663859327
transform -1 0 9476 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1663859327
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1663859327
transform -1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1663859327
transform -1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1663859327
transform -1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1663859327
transform -1 0 4324 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1663859327
transform -1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1663859327
transform 1 0 6716 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1663859327
transform -1 0 6900 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1663859327
transform 1 0 3680 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1663859327
transform 1 0 1196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1663859327
transform 1 0 9016 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1663859327
transform -1 0 10120 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1663859327
transform -1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1663859327
transform -1 0 6072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1663859327
transform -1 0 10120 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  one_buffer $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform -1 0 6072 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output6
timestamp 1663859327
transform -1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output7
timestamp 1663859327
transform 1 0 6624 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output8
timestamp 1663859327
transform -1 0 8188 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output9
timestamp 1663859327
transform 1 0 6072 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output10
timestamp 1663859327
transform -1 0 6164 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output11
timestamp 1663859327
transform -1 0 8188 0 -1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output12
timestamp 1663859327
transform -1 0 10120 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output13
timestamp 1663859327
transform 1 0 6164 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output14
timestamp 1663859327
transform 1 0 6072 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output15
timestamp 1663859327
transform 1 0 8096 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output16
timestamp 1663859327
transform -1 0 10120 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output17
timestamp 1663859327
transform -1 0 8648 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output18
timestamp 1663859327
transform -1 0 8096 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output19
timestamp 1663859327
transform -1 0 3496 0 -1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output20
timestamp 1663859327
transform -1 0 3956 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output21
timestamp 1663859327
transform 1 0 4048 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output22
timestamp 1663859327
transform -1 0 3496 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_16  serial_clock_out_buffer
timestamp 1663859327
transform 1 0 3312 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  serial_load_out_buffer
timestamp 1663859327
transform 1 0 3312 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__macro_sparecell  spare_cell $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1663859327
transform 1 0 7452 0 1 2720
box -38 -48 2706 592
use sky130_fd_sc_hd__buf_16  zero_buffer
timestamp 1663859327
transform -1 0 6164 0 -1 2720
box -38 -48 2062 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 496 2880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 496 7880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1180 10000 1500 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4560 10000 4880 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7940 10000 8260 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 11320 10000 11640 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3560 496 3880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8560 496 8880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2228 10000 2548 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 5608 10000 5928 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 8988 10000 9308 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 5060 496 5380 12016 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2870 10000 3190 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 6250 10000 6570 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9630 10000 9950 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6060 496 6380 12016 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3918 10000 4238 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 7298 10000 7618 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 10678 10000 10998 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
