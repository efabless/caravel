magic
tech sky130A
magscale 1 2
timestamp 1506572754
<< checkpaint >>
rect -4476 -4198 636864 956856
<< isosubstrate >>
rect 50674 930615 55576 935630
rect 110775 930502 115563 935668
rect 190632 930600 195676 935619
rect 230738 930793 235564 935619
rect 290688 930538 295611 935711
rect 350643 930793 355711 935595
rect 410680 930649 415627 935619
rect 470693 930383 475785 935692
rect 550682 930649 555726 935644
rect 1780 899622 6787 904630
rect 625545 889766 630410 894592
rect 625448 799518 630352 804614
rect 1906 729809 6781 734756
rect 625540 713762 630366 718588
rect 1780 685644 6726 690832
rect 625448 669636 630410 674617
rect 1930 641605 6817 646672
rect 625516 623658 630366 628653
rect 1869 599739 6780 604711
rect 625377 577598 630384 582636
rect 1810 553536 6862 558739
rect 625347 533620 630354 538718
rect 1930 513531 6817 518719
rect 625407 485691 630384 490637
rect 1930 471604 6877 476823
rect 1870 341691 6787 346668
rect 625498 311678 630414 316746
rect 1810 299703 6817 304680
rect 625395 263724 630390 268623
rect 1870 253764 6666 258621
rect 625540 219734 630294 224609
rect 2021 211717 6757 216724
rect 163965 179571 185037 181815
rect 237194 179822 308640 184521
rect 625506 175768 630294 180652
rect 1882 167660 6757 172728
rect 1858 125455 6781 130668
rect 625371 129591 630429 134572
rect 625429 85751 630332 90770
rect 625560 39752 630379 44648
rect 136275 4720 141007 8871
<< metal3 >>
rect 533387 954354 538193 955596
rect 533387 952770 533467 954354
rect 538091 952770 538193 954354
rect 533387 952680 538193 952770
rect 543368 954354 548174 955596
rect 543368 952770 543448 954354
rect 548072 952770 548174 954354
rect 543368 952680 548174 952770
rect 609647 911040 628047 911068
rect 609647 910816 609696 911040
rect 610240 910816 627064 911040
rect 628008 910816 628047 911040
rect 609647 910788 628047 910816
rect 610600 910496 626860 910524
rect 610600 910272 610656 910496
rect 611200 910272 625864 910496
rect 626808 910272 626860 910496
rect 610600 910244 626860 910272
rect 616360 909952 625660 909980
rect 616360 909728 616416 909952
rect 616960 909728 624664 909952
rect 625608 909728 625660 909952
rect 616360 909700 625660 909728
rect 615400 909408 624460 909436
rect 615400 909184 615456 909408
rect 616000 909184 623464 909408
rect 624408 909184 624460 909408
rect 615400 909156 624460 909184
rect 614450 908864 623260 908892
rect 614450 908640 614496 908864
rect 615040 908640 622264 908864
rect 623208 908640 623260 908864
rect 614450 908612 623260 908640
rect 613460 908320 622060 908348
rect 613460 908096 613536 908320
rect 614080 908096 621064 908320
rect 622008 908096 622060 908320
rect 613460 908068 622060 908096
rect 612500 907776 620860 907804
rect 612500 907552 612576 907776
rect 613120 907552 619864 907776
rect 620808 907552 620860 907776
rect 612500 907524 620860 907552
rect 611560 907232 619660 907260
rect 611560 907008 611616 907232
rect 612160 907008 618664 907232
rect 619608 907008 619660 907232
rect 611560 906980 619660 907008
rect 4573 906144 22973 906172
rect 4573 905920 4612 906144
rect 5556 905920 22380 906144
rect 22924 905920 22973 906144
rect 4573 905892 22973 905920
rect 5760 905600 22020 905628
rect 5760 905376 5812 905600
rect 6756 905376 21420 905600
rect 21964 905376 22020 905600
rect 5760 905348 22020 905376
rect 6960 905056 16260 905084
rect 6960 904832 7012 905056
rect 7956 904832 15660 905056
rect 16204 904832 16260 905056
rect 6960 904804 16260 904832
rect 8160 904512 17220 904540
rect 8160 904288 8212 904512
rect 9156 904288 16620 904512
rect 17164 904288 17220 904512
rect 8160 904260 17220 904288
rect 9360 903968 18170 903996
rect 9360 903744 9412 903968
rect 10356 903744 17580 903968
rect 18124 903744 18170 903968
rect 9360 903716 18170 903744
rect 10560 903424 19160 903452
rect 10560 903200 10612 903424
rect 11556 903200 18540 903424
rect 19084 903200 19160 903424
rect 10560 903172 19160 903200
rect 11760 902880 20120 902908
rect 11760 902656 11812 902880
rect 12756 902656 19500 902880
rect 20044 902656 20120 902880
rect 11760 902628 20120 902656
rect 12960 902336 21060 902364
rect 12960 902112 13012 902336
rect 13956 902112 20460 902336
rect 21004 902112 21060 902336
rect 12960 902084 21060 902112
rect 609647 896352 628047 896380
rect 609647 896128 609696 896352
rect 610240 896128 627064 896352
rect 628008 896128 628047 896352
rect 609647 896100 628047 896128
rect 610600 895808 626860 895836
rect 610600 895584 610656 895808
rect 611200 895584 625864 895808
rect 626808 895584 626860 895808
rect 610600 895556 626860 895584
rect 616360 895264 625660 895292
rect 616360 895040 616416 895264
rect 616960 895040 624664 895264
rect 625608 895040 625660 895264
rect 616360 895012 625660 895040
rect 615400 894720 624460 894748
rect 615400 894496 615456 894720
rect 616000 894496 623464 894720
rect 624408 894496 624460 894720
rect 615400 894468 624460 894496
rect 614450 894176 623260 894204
rect 614450 893952 614496 894176
rect 615040 893952 622264 894176
rect 623208 893952 623260 894176
rect 614450 893924 623260 893952
rect 613460 893632 622060 893660
rect 613460 893408 613536 893632
rect 614080 893408 621064 893632
rect 622008 893408 622060 893632
rect 613460 893380 622060 893408
rect 612500 893088 620860 893116
rect 612500 892864 612576 893088
rect 613120 892864 619864 893088
rect 620808 892864 620860 893088
rect 612500 892836 620860 892864
rect 611560 892544 619660 892572
rect 611560 892320 611616 892544
rect 612160 892320 618664 892544
rect 619608 892320 619660 892544
rect 611560 892292 619660 892320
rect 4573 891456 22973 891484
rect 4573 891232 4612 891456
rect 5556 891232 22380 891456
rect 22924 891232 22973 891456
rect 4573 891204 22973 891232
rect 5760 890912 22020 890940
rect 5760 890688 5812 890912
rect 6756 890688 21420 890912
rect 21964 890688 22020 890912
rect 5760 890660 22020 890688
rect 6960 890368 16260 890396
rect 6960 890144 7012 890368
rect 7956 890144 15660 890368
rect 16204 890144 16260 890368
rect 6960 890116 16260 890144
rect 8160 889824 17220 889852
rect 8160 889600 8212 889824
rect 9156 889600 16620 889824
rect 17164 889600 17220 889824
rect 8160 889572 17220 889600
rect 9360 889280 18170 889308
rect 9360 889056 9412 889280
rect 10356 889056 17580 889280
rect 18124 889056 18170 889280
rect 9360 889028 18170 889056
rect 10560 888736 19160 888764
rect 10560 888512 10612 888736
rect 11556 888512 18540 888736
rect 19084 888512 19160 888736
rect 10560 888484 19160 888512
rect 11760 888192 20120 888220
rect 11760 887968 11812 888192
rect 12756 887968 19500 888192
rect 20044 887968 20120 888192
rect 11760 887940 20120 887968
rect 12960 887648 21060 887676
rect 12960 887424 13012 887648
rect 13956 887424 20460 887648
rect 21004 887424 21060 887648
rect 12960 887396 21060 887424
rect 609647 884928 628047 884956
rect -3216 884758 1182 884840
rect -3216 880134 -1777 884758
rect 1087 880134 1182 884758
rect 609647 884704 609696 884928
rect 610240 884704 627064 884928
rect 628008 884704 628047 884928
rect 609647 884676 628047 884704
rect 610600 884384 626860 884412
rect 610600 884160 610656 884384
rect 611200 884160 625864 884384
rect 626808 884160 626860 884384
rect 610600 884132 626860 884160
rect 616360 883840 625660 883868
rect 616360 883616 616416 883840
rect 616960 883616 624664 883840
rect 625608 883616 625660 883840
rect 616360 883588 625660 883616
rect 615400 883296 624460 883324
rect 615400 883072 615456 883296
rect 616000 883072 623464 883296
rect 624408 883072 624460 883296
rect 615400 883044 624460 883072
rect 614450 882752 623260 882780
rect 614450 882528 614496 882752
rect 615040 882528 622264 882752
rect 623208 882528 623260 882752
rect 614450 882500 623260 882528
rect 613460 882208 622060 882236
rect 613460 881984 613536 882208
rect 614080 881984 621064 882208
rect 622008 881984 622060 882208
rect 613460 881956 622060 881984
rect 612500 881664 620860 881692
rect 612500 881440 612576 881664
rect 613120 881440 619864 881664
rect 620808 881440 620860 881664
rect 612500 881412 620860 881440
rect 611560 881120 619660 881148
rect 611560 880896 611616 881120
rect 612160 880896 618664 881120
rect 619608 880896 619660 881120
rect 611560 880868 619660 880896
rect -3216 880051 1182 880134
rect 631206 880318 635604 880400
rect -2200 879648 1182 879730
rect -2200 875184 -1777 879648
rect 1087 875184 1182 879648
rect 4573 878400 22973 878428
rect 4573 878176 4612 878400
rect 5556 878176 22380 878400
rect 22924 878176 22973 878400
rect 4573 878148 22973 878176
rect 5760 877856 22020 877884
rect 5760 877632 5812 877856
rect 6756 877632 21420 877856
rect 21964 877632 22020 877856
rect 5760 877604 22020 877632
rect 6960 877312 16260 877340
rect 6960 877088 7012 877312
rect 7956 877088 15660 877312
rect 16204 877088 16260 877312
rect 6960 877060 16260 877088
rect 8160 876768 17220 876796
rect 8160 876544 8212 876768
rect 9156 876544 16620 876768
rect 17164 876544 17220 876768
rect 8160 876516 17220 876544
rect 9360 876224 18170 876252
rect 9360 876000 9412 876224
rect 10356 876000 17580 876224
rect 18124 876000 18170 876224
rect 9360 875972 18170 876000
rect 10560 875680 19160 875708
rect 10560 875456 10612 875680
rect 11556 875456 18540 875680
rect 19084 875456 19160 875680
rect 631206 875694 631301 880318
rect 634165 875694 635604 880318
rect 631206 875611 635604 875694
rect 10560 875428 19160 875456
rect -2200 875120 1182 875184
rect 631206 875208 635204 875290
rect 11760 875136 20120 875164
rect 11760 874912 11812 875136
rect 12756 874912 19500 875136
rect 20044 874912 20120 875136
rect 11760 874884 20120 874912
rect -3216 874718 1182 874800
rect -3216 870094 -1777 874718
rect 1087 870094 1182 874718
rect 12960 874592 21060 874620
rect 12960 874368 13012 874592
rect 13956 874368 20460 874592
rect 21004 874368 21060 874592
rect 12960 874340 21060 874368
rect 609647 871872 628047 871900
rect 609647 871648 609696 871872
rect 610240 871648 627064 871872
rect 628008 871648 628047 871872
rect 609647 871620 628047 871648
rect 610600 871328 626860 871356
rect 610600 871104 610656 871328
rect 611200 871104 625864 871328
rect 626808 871104 626860 871328
rect 610600 871076 626860 871104
rect 616360 870784 625660 870812
rect 616360 870560 616416 870784
rect 616960 870560 624664 870784
rect 625608 870560 625660 870784
rect 631206 870744 631301 875208
rect 634165 870744 635204 875208
rect 631206 870669 635204 870744
rect 616360 870532 625660 870560
rect -3216 870011 1182 870094
rect 615400 870240 624460 870268
rect 615400 870016 615456 870240
rect 616000 870016 623464 870240
rect 624408 870016 624460 870240
rect 615400 869988 624460 870016
rect 631206 870267 635604 870349
rect 614450 869696 623260 869724
rect 614450 869472 614496 869696
rect 615040 869472 622264 869696
rect 623208 869472 623260 869696
rect 614450 869444 623260 869472
rect 613460 869152 622060 869180
rect 613460 868928 613536 869152
rect 614080 868928 621064 869152
rect 622008 868928 622060 869152
rect 613460 868900 622060 868928
rect 612500 868608 620860 868636
rect 612500 868384 612576 868608
rect 613120 868384 619864 868608
rect 620808 868384 620860 868608
rect 612500 868356 620860 868384
rect 611560 868064 619660 868092
rect 611560 867840 611616 868064
rect 612160 867840 618664 868064
rect 619608 867840 619660 868064
rect 611560 867812 619660 867840
rect 631206 865643 631301 870267
rect 634165 865643 635604 870267
rect 631206 865560 635604 865643
rect 4573 865344 22973 865372
rect 4573 865120 4612 865344
rect 5556 865120 22380 865344
rect 22924 865120 22973 865344
rect 4573 865092 22973 865120
rect 5760 864800 22020 864828
rect 5760 864576 5812 864800
rect 6756 864576 21420 864800
rect 21964 864576 22020 864800
rect 5760 864548 22020 864576
rect 6960 864256 16260 864284
rect 6960 864032 7012 864256
rect 7956 864032 15660 864256
rect 16204 864032 16260 864256
rect 6960 864004 16260 864032
rect 8160 863712 17220 863740
rect 8160 863488 8212 863712
rect 9156 863488 16620 863712
rect 17164 863488 17220 863712
rect 8160 863460 17220 863488
rect 9360 863168 18170 863196
rect 9360 862944 9412 863168
rect 10356 862944 17580 863168
rect 18124 862944 18170 863168
rect 9360 862916 18170 862944
rect 10560 862624 19160 862652
rect 10560 862400 10612 862624
rect 11556 862400 18540 862624
rect 19084 862400 19160 862624
rect 10560 862372 19160 862400
rect 11760 862080 20120 862108
rect 11760 861856 11812 862080
rect 12756 861856 19500 862080
rect 20044 861856 20120 862080
rect 11760 861828 20120 861856
rect 12960 861536 21060 861564
rect 12960 861312 13012 861536
rect 13956 861312 20460 861536
rect 21004 861312 21060 861536
rect 12960 861284 21060 861312
rect 609647 858816 628047 858844
rect 609647 858592 609696 858816
rect 610240 858592 627064 858816
rect 628008 858592 628047 858816
rect 609647 858564 628047 858592
rect 610600 858272 626860 858300
rect 610600 858048 610656 858272
rect 611200 858048 625864 858272
rect 626808 858048 626860 858272
rect 610600 858020 626860 858048
rect 616360 857728 625660 857756
rect 616360 857504 616416 857728
rect 616960 857504 624664 857728
rect 625608 857504 625660 857728
rect 616360 857476 625660 857504
rect 615400 857184 624460 857212
rect 615400 856960 615456 857184
rect 616000 856960 623464 857184
rect 624408 856960 624460 857184
rect 615400 856932 624460 856960
rect 614450 856640 623260 856668
rect 614450 856416 614496 856640
rect 615040 856416 622264 856640
rect 623208 856416 623260 856640
rect 614450 856388 623260 856416
rect 613460 856096 622060 856124
rect 613460 855872 613536 856096
rect 614080 855872 621064 856096
rect 622008 855872 622060 856096
rect 613460 855844 622060 855872
rect 612500 855552 620860 855580
rect 612500 855328 612576 855552
rect 613120 855328 619864 855552
rect 620808 855328 620860 855552
rect 612500 855300 620860 855328
rect 611560 855008 619660 855036
rect 611560 854784 611616 855008
rect 612160 854784 618664 855008
rect 619608 854784 619660 855008
rect 611560 854756 619660 854784
rect 4573 852288 22973 852316
rect 4573 852064 4612 852288
rect 5556 852064 22380 852288
rect 22924 852064 22973 852288
rect 4573 852036 22973 852064
rect 5760 851744 22020 851772
rect 5760 851520 5812 851744
rect 6756 851520 21420 851744
rect 21964 851520 22020 851744
rect 5760 851492 22020 851520
rect 6960 851200 16260 851228
rect 6960 850976 7012 851200
rect 7956 850976 15660 851200
rect 16204 850976 16260 851200
rect 6960 850948 16260 850976
rect 8160 850656 17220 850684
rect 8160 850432 8212 850656
rect 9156 850432 16620 850656
rect 17164 850432 17220 850656
rect 8160 850404 17220 850432
rect 9360 850112 18170 850140
rect 9360 849888 9412 850112
rect 10356 849888 17580 850112
rect 18124 849888 18170 850112
rect 9360 849860 18170 849888
rect 10560 849568 19160 849596
rect 10560 849344 10612 849568
rect 11556 849344 18540 849568
rect 19084 849344 19160 849568
rect 10560 849316 19160 849344
rect 11760 849024 20120 849052
rect 11760 848800 11812 849024
rect 12756 848800 19500 849024
rect 20044 848800 20120 849024
rect 11760 848772 20120 848800
rect 12960 848480 21060 848508
rect 12960 848256 13012 848480
rect 13956 848256 20460 848480
rect 21004 848256 21060 848480
rect 12960 848228 21060 848256
rect 609647 845760 628047 845788
rect 609647 845536 609696 845760
rect 610240 845536 627064 845760
rect 628008 845536 628047 845760
rect 609647 845508 628047 845536
rect 610600 845216 626860 845244
rect 610600 844992 610656 845216
rect 611200 844992 625864 845216
rect 626808 844992 626860 845216
rect 610600 844964 626860 844992
rect 616360 844672 625660 844700
rect 616360 844448 616416 844672
rect 616960 844448 624664 844672
rect 625608 844448 625660 844672
rect 616360 844420 625660 844448
rect 615400 844128 624460 844156
rect 615400 843904 615456 844128
rect 616000 843904 623464 844128
rect 624408 843904 624460 844128
rect 615400 843876 624460 843904
rect 614450 843584 623260 843612
rect 614450 843360 614496 843584
rect 615040 843360 622264 843584
rect 623208 843360 623260 843584
rect 614450 843332 623260 843360
rect 613460 843040 622060 843068
rect 613460 842816 613536 843040
rect 614080 842816 621064 843040
rect 622008 842816 622060 843040
rect 613460 842788 622060 842816
rect 612500 842496 620860 842524
rect 612500 842272 612576 842496
rect 613120 842272 619864 842496
rect 620808 842272 620860 842496
rect 612500 842244 620860 842272
rect 611560 841952 619660 841980
rect 611560 841728 611616 841952
rect 612160 841728 618664 841952
rect 619608 841728 619660 841952
rect 611560 841700 619660 841728
rect 4573 839232 22973 839260
rect 4573 839008 4612 839232
rect 5556 839008 22380 839232
rect 22924 839008 22973 839232
rect 4573 838980 22973 839008
rect 5760 838688 22020 838716
rect 5760 838464 5812 838688
rect 6756 838464 21420 838688
rect 21964 838464 22020 838688
rect 5760 838436 22020 838464
rect 6960 838144 16260 838172
rect 6960 837920 7012 838144
rect 7956 837920 15660 838144
rect 16204 837920 16260 838144
rect 6960 837892 16260 837920
rect 8160 837600 17220 837628
rect 8160 837376 8212 837600
rect 9156 837376 16620 837600
rect 17164 837376 17220 837600
rect 8160 837348 17220 837376
rect 9360 837056 18170 837084
rect 9360 836832 9412 837056
rect 10356 836832 17580 837056
rect 18124 836832 18170 837056
rect 9360 836804 18170 836832
rect 10560 836512 19160 836540
rect 10560 836288 10612 836512
rect 11556 836288 18540 836512
rect 19084 836288 19160 836512
rect 10560 836260 19160 836288
rect 11760 835968 20120 835996
rect 11760 835744 11812 835968
rect 12756 835744 19500 835968
rect 20044 835744 20120 835968
rect 11760 835716 20120 835744
rect 12960 835424 21060 835452
rect 12960 835200 13012 835424
rect 13956 835200 20460 835424
rect 21004 835200 21060 835424
rect 12960 835172 21060 835200
rect 609647 832704 628047 832732
rect 609647 832480 609696 832704
rect 610240 832480 627064 832704
rect 628008 832480 628047 832704
rect 609647 832452 628047 832480
rect 610600 832160 626860 832188
rect 610600 831936 610656 832160
rect 611200 831936 625864 832160
rect 626808 831936 626860 832160
rect 610600 831908 626860 831936
rect 616360 831616 625660 831644
rect 616360 831392 616416 831616
rect 616960 831392 624664 831616
rect 625608 831392 625660 831616
rect 616360 831364 625660 831392
rect 615400 831072 624460 831100
rect 615400 830848 615456 831072
rect 616000 830848 623464 831072
rect 624408 830848 624460 831072
rect 615400 830820 624460 830848
rect 614450 830528 623260 830556
rect 614450 830304 614496 830528
rect 615040 830304 622264 830528
rect 623208 830304 623260 830528
rect 614450 830276 623260 830304
rect 613460 829984 622060 830012
rect 613460 829760 613536 829984
rect 614080 829760 621064 829984
rect 622008 829760 622060 829984
rect 613460 829732 622060 829760
rect 612500 829440 620860 829468
rect 612500 829216 612576 829440
rect 613120 829216 619864 829440
rect 620808 829216 620860 829440
rect 612500 829188 620860 829216
rect 611560 828896 619660 828924
rect 611560 828672 611616 828896
rect 612160 828672 618664 828896
rect 619608 828672 619660 828896
rect 611560 828644 619660 828672
rect 4573 826176 22973 826204
rect 4573 825952 4612 826176
rect 5556 825952 22380 826176
rect 22924 825952 22973 826176
rect 4573 825924 22973 825952
rect 5760 825632 22020 825660
rect 5760 825408 5812 825632
rect 6756 825408 21420 825632
rect 21964 825408 22020 825632
rect 5760 825380 22020 825408
rect 6960 825088 16260 825116
rect 6960 824864 7012 825088
rect 7956 824864 15660 825088
rect 16204 824864 16260 825088
rect 6960 824836 16260 824864
rect 8160 824544 17220 824572
rect 8160 824320 8212 824544
rect 9156 824320 16620 824544
rect 17164 824320 17220 824544
rect 8160 824292 17220 824320
rect 9360 824000 18170 824028
rect 9360 823776 9412 824000
rect 10356 823776 17580 824000
rect 18124 823776 18170 824000
rect 9360 823748 18170 823776
rect 10560 823456 19160 823484
rect 10560 823232 10612 823456
rect 11556 823232 18540 823456
rect 19084 823232 19160 823456
rect 10560 823204 19160 823232
rect 11760 822912 20120 822940
rect 11760 822688 11812 822912
rect 12756 822688 19500 822912
rect 20044 822688 20120 822912
rect 11760 822660 20120 822688
rect 12960 822368 21060 822396
rect 12960 822144 13012 822368
rect 13956 822144 20460 822368
rect 21004 822144 21060 822368
rect 12960 822116 21060 822144
rect 609647 819648 628047 819676
rect 609647 819424 609696 819648
rect 610240 819424 627064 819648
rect 628008 819424 628047 819648
rect 609647 819396 628047 819424
rect 610600 819104 626860 819132
rect 610600 818880 610656 819104
rect 611200 818880 625864 819104
rect 626808 818880 626860 819104
rect 610600 818852 626860 818880
rect 616360 818560 625660 818588
rect 616360 818336 616416 818560
rect 616960 818336 624664 818560
rect 625608 818336 625660 818560
rect 616360 818308 625660 818336
rect 615400 818016 624460 818044
rect 615400 817792 615456 818016
rect 616000 817792 623464 818016
rect 624408 817792 624460 818016
rect 615400 817764 624460 817792
rect 614450 817472 623260 817500
rect 614450 817248 614496 817472
rect 615040 817248 622264 817472
rect 623208 817248 623260 817472
rect 614450 817220 623260 817248
rect 613460 816928 622060 816956
rect 613460 816704 613536 816928
rect 614080 816704 621064 816928
rect 622008 816704 622060 816928
rect 613460 816676 622060 816704
rect 612500 816384 620860 816412
rect 612500 816160 612576 816384
rect 613120 816160 619864 816384
rect 620808 816160 620860 816384
rect 612500 816132 620860 816160
rect 611560 815840 619660 815868
rect 611560 815616 611616 815840
rect 612160 815616 618664 815840
rect 619608 815616 619660 815840
rect 611560 815588 619660 815616
rect 4573 813120 22973 813148
rect 4573 812896 4612 813120
rect 5556 812896 22380 813120
rect 22924 812896 22973 813120
rect 4573 812868 22973 812896
rect 5760 812576 22020 812604
rect 5760 812352 5812 812576
rect 6756 812352 21420 812576
rect 21964 812352 22020 812576
rect 5760 812324 22020 812352
rect 6960 812032 16260 812060
rect 6960 811808 7012 812032
rect 7956 811808 15660 812032
rect 16204 811808 16260 812032
rect 6960 811780 16260 811808
rect 8160 811488 17220 811516
rect 8160 811264 8212 811488
rect 9156 811264 16620 811488
rect 17164 811264 17220 811488
rect 8160 811236 17220 811264
rect 9360 810944 18170 810972
rect 9360 810720 9412 810944
rect 10356 810720 17580 810944
rect 18124 810720 18170 810944
rect 9360 810692 18170 810720
rect 10560 810400 19160 810428
rect 10560 810176 10612 810400
rect 11556 810176 18540 810400
rect 19084 810176 19160 810400
rect 10560 810148 19160 810176
rect 11760 809856 20120 809884
rect 11760 809632 11812 809856
rect 12756 809632 19500 809856
rect 20044 809632 20120 809856
rect 11760 809604 20120 809632
rect 12960 809312 21060 809340
rect 12960 809088 13012 809312
rect 13956 809088 20460 809312
rect 21004 809088 21060 809312
rect 12960 809060 21060 809088
rect 609647 806592 628047 806620
rect 609647 806368 609696 806592
rect 610240 806368 627064 806592
rect 628008 806368 628047 806592
rect 609647 806340 628047 806368
rect 610600 806048 626860 806076
rect 610600 805824 610656 806048
rect 611200 805824 625864 806048
rect 626808 805824 626860 806048
rect 610600 805796 626860 805824
rect 616360 805504 625660 805532
rect 616360 805280 616416 805504
rect 616960 805280 624664 805504
rect 625608 805280 625660 805504
rect 616360 805252 625660 805280
rect 615400 804960 624460 804988
rect 615400 804736 615456 804960
rect 616000 804736 623464 804960
rect 624408 804736 624460 804960
rect 615400 804708 624460 804736
rect 614450 804416 623260 804444
rect 614450 804192 614496 804416
rect 615040 804192 622264 804416
rect 623208 804192 623260 804416
rect 614450 804164 623260 804192
rect 613460 803872 622060 803900
rect 613460 803648 613536 803872
rect 614080 803648 621064 803872
rect 622008 803648 622060 803872
rect 613460 803620 622060 803648
rect 612500 803328 620860 803356
rect 612500 803104 612576 803328
rect 613120 803104 619864 803328
rect 620808 803104 620860 803328
rect 612500 803076 620860 803104
rect 611560 802784 619660 802812
rect 611560 802560 611616 802784
rect 612160 802560 618664 802784
rect 619608 802560 619660 802784
rect 611560 802532 619660 802560
rect -3216 800276 1182 800358
rect -3216 795652 -1777 800276
rect 1087 795652 1182 800276
rect 4573 800064 22973 800092
rect 4573 799840 4612 800064
rect 5556 799840 22380 800064
rect 22924 799840 22973 800064
rect 4573 799812 22973 799840
rect 5760 799520 22020 799548
rect 5760 799296 5812 799520
rect 6756 799296 21420 799520
rect 21964 799296 22020 799520
rect 5760 799268 22020 799296
rect 6960 798976 16260 799004
rect 6960 798752 7012 798976
rect 7956 798752 15660 798976
rect 16204 798752 16260 798976
rect 6960 798724 16260 798752
rect 8160 798432 17220 798460
rect 8160 798208 8212 798432
rect 9156 798208 16620 798432
rect 17164 798208 17220 798432
rect 8160 798180 17220 798208
rect 9360 797888 18170 797916
rect 9360 797664 9412 797888
rect 10356 797664 17580 797888
rect 18124 797664 18170 797888
rect 9360 797636 18170 797664
rect 10560 797344 19160 797372
rect 10560 797120 10612 797344
rect 11556 797120 18540 797344
rect 19084 797120 19160 797344
rect 10560 797092 19160 797120
rect 11760 796800 20120 796828
rect 11760 796576 11812 796800
rect 12756 796576 19500 796800
rect 20044 796576 20120 796800
rect 11760 796548 20120 796576
rect 12960 796256 21060 796284
rect 12960 796032 13012 796256
rect 13956 796032 20460 796256
rect 21004 796032 21060 796256
rect 12960 796004 21060 796032
rect -3216 795569 1182 795652
rect 609647 793536 628047 793564
rect 609647 793312 609696 793536
rect 610240 793312 627064 793536
rect 628008 793312 628047 793536
rect 609647 793284 628047 793312
rect 610600 792992 626860 793020
rect 610600 792768 610656 792992
rect 611200 792768 625864 792992
rect 626808 792768 626860 792992
rect 610600 792740 626860 792768
rect 616360 792448 625660 792476
rect 616360 792224 616416 792448
rect 616960 792224 624664 792448
rect 625608 792224 625660 792448
rect 616360 792196 625660 792224
rect 615400 791904 624460 791932
rect 615400 791680 615456 791904
rect 616000 791680 623464 791904
rect 624408 791680 624460 791904
rect 615400 791652 624460 791680
rect 614450 791360 623260 791388
rect 614450 791136 614496 791360
rect 615040 791136 622264 791360
rect 623208 791136 623260 791360
rect 614450 791108 623260 791136
rect 631206 791119 635604 791201
rect 613460 790816 622060 790844
rect 613460 790592 613536 790816
rect 614080 790592 621064 790816
rect 622008 790592 622060 790816
rect 613460 790564 622060 790592
rect -3216 790297 1182 790379
rect -3216 785673 -1777 790297
rect 1087 785673 1182 790297
rect 612500 790272 620860 790300
rect 612500 790048 612576 790272
rect 613120 790048 619864 790272
rect 620808 790048 620860 790272
rect 612500 790020 620860 790048
rect 611560 789728 619660 789756
rect 611560 789504 611616 789728
rect 612160 789504 618664 789728
rect 619608 789504 619660 789728
rect 611560 789476 619660 789504
rect 4573 787008 22973 787036
rect 4573 786784 4612 787008
rect 5556 786784 22380 787008
rect 22924 786784 22973 787008
rect 4573 786756 22973 786784
rect 631206 786495 631301 791119
rect 634165 786495 635604 791119
rect 5760 786464 22020 786492
rect 5760 786240 5812 786464
rect 6756 786240 21420 786464
rect 21964 786240 22020 786464
rect 631206 786412 635604 786495
rect 5760 786212 22020 786240
rect -3216 785590 1182 785673
rect 6960 785920 16260 785948
rect 6960 785696 7012 785920
rect 7956 785696 15660 785920
rect 16204 785696 16260 785920
rect 6960 785668 16260 785696
rect 8160 785376 17220 785404
rect 8160 785152 8212 785376
rect 9156 785152 16620 785376
rect 17164 785152 17220 785376
rect 8160 785124 17220 785152
rect 9360 784832 18170 784860
rect 9360 784608 9412 784832
rect 10356 784608 17580 784832
rect 18124 784608 18170 784832
rect 9360 784580 18170 784608
rect 10560 784288 19160 784316
rect 10560 784064 10612 784288
rect 11556 784064 18540 784288
rect 19084 784064 19160 784288
rect 10560 784036 19160 784064
rect 11760 783744 20120 783772
rect 11760 783520 11812 783744
rect 12756 783520 19500 783744
rect 20044 783520 20120 783744
rect 11760 783492 20120 783520
rect 12960 783200 21060 783228
rect 12960 782976 13012 783200
rect 13956 782976 20460 783200
rect 21004 782976 21060 783200
rect 12960 782948 21060 782976
rect 631206 781136 635604 781218
rect 609647 780480 628047 780508
rect 609647 780256 609696 780480
rect 610240 780256 627064 780480
rect 628008 780256 628047 780480
rect 609647 780228 628047 780256
rect 610600 779936 626860 779964
rect 610600 779712 610656 779936
rect 611200 779712 625864 779936
rect 626808 779712 626860 779936
rect 610600 779684 626860 779712
rect 616360 779392 625660 779420
rect 616360 779168 616416 779392
rect 616960 779168 624664 779392
rect 625608 779168 625660 779392
rect 616360 779140 625660 779168
rect 615400 778848 624460 778876
rect 615400 778624 615456 778848
rect 616000 778624 623464 778848
rect 624408 778624 624460 778848
rect 615400 778596 624460 778624
rect 614450 778304 623260 778332
rect 614450 778080 614496 778304
rect 615040 778080 622264 778304
rect 623208 778080 623260 778304
rect 614450 778052 623260 778080
rect 613460 777760 622060 777788
rect 613460 777536 613536 777760
rect 614080 777536 621064 777760
rect 622008 777536 622060 777760
rect 613460 777508 622060 777536
rect 612500 777216 620860 777244
rect 612500 776992 612576 777216
rect 613120 776992 619864 777216
rect 620808 776992 620860 777216
rect 612500 776964 620860 776992
rect 611560 776672 619660 776700
rect 611560 776448 611616 776672
rect 612160 776448 618664 776672
rect 619608 776448 619660 776672
rect 611560 776420 619660 776448
rect 631206 776512 631301 781136
rect 634165 776512 635604 781136
rect 631206 776429 635604 776512
rect 4573 773952 22973 773980
rect 4573 773728 4612 773952
rect 5556 773728 22380 773952
rect 22924 773728 22973 773952
rect 4573 773700 22973 773728
rect 5760 773408 22020 773436
rect 5760 773184 5812 773408
rect 6756 773184 21420 773408
rect 21964 773184 22020 773408
rect 5760 773156 22020 773184
rect 6960 772864 16260 772892
rect 6960 772640 7012 772864
rect 7956 772640 15660 772864
rect 16204 772640 16260 772864
rect 6960 772612 16260 772640
rect 8160 772320 17220 772348
rect 8160 772096 8212 772320
rect 9156 772096 16620 772320
rect 17164 772096 17220 772320
rect 8160 772068 17220 772096
rect 9360 771776 18170 771804
rect 9360 771552 9412 771776
rect 10356 771552 17580 771776
rect 18124 771552 18170 771776
rect 9360 771524 18170 771552
rect 10560 771232 19160 771260
rect 10560 771008 10612 771232
rect 11556 771008 18540 771232
rect 19084 771008 19160 771232
rect 10560 770980 19160 771008
rect 11760 770688 20120 770716
rect 11760 770464 11812 770688
rect 12756 770464 19500 770688
rect 20044 770464 20120 770688
rect 11760 770436 20120 770464
rect 12960 770144 21060 770172
rect 12960 769920 13012 770144
rect 13956 769920 20460 770144
rect 21004 769920 21060 770144
rect 12960 769892 21060 769920
rect 609647 767424 628047 767452
rect 609647 767200 609696 767424
rect 610240 767200 627064 767424
rect 628008 767200 628047 767424
rect 609647 767172 628047 767200
rect 610600 766880 626860 766908
rect 610600 766656 610656 766880
rect 611200 766656 625864 766880
rect 626808 766656 626860 766880
rect 610600 766628 626860 766656
rect 616360 766336 625660 766364
rect 616360 766112 616416 766336
rect 616960 766112 624664 766336
rect 625608 766112 625660 766336
rect 616360 766084 625660 766112
rect 615400 765792 624460 765820
rect 615400 765568 615456 765792
rect 616000 765568 623464 765792
rect 624408 765568 624460 765792
rect 615400 765540 624460 765568
rect 614450 765248 623260 765276
rect 614450 765024 614496 765248
rect 615040 765024 622264 765248
rect 623208 765024 623260 765248
rect 614450 764996 623260 765024
rect 613460 764704 622060 764732
rect 613460 764480 613536 764704
rect 614080 764480 621064 764704
rect 622008 764480 622060 764704
rect 613460 764452 622060 764480
rect 612500 764160 620860 764188
rect 612500 763936 612576 764160
rect 613120 763936 619864 764160
rect 620808 763936 620860 764160
rect 612500 763908 620860 763936
rect 611560 763616 619660 763644
rect 611560 763392 611616 763616
rect 612160 763392 618664 763616
rect 619608 763392 619660 763616
rect 611560 763364 619660 763392
rect 4573 760896 22973 760924
rect 4573 760672 4612 760896
rect 5556 760672 22380 760896
rect 22924 760672 22973 760896
rect 4573 760644 22973 760672
rect 5760 760352 22020 760380
rect 5760 760128 5812 760352
rect 6756 760128 21420 760352
rect 21964 760128 22020 760352
rect 5760 760100 22020 760128
rect 6960 759808 16260 759836
rect 6960 759584 7012 759808
rect 7956 759584 15660 759808
rect 16204 759584 16260 759808
rect 6960 759556 16260 759584
rect 8160 759264 17220 759292
rect 8160 759040 8212 759264
rect 9156 759040 16620 759264
rect 17164 759040 17220 759264
rect 8160 759012 17220 759040
rect 9360 758720 18170 758748
rect 9360 758496 9412 758720
rect 10356 758496 17580 758720
rect 18124 758496 18170 758720
rect 9360 758468 18170 758496
rect 10560 758176 19160 758204
rect 10560 757952 10612 758176
rect 11556 757952 18540 758176
rect 19084 757952 19160 758176
rect 10560 757924 19160 757952
rect 11760 757632 20120 757660
rect 11760 757408 11812 757632
rect 12756 757408 19500 757632
rect 20044 757408 20120 757632
rect 11760 757380 20120 757408
rect 12960 757088 21060 757116
rect 12960 756864 13012 757088
rect 13956 756864 20460 757088
rect 21004 756864 21060 757088
rect 12960 756836 21060 756864
rect 609647 754368 628047 754396
rect 609647 754144 609696 754368
rect 610240 754144 627064 754368
rect 628008 754144 628047 754368
rect 609647 754116 628047 754144
rect 610600 753824 626860 753852
rect 610600 753600 610656 753824
rect 611200 753600 625864 753824
rect 626808 753600 626860 753824
rect 610600 753572 626860 753600
rect 616360 753280 625660 753308
rect 616360 753056 616416 753280
rect 616960 753056 624664 753280
rect 625608 753056 625660 753280
rect 616360 753028 625660 753056
rect 615400 752736 624460 752764
rect 615400 752512 615456 752736
rect 616000 752512 623464 752736
rect 624408 752512 624460 752736
rect 615400 752484 624460 752512
rect 614450 752192 623260 752220
rect 614450 751968 614496 752192
rect 615040 751968 622264 752192
rect 623208 751968 623260 752192
rect 614450 751940 623260 751968
rect 613460 751648 622060 751676
rect 613460 751424 613536 751648
rect 614080 751424 621064 751648
rect 622008 751424 622060 751648
rect 613460 751396 622060 751424
rect 612500 751104 620860 751132
rect 612500 750880 612576 751104
rect 613120 750880 619864 751104
rect 620808 750880 620860 751104
rect 612500 750852 620860 750880
rect 611560 750560 619660 750588
rect 611560 750336 611616 750560
rect 612160 750336 618664 750560
rect 619608 750336 619660 750560
rect 611560 750308 619660 750336
rect 4573 747840 22973 747868
rect 4573 747616 4612 747840
rect 5556 747616 22380 747840
rect 22924 747616 22973 747840
rect 4573 747588 22973 747616
rect 5760 747296 22020 747324
rect 5760 747072 5812 747296
rect 6756 747072 21420 747296
rect 21964 747072 22020 747296
rect 5760 747044 22020 747072
rect 6960 746752 16260 746780
rect 6960 746528 7012 746752
rect 7956 746528 15660 746752
rect 16204 746528 16260 746752
rect 6960 746500 16260 746528
rect 8160 746208 17220 746236
rect 8160 745984 8212 746208
rect 9156 745984 16620 746208
rect 17164 745984 17220 746208
rect 8160 745956 17220 745984
rect 9360 745664 18170 745692
rect 9360 745440 9412 745664
rect 10356 745440 17580 745664
rect 18124 745440 18170 745664
rect 9360 745412 18170 745440
rect 10560 745120 19160 745148
rect 10560 744896 10612 745120
rect 11556 744896 18540 745120
rect 19084 744896 19160 745120
rect 10560 744868 19160 744896
rect 11760 744576 20120 744604
rect 11760 744352 11812 744576
rect 12756 744352 19500 744576
rect 20044 744352 20120 744576
rect 11760 744324 20120 744352
rect 12960 744032 21060 744060
rect 12960 743808 13012 744032
rect 13956 743808 20460 744032
rect 21004 743808 21060 744032
rect 12960 743780 21060 743808
rect 609647 741312 628047 741340
rect 609647 741088 609696 741312
rect 610240 741088 627064 741312
rect 628008 741088 628047 741312
rect 609647 741060 628047 741088
rect 610600 740768 626860 740796
rect 610600 740544 610656 740768
rect 611200 740544 625864 740768
rect 626808 740544 626860 740768
rect 610600 740516 626860 740544
rect 616360 740224 625660 740252
rect 616360 740000 616416 740224
rect 616960 740000 624664 740224
rect 625608 740000 625660 740224
rect 616360 739972 625660 740000
rect 615400 739680 624460 739708
rect 615400 739456 615456 739680
rect 616000 739456 623464 739680
rect 624408 739456 624460 739680
rect 615400 739428 624460 739456
rect 614450 739136 623260 739164
rect 614450 738912 614496 739136
rect 615040 738912 622264 739136
rect 623208 738912 623260 739136
rect 614450 738884 623260 738912
rect 613460 738592 622060 738620
rect 613460 738368 613536 738592
rect 614080 738368 621064 738592
rect 622008 738368 622060 738592
rect 613460 738340 622060 738368
rect 612500 738048 620860 738076
rect 612500 737824 612576 738048
rect 613120 737824 619864 738048
rect 620808 737824 620860 738048
rect 612500 737796 620860 737824
rect 611560 737504 619660 737532
rect 611560 737280 611616 737504
rect 612160 737280 618664 737504
rect 619608 737280 619660 737504
rect 611560 737252 619660 737280
rect 4573 736416 22973 736444
rect 4573 736192 4612 736416
rect 5556 736192 22380 736416
rect 22924 736192 22973 736416
rect 4573 736164 22973 736192
rect 5760 735872 22020 735900
rect 5760 735648 5812 735872
rect 6756 735648 21420 735872
rect 21964 735648 22020 735872
rect 5760 735620 22020 735648
rect 6960 735328 16260 735356
rect 6960 735104 7012 735328
rect 7956 735104 15660 735328
rect 16204 735104 16260 735328
rect 6960 735076 16260 735104
rect 8160 734784 17220 734812
rect 8160 734560 8212 734784
rect 9156 734560 16620 734784
rect 17164 734560 17220 734784
rect 8160 734532 17220 734560
rect 9360 734240 18170 734268
rect 9360 734016 9412 734240
rect 10356 734016 17580 734240
rect 18124 734016 18170 734240
rect 9360 733988 18170 734016
rect 10560 733696 19160 733724
rect 10560 733472 10612 733696
rect 11556 733472 18540 733696
rect 19084 733472 19160 733696
rect 10560 733444 19160 733472
rect 11760 733152 20120 733180
rect 11760 732928 11812 733152
rect 12756 732928 19500 733152
rect 20044 732928 20120 733152
rect 11760 732900 20120 732928
rect 12960 732608 21060 732636
rect 12960 732384 13012 732608
rect 13956 732384 20460 732608
rect 21004 732384 21060 732608
rect 12960 732356 21060 732384
rect 609647 728256 628047 728284
rect 609647 728032 609696 728256
rect 610240 728032 627064 728256
rect 628008 728032 628047 728256
rect 609647 728004 628047 728032
rect 610600 727712 626860 727740
rect 610600 727488 610656 727712
rect 611200 727488 625864 727712
rect 626808 727488 626860 727712
rect 610600 727460 626860 727488
rect 616360 727168 625660 727196
rect 616360 726944 616416 727168
rect 616960 726944 624664 727168
rect 625608 726944 625660 727168
rect 616360 726916 625660 726944
rect 615400 726624 624460 726652
rect 615400 726400 615456 726624
rect 616000 726400 623464 726624
rect 624408 726400 624460 726624
rect 615400 726372 624460 726400
rect 614450 726080 623260 726108
rect 614450 725856 614496 726080
rect 615040 725856 622264 726080
rect 623208 725856 623260 726080
rect 614450 725828 623260 725856
rect 613460 725536 622060 725564
rect 613460 725312 613536 725536
rect 614080 725312 621064 725536
rect 622008 725312 622060 725536
rect 613460 725284 622060 725312
rect 612500 724992 620860 725020
rect 612500 724768 612576 724992
rect 613120 724768 619864 724992
rect 620808 724768 620860 724992
rect 612500 724740 620860 724768
rect 611560 724448 619660 724476
rect 611560 724224 611616 724448
rect 612160 724224 618664 724448
rect 619608 724224 619660 724448
rect 611560 724196 619660 724224
rect 4573 721728 22973 721756
rect 4573 721504 4612 721728
rect 5556 721504 22380 721728
rect 22924 721504 22973 721728
rect 4573 721476 22973 721504
rect 5760 721184 22020 721212
rect 5760 720960 5812 721184
rect 6756 720960 21420 721184
rect 21964 720960 22020 721184
rect 5760 720932 22020 720960
rect 6960 720640 16260 720668
rect 6960 720416 7012 720640
rect 7956 720416 15660 720640
rect 16204 720416 16260 720640
rect 6960 720388 16260 720416
rect 8160 720096 17220 720124
rect 8160 719872 8212 720096
rect 9156 719872 16620 720096
rect 17164 719872 17220 720096
rect 8160 719844 17220 719872
rect 9360 719552 18170 719580
rect 9360 719328 9412 719552
rect 10356 719328 17580 719552
rect 18124 719328 18170 719552
rect 9360 719300 18170 719328
rect 10560 719008 19160 719036
rect 10560 718784 10612 719008
rect 11556 718784 18540 719008
rect 19084 718784 19160 719008
rect 10560 718756 19160 718784
rect 11760 718464 20120 718492
rect 11760 718240 11812 718464
rect 12756 718240 19500 718464
rect 20044 718240 20120 718464
rect 11760 718212 20120 718240
rect 12960 717920 21060 717948
rect 12960 717696 13012 717920
rect 13956 717696 20460 717920
rect 21004 717696 21060 717920
rect 12960 717668 21060 717696
rect 609647 713568 628047 713596
rect 609647 713344 609696 713568
rect 610240 713344 627064 713568
rect 628008 713344 628047 713568
rect 609647 713316 628047 713344
rect 610600 713024 626860 713052
rect 610600 712800 610656 713024
rect 611200 712800 625864 713024
rect 626808 712800 626860 713024
rect 610600 712772 626860 712800
rect 616360 712480 625660 712508
rect 616360 712256 616416 712480
rect 616960 712256 624664 712480
rect 625608 712256 625660 712480
rect 616360 712228 625660 712256
rect 615400 711936 624460 711964
rect 615400 711712 615456 711936
rect 616000 711712 623464 711936
rect 624408 711712 624460 711936
rect 615400 711684 624460 711712
rect 614450 711392 623260 711420
rect 614450 711168 614496 711392
rect 615040 711168 622264 711392
rect 623208 711168 623260 711392
rect 614450 711140 623260 711168
rect 613460 710848 622060 710876
rect 613460 710624 613536 710848
rect 614080 710624 621064 710848
rect 622008 710624 622060 710848
rect 613460 710596 622060 710624
rect 612500 710304 620860 710332
rect 612500 710080 612576 710304
rect 613120 710080 619864 710304
rect 620808 710080 620860 710304
rect 612500 710052 620860 710080
rect 611560 709760 619660 709788
rect 611560 709536 611616 709760
rect 612160 709536 618664 709760
rect 619608 709536 619660 709760
rect 611560 709508 619660 709536
rect 4573 708672 22973 708700
rect 4573 708448 4612 708672
rect 5556 708448 22380 708672
rect 22924 708448 22973 708672
rect 4573 708420 22973 708448
rect 5760 708128 22020 708156
rect 5760 707904 5812 708128
rect 6756 707904 21420 708128
rect 21964 707904 22020 708128
rect 5760 707876 22020 707904
rect 6960 707584 16260 707612
rect 6960 707360 7012 707584
rect 7956 707360 15660 707584
rect 16204 707360 16260 707584
rect 6960 707332 16260 707360
rect 8160 707040 17220 707068
rect 8160 706816 8212 707040
rect 9156 706816 16620 707040
rect 17164 706816 17220 707040
rect 8160 706788 17220 706816
rect 9360 706496 18170 706524
rect 9360 706272 9412 706496
rect 10356 706272 17580 706496
rect 18124 706272 18170 706496
rect 9360 706244 18170 706272
rect 10560 705952 19160 705980
rect 10560 705728 10612 705952
rect 11556 705728 18540 705952
rect 19084 705728 19160 705952
rect 10560 705700 19160 705728
rect 11760 705408 20120 705436
rect 11760 705184 11812 705408
rect 12756 705184 19500 705408
rect 20044 705184 20120 705408
rect 11760 705156 20120 705184
rect 12960 704864 21060 704892
rect 12960 704640 13012 704864
rect 13956 704640 20460 704864
rect 21004 704640 21060 704864
rect 12960 704612 21060 704640
rect 609647 702144 628047 702172
rect 609647 701920 609696 702144
rect 610240 701920 627064 702144
rect 628008 701920 628047 702144
rect 609647 701892 628047 701920
rect 610600 701600 626860 701628
rect 610600 701376 610656 701600
rect 611200 701376 625864 701600
rect 626808 701376 626860 701600
rect 610600 701348 626860 701376
rect 616360 701056 625660 701084
rect 616360 700832 616416 701056
rect 616960 700832 624664 701056
rect 625608 700832 625660 701056
rect 616360 700804 625660 700832
rect 615400 700512 624460 700540
rect 615400 700288 615456 700512
rect 616000 700288 623464 700512
rect 624408 700288 624460 700512
rect 615400 700260 624460 700288
rect 614450 699968 623260 699996
rect 614450 699744 614496 699968
rect 615040 699744 622264 699968
rect 623208 699744 623260 699968
rect 614450 699716 623260 699744
rect 613460 699424 622060 699452
rect 613460 699200 613536 699424
rect 614080 699200 621064 699424
rect 622008 699200 622060 699424
rect 613460 699172 622060 699200
rect 612500 698880 620860 698908
rect 612500 698656 612576 698880
rect 613120 698656 619864 698880
rect 620808 698656 620860 698880
rect 612500 698628 620860 698656
rect 611560 698336 619660 698364
rect 611560 698112 611616 698336
rect 612160 698112 618664 698336
rect 619608 698112 619660 698336
rect 611560 698084 619660 698112
rect 4573 692352 22973 692380
rect 4573 692128 4612 692352
rect 5556 692128 22380 692352
rect 22924 692128 22973 692352
rect 4573 692100 22973 692128
rect 5760 691808 22020 691836
rect 5760 691584 5812 691808
rect 6756 691584 21420 691808
rect 21964 691584 22020 691808
rect 5760 691556 22020 691584
rect 6960 691264 16260 691292
rect 6960 691040 7012 691264
rect 7956 691040 15660 691264
rect 16204 691040 16260 691264
rect 6960 691012 16260 691040
rect 8160 690720 17220 690748
rect 8160 690496 8212 690720
rect 9156 690496 16620 690720
rect 17164 690496 17220 690720
rect 8160 690468 17220 690496
rect 9360 690176 18170 690204
rect 9360 689952 9412 690176
rect 10356 689952 17580 690176
rect 18124 689952 18170 690176
rect 9360 689924 18170 689952
rect 10560 689632 19160 689660
rect 10560 689408 10612 689632
rect 11556 689408 18540 689632
rect 19084 689408 19160 689632
rect 10560 689380 19160 689408
rect 11760 689088 20120 689116
rect 11760 688864 11812 689088
rect 12756 688864 19500 689088
rect 20044 688864 20120 689088
rect 11760 688836 20120 688864
rect 609647 689088 628047 689116
rect 609647 688864 609696 689088
rect 610240 688864 627064 689088
rect 628008 688864 628047 689088
rect 609647 688836 628047 688864
rect 12960 688544 21060 688572
rect 12960 688320 13012 688544
rect 13956 688320 20460 688544
rect 21004 688320 21060 688544
rect 12960 688292 21060 688320
rect 610600 688544 626860 688572
rect 610600 688320 610656 688544
rect 611200 688320 625864 688544
rect 626808 688320 626860 688544
rect 610600 688292 626860 688320
rect 616360 688000 625660 688028
rect 616360 687776 616416 688000
rect 616960 687776 624664 688000
rect 625608 687776 625660 688000
rect 616360 687748 625660 687776
rect 615400 687456 624460 687484
rect 615400 687232 615456 687456
rect 616000 687232 623464 687456
rect 624408 687232 624460 687456
rect 615400 687204 624460 687232
rect 614450 686912 623260 686940
rect 614450 686688 614496 686912
rect 615040 686688 622264 686912
rect 623208 686688 623260 686912
rect 614450 686660 623260 686688
rect 613460 686368 622060 686396
rect 613460 686144 613536 686368
rect 614080 686144 621064 686368
rect 622008 686144 622060 686368
rect 613460 686116 622060 686144
rect 612500 685824 620860 685852
rect 612500 685600 612576 685824
rect 613120 685600 619864 685824
rect 620808 685600 620860 685824
rect 612500 685572 620860 685600
rect 611560 685280 619660 685308
rect 611560 685056 611616 685280
rect 612160 685056 618664 685280
rect 619608 685056 619660 685280
rect 611560 685028 619660 685056
rect 4573 682560 22973 682588
rect 4573 682336 4612 682560
rect 5556 682336 22380 682560
rect 22924 682336 22973 682560
rect 4573 682308 22973 682336
rect 5760 682016 22020 682044
rect 5760 681792 5812 682016
rect 6756 681792 21420 682016
rect 21964 681792 22020 682016
rect 5760 681764 22020 681792
rect 6960 681472 16260 681500
rect 6960 681248 7012 681472
rect 7956 681248 15660 681472
rect 16204 681248 16260 681472
rect 6960 681220 16260 681248
rect 8160 680928 17220 680956
rect 8160 680704 8212 680928
rect 9156 680704 16620 680928
rect 17164 680704 17220 680928
rect 8160 680676 17220 680704
rect 9360 680384 18170 680412
rect 9360 680160 9412 680384
rect 10356 680160 17580 680384
rect 18124 680160 18170 680384
rect 9360 680132 18170 680160
rect 10560 679840 19160 679868
rect 10560 679616 10612 679840
rect 11556 679616 18540 679840
rect 19084 679616 19160 679840
rect 10560 679588 19160 679616
rect 11760 679296 20120 679324
rect 11760 679072 11812 679296
rect 12756 679072 19500 679296
rect 20044 679072 20120 679296
rect 11760 679044 20120 679072
rect 12960 678752 21060 678780
rect 12960 678528 13012 678752
rect 13956 678528 20460 678752
rect 21004 678528 21060 678752
rect 12960 678500 21060 678528
rect 609647 676032 628047 676060
rect 609647 675808 609696 676032
rect 610240 675808 627064 676032
rect 628008 675808 628047 676032
rect 609647 675780 628047 675808
rect 610600 675488 626860 675516
rect 610600 675264 610656 675488
rect 611200 675264 625864 675488
rect 626808 675264 626860 675488
rect 610600 675236 626860 675264
rect 616360 674944 625660 674972
rect 616360 674720 616416 674944
rect 616960 674720 624664 674944
rect 625608 674720 625660 674944
rect 616360 674692 625660 674720
rect 615400 674400 624460 674428
rect 615400 674176 615456 674400
rect 616000 674176 623464 674400
rect 624408 674176 624460 674400
rect 615400 674148 624460 674176
rect 614450 673856 623260 673884
rect 614450 673632 614496 673856
rect 615040 673632 622264 673856
rect 623208 673632 623260 673856
rect 614450 673604 623260 673632
rect 613460 673312 622060 673340
rect 613460 673088 613536 673312
rect 614080 673088 621064 673312
rect 622008 673088 622060 673312
rect 613460 673060 622060 673088
rect 612500 672768 620860 672796
rect 612500 672544 612576 672768
rect 613120 672544 619864 672768
rect 620808 672544 620860 672768
rect 612500 672516 620860 672544
rect 611560 672224 619660 672252
rect 611560 672000 611616 672224
rect 612160 672000 618664 672224
rect 619608 672000 619660 672224
rect 611560 671972 619660 672000
rect 4573 669504 22973 669532
rect 4573 669280 4612 669504
rect 5556 669280 22380 669504
rect 22924 669280 22973 669504
rect 4573 669252 22973 669280
rect 5760 668960 22020 668988
rect 5760 668736 5812 668960
rect 6756 668736 21420 668960
rect 21964 668736 22020 668960
rect 5760 668708 22020 668736
rect 6960 668416 16260 668444
rect 6960 668192 7012 668416
rect 7956 668192 15660 668416
rect 16204 668192 16260 668416
rect 6960 668164 16260 668192
rect 8160 667872 17220 667900
rect 8160 667648 8212 667872
rect 9156 667648 16620 667872
rect 17164 667648 17220 667872
rect 8160 667620 17220 667648
rect 9360 667328 18170 667356
rect 9360 667104 9412 667328
rect 10356 667104 17580 667328
rect 18124 667104 18170 667328
rect 9360 667076 18170 667104
rect 10560 666784 19160 666812
rect 10560 666560 10612 666784
rect 11556 666560 18540 666784
rect 19084 666560 19160 666784
rect 10560 666532 19160 666560
rect 11760 666240 20120 666268
rect 11760 666016 11812 666240
rect 12756 666016 19500 666240
rect 20044 666016 20120 666240
rect 11760 665988 20120 666016
rect 12960 665696 21060 665724
rect 12960 665472 13012 665696
rect 13956 665472 20460 665696
rect 21004 665472 21060 665696
rect 12960 665444 21060 665472
rect 609647 662976 628047 663004
rect 609647 662752 609696 662976
rect 610240 662752 627064 662976
rect 628008 662752 628047 662976
rect 609647 662724 628047 662752
rect 610600 662432 626860 662460
rect 610600 662208 610656 662432
rect 611200 662208 625864 662432
rect 626808 662208 626860 662432
rect 610600 662180 626860 662208
rect 616360 661888 625660 661916
rect 616360 661664 616416 661888
rect 616960 661664 624664 661888
rect 625608 661664 625660 661888
rect 616360 661636 625660 661664
rect 615400 661344 624460 661372
rect 615400 661120 615456 661344
rect 616000 661120 623464 661344
rect 624408 661120 624460 661344
rect 615400 661092 624460 661120
rect 614450 660800 623260 660828
rect 614450 660576 614496 660800
rect 615040 660576 622264 660800
rect 623208 660576 623260 660800
rect 614450 660548 623260 660576
rect 613460 660256 622060 660284
rect 613460 660032 613536 660256
rect 614080 660032 621064 660256
rect 622008 660032 622060 660256
rect 613460 660004 622060 660032
rect 612500 659712 620860 659740
rect 612500 659488 612576 659712
rect 613120 659488 619864 659712
rect 620808 659488 620860 659712
rect 612500 659460 620860 659488
rect 611560 659168 619660 659196
rect 611560 658944 611616 659168
rect 612160 658944 618664 659168
rect 619608 658944 619660 659168
rect 611560 658916 619660 658944
rect 4573 656448 22973 656476
rect 4573 656224 4612 656448
rect 5556 656224 22380 656448
rect 22924 656224 22973 656448
rect 4573 656196 22973 656224
rect 5760 655904 22020 655932
rect 5760 655680 5812 655904
rect 6756 655680 21420 655904
rect 21964 655680 22020 655904
rect 5760 655652 22020 655680
rect 6960 655360 16260 655388
rect 6960 655136 7012 655360
rect 7956 655136 15660 655360
rect 16204 655136 16260 655360
rect 6960 655108 16260 655136
rect 8160 654816 17220 654844
rect 8160 654592 8212 654816
rect 9156 654592 16620 654816
rect 17164 654592 17220 654816
rect 8160 654564 17220 654592
rect 9360 654272 18170 654300
rect 9360 654048 9412 654272
rect 10356 654048 17580 654272
rect 18124 654048 18170 654272
rect 9360 654020 18170 654048
rect 10560 653728 19160 653756
rect 10560 653504 10612 653728
rect 11556 653504 18540 653728
rect 19084 653504 19160 653728
rect 10560 653476 19160 653504
rect 11760 653184 20120 653212
rect 11760 652960 11812 653184
rect 12756 652960 19500 653184
rect 20044 652960 20120 653184
rect 11760 652932 20120 652960
rect 12960 652640 21060 652668
rect 12960 652416 13012 652640
rect 13956 652416 20460 652640
rect 21004 652416 21060 652640
rect 12960 652388 21060 652416
rect 609647 649920 628047 649948
rect 609647 649696 609696 649920
rect 610240 649696 627064 649920
rect 628008 649696 628047 649920
rect 609647 649668 628047 649696
rect 610600 649376 626860 649404
rect 610600 649152 610656 649376
rect 611200 649152 625864 649376
rect 626808 649152 626860 649376
rect 610600 649124 626860 649152
rect 616360 648832 625660 648860
rect 616360 648608 616416 648832
rect 616960 648608 624664 648832
rect 625608 648608 625660 648832
rect 616360 648580 625660 648608
rect 615400 648288 624460 648316
rect 615400 648064 615456 648288
rect 616000 648064 623464 648288
rect 624408 648064 624460 648288
rect 615400 648036 624460 648064
rect 614450 647744 623260 647772
rect 614450 647520 614496 647744
rect 615040 647520 622264 647744
rect 623208 647520 623260 647744
rect 614450 647492 623260 647520
rect 613460 647200 622060 647228
rect 613460 646976 613536 647200
rect 614080 646976 621064 647200
rect 622008 646976 622060 647200
rect 613460 646948 622060 646976
rect 612500 646656 620860 646684
rect 612500 646432 612576 646656
rect 613120 646432 619864 646656
rect 620808 646432 620860 646656
rect 612500 646404 620860 646432
rect 611560 646112 619660 646140
rect 611560 645888 611616 646112
rect 612160 645888 618664 646112
rect 619608 645888 619660 646112
rect 611560 645860 619660 645888
rect 4573 641760 22973 641788
rect 4573 641536 4612 641760
rect 5556 641536 22380 641760
rect 22924 641536 22973 641760
rect 4573 641508 22973 641536
rect 5760 641216 22020 641244
rect 5760 640992 5812 641216
rect 6756 640992 21420 641216
rect 21964 640992 22020 641216
rect 5760 640964 22020 640992
rect 6960 640672 16260 640700
rect 6960 640448 7012 640672
rect 7956 640448 15660 640672
rect 16204 640448 16260 640672
rect 6960 640420 16260 640448
rect 8160 640128 17220 640156
rect 8160 639904 8212 640128
rect 9156 639904 16620 640128
rect 17164 639904 17220 640128
rect 8160 639876 17220 639904
rect 9360 639584 18170 639612
rect 9360 639360 9412 639584
rect 10356 639360 17580 639584
rect 18124 639360 18170 639584
rect 9360 639332 18170 639360
rect 10560 639040 19160 639068
rect 10560 638816 10612 639040
rect 11556 638816 18540 639040
rect 19084 638816 19160 639040
rect 10560 638788 19160 638816
rect 11760 638496 20120 638524
rect 11760 638272 11812 638496
rect 12756 638272 19500 638496
rect 20044 638272 20120 638496
rect 11760 638244 20120 638272
rect 12960 637952 21060 637980
rect 12960 637728 13012 637952
rect 13956 637728 20460 637952
rect 21004 637728 21060 637952
rect 12960 637700 21060 637728
rect 609647 636864 628047 636892
rect 609647 636640 609696 636864
rect 610240 636640 627064 636864
rect 628008 636640 628047 636864
rect 609647 636612 628047 636640
rect 610600 636320 626860 636348
rect 610600 636096 610656 636320
rect 611200 636096 625864 636320
rect 626808 636096 626860 636320
rect 610600 636068 626860 636096
rect 616360 635776 625660 635804
rect 616360 635552 616416 635776
rect 616960 635552 624664 635776
rect 625608 635552 625660 635776
rect 616360 635524 625660 635552
rect 615400 635232 624460 635260
rect 615400 635008 615456 635232
rect 616000 635008 623464 635232
rect 624408 635008 624460 635232
rect 615400 634980 624460 635008
rect 614450 634688 623260 634716
rect 614450 634464 614496 634688
rect 615040 634464 622264 634688
rect 623208 634464 623260 634688
rect 614450 634436 623260 634464
rect 613460 634144 622060 634172
rect 613460 633920 613536 634144
rect 614080 633920 621064 634144
rect 622008 633920 622060 634144
rect 613460 633892 622060 633920
rect 612500 633600 620860 633628
rect 612500 633376 612576 633600
rect 613120 633376 619864 633600
rect 620808 633376 620860 633600
rect 612500 633348 620860 633376
rect 611560 633056 619660 633084
rect 611560 632832 611616 633056
rect 612160 632832 618664 633056
rect 619608 632832 619660 633056
rect 611560 632804 619660 632832
rect 4573 630336 22973 630364
rect 4573 630112 4612 630336
rect 5556 630112 22380 630336
rect 22924 630112 22973 630336
rect 4573 630084 22973 630112
rect 5760 629792 22020 629820
rect 5760 629568 5812 629792
rect 6756 629568 21420 629792
rect 21964 629568 22020 629792
rect 5760 629540 22020 629568
rect 6960 629248 16260 629276
rect 6960 629024 7012 629248
rect 7956 629024 15660 629248
rect 16204 629024 16260 629248
rect 6960 628996 16260 629024
rect 8160 628704 17220 628732
rect 8160 628480 8212 628704
rect 9156 628480 16620 628704
rect 17164 628480 17220 628704
rect 8160 628452 17220 628480
rect 9360 628160 18170 628188
rect 9360 627936 9412 628160
rect 10356 627936 17580 628160
rect 18124 627936 18170 628160
rect 9360 627908 18170 627936
rect 10560 627616 19160 627644
rect 10560 627392 10612 627616
rect 11556 627392 18540 627616
rect 19084 627392 19160 627616
rect 10560 627364 19160 627392
rect 11760 627072 20120 627100
rect 11760 626848 11812 627072
rect 12756 626848 19500 627072
rect 20044 626848 20120 627072
rect 11760 626820 20120 626848
rect 12960 626528 21060 626556
rect 12960 626304 13012 626528
rect 13956 626304 20460 626528
rect 21004 626304 21060 626528
rect 12960 626276 21060 626304
rect 609647 623808 628047 623836
rect 609647 623584 609696 623808
rect 610240 623584 627064 623808
rect 628008 623584 628047 623808
rect 609647 623556 628047 623584
rect 610600 623264 626860 623292
rect 610600 623040 610656 623264
rect 611200 623040 625864 623264
rect 626808 623040 626860 623264
rect 610600 623012 626860 623040
rect 616360 622720 625660 622748
rect 616360 622496 616416 622720
rect 616960 622496 624664 622720
rect 625608 622496 625660 622720
rect 616360 622468 625660 622496
rect 615400 622176 624460 622204
rect 615400 621952 615456 622176
rect 616000 621952 623464 622176
rect 624408 621952 624460 622176
rect 615400 621924 624460 621952
rect 614450 621632 623260 621660
rect 614450 621408 614496 621632
rect 615040 621408 622264 621632
rect 623208 621408 623260 621632
rect 614450 621380 623260 621408
rect 613460 621088 622060 621116
rect 613460 620864 613536 621088
rect 614080 620864 621064 621088
rect 622008 620864 622060 621088
rect 613460 620836 622060 620864
rect 612500 620544 620860 620572
rect 612500 620320 612576 620544
rect 613120 620320 619864 620544
rect 620808 620320 620860 620544
rect 612500 620292 620860 620320
rect 611560 620000 619660 620028
rect 611560 619776 611616 620000
rect 612160 619776 618664 620000
rect 619608 619776 619660 620000
rect 611560 619748 619660 619776
rect 4573 617280 22973 617308
rect 4573 617056 4612 617280
rect 5556 617056 22380 617280
rect 22924 617056 22973 617280
rect 4573 617028 22973 617056
rect 5760 616736 22020 616764
rect 5760 616512 5812 616736
rect 6756 616512 21420 616736
rect 21964 616512 22020 616736
rect 5760 616484 22020 616512
rect 6960 616192 16260 616220
rect 6960 615968 7012 616192
rect 7956 615968 15660 616192
rect 16204 615968 16260 616192
rect 6960 615940 16260 615968
rect 8160 615648 17220 615676
rect 8160 615424 8212 615648
rect 9156 615424 16620 615648
rect 17164 615424 17220 615648
rect 8160 615396 17220 615424
rect 9360 615104 18170 615132
rect 9360 614880 9412 615104
rect 10356 614880 17580 615104
rect 18124 614880 18170 615104
rect 9360 614852 18170 614880
rect 10560 614560 19160 614588
rect 10560 614336 10612 614560
rect 11556 614336 18540 614560
rect 19084 614336 19160 614560
rect 10560 614308 19160 614336
rect 11760 614016 20120 614044
rect 11760 613792 11812 614016
rect 12756 613792 19500 614016
rect 20044 613792 20120 614016
rect 11760 613764 20120 613792
rect 12960 613472 21060 613500
rect 12960 613248 13012 613472
rect 13956 613248 20460 613472
rect 21004 613248 21060 613472
rect 12960 613220 21060 613248
rect 609647 610752 628047 610780
rect 609647 610528 609696 610752
rect 610240 610528 627064 610752
rect 628008 610528 628047 610752
rect 609647 610500 628047 610528
rect 610600 610208 626860 610236
rect 610600 609984 610656 610208
rect 611200 609984 625864 610208
rect 626808 609984 626860 610208
rect 610600 609956 626860 609984
rect 616360 609664 625660 609692
rect 616360 609440 616416 609664
rect 616960 609440 624664 609664
rect 625608 609440 625660 609664
rect 616360 609412 625660 609440
rect 615400 609120 624460 609148
rect 615400 608896 615456 609120
rect 616000 608896 623464 609120
rect 624408 608896 624460 609120
rect 615400 608868 624460 608896
rect 614450 608576 623260 608604
rect 614450 608352 614496 608576
rect 615040 608352 622264 608576
rect 623208 608352 623260 608576
rect 614450 608324 623260 608352
rect 613460 608032 622060 608060
rect 613460 607808 613536 608032
rect 614080 607808 621064 608032
rect 622008 607808 622060 608032
rect 613460 607780 622060 607808
rect 612500 607488 620860 607516
rect 612500 607264 612576 607488
rect 613120 607264 619864 607488
rect 620808 607264 620860 607488
rect 612500 607236 620860 607264
rect 611560 606944 619660 606972
rect 611560 606720 611616 606944
rect 612160 606720 618664 606944
rect 619608 606720 619660 606944
rect 611560 606692 619660 606720
rect 4573 606400 22973 606428
rect 4573 606176 4612 606400
rect 5556 606176 22380 606400
rect 22924 606176 22973 606400
rect 4573 606148 22973 606176
rect 5760 605856 22020 605884
rect 5760 605632 5812 605856
rect 6756 605632 21420 605856
rect 21964 605632 22020 605856
rect 5760 605604 22020 605632
rect 6960 605312 16260 605340
rect 6960 605088 7012 605312
rect 7956 605088 15660 605312
rect 16204 605088 16260 605312
rect 6960 605060 16260 605088
rect 8160 604768 17220 604796
rect 8160 604544 8212 604768
rect 9156 604544 16620 604768
rect 17164 604544 17220 604768
rect 8160 604516 17220 604544
rect 9360 604224 18170 604252
rect 9360 604000 9412 604224
rect 10356 604000 17580 604224
rect 18124 604000 18170 604224
rect 9360 603972 18170 604000
rect 10560 603680 19160 603708
rect 10560 603456 10612 603680
rect 11556 603456 18540 603680
rect 19084 603456 19160 603680
rect 10560 603428 19160 603456
rect 11760 603136 20120 603164
rect 11760 602912 11812 603136
rect 12756 602912 19500 603136
rect 20044 602912 20120 603136
rect 11760 602884 20120 602912
rect 12960 602592 21060 602620
rect 12960 602368 13012 602592
rect 13956 602368 20460 602592
rect 21004 602368 21060 602592
rect 12960 602340 21060 602368
rect 609647 597696 628047 597724
rect 609647 597472 609696 597696
rect 610240 597472 627064 597696
rect 628008 597472 628047 597696
rect 609647 597444 628047 597472
rect 610600 597152 626860 597180
rect 610600 596928 610656 597152
rect 611200 596928 625864 597152
rect 626808 596928 626860 597152
rect 610600 596900 626860 596928
rect 616360 596608 625660 596636
rect 616360 596384 616416 596608
rect 616960 596384 624664 596608
rect 625608 596384 625660 596608
rect 616360 596356 625660 596384
rect 615400 596064 624460 596092
rect 615400 595840 615456 596064
rect 616000 595840 623464 596064
rect 624408 595840 624460 596064
rect 615400 595812 624460 595840
rect 614450 595520 623260 595548
rect 614450 595296 614496 595520
rect 615040 595296 622264 595520
rect 623208 595296 623260 595520
rect 614450 595268 623260 595296
rect 613460 594976 622060 595004
rect 613460 594752 613536 594976
rect 614080 594752 621064 594976
rect 622008 594752 622060 594976
rect 613460 594724 622060 594752
rect 612500 594432 620860 594460
rect 612500 594208 612576 594432
rect 613120 594208 619864 594432
rect 620808 594208 620860 594432
rect 612500 594180 620860 594208
rect 611560 593888 619660 593916
rect 611560 593664 611616 593888
rect 612160 593664 618664 593888
rect 619608 593664 619660 593888
rect 611560 593636 619660 593664
rect 4573 591168 22973 591196
rect 4573 590944 4612 591168
rect 5556 590944 22380 591168
rect 22924 590944 22973 591168
rect 4573 590916 22973 590944
rect 5760 590624 22020 590652
rect 5760 590400 5812 590624
rect 6756 590400 21420 590624
rect 21964 590400 22020 590624
rect 5760 590372 22020 590400
rect 6960 590080 16260 590108
rect 6960 589856 7012 590080
rect 7956 589856 15660 590080
rect 16204 589856 16260 590080
rect 6960 589828 16260 589856
rect 8160 589536 17220 589564
rect 8160 589312 8212 589536
rect 9156 589312 16620 589536
rect 17164 589312 17220 589536
rect 8160 589284 17220 589312
rect 9360 588992 18170 589020
rect 9360 588768 9412 588992
rect 10356 588768 17580 588992
rect 18124 588768 18170 588992
rect 9360 588740 18170 588768
rect 10560 588448 19160 588476
rect 10560 588224 10612 588448
rect 11556 588224 18540 588448
rect 19084 588224 19160 588448
rect 10560 588196 19160 588224
rect 11760 587904 20120 587932
rect 11760 587680 11812 587904
rect 12756 587680 19500 587904
rect 20044 587680 20120 587904
rect 11760 587652 20120 587680
rect 12960 587360 21060 587388
rect 12960 587136 13012 587360
rect 13956 587136 20460 587360
rect 21004 587136 21060 587360
rect 12960 587108 21060 587136
rect 609647 584640 628047 584668
rect 609647 584416 609696 584640
rect 610240 584416 627064 584640
rect 628008 584416 628047 584640
rect 609647 584388 628047 584416
rect 610600 584096 626860 584124
rect 610600 583872 610656 584096
rect 611200 583872 625864 584096
rect 626808 583872 626860 584096
rect 610600 583844 626860 583872
rect 616360 583552 625660 583580
rect 616360 583328 616416 583552
rect 616960 583328 624664 583552
rect 625608 583328 625660 583552
rect 616360 583300 625660 583328
rect 615400 583008 624460 583036
rect 615400 582784 615456 583008
rect 616000 582784 623464 583008
rect 624408 582784 624460 583008
rect 615400 582756 624460 582784
rect 614450 582464 623260 582492
rect 614450 582240 614496 582464
rect 615040 582240 622264 582464
rect 623208 582240 623260 582464
rect 614450 582212 623260 582240
rect 613460 581920 622060 581948
rect 613460 581696 613536 581920
rect 614080 581696 621064 581920
rect 622008 581696 622060 581920
rect 613460 581668 622060 581696
rect 612500 581376 620860 581404
rect 612500 581152 612576 581376
rect 613120 581152 619864 581376
rect 620808 581152 620860 581376
rect 612500 581124 620860 581152
rect 611560 580832 619660 580860
rect 611560 580608 611616 580832
rect 612160 580608 618664 580832
rect 619608 580608 619660 580832
rect 611560 580580 619660 580608
rect 4573 578112 22973 578140
rect 4573 577888 4612 578112
rect 5556 577888 22380 578112
rect 22924 577888 22973 578112
rect 4573 577860 22973 577888
rect 5760 577568 22020 577596
rect 5760 577344 5812 577568
rect 6756 577344 21420 577568
rect 21964 577344 22020 577568
rect 5760 577316 22020 577344
rect 6960 577024 16260 577052
rect 6960 576800 7012 577024
rect 7956 576800 15660 577024
rect 16204 576800 16260 577024
rect 6960 576772 16260 576800
rect 8160 576480 17220 576508
rect 8160 576256 8212 576480
rect 9156 576256 16620 576480
rect 17164 576256 17220 576480
rect 8160 576228 17220 576256
rect 9360 575936 18170 575964
rect 9360 575712 9412 575936
rect 10356 575712 17580 575936
rect 18124 575712 18170 575936
rect 9360 575684 18170 575712
rect 10560 575392 19160 575420
rect 10560 575168 10612 575392
rect 11556 575168 18540 575392
rect 19084 575168 19160 575392
rect 10560 575140 19160 575168
rect 11760 574848 20120 574876
rect 11760 574624 11812 574848
rect 12756 574624 19500 574848
rect 20044 574624 20120 574848
rect 11760 574596 20120 574624
rect 12960 574304 21060 574332
rect 12960 574080 13012 574304
rect 13956 574080 20460 574304
rect 21004 574080 21060 574304
rect 12960 574052 21060 574080
rect 609647 571584 628047 571612
rect 609647 571360 609696 571584
rect 610240 571360 627064 571584
rect 628008 571360 628047 571584
rect 609647 571332 628047 571360
rect 610600 571040 626860 571068
rect 610600 570816 610656 571040
rect 611200 570816 625864 571040
rect 626808 570816 626860 571040
rect 610600 570788 626860 570816
rect 616360 570496 625660 570524
rect 616360 570272 616416 570496
rect 616960 570272 624664 570496
rect 625608 570272 625660 570496
rect 616360 570244 625660 570272
rect 615400 569952 624460 569980
rect 615400 569728 615456 569952
rect 616000 569728 623464 569952
rect 624408 569728 624460 569952
rect 615400 569700 624460 569728
rect 614450 569408 623260 569436
rect 614450 569184 614496 569408
rect 615040 569184 622264 569408
rect 623208 569184 623260 569408
rect 614450 569156 623260 569184
rect 613460 568864 622060 568892
rect 613460 568640 613536 568864
rect 614080 568640 621064 568864
rect 622008 568640 622060 568864
rect 613460 568612 622060 568640
rect 612500 568320 620860 568348
rect 612500 568096 612576 568320
rect 613120 568096 619864 568320
rect 620808 568096 620860 568320
rect 612500 568068 620860 568096
rect 611560 567776 619660 567804
rect 611560 567552 611616 567776
rect 612160 567552 618664 567776
rect 619608 567552 619660 567776
rect 611560 567524 619660 567552
rect 4573 567232 22973 567260
rect 4573 567008 4612 567232
rect 5556 567008 22380 567232
rect 22924 567008 22973 567232
rect 4573 566980 22973 567008
rect 5760 566688 22020 566716
rect 5760 566464 5812 566688
rect 6756 566464 21420 566688
rect 21964 566464 22020 566688
rect 5760 566436 22020 566464
rect 6960 566144 16260 566172
rect 6960 565920 7012 566144
rect 7956 565920 15660 566144
rect 16204 565920 16260 566144
rect 6960 565892 16260 565920
rect 8160 565600 17220 565628
rect 8160 565376 8212 565600
rect 9156 565376 16620 565600
rect 17164 565376 17220 565600
rect 8160 565348 17220 565376
rect 9360 565056 18170 565084
rect 9360 564832 9412 565056
rect 10356 564832 17580 565056
rect 18124 564832 18170 565056
rect 9360 564804 18170 564832
rect 10560 564512 19160 564540
rect 10560 564288 10612 564512
rect 11556 564288 18540 564512
rect 19084 564288 19160 564512
rect 10560 564260 19160 564288
rect 11760 563968 20120 563996
rect 11760 563744 11812 563968
rect 12756 563744 19500 563968
rect 20044 563744 20120 563968
rect 11760 563716 20120 563744
rect 12960 563424 21060 563452
rect 12960 563200 13012 563424
rect 13956 563200 20460 563424
rect 21004 563200 21060 563424
rect 12960 563172 21060 563200
rect 609647 558528 628047 558556
rect 609647 558304 609696 558528
rect 610240 558304 627064 558528
rect 628008 558304 628047 558528
rect 609647 558276 628047 558304
rect 610600 557984 626860 558012
rect 610600 557760 610656 557984
rect 611200 557760 625864 557984
rect 626808 557760 626860 557984
rect 610600 557732 626860 557760
rect 616360 557440 625660 557468
rect 616360 557216 616416 557440
rect 616960 557216 624664 557440
rect 625608 557216 625660 557440
rect 616360 557188 625660 557216
rect 615400 556896 624460 556924
rect 615400 556672 615456 556896
rect 616000 556672 623464 556896
rect 624408 556672 624460 556896
rect 615400 556644 624460 556672
rect 614450 556352 623260 556380
rect 614450 556128 614496 556352
rect 615040 556128 622264 556352
rect 623208 556128 623260 556352
rect 614450 556100 623260 556128
rect 613460 555808 622060 555836
rect 613460 555584 613536 555808
rect 614080 555584 621064 555808
rect 622008 555584 622060 555808
rect 613460 555556 622060 555584
rect 612500 555264 620860 555292
rect 612500 555040 612576 555264
rect 613120 555040 619864 555264
rect 620808 555040 620860 555264
rect 612500 555012 620860 555040
rect 611560 554720 619660 554748
rect 611560 554496 611616 554720
rect 612160 554496 618664 554720
rect 619608 554496 619660 554720
rect 611560 554468 619660 554496
rect 4573 552000 22973 552028
rect 4573 551776 4612 552000
rect 5556 551776 22380 552000
rect 22924 551776 22973 552000
rect 4573 551748 22973 551776
rect 5760 551456 22020 551484
rect 5760 551232 5812 551456
rect 6756 551232 21420 551456
rect 21964 551232 22020 551456
rect 5760 551204 22020 551232
rect 6960 550912 16260 550940
rect 6960 550688 7012 550912
rect 7956 550688 15660 550912
rect 16204 550688 16260 550912
rect 6960 550660 16260 550688
rect 8160 550368 17220 550396
rect 8160 550144 8212 550368
rect 9156 550144 16620 550368
rect 17164 550144 17220 550368
rect 8160 550116 17220 550144
rect 9360 549824 18170 549852
rect 9360 549600 9412 549824
rect 10356 549600 17580 549824
rect 18124 549600 18170 549824
rect 9360 549572 18170 549600
rect 10560 549280 19160 549308
rect 10560 549056 10612 549280
rect 11556 549056 18540 549280
rect 19084 549056 19160 549280
rect 10560 549028 19160 549056
rect 11760 548736 20120 548764
rect 11760 548512 11812 548736
rect 12756 548512 19500 548736
rect 20044 548512 20120 548736
rect 11760 548484 20120 548512
rect 12960 548192 21060 548220
rect 12960 547968 13012 548192
rect 13956 547968 20460 548192
rect 21004 547968 21060 548192
rect 12960 547940 21060 547968
rect 614450 543296 623260 543324
rect 614450 543072 614496 543296
rect 615040 543072 622264 543296
rect 623208 543072 623260 543296
rect 614450 543044 623260 543072
rect 613460 542752 622060 542780
rect 613460 542528 613536 542752
rect 614080 542528 621064 542752
rect 622008 542528 622060 542752
rect 613460 542500 622060 542528
rect 612500 542208 620860 542236
rect 612500 541984 612576 542208
rect 613120 541984 619864 542208
rect 620808 541984 620860 542208
rect 612500 541956 620860 541984
rect 611560 541664 619660 541692
rect 611560 541440 611616 541664
rect 612160 541440 618664 541664
rect 619608 541440 619660 541664
rect 611560 541412 619660 541440
rect 4573 538944 22973 538972
rect 4573 538720 4612 538944
rect 5556 538720 22380 538944
rect 22924 538720 22973 538944
rect 4573 538692 22973 538720
rect 5760 538400 22020 538428
rect 5760 538176 5812 538400
rect 6756 538176 21420 538400
rect 21964 538176 22020 538400
rect 5760 538148 22020 538176
rect 6960 537856 16260 537884
rect 6960 537632 7012 537856
rect 7956 537632 15660 537856
rect 16204 537632 16260 537856
rect 6960 537604 16260 537632
rect 8160 537312 17220 537340
rect 8160 537088 8212 537312
rect 9156 537088 16620 537312
rect 17164 537088 17220 537312
rect 8160 537060 17220 537088
rect 9360 536768 18170 536796
rect 9360 536544 9412 536768
rect 10356 536544 17580 536768
rect 18124 536544 18170 536768
rect 9360 536516 18170 536544
rect 10560 536224 19160 536252
rect 10560 536000 10612 536224
rect 11556 536000 18540 536224
rect 19084 536000 19160 536224
rect 10560 535972 19160 536000
rect 11760 535680 20120 535708
rect 11760 535456 11812 535680
rect 12756 535456 19500 535680
rect 20044 535456 20120 535680
rect 11760 535428 20120 535456
rect 12960 535136 21060 535164
rect 12960 534912 13012 535136
rect 13956 534912 20460 535136
rect 21004 534912 21060 535136
rect 12960 534884 21060 534912
rect 609647 530784 628047 530812
rect 609647 530560 609696 530784
rect 610240 530560 627064 530784
rect 628008 530560 628047 530784
rect 609647 530532 628047 530560
rect 610600 530240 626860 530268
rect 610600 530016 610656 530240
rect 611200 530016 625864 530240
rect 626808 530016 626860 530240
rect 610600 529988 626860 530016
rect 616360 529696 625660 529724
rect 616360 529472 616416 529696
rect 616960 529472 624664 529696
rect 625608 529472 625660 529696
rect 616360 529444 625660 529472
rect 615400 529152 624460 529180
rect 615400 528928 615456 529152
rect 616000 528928 623464 529152
rect 624408 528928 624460 529152
rect 615400 528900 624460 528928
rect 614450 528608 623260 528636
rect 614450 528384 614496 528608
rect 615040 528384 622264 528608
rect 623208 528384 623260 528608
rect 614450 528356 623260 528384
rect 613460 528064 622060 528092
rect 613460 527840 613536 528064
rect 614080 527840 621064 528064
rect 622008 527840 622060 528064
rect 613460 527812 622060 527840
rect 612500 527520 620860 527548
rect 612500 527296 612576 527520
rect 613120 527296 619864 527520
rect 620808 527296 620860 527520
rect 612500 527268 620860 527296
rect 611560 526976 619660 527004
rect 611560 526752 611616 526976
rect 612160 526752 618664 526976
rect 619608 526752 619660 526976
rect 611560 526724 619660 526752
rect 4573 525888 22973 525916
rect 4573 525664 4612 525888
rect 5556 525664 22380 525888
rect 22924 525664 22973 525888
rect 4573 525636 22973 525664
rect 5760 525344 22020 525372
rect 5760 525120 5812 525344
rect 6756 525120 21420 525344
rect 21964 525120 22020 525344
rect 5760 525092 22020 525120
rect 6960 524800 16260 524828
rect 6960 524576 7012 524800
rect 7956 524576 15660 524800
rect 16204 524576 16260 524800
rect 6960 524548 16260 524576
rect 8160 524256 17220 524284
rect 8160 524032 8212 524256
rect 9156 524032 16620 524256
rect 17164 524032 17220 524256
rect 8160 524004 17220 524032
rect 9360 523712 18170 523740
rect 9360 523488 9412 523712
rect 10356 523488 17580 523712
rect 18124 523488 18170 523712
rect 9360 523460 18170 523488
rect 10560 523168 19160 523196
rect 10560 522944 10612 523168
rect 11556 522944 18540 523168
rect 19084 522944 19160 523168
rect 10560 522916 19160 522944
rect 11760 522624 20120 522652
rect 11760 522400 11812 522624
rect 12756 522400 19500 522624
rect 20044 522400 20120 522624
rect 11760 522372 20120 522400
rect 12960 522080 21060 522108
rect 12960 521856 13012 522080
rect 13956 521856 20460 522080
rect 21004 521856 21060 522080
rect 12960 521828 21060 521856
rect 609647 517728 628047 517756
rect 609647 517504 609696 517728
rect 610240 517504 627064 517728
rect 628008 517504 628047 517728
rect 609647 517476 628047 517504
rect 610600 517184 626860 517212
rect 610600 516960 610656 517184
rect 611200 516960 625864 517184
rect 626808 516960 626860 517184
rect 610600 516932 626860 516960
rect 616360 516640 625660 516668
rect 616360 516416 616416 516640
rect 616960 516416 624664 516640
rect 625608 516416 625660 516640
rect 616360 516388 625660 516416
rect 615400 516096 624460 516124
rect 615400 515872 615456 516096
rect 616000 515872 623464 516096
rect 624408 515872 624460 516096
rect 615400 515844 624460 515872
rect 614450 515552 623260 515580
rect 614450 515328 614496 515552
rect 615040 515328 622264 515552
rect 623208 515328 623260 515552
rect 614450 515300 623260 515328
rect 613460 515008 622060 515036
rect 613460 514784 613536 515008
rect 614080 514784 621064 515008
rect 622008 514784 622060 515008
rect 613460 514756 622060 514784
rect 612500 514464 620860 514492
rect 612500 514240 612576 514464
rect 613120 514240 619864 514464
rect 620808 514240 620860 514464
rect 612500 514212 620860 514240
rect 611560 513920 619660 513948
rect 611560 513696 611616 513920
rect 612160 513696 618664 513920
rect 619608 513696 619660 513920
rect 611560 513668 619660 513696
rect 4573 512832 22973 512860
rect 4573 512608 4612 512832
rect 5556 512608 22380 512832
rect 22924 512608 22973 512832
rect 4573 512580 22973 512608
rect 5760 512288 22020 512316
rect 5760 512064 5812 512288
rect 6756 512064 21420 512288
rect 21964 512064 22020 512288
rect 5760 512036 22020 512064
rect 6960 511744 16260 511772
rect 6960 511520 7012 511744
rect 7956 511520 15660 511744
rect 16204 511520 16260 511744
rect 6960 511492 16260 511520
rect 8160 511200 17220 511228
rect 8160 510976 8212 511200
rect 9156 510976 16620 511200
rect 17164 510976 17220 511200
rect 8160 510948 17220 510976
rect 9360 510656 18170 510684
rect 9360 510432 9412 510656
rect 10356 510432 17580 510656
rect 18124 510432 18170 510656
rect 9360 510404 18170 510432
rect 10560 510112 19160 510140
rect 10560 509888 10612 510112
rect 11556 509888 18540 510112
rect 19084 509888 19160 510112
rect 10560 509860 19160 509888
rect 11760 509568 20120 509596
rect 11760 509344 11812 509568
rect 12756 509344 19500 509568
rect 20044 509344 20120 509568
rect 11760 509316 20120 509344
rect 12960 509024 21060 509052
rect 12960 508800 13012 509024
rect 13956 508800 20460 509024
rect 21004 508800 21060 509024
rect 12960 508772 21060 508800
rect 609647 504672 628047 504700
rect 609647 504448 609696 504672
rect 610240 504448 627064 504672
rect 628008 504448 628047 504672
rect 609647 504420 628047 504448
rect 610600 504128 626860 504156
rect 610600 503904 610656 504128
rect 611200 503904 625864 504128
rect 626808 503904 626860 504128
rect 610600 503876 626860 503904
rect 616360 503584 625660 503612
rect 616360 503360 616416 503584
rect 616960 503360 624664 503584
rect 625608 503360 625660 503584
rect 616360 503332 625660 503360
rect 615400 503040 624460 503068
rect 615400 502816 615456 503040
rect 616000 502816 623464 503040
rect 624408 502816 624460 503040
rect 615400 502788 624460 502816
rect 614450 502496 623260 502524
rect 614450 502272 614496 502496
rect 615040 502272 622264 502496
rect 623208 502272 623260 502496
rect 614450 502244 623260 502272
rect 613460 501952 622060 501980
rect 613460 501728 613536 501952
rect 614080 501728 621064 501952
rect 622008 501728 622060 501952
rect 613460 501700 622060 501728
rect 612500 501408 620860 501436
rect 612500 501184 612576 501408
rect 613120 501184 619864 501408
rect 620808 501184 620860 501408
rect 612500 501156 620860 501184
rect 611560 500864 619660 500892
rect 611560 500640 611616 500864
rect 612160 500640 618664 500864
rect 619608 500640 619660 500864
rect 611560 500612 619660 500640
rect 4573 499776 22973 499804
rect 4573 499552 4612 499776
rect 5556 499552 22380 499776
rect 22924 499552 22973 499776
rect 4573 499524 22973 499552
rect 5760 499232 22020 499260
rect 5760 499008 5812 499232
rect 6756 499008 21420 499232
rect 21964 499008 22020 499232
rect 5760 498980 22020 499008
rect 6960 498688 16260 498716
rect 6960 498464 7012 498688
rect 7956 498464 15660 498688
rect 16204 498464 16260 498688
rect 6960 498436 16260 498464
rect 8160 498144 17220 498172
rect 8160 497920 8212 498144
rect 9156 497920 16620 498144
rect 17164 497920 17220 498144
rect 8160 497892 17220 497920
rect 9360 497600 18170 497628
rect 9360 497376 9412 497600
rect 10356 497376 17580 497600
rect 18124 497376 18170 497600
rect 9360 497348 18170 497376
rect 10560 497056 19160 497084
rect 10560 496832 10612 497056
rect 11556 496832 18540 497056
rect 19084 496832 19160 497056
rect 10560 496804 19160 496832
rect 11760 496512 20120 496540
rect 11760 496288 11812 496512
rect 12756 496288 19500 496512
rect 20044 496288 20120 496512
rect 11760 496260 20120 496288
rect 12960 495968 21060 495996
rect 12960 495744 13012 495968
rect 13956 495744 20460 495968
rect 21004 495744 21060 495968
rect 12960 495716 21060 495744
rect 609647 491616 628047 491644
rect 609647 491392 609696 491616
rect 610240 491392 627064 491616
rect 628008 491392 628047 491616
rect 609647 491364 628047 491392
rect 610600 491072 626860 491100
rect 610600 490848 610656 491072
rect 611200 490848 625864 491072
rect 626808 490848 626860 491072
rect 610600 490820 626860 490848
rect 616360 490528 625660 490556
rect 616360 490304 616416 490528
rect 616960 490304 624664 490528
rect 625608 490304 625660 490528
rect 616360 490276 625660 490304
rect 615400 489984 624460 490012
rect 615400 489760 615456 489984
rect 616000 489760 623464 489984
rect 624408 489760 624460 489984
rect 615400 489732 624460 489760
rect 614450 489440 623260 489468
rect 614450 489216 614496 489440
rect 615040 489216 622264 489440
rect 623208 489216 623260 489440
rect 614450 489188 623260 489216
rect 613460 488896 622060 488924
rect 613460 488672 613536 488896
rect 614080 488672 621064 488896
rect 622008 488672 622060 488896
rect 613460 488644 622060 488672
rect 612500 488352 620860 488380
rect 612500 488128 612576 488352
rect 613120 488128 619864 488352
rect 620808 488128 620860 488352
rect 612500 488100 620860 488128
rect 611560 487808 619660 487836
rect 611560 487584 611616 487808
rect 612160 487584 618664 487808
rect 619608 487584 619660 487808
rect 611560 487556 619660 487584
rect 4573 486720 22973 486748
rect 4573 486496 4612 486720
rect 5556 486496 22380 486720
rect 22924 486496 22973 486720
rect 4573 486468 22973 486496
rect 5760 486176 22020 486204
rect 5760 485952 5812 486176
rect 6756 485952 21420 486176
rect 21964 485952 22020 486176
rect 5760 485924 22020 485952
rect 6960 485632 16260 485660
rect 6960 485408 7012 485632
rect 7956 485408 15660 485632
rect 16204 485408 16260 485632
rect 6960 485380 16260 485408
rect 8160 485088 17220 485116
rect 8160 484864 8212 485088
rect 9156 484864 16620 485088
rect 17164 484864 17220 485088
rect 8160 484836 17220 484864
rect 9360 484544 18170 484572
rect 9360 484320 9412 484544
rect 10356 484320 17580 484544
rect 18124 484320 18170 484544
rect 9360 484292 18170 484320
rect 10560 484000 19160 484028
rect 10560 483776 10612 484000
rect 11556 483776 18540 484000
rect 19084 483776 19160 484000
rect 10560 483748 19160 483776
rect 11760 483456 20120 483484
rect 11760 483232 11812 483456
rect 12756 483232 19500 483456
rect 20044 483232 20120 483456
rect 11760 483204 20120 483232
rect 12960 482912 21060 482940
rect 12960 482688 13012 482912
rect 13956 482688 20460 482912
rect 21004 482688 21060 482912
rect 12960 482660 21060 482688
rect 609647 476928 628047 476956
rect 609647 476704 609696 476928
rect 610240 476704 627064 476928
rect 628008 476704 628047 476928
rect 609647 476676 628047 476704
rect 631206 476519 635604 476601
rect 610600 476384 626860 476412
rect 610600 476160 610656 476384
rect 611200 476160 625864 476384
rect 626808 476160 626860 476384
rect 610600 476132 626860 476160
rect 616360 475840 625660 475868
rect 616360 475616 616416 475840
rect 616960 475616 624664 475840
rect 625608 475616 625660 475840
rect 616360 475588 625660 475616
rect 615400 475296 624460 475324
rect 615400 475072 615456 475296
rect 616000 475072 623464 475296
rect 624408 475072 624460 475296
rect 615400 475044 624460 475072
rect 614450 474752 623260 474780
rect 614450 474528 614496 474752
rect 615040 474528 622264 474752
rect 623208 474528 623260 474752
rect 614450 474500 623260 474528
rect 613460 474208 622060 474236
rect 613460 473984 613536 474208
rect 614080 473984 621064 474208
rect 622008 473984 622060 474208
rect 613460 473956 622060 473984
rect 612500 473664 620860 473692
rect 612500 473440 612576 473664
rect 613120 473440 619864 473664
rect 620808 473440 620860 473664
rect 612500 473412 620860 473440
rect 611560 473120 619660 473148
rect 611560 472896 611616 473120
rect 612160 472896 618664 473120
rect 619608 472896 619660 473120
rect 611560 472868 619660 472896
rect 631206 471895 631301 476519
rect 634165 471895 635604 476519
rect 631206 471812 635604 471895
rect 4573 471488 22973 471516
rect 4573 471264 4612 471488
rect 5556 471264 22380 471488
rect 22924 471264 22973 471488
rect 4573 471236 22973 471264
rect 5760 470944 22020 470972
rect 5760 470720 5812 470944
rect 6756 470720 21420 470944
rect 21964 470720 22020 470944
rect 5760 470692 22020 470720
rect 6960 470400 16260 470428
rect 6960 470176 7012 470400
rect 7956 470176 15660 470400
rect 16204 470176 16260 470400
rect 6960 470148 16260 470176
rect 8160 469856 17220 469884
rect 8160 469632 8212 469856
rect 9156 469632 16620 469856
rect 17164 469632 17220 469856
rect 8160 469604 17220 469632
rect 9360 469312 18170 469340
rect 9360 469088 9412 469312
rect 10356 469088 17580 469312
rect 18124 469088 18170 469312
rect 9360 469060 18170 469088
rect 10560 468768 19160 468796
rect 10560 468544 10612 468768
rect 11556 468544 18540 468768
rect 19084 468544 19160 468768
rect 10560 468516 19160 468544
rect 11760 468224 20120 468252
rect 11760 468000 11812 468224
rect 12756 468000 19500 468224
rect 20044 468000 20120 468224
rect 11760 467972 20120 468000
rect 12960 467680 21060 467708
rect 12960 467456 13012 467680
rect 13956 467456 20460 467680
rect 21004 467456 21060 467680
rect 12960 467428 21060 467456
rect 631206 466536 635604 466618
rect 609647 463872 628047 463900
rect 609647 463648 609696 463872
rect 610240 463648 627064 463872
rect 628008 463648 628047 463872
rect 609647 463620 628047 463648
rect 610600 463328 626860 463356
rect 610600 463104 610656 463328
rect 611200 463104 625864 463328
rect 626808 463104 626860 463328
rect 610600 463076 626860 463104
rect 616360 462784 625660 462812
rect 616360 462560 616416 462784
rect 616960 462560 624664 462784
rect 625608 462560 625660 462784
rect 616360 462532 625660 462560
rect 615400 462240 624460 462268
rect 615400 462016 615456 462240
rect 616000 462016 623464 462240
rect 624408 462016 624460 462240
rect 615400 461988 624460 462016
rect 631206 461912 631301 466536
rect 634165 461912 635604 466536
rect 631206 461829 635604 461912
rect 614450 461696 623260 461724
rect 614450 461472 614496 461696
rect 615040 461472 622264 461696
rect 623208 461472 623260 461696
rect 614450 461444 623260 461472
rect 613460 461152 622060 461180
rect 613460 460928 613536 461152
rect 614080 460928 621064 461152
rect 622008 460928 622060 461152
rect 613460 460900 622060 460928
rect 4573 460608 22973 460636
rect 4573 460384 4612 460608
rect 5556 460384 22380 460608
rect 22924 460384 22973 460608
rect 4573 460356 22973 460384
rect 612500 460608 620860 460636
rect 612500 460384 612576 460608
rect 613120 460384 619864 460608
rect 620808 460384 620860 460608
rect 612500 460356 620860 460384
rect 5760 460064 22020 460092
rect 5760 459840 5812 460064
rect 6756 459840 21420 460064
rect 21964 459840 22020 460064
rect 5760 459812 22020 459840
rect 611560 460064 619660 460092
rect 611560 459840 611616 460064
rect 612160 459840 618664 460064
rect 619608 459840 619660 460064
rect 611560 459812 619660 459840
rect 6960 459520 16260 459548
rect 6960 459296 7012 459520
rect 7956 459296 15660 459520
rect 16204 459296 16260 459520
rect 6960 459268 16260 459296
rect 8160 458976 17220 459004
rect 8160 458752 8212 458976
rect 9156 458752 16620 458976
rect 17164 458752 17220 458976
rect 8160 458724 17220 458752
rect 9360 458432 18170 458460
rect 9360 458208 9412 458432
rect 10356 458208 17580 458432
rect 18124 458208 18170 458432
rect 9360 458180 18170 458208
rect 10560 457888 19160 457916
rect 10560 457664 10612 457888
rect 11556 457664 18540 457888
rect 19084 457664 19160 457888
rect 10560 457636 19160 457664
rect 11760 457344 20120 457372
rect 11760 457120 11812 457344
rect 12756 457120 19500 457344
rect 20044 457120 20120 457344
rect 11760 457092 20120 457120
rect 12960 456800 21060 456828
rect 12960 456576 13012 456800
rect 13956 456576 20460 456800
rect 21004 456576 21060 456800
rect 12960 456548 21060 456576
rect -3216 455676 1182 455758
rect -3216 451052 -1777 455676
rect 1087 451052 1182 455676
rect -3216 450969 1182 451052
rect 609647 450816 628047 450844
rect 609647 450592 609696 450816
rect 610240 450592 627064 450816
rect 628008 450592 628047 450816
rect 609647 450564 628047 450592
rect 610600 450272 626860 450300
rect 610600 450048 610656 450272
rect 611200 450048 625864 450272
rect 626808 450048 626860 450272
rect 610600 450020 626860 450048
rect 616360 449728 625660 449756
rect 616360 449504 616416 449728
rect 616960 449504 624664 449728
rect 625608 449504 625660 449728
rect 616360 449476 625660 449504
rect 615400 449184 624460 449212
rect 615400 448960 615456 449184
rect 616000 448960 623464 449184
rect 624408 448960 624460 449184
rect 615400 448932 624460 448960
rect 614450 448640 623260 448668
rect 614450 448416 614496 448640
rect 615040 448416 622264 448640
rect 623208 448416 623260 448640
rect 614450 448388 623260 448416
rect 613460 448096 622060 448124
rect 613460 447872 613536 448096
rect 614080 447872 621064 448096
rect 622008 447872 622060 448096
rect 613460 447844 622060 447872
rect 4573 447552 22973 447580
rect 4573 447328 4612 447552
rect 5556 447328 22380 447552
rect 22924 447328 22973 447552
rect 4573 447300 22973 447328
rect 612500 447552 620860 447580
rect 612500 447328 612576 447552
rect 613120 447328 619864 447552
rect 620808 447328 620860 447552
rect 612500 447300 620860 447328
rect 5760 447008 22020 447036
rect 5760 446784 5812 447008
rect 6756 446784 21420 447008
rect 21964 446784 22020 447008
rect 5760 446756 22020 446784
rect 611560 447008 619660 447036
rect 611560 446784 611616 447008
rect 612160 446784 618664 447008
rect 619608 446784 619660 447008
rect 611560 446756 619660 446784
rect 6960 446464 16260 446492
rect 6960 446240 7012 446464
rect 7956 446240 15660 446464
rect 16204 446240 16260 446464
rect 6960 446212 16260 446240
rect 8160 445920 17220 445948
rect -3216 445697 1182 445779
rect -3216 441073 -1777 445697
rect 1087 441073 1182 445697
rect 8160 445696 8212 445920
rect 9156 445696 16620 445920
rect 17164 445696 17220 445920
rect 8160 445668 17220 445696
rect 9360 445376 18170 445404
rect 9360 445152 9412 445376
rect 10356 445152 17580 445376
rect 18124 445152 18170 445376
rect 9360 445124 18170 445152
rect 10560 444832 19160 444860
rect 10560 444608 10612 444832
rect 11556 444608 18540 444832
rect 19084 444608 19160 444832
rect 10560 444580 19160 444608
rect 11760 444288 20120 444316
rect 11760 444064 11812 444288
rect 12756 444064 19500 444288
rect 20044 444064 20120 444288
rect 11760 444036 20120 444064
rect 12960 443744 21060 443772
rect 12960 443520 13012 443744
rect 13956 443520 20460 443744
rect 21004 443520 21060 443744
rect 12960 443492 21060 443520
rect -3216 440990 1182 441073
rect 609647 437760 628047 437788
rect 609647 437536 609696 437760
rect 610240 437536 627064 437760
rect 628008 437536 628047 437760
rect 609647 437508 628047 437536
rect 610600 437216 626860 437244
rect 610600 436992 610656 437216
rect 611200 436992 625864 437216
rect 626808 436992 626860 437216
rect 610600 436964 626860 436992
rect 616360 436672 625660 436700
rect 616360 436448 616416 436672
rect 616960 436448 624664 436672
rect 625608 436448 625660 436672
rect 616360 436420 625660 436448
rect 615400 436128 624460 436156
rect 615400 435904 615456 436128
rect 616000 435904 623464 436128
rect 624408 435904 624460 436128
rect 615400 435876 624460 435904
rect 614450 435584 623260 435612
rect 614450 435360 614496 435584
rect 615040 435360 622264 435584
rect 623208 435360 623260 435584
rect 614450 435332 623260 435360
rect 613460 435040 622060 435068
rect 613460 434816 613536 435040
rect 614080 434816 621064 435040
rect 622008 434816 622060 435040
rect 613460 434788 622060 434816
rect 4573 434496 22973 434524
rect 4573 434272 4612 434496
rect 5556 434272 22380 434496
rect 22924 434272 22973 434496
rect 4573 434244 22973 434272
rect 612500 434496 620860 434524
rect 612500 434272 612576 434496
rect 613120 434272 619864 434496
rect 620808 434272 620860 434496
rect 612500 434244 620860 434272
rect 5760 433952 22020 433980
rect 5760 433728 5812 433952
rect 6756 433728 21420 433952
rect 21964 433728 22020 433952
rect 5760 433700 22020 433728
rect 611560 433952 619660 433980
rect 611560 433728 611616 433952
rect 612160 433728 618664 433952
rect 619608 433728 619660 433952
rect 611560 433700 619660 433728
rect 6960 433408 16260 433436
rect 6960 433184 7012 433408
rect 7956 433184 15660 433408
rect 16204 433184 16260 433408
rect 6960 433156 16260 433184
rect 8160 432864 17220 432892
rect 8160 432640 8212 432864
rect 9156 432640 16620 432864
rect 17164 432640 17220 432864
rect 8160 432612 17220 432640
rect 631206 432518 635604 432600
rect 9360 432320 18170 432348
rect 9360 432096 9412 432320
rect 10356 432096 17580 432320
rect 18124 432096 18170 432320
rect 9360 432068 18170 432096
rect 10560 431776 19160 431804
rect 10560 431552 10612 431776
rect 11556 431552 18540 431776
rect 19084 431552 19160 431776
rect 10560 431524 19160 431552
rect 11760 431232 20120 431260
rect 11760 431008 11812 431232
rect 12756 431008 19500 431232
rect 20044 431008 20120 431232
rect 11760 430980 20120 431008
rect 12960 430688 21060 430716
rect 12960 430464 13012 430688
rect 13956 430464 20460 430688
rect 21004 430464 21060 430688
rect 12960 430436 21060 430464
rect 631206 427894 631301 432518
rect 634165 427894 635604 432518
rect 631206 427811 635604 427894
rect 631206 427408 635204 427490
rect 609647 424704 628047 424732
rect 609647 424480 609696 424704
rect 610240 424480 627064 424704
rect 628008 424480 628047 424704
rect 609647 424452 628047 424480
rect 610600 424160 626860 424188
rect 610600 423936 610656 424160
rect 611200 423936 625864 424160
rect 626808 423936 626860 424160
rect 610600 423908 626860 423936
rect 616360 423616 625660 423644
rect 616360 423392 616416 423616
rect 616960 423392 624664 423616
rect 625608 423392 625660 423616
rect 616360 423364 625660 423392
rect 615400 423072 624460 423100
rect 615400 422848 615456 423072
rect 616000 422848 623464 423072
rect 624408 422848 624460 423072
rect 631206 422944 631301 427408
rect 634165 422944 635204 427408
rect 631206 422869 635204 422944
rect 615400 422820 624460 422848
rect 614450 422528 623260 422556
rect 614450 422304 614496 422528
rect 615040 422304 622264 422528
rect 623208 422304 623260 422528
rect 614450 422276 623260 422304
rect 631206 422467 635604 422549
rect 613460 421984 622060 422012
rect 613460 421760 613536 421984
rect 614080 421760 621064 421984
rect 622008 421760 622060 421984
rect 613460 421732 622060 421760
rect 4573 421440 22973 421468
rect 4573 421216 4612 421440
rect 5556 421216 22380 421440
rect 22924 421216 22973 421440
rect 4573 421188 22973 421216
rect 612500 421440 620860 421468
rect 612500 421216 612576 421440
rect 613120 421216 619864 421440
rect 620808 421216 620860 421440
rect 612500 421188 620860 421216
rect 5760 420896 22020 420924
rect 5760 420672 5812 420896
rect 6756 420672 21420 420896
rect 21964 420672 22020 420896
rect 5760 420644 22020 420672
rect 611560 420896 619660 420924
rect 611560 420672 611616 420896
rect 612160 420672 618664 420896
rect 619608 420672 619660 420896
rect 611560 420644 619660 420672
rect 6960 420352 16260 420380
rect 6960 420128 7012 420352
rect 7956 420128 15660 420352
rect 16204 420128 16260 420352
rect 6960 420100 16260 420128
rect 8160 419808 17220 419836
rect 8160 419584 8212 419808
rect 9156 419584 16620 419808
rect 17164 419584 17220 419808
rect 8160 419556 17220 419584
rect 9360 419264 18170 419292
rect 9360 419040 9412 419264
rect 10356 419040 17580 419264
rect 18124 419040 18170 419264
rect 9360 419012 18170 419040
rect 10560 418720 19160 418748
rect 10560 418496 10612 418720
rect 11556 418496 18540 418720
rect 19084 418496 19160 418720
rect 10560 418468 19160 418496
rect 11760 418176 20120 418204
rect 11760 417952 11812 418176
rect 12756 417952 19500 418176
rect 20044 417952 20120 418176
rect 11760 417924 20120 417952
rect 631206 417843 631301 422467
rect 634165 417843 635604 422467
rect 631206 417760 635604 417843
rect 12960 417632 21060 417660
rect 12960 417408 13012 417632
rect 13956 417408 20460 417632
rect 21004 417408 21060 417632
rect 12960 417380 21060 417408
rect -3216 413558 1182 413640
rect -3216 408934 -1777 413558
rect 1087 408934 1182 413558
rect 609647 411648 628047 411676
rect 609647 411424 609696 411648
rect 610240 411424 627064 411648
rect 628008 411424 628047 411648
rect 609647 411396 628047 411424
rect 610600 411104 626860 411132
rect 610600 410880 610656 411104
rect 611200 410880 625864 411104
rect 626808 410880 626860 411104
rect 610600 410852 626860 410880
rect 616360 410560 625660 410588
rect 616360 410336 616416 410560
rect 616960 410336 624664 410560
rect 625608 410336 625660 410560
rect 616360 410308 625660 410336
rect 615400 410016 624460 410044
rect 615400 409792 615456 410016
rect 616000 409792 623464 410016
rect 624408 409792 624460 410016
rect 615400 409764 624460 409792
rect 614450 409472 623260 409500
rect 614450 409248 614496 409472
rect 615040 409248 622264 409472
rect 623208 409248 623260 409472
rect 614450 409220 623260 409248
rect -3216 408851 1182 408934
rect 613460 408928 622060 408956
rect 613460 408704 613536 408928
rect 614080 408704 621064 408928
rect 622008 408704 622060 408928
rect 613460 408676 622060 408704
rect -2216 408448 1182 408530
rect -2216 403984 -1777 408448
rect 1087 403984 1182 408448
rect 4573 408384 22973 408412
rect 4573 408160 4612 408384
rect 5556 408160 22380 408384
rect 22924 408160 22973 408384
rect 4573 408132 22973 408160
rect 612500 408384 620860 408412
rect 612500 408160 612576 408384
rect 613120 408160 619864 408384
rect 620808 408160 620860 408384
rect 612500 408132 620860 408160
rect 5760 407840 22020 407868
rect 5760 407616 5812 407840
rect 6756 407616 21420 407840
rect 21964 407616 22020 407840
rect 5760 407588 22020 407616
rect 611560 407840 619660 407868
rect 611560 407616 611616 407840
rect 612160 407616 618664 407840
rect 619608 407616 619660 407840
rect 611560 407588 619660 407616
rect 6960 407296 16260 407324
rect 6960 407072 7012 407296
rect 7956 407072 15660 407296
rect 16204 407072 16260 407296
rect 6960 407044 16260 407072
rect 8160 406752 17220 406780
rect 8160 406528 8212 406752
rect 9156 406528 16620 406752
rect 17164 406528 17220 406752
rect 8160 406500 17220 406528
rect 9360 406208 18170 406236
rect 9360 405984 9412 406208
rect 10356 405984 17580 406208
rect 18124 405984 18170 406208
rect 9360 405956 18170 405984
rect 10560 405664 19160 405692
rect 10560 405440 10612 405664
rect 11556 405440 18540 405664
rect 19084 405440 19160 405664
rect 10560 405412 19160 405440
rect 11760 405120 20120 405148
rect 11760 404896 11812 405120
rect 12756 404896 19500 405120
rect 20044 404896 20120 405120
rect 11760 404868 20120 404896
rect 12960 404576 21060 404604
rect 12960 404352 13012 404576
rect 13956 404352 20460 404576
rect 21004 404352 21060 404576
rect 12960 404324 21060 404352
rect -2216 403920 1182 403984
rect -3216 403518 1182 403600
rect -3216 398894 -1777 403518
rect 1087 398894 1182 403518
rect -3216 398811 1182 398894
rect 609647 398592 628047 398620
rect 609647 398368 609696 398592
rect 610240 398368 627064 398592
rect 628008 398368 628047 398592
rect 609647 398340 628047 398368
rect 610600 398048 626860 398076
rect 610600 397824 610656 398048
rect 611200 397824 625864 398048
rect 626808 397824 626860 398048
rect 610600 397796 626860 397824
rect 616360 397504 625660 397532
rect 616360 397280 616416 397504
rect 616960 397280 624664 397504
rect 625608 397280 625660 397504
rect 616360 397252 625660 397280
rect 615400 396960 624460 396988
rect 615400 396736 615456 396960
rect 616000 396736 623464 396960
rect 624408 396736 624460 396960
rect 615400 396708 624460 396736
rect 614450 396416 623260 396444
rect 614450 396192 614496 396416
rect 615040 396192 622264 396416
rect 623208 396192 623260 396416
rect 614450 396164 623260 396192
rect 613460 395872 622060 395900
rect 613460 395648 613536 395872
rect 614080 395648 621064 395872
rect 622008 395648 622060 395872
rect 613460 395620 622060 395648
rect 4573 395328 22973 395356
rect 4573 395104 4612 395328
rect 5556 395104 22380 395328
rect 22924 395104 22973 395328
rect 4573 395076 22973 395104
rect 612500 395328 620860 395356
rect 612500 395104 612576 395328
rect 613120 395104 619864 395328
rect 620808 395104 620860 395328
rect 612500 395076 620860 395104
rect 5760 394784 22020 394812
rect 5760 394560 5812 394784
rect 6756 394560 21420 394784
rect 21964 394560 22020 394784
rect 5760 394532 22020 394560
rect 611560 394784 619660 394812
rect 611560 394560 611616 394784
rect 612160 394560 618664 394784
rect 619608 394560 619660 394784
rect 611560 394532 619660 394560
rect 6960 394240 16260 394268
rect 6960 394016 7012 394240
rect 7956 394016 15660 394240
rect 16204 394016 16260 394240
rect 6960 393988 16260 394016
rect 8160 393696 17220 393724
rect 8160 393472 8212 393696
rect 9156 393472 16620 393696
rect 17164 393472 17220 393696
rect 8160 393444 17220 393472
rect 9360 393152 18170 393180
rect 9360 392928 9412 393152
rect 10356 392928 17580 393152
rect 18124 392928 18170 393152
rect 9360 392900 18170 392928
rect 10560 392608 19160 392636
rect 10560 392384 10612 392608
rect 11556 392384 18540 392608
rect 19084 392384 19160 392608
rect 10560 392356 19160 392384
rect 11760 392064 20120 392092
rect 11760 391840 11812 392064
rect 12756 391840 19500 392064
rect 20044 391840 20120 392064
rect 11760 391812 20120 391840
rect 12960 391520 21060 391548
rect 12960 391296 13012 391520
rect 13956 391296 20460 391520
rect 21004 391296 21060 391520
rect 12960 391268 21060 391296
rect 631206 388327 635604 388409
rect 609647 385536 628047 385564
rect 609647 385312 609696 385536
rect 610240 385312 627064 385536
rect 628008 385312 628047 385536
rect 609647 385284 628047 385312
rect 610600 384992 626860 385020
rect 610600 384768 610656 384992
rect 611200 384768 625864 384992
rect 626808 384768 626860 384992
rect 610600 384740 626860 384768
rect 616360 384448 625660 384476
rect 616360 384224 616416 384448
rect 616960 384224 624664 384448
rect 625608 384224 625660 384448
rect 616360 384196 625660 384224
rect 615400 383904 624460 383932
rect 615400 383680 615456 383904
rect 616000 383680 623464 383904
rect 624408 383680 624460 383904
rect 615400 383652 624460 383680
rect 631206 383703 631301 388327
rect 634165 383703 635604 388327
rect 631206 383620 635604 383703
rect 614450 383360 623260 383388
rect 614450 383136 614496 383360
rect 615040 383136 622264 383360
rect 623208 383136 623260 383360
rect 614450 383108 623260 383136
rect 613460 382816 622060 382844
rect 613460 382592 613536 382816
rect 614080 382592 621064 382816
rect 622008 382592 622060 382816
rect 613460 382564 622060 382592
rect 4573 382272 22973 382300
rect 4573 382048 4612 382272
rect 5556 382048 22380 382272
rect 22924 382048 22973 382272
rect 4573 382020 22973 382048
rect 612500 382272 620860 382300
rect 612500 382048 612576 382272
rect 613120 382048 619864 382272
rect 620808 382048 620860 382272
rect 612500 382020 620860 382048
rect 5760 381728 22020 381756
rect 5760 381504 5812 381728
rect 6756 381504 21420 381728
rect 21964 381504 22020 381728
rect 5760 381476 22020 381504
rect 611560 381728 619660 381756
rect 611560 381504 611616 381728
rect 612160 381504 618664 381728
rect 619608 381504 619660 381728
rect 611560 381476 619660 381504
rect 6960 381184 16260 381212
rect 6960 380960 7012 381184
rect 7956 380960 15660 381184
rect 16204 380960 16260 381184
rect 6960 380932 16260 380960
rect 8160 380640 17220 380668
rect 8160 380416 8212 380640
rect 9156 380416 16620 380640
rect 17164 380416 17220 380640
rect 8160 380388 17220 380416
rect 9360 380096 18170 380124
rect 9360 379872 9412 380096
rect 10356 379872 17580 380096
rect 18124 379872 18170 380096
rect 9360 379844 18170 379872
rect 10560 379552 19160 379580
rect 10560 379328 10612 379552
rect 11556 379328 18540 379552
rect 19084 379328 19160 379552
rect 10560 379300 19160 379328
rect 11760 379008 20120 379036
rect 11760 378784 11812 379008
rect 12756 378784 19500 379008
rect 20044 378784 20120 379008
rect 11760 378756 20120 378784
rect 12960 378464 21060 378492
rect 12960 378240 13012 378464
rect 13956 378240 20460 378464
rect 21004 378240 21060 378464
rect 12960 378212 21060 378240
rect 631206 378344 635604 378426
rect 631206 373720 631301 378344
rect 634165 373720 635604 378344
rect 631206 373637 635604 373720
rect 4573 369216 22973 369244
rect 4573 368992 4612 369216
rect 5556 368992 22380 369216
rect 22924 368992 22973 369216
rect 4573 368964 22973 368992
rect 609647 369216 628047 369244
rect 609647 368992 609696 369216
rect 610240 368992 627064 369216
rect 628008 368992 628047 369216
rect 609647 368964 628047 368992
rect 5760 368672 22020 368700
rect 5760 368448 5812 368672
rect 6756 368448 21420 368672
rect 21964 368448 22020 368672
rect 5760 368420 22020 368448
rect 610600 368672 626860 368700
rect 610600 368448 610656 368672
rect 611200 368448 625864 368672
rect 626808 368448 626860 368672
rect 610600 368420 626860 368448
rect 6960 368128 16260 368156
rect 6960 367904 7012 368128
rect 7956 367904 15660 368128
rect 16204 367904 16260 368128
rect 6960 367876 16260 367904
rect 616360 368128 625660 368156
rect 616360 367904 616416 368128
rect 616960 367904 624664 368128
rect 625608 367904 625660 368128
rect 616360 367876 625660 367904
rect 8160 367584 17220 367612
rect 8160 367360 8212 367584
rect 9156 367360 16620 367584
rect 17164 367360 17220 367584
rect 8160 367332 17220 367360
rect 615400 367584 624460 367612
rect 615400 367360 615456 367584
rect 616000 367360 623464 367584
rect 624408 367360 624460 367584
rect 615400 367332 624460 367360
rect 9360 367040 18170 367068
rect 9360 366816 9412 367040
rect 10356 366816 17580 367040
rect 18124 366816 18170 367040
rect 9360 366788 18170 366816
rect 614450 367040 623260 367068
rect 614450 366816 614496 367040
rect 615040 366816 622264 367040
rect 623208 366816 623260 367040
rect 614450 366788 623260 366816
rect 10560 366496 19160 366524
rect 10560 366272 10612 366496
rect 11556 366272 18540 366496
rect 19084 366272 19160 366496
rect 10560 366244 19160 366272
rect 613460 366496 622060 366524
rect 613460 366272 613536 366496
rect 614080 366272 621064 366496
rect 622008 366272 622060 366496
rect 613460 366244 622060 366272
rect 11760 365952 20120 365980
rect 11760 365728 11812 365952
rect 12756 365728 19500 365952
rect 20044 365728 20120 365952
rect 11760 365700 20120 365728
rect 612500 365952 620860 365980
rect 612500 365728 612576 365952
rect 613120 365728 619864 365952
rect 620808 365728 620860 365952
rect 612500 365700 620860 365728
rect 12960 365408 21060 365436
rect 12960 365184 13012 365408
rect 13956 365184 20460 365408
rect 21004 365184 21060 365408
rect 12960 365156 21060 365184
rect 611560 365408 619660 365436
rect 611560 365184 611616 365408
rect 612160 365184 618664 365408
rect 619608 365184 619660 365408
rect 611560 365156 619660 365184
rect 4573 356160 22973 356188
rect 4573 355936 4612 356160
rect 5556 355936 22380 356160
rect 22924 355936 22973 356160
rect 4573 355908 22973 355936
rect 609647 356160 628047 356188
rect 609647 355936 609696 356160
rect 610240 355936 627064 356160
rect 628008 355936 628047 356160
rect 609647 355908 628047 355936
rect 5760 355616 22020 355644
rect 5760 355392 5812 355616
rect 6756 355392 21420 355616
rect 21964 355392 22020 355616
rect 5760 355364 22020 355392
rect 610600 355616 626860 355644
rect 610600 355392 610656 355616
rect 611200 355392 625864 355616
rect 626808 355392 626860 355616
rect 610600 355364 626860 355392
rect 6960 355072 16260 355100
rect 6960 354848 7012 355072
rect 7956 354848 15660 355072
rect 16204 354848 16260 355072
rect 6960 354820 16260 354848
rect 616360 355072 625660 355100
rect 616360 354848 616416 355072
rect 616960 354848 624664 355072
rect 625608 354848 625660 355072
rect 616360 354820 625660 354848
rect 8160 354528 17220 354556
rect 8160 354304 8212 354528
rect 9156 354304 16620 354528
rect 17164 354304 17220 354528
rect 8160 354276 17220 354304
rect 615400 354528 624460 354556
rect 615400 354304 615456 354528
rect 616000 354304 623464 354528
rect 624408 354304 624460 354528
rect 615400 354276 624460 354304
rect 9360 353984 18170 354012
rect 9360 353760 9412 353984
rect 10356 353760 17580 353984
rect 18124 353760 18170 353984
rect 9360 353732 18170 353760
rect 614450 353984 623260 354012
rect 614450 353760 614496 353984
rect 615040 353760 622264 353984
rect 623208 353760 623260 353984
rect 614450 353732 623260 353760
rect 10560 353440 19160 353468
rect 10560 353216 10612 353440
rect 11556 353216 18540 353440
rect 19084 353216 19160 353440
rect 10560 353188 19160 353216
rect 613460 353440 622060 353468
rect 613460 353216 613536 353440
rect 614080 353216 621064 353440
rect 622008 353216 622060 353440
rect 613460 353188 622060 353216
rect 11760 352896 20120 352924
rect 11760 352672 11812 352896
rect 12756 352672 19500 352896
rect 20044 352672 20120 352896
rect 11760 352644 20120 352672
rect 612500 352896 620860 352924
rect 612500 352672 612576 352896
rect 613120 352672 619864 352896
rect 620808 352672 620860 352896
rect 612500 352644 620860 352672
rect 12960 352352 21060 352380
rect 12960 352128 13012 352352
rect 13956 352128 20460 352352
rect 21004 352128 21060 352352
rect 12960 352100 21060 352128
rect 611560 352352 619660 352380
rect 611560 352128 611616 352352
rect 612160 352128 618664 352352
rect 619608 352128 619660 352352
rect 611560 352100 619660 352128
rect 609647 343104 628047 343132
rect 609647 342880 609696 343104
rect 610240 342880 627064 343104
rect 628008 342880 628047 343104
rect 609647 342852 628047 342880
rect 610600 342560 626860 342588
rect 610600 342336 610656 342560
rect 611200 342336 625864 342560
rect 626808 342336 626860 342560
rect 610600 342308 626860 342336
rect 616360 342016 625660 342044
rect 616360 341792 616416 342016
rect 616960 341792 624664 342016
rect 625608 341792 625660 342016
rect 616360 341764 625660 341792
rect 615400 341472 624460 341500
rect 615400 341248 615456 341472
rect 616000 341248 623464 341472
rect 624408 341248 624460 341472
rect 615400 341220 624460 341248
rect 4573 340928 22973 340956
rect 4573 340704 4612 340928
rect 5556 340704 22380 340928
rect 22924 340704 22973 340928
rect 4573 340676 22973 340704
rect 614450 340928 623260 340956
rect 614450 340704 614496 340928
rect 615040 340704 622264 340928
rect 623208 340704 623260 340928
rect 614450 340676 623260 340704
rect 5760 340384 22020 340412
rect 5760 340160 5812 340384
rect 6756 340160 21420 340384
rect 21964 340160 22020 340384
rect 5760 340132 22020 340160
rect 613460 340384 622060 340412
rect 613460 340160 613536 340384
rect 614080 340160 621064 340384
rect 622008 340160 622060 340384
rect 613460 340132 622060 340160
rect 6960 339840 16260 339868
rect 6960 339616 7012 339840
rect 7956 339616 15660 339840
rect 16204 339616 16260 339840
rect 6960 339588 16260 339616
rect 612500 339840 620860 339868
rect 612500 339616 612576 339840
rect 613120 339616 619864 339840
rect 620808 339616 620860 339840
rect 612500 339588 620860 339616
rect 8160 339296 17220 339324
rect 8160 339072 8212 339296
rect 9156 339072 16620 339296
rect 17164 339072 17220 339296
rect 8160 339044 17220 339072
rect 611560 339296 619660 339324
rect 611560 339072 611616 339296
rect 612160 339072 618664 339296
rect 619608 339072 619660 339296
rect 611560 339044 619660 339072
rect 9360 338752 18170 338780
rect 9360 338528 9412 338752
rect 10356 338528 17580 338752
rect 18124 338528 18170 338752
rect 9360 338500 18170 338528
rect 10560 338208 19160 338236
rect 10560 337984 10612 338208
rect 11556 337984 18540 338208
rect 19084 337984 19160 338208
rect 10560 337956 19160 337984
rect 11760 337664 20120 337692
rect 11760 337440 11812 337664
rect 12756 337440 19500 337664
rect 20044 337440 20120 337664
rect 11760 337412 20120 337440
rect 12960 337120 21060 337148
rect 12960 336896 13012 337120
rect 13956 336896 20460 337120
rect 21004 336896 21060 337120
rect 12960 336868 21060 336896
rect 4573 330048 22973 330076
rect 4573 329824 4612 330048
rect 5556 329824 22380 330048
rect 22924 329824 22973 330048
rect 4573 329796 22973 329824
rect 609647 330048 628047 330076
rect 609647 329824 609696 330048
rect 610240 329824 627064 330048
rect 628008 329824 628047 330048
rect 609647 329796 628047 329824
rect 5760 329504 22020 329532
rect 5760 329280 5812 329504
rect 6756 329280 21420 329504
rect 21964 329280 22020 329504
rect 5760 329252 22020 329280
rect 610600 329504 626860 329532
rect 610600 329280 610656 329504
rect 611200 329280 625864 329504
rect 626808 329280 626860 329504
rect 610600 329252 626860 329280
rect 6960 328960 16260 328988
rect 6960 328736 7012 328960
rect 7956 328736 15660 328960
rect 16204 328736 16260 328960
rect 6960 328708 16260 328736
rect 616360 328960 625660 328988
rect 616360 328736 616416 328960
rect 616960 328736 624664 328960
rect 625608 328736 625660 328960
rect 616360 328708 625660 328736
rect 8160 328416 17220 328444
rect 8160 328192 8212 328416
rect 9156 328192 16620 328416
rect 17164 328192 17220 328416
rect 8160 328164 17220 328192
rect 615400 328416 624460 328444
rect 615400 328192 615456 328416
rect 616000 328192 623464 328416
rect 624408 328192 624460 328416
rect 615400 328164 624460 328192
rect 9360 327872 18170 327900
rect 9360 327648 9412 327872
rect 10356 327648 17580 327872
rect 18124 327648 18170 327872
rect 9360 327620 18170 327648
rect 614450 327872 623260 327900
rect 614450 327648 614496 327872
rect 615040 327648 622264 327872
rect 623208 327648 623260 327872
rect 614450 327620 623260 327648
rect 10560 327328 19160 327356
rect 10560 327104 10612 327328
rect 11556 327104 18540 327328
rect 19084 327104 19160 327328
rect 10560 327076 19160 327104
rect 613460 327328 622060 327356
rect 613460 327104 613536 327328
rect 614080 327104 621064 327328
rect 622008 327104 622060 327328
rect 613460 327076 622060 327104
rect 11760 326784 20120 326812
rect 11760 326560 11812 326784
rect 12756 326560 19500 326784
rect 20044 326560 20120 326784
rect 11760 326532 20120 326560
rect 612500 326784 620860 326812
rect 612500 326560 612576 326784
rect 613120 326560 619864 326784
rect 620808 326560 620860 326784
rect 612500 326532 620860 326560
rect 12960 326240 21060 326268
rect 12960 326016 13012 326240
rect 13956 326016 20460 326240
rect 21004 326016 21060 326240
rect 12960 325988 21060 326016
rect 611560 326240 619660 326268
rect 611560 326016 611616 326240
rect 612160 326016 618664 326240
rect 619608 326016 619660 326240
rect 611560 325988 619660 326016
rect 609647 318624 628047 318652
rect 609647 318400 609696 318624
rect 610240 318400 627064 318624
rect 628008 318400 628047 318624
rect 609647 318372 628047 318400
rect 610600 318080 626860 318108
rect 610600 317856 610656 318080
rect 611200 317856 625864 318080
rect 626808 317856 626860 318080
rect 610600 317828 626860 317856
rect 616360 317536 625660 317564
rect 616360 317312 616416 317536
rect 616960 317312 624664 317536
rect 625608 317312 625660 317536
rect 616360 317284 625660 317312
rect 4573 316992 22973 317020
rect 4573 316768 4612 316992
rect 5556 316768 22380 316992
rect 22924 316768 22973 316992
rect 4573 316740 22973 316768
rect 615400 316992 624460 317020
rect 615400 316768 615456 316992
rect 616000 316768 623464 316992
rect 624408 316768 624460 316992
rect 615400 316740 624460 316768
rect 5760 316448 22020 316476
rect 5760 316224 5812 316448
rect 6756 316224 21420 316448
rect 21964 316224 22020 316448
rect 5760 316196 22020 316224
rect 614450 316448 623260 316476
rect 614450 316224 614496 316448
rect 615040 316224 622264 316448
rect 623208 316224 623260 316448
rect 614450 316196 623260 316224
rect 6960 315904 16260 315932
rect 6960 315680 7012 315904
rect 7956 315680 15660 315904
rect 16204 315680 16260 315904
rect 6960 315652 16260 315680
rect 613460 315904 622060 315932
rect 613460 315680 613536 315904
rect 614080 315680 621064 315904
rect 622008 315680 622060 315904
rect 613460 315652 622060 315680
rect 8160 315360 17220 315388
rect 8160 315136 8212 315360
rect 9156 315136 16620 315360
rect 17164 315136 17220 315360
rect 8160 315108 17220 315136
rect 612500 315360 620860 315388
rect 612500 315136 612576 315360
rect 613120 315136 619864 315360
rect 620808 315136 620860 315360
rect 612500 315108 620860 315136
rect 9360 314816 18170 314844
rect 9360 314592 9412 314816
rect 10356 314592 17580 314816
rect 18124 314592 18170 314816
rect 9360 314564 18170 314592
rect 611560 314816 619660 314844
rect 611560 314592 611616 314816
rect 612160 314592 618664 314816
rect 619608 314592 619660 314816
rect 611560 314564 619660 314592
rect 10560 314272 19160 314300
rect 10560 314048 10612 314272
rect 11556 314048 18540 314272
rect 19084 314048 19160 314272
rect 10560 314020 19160 314048
rect 11760 313728 20120 313756
rect 11760 313504 11812 313728
rect 12756 313504 19500 313728
rect 20044 313504 20120 313728
rect 11760 313476 20120 313504
rect 12960 313184 21060 313212
rect 12960 312960 13012 313184
rect 13956 312960 20460 313184
rect 21004 312960 21060 313184
rect 12960 312932 21060 312960
rect 4573 306112 22973 306140
rect 4573 305888 4612 306112
rect 5556 305888 22380 306112
rect 22924 305888 22973 306112
rect 4573 305860 22973 305888
rect 5760 305568 22020 305596
rect 5760 305344 5812 305568
rect 6756 305344 21420 305568
rect 21964 305344 22020 305568
rect 5760 305316 22020 305344
rect 6960 305024 16260 305052
rect 6960 304800 7012 305024
rect 7956 304800 15660 305024
rect 16204 304800 16260 305024
rect 6960 304772 16260 304800
rect 8160 304480 17220 304508
rect 8160 304256 8212 304480
rect 9156 304256 16620 304480
rect 17164 304256 17220 304480
rect 8160 304228 17220 304256
rect 9360 303936 18170 303964
rect 9360 303712 9412 303936
rect 10356 303712 17580 303936
rect 18124 303712 18170 303936
rect 9360 303684 18170 303712
rect 609647 303936 628047 303964
rect 609647 303712 609696 303936
rect 610240 303712 627064 303936
rect 628008 303712 628047 303936
rect 609647 303684 628047 303712
rect 10560 303392 19160 303420
rect 10560 303168 10612 303392
rect 11556 303168 18540 303392
rect 19084 303168 19160 303392
rect 10560 303140 19160 303168
rect 610600 303392 626860 303420
rect 610600 303168 610656 303392
rect 611200 303168 625864 303392
rect 626808 303168 626860 303392
rect 610600 303140 626860 303168
rect 11760 302848 20120 302876
rect 11760 302624 11812 302848
rect 12756 302624 19500 302848
rect 20044 302624 20120 302848
rect 11760 302596 20120 302624
rect 616360 302848 625660 302876
rect 616360 302624 616416 302848
rect 616960 302624 624664 302848
rect 625608 302624 625660 302848
rect 616360 302596 625660 302624
rect 12960 302304 21060 302332
rect 12960 302080 13012 302304
rect 13956 302080 20460 302304
rect 21004 302080 21060 302304
rect 12960 302052 21060 302080
rect 615400 302304 624460 302332
rect 615400 302080 615456 302304
rect 616000 302080 623464 302304
rect 624408 302080 624460 302304
rect 615400 302052 624460 302080
rect 614450 301760 623260 301788
rect 614450 301536 614496 301760
rect 615040 301536 622264 301760
rect 623208 301536 623260 301760
rect 614450 301508 623260 301536
rect 613460 301216 622060 301244
rect 613460 300992 613536 301216
rect 614080 300992 621064 301216
rect 622008 300992 622060 301216
rect 613460 300964 622060 300992
rect 612500 300672 620860 300700
rect 612500 300448 612576 300672
rect 613120 300448 619864 300672
rect 620808 300448 620860 300672
rect 612500 300420 620860 300448
rect 611560 300128 619660 300156
rect 611560 299904 611616 300128
rect 612160 299904 618664 300128
rect 619608 299904 619660 300128
rect 611560 299876 619660 299904
rect 4573 290880 22973 290908
rect 4573 290656 4612 290880
rect 5556 290656 22380 290880
rect 22924 290656 22973 290880
rect 4573 290628 22973 290656
rect 609647 290880 628047 290908
rect 609647 290656 609696 290880
rect 610240 290656 627064 290880
rect 628008 290656 628047 290880
rect 609647 290628 628047 290656
rect 5760 290336 22020 290364
rect 5760 290112 5812 290336
rect 6756 290112 21420 290336
rect 21964 290112 22020 290336
rect 5760 290084 22020 290112
rect 610600 290336 626860 290364
rect 610600 290112 610656 290336
rect 611200 290112 625864 290336
rect 626808 290112 626860 290336
rect 610600 290084 626860 290112
rect 6960 289792 16260 289820
rect 6960 289568 7012 289792
rect 7956 289568 15660 289792
rect 16204 289568 16260 289792
rect 6960 289540 16260 289568
rect 616360 289792 625660 289820
rect 616360 289568 616416 289792
rect 616960 289568 624664 289792
rect 625608 289568 625660 289792
rect 616360 289540 625660 289568
rect 8160 289248 17220 289276
rect 8160 289024 8212 289248
rect 9156 289024 16620 289248
rect 17164 289024 17220 289248
rect 8160 288996 17220 289024
rect 615400 289248 624460 289276
rect 615400 289024 615456 289248
rect 616000 289024 623464 289248
rect 624408 289024 624460 289248
rect 615400 288996 624460 289024
rect 9360 288704 18170 288732
rect 9360 288480 9412 288704
rect 10356 288480 17580 288704
rect 18124 288480 18170 288704
rect 9360 288452 18170 288480
rect 614450 288704 623260 288732
rect 614450 288480 614496 288704
rect 615040 288480 622264 288704
rect 623208 288480 623260 288704
rect 614450 288452 623260 288480
rect 10560 288160 19160 288188
rect 10560 287936 10612 288160
rect 11556 287936 18540 288160
rect 19084 287936 19160 288160
rect 10560 287908 19160 287936
rect 613460 288160 622060 288188
rect 613460 287936 613536 288160
rect 614080 287936 621064 288160
rect 622008 287936 622060 288160
rect 613460 287908 622060 287936
rect 11760 287616 20120 287644
rect 11760 287392 11812 287616
rect 12756 287392 19500 287616
rect 20044 287392 20120 287616
rect 11760 287364 20120 287392
rect 612500 287616 620860 287644
rect 612500 287392 612576 287616
rect 613120 287392 619864 287616
rect 620808 287392 620860 287616
rect 612500 287364 620860 287392
rect 12960 287072 21060 287100
rect 12960 286848 13012 287072
rect 13956 286848 20460 287072
rect 21004 286848 21060 287072
rect 12960 286820 21060 286848
rect 611560 287072 619660 287100
rect 611560 286848 611616 287072
rect 612160 286848 618664 287072
rect 619608 286848 619660 287072
rect 611560 286820 619660 286848
rect 4573 277824 22973 277852
rect 4573 277600 4612 277824
rect 5556 277600 22380 277824
rect 22924 277600 22973 277824
rect 4573 277572 22973 277600
rect 609647 277824 628047 277852
rect 609647 277600 609696 277824
rect 610240 277600 627064 277824
rect 628008 277600 628047 277824
rect 609647 277572 628047 277600
rect 5760 277280 22020 277308
rect 5760 277056 5812 277280
rect 6756 277056 21420 277280
rect 21964 277056 22020 277280
rect 5760 277028 22020 277056
rect 610600 277280 626860 277308
rect 610600 277056 610656 277280
rect 611200 277056 625864 277280
rect 626808 277056 626860 277280
rect 610600 277028 626860 277056
rect 6960 276736 16260 276764
rect 6960 276512 7012 276736
rect 7956 276512 15660 276736
rect 16204 276512 16260 276736
rect 6960 276484 16260 276512
rect 616360 276736 625660 276764
rect 616360 276512 616416 276736
rect 616960 276512 624664 276736
rect 625608 276512 625660 276736
rect 616360 276484 625660 276512
rect 8160 276192 17220 276220
rect 8160 275968 8212 276192
rect 9156 275968 16620 276192
rect 17164 275968 17220 276192
rect 8160 275940 17220 275968
rect 615400 276192 624460 276220
rect 615400 275968 615456 276192
rect 616000 275968 623464 276192
rect 624408 275968 624460 276192
rect 615400 275940 624460 275968
rect 9360 275648 18170 275676
rect 9360 275424 9412 275648
rect 10356 275424 17580 275648
rect 18124 275424 18170 275648
rect 9360 275396 18170 275424
rect 614450 275648 623260 275676
rect 614450 275424 614496 275648
rect 615040 275424 622264 275648
rect 623208 275424 623260 275648
rect 614450 275396 623260 275424
rect 10560 275104 19160 275132
rect 10560 274880 10612 275104
rect 11556 274880 18540 275104
rect 19084 274880 19160 275104
rect 10560 274852 19160 274880
rect 613460 275104 622060 275132
rect 613460 274880 613536 275104
rect 614080 274880 621064 275104
rect 622008 274880 622060 275104
rect 613460 274852 622060 274880
rect 11760 274560 20120 274588
rect 11760 274336 11812 274560
rect 12756 274336 19500 274560
rect 20044 274336 20120 274560
rect 11760 274308 20120 274336
rect 612500 274560 620860 274588
rect 612500 274336 612576 274560
rect 613120 274336 619864 274560
rect 620808 274336 620860 274560
rect 612500 274308 620860 274336
rect 12960 274016 21060 274044
rect 12960 273792 13012 274016
rect 13956 273792 20460 274016
rect 21004 273792 21060 274016
rect 12960 273764 21060 273792
rect 611560 274016 619660 274044
rect 611560 273792 611616 274016
rect 612160 273792 618664 274016
rect 619608 273792 619660 274016
rect 611560 273764 619660 273792
rect 4573 266944 22973 266972
rect 4573 266720 4612 266944
rect 5556 266720 22380 266944
rect 22924 266720 22973 266944
rect 4573 266692 22973 266720
rect 5760 266400 22020 266428
rect 5760 266176 5812 266400
rect 6756 266176 21420 266400
rect 21964 266176 22020 266400
rect 5760 266148 22020 266176
rect 6960 265856 16260 265884
rect 6960 265632 7012 265856
rect 7956 265632 15660 265856
rect 16204 265632 16260 265856
rect 6960 265604 16260 265632
rect 8160 265312 17220 265340
rect 8160 265088 8212 265312
rect 9156 265088 16620 265312
rect 17164 265088 17220 265312
rect 8160 265060 17220 265088
rect 9360 264768 18170 264796
rect 9360 264544 9412 264768
rect 10356 264544 17580 264768
rect 18124 264544 18170 264768
rect 9360 264516 18170 264544
rect 10560 264224 19160 264252
rect 10560 264000 10612 264224
rect 11556 264000 18540 264224
rect 19084 264000 19160 264224
rect 10560 263972 19160 264000
rect 11760 263680 20120 263708
rect 11760 263456 11812 263680
rect 12756 263456 19500 263680
rect 20044 263456 20120 263680
rect 11760 263428 20120 263456
rect 12960 263136 21060 263164
rect 12960 262912 13012 263136
rect 13956 262912 20460 263136
rect 21004 262912 21060 263136
rect 12960 262884 21060 262912
rect 609647 263136 628047 263164
rect 609647 262912 609696 263136
rect 610240 262912 627064 263136
rect 628008 262912 628047 263136
rect 609647 262884 628047 262912
rect 610600 262592 626860 262620
rect 610600 262368 610656 262592
rect 611200 262368 625864 262592
rect 626808 262368 626860 262592
rect 610600 262340 626860 262368
rect 616360 262048 625660 262076
rect 616360 261824 616416 262048
rect 616960 261824 624664 262048
rect 625608 261824 625660 262048
rect 616360 261796 625660 261824
rect 615400 261504 624460 261532
rect 615400 261280 615456 261504
rect 616000 261280 623464 261504
rect 624408 261280 624460 261504
rect 615400 261252 624460 261280
rect 614450 260960 623260 260988
rect 614450 260736 614496 260960
rect 615040 260736 622264 260960
rect 623208 260736 623260 260960
rect 614450 260708 623260 260736
rect 613460 260416 622060 260444
rect 613460 260192 613536 260416
rect 614080 260192 621064 260416
rect 622008 260192 622060 260416
rect 613460 260164 622060 260192
rect 612500 259872 620860 259900
rect 612500 259648 612576 259872
rect 613120 259648 619864 259872
rect 620808 259648 620860 259872
rect 612500 259620 620860 259648
rect 611560 259328 619660 259356
rect 611560 259104 611616 259328
rect 612160 259104 618664 259328
rect 619608 259104 619660 259328
rect 611560 259076 619660 259104
rect 4573 251712 22973 251740
rect 4573 251488 4612 251712
rect 5556 251488 22380 251712
rect 22924 251488 22973 251712
rect 4573 251460 22973 251488
rect 609647 251712 628047 251740
rect 609647 251488 609696 251712
rect 610240 251488 627064 251712
rect 628008 251488 628047 251712
rect 609647 251460 628047 251488
rect 5760 251168 22020 251196
rect 5760 250944 5812 251168
rect 6756 250944 21420 251168
rect 21964 250944 22020 251168
rect 5760 250916 22020 250944
rect 610600 251168 626860 251196
rect 610600 250944 610656 251168
rect 611200 250944 625864 251168
rect 626808 250944 626860 251168
rect 610600 250916 626860 250944
rect 6960 250624 16260 250652
rect 6960 250400 7012 250624
rect 7956 250400 15660 250624
rect 16204 250400 16260 250624
rect 6960 250372 16260 250400
rect 616360 250624 625660 250652
rect 616360 250400 616416 250624
rect 616960 250400 624664 250624
rect 625608 250400 625660 250624
rect 616360 250372 625660 250400
rect 8160 250080 17220 250108
rect 8160 249856 8212 250080
rect 9156 249856 16620 250080
rect 17164 249856 17220 250080
rect 8160 249828 17220 249856
rect 615400 250080 624460 250108
rect 615400 249856 615456 250080
rect 616000 249856 623464 250080
rect 624408 249856 624460 250080
rect 615400 249828 624460 249856
rect 9360 249536 18170 249564
rect 9360 249312 9412 249536
rect 10356 249312 17580 249536
rect 18124 249312 18170 249536
rect 9360 249284 18170 249312
rect 614450 249536 623260 249564
rect 614450 249312 614496 249536
rect 615040 249312 622264 249536
rect 623208 249312 623260 249536
rect 614450 249284 623260 249312
rect 10560 248992 19160 249020
rect 10560 248768 10612 248992
rect 11556 248768 18540 248992
rect 19084 248768 19160 248992
rect 10560 248740 19160 248768
rect 613460 248992 622060 249020
rect 613460 248768 613536 248992
rect 614080 248768 621064 248992
rect 622008 248768 622060 248992
rect 613460 248740 622060 248768
rect 11760 248448 20120 248476
rect 11760 248224 11812 248448
rect 12756 248224 19500 248448
rect 20044 248224 20120 248448
rect 11760 248196 20120 248224
rect 612500 248448 620860 248476
rect 612500 248224 612576 248448
rect 613120 248224 619864 248448
rect 620808 248224 620860 248448
rect 612500 248196 620860 248224
rect 12960 247904 21060 247932
rect 12960 247680 13012 247904
rect 13956 247680 20460 247904
rect 21004 247680 21060 247904
rect 12960 247652 21060 247680
rect 611560 247904 619660 247932
rect 611560 247680 611616 247904
rect 612160 247680 618664 247904
rect 619608 247680 619660 247904
rect 611560 247652 619660 247680
rect 4573 238656 22973 238684
rect 4573 238432 4612 238656
rect 5556 238432 22380 238656
rect 22924 238432 22973 238656
rect 4573 238404 22973 238432
rect 609647 238656 628047 238684
rect 609647 238432 609696 238656
rect 610240 238432 627064 238656
rect 628008 238432 628047 238656
rect 609647 238404 628047 238432
rect 5760 238112 22020 238140
rect 5760 237888 5812 238112
rect 6756 237888 21420 238112
rect 21964 237888 22020 238112
rect 5760 237860 22020 237888
rect 610600 238112 626860 238140
rect 610600 237888 610656 238112
rect 611200 237888 625864 238112
rect 626808 237888 626860 238112
rect 610600 237860 626860 237888
rect 6960 237568 16260 237596
rect 6960 237344 7012 237568
rect 7956 237344 15660 237568
rect 16204 237344 16260 237568
rect 6960 237316 16260 237344
rect 616360 237568 625660 237596
rect 616360 237344 616416 237568
rect 616960 237344 624664 237568
rect 625608 237344 625660 237568
rect 616360 237316 625660 237344
rect 8160 237024 17220 237052
rect 8160 236800 8212 237024
rect 9156 236800 16620 237024
rect 17164 236800 17220 237024
rect 8160 236772 17220 236800
rect 615400 237024 624460 237052
rect 615400 236800 615456 237024
rect 616000 236800 623464 237024
rect 624408 236800 624460 237024
rect 615400 236772 624460 236800
rect 9360 236480 18170 236508
rect 9360 236256 9412 236480
rect 10356 236256 17580 236480
rect 18124 236256 18170 236480
rect 9360 236228 18170 236256
rect 614450 236480 623260 236508
rect 614450 236256 614496 236480
rect 615040 236256 622264 236480
rect 623208 236256 623260 236480
rect 614450 236228 623260 236256
rect 10560 235936 19160 235964
rect 10560 235712 10612 235936
rect 11556 235712 18540 235936
rect 19084 235712 19160 235936
rect 10560 235684 19160 235712
rect 613460 235936 622060 235964
rect 613460 235712 613536 235936
rect 614080 235712 621064 235936
rect 622008 235712 622060 235936
rect 613460 235684 622060 235712
rect 11760 235392 20120 235420
rect 11760 235168 11812 235392
rect 12756 235168 19500 235392
rect 20044 235168 20120 235392
rect 11760 235140 20120 235168
rect 612500 235392 620860 235420
rect 612500 235168 612576 235392
rect 613120 235168 619864 235392
rect 620808 235168 620860 235392
rect 612500 235140 620860 235168
rect 12960 234848 21060 234876
rect 12960 234624 13012 234848
rect 13956 234624 20460 234848
rect 21004 234624 21060 234848
rect 12960 234596 21060 234624
rect 611560 234848 619660 234876
rect 611560 234624 611616 234848
rect 612160 234624 618664 234848
rect 619608 234624 619660 234848
rect 611560 234596 619660 234624
rect 4573 225600 22973 225628
rect 4573 225376 4612 225600
rect 5556 225376 22380 225600
rect 22924 225376 22973 225600
rect 4573 225348 22973 225376
rect 609647 225600 628047 225628
rect 609647 225376 609696 225600
rect 610240 225376 627064 225600
rect 628008 225376 628047 225600
rect 609647 225348 628047 225376
rect 5760 225056 22020 225084
rect 5760 224832 5812 225056
rect 6756 224832 21420 225056
rect 21964 224832 22020 225056
rect 5760 224804 22020 224832
rect 610600 225056 626860 225084
rect 610600 224832 610656 225056
rect 611200 224832 625864 225056
rect 626808 224832 626860 225056
rect 610600 224804 626860 224832
rect 6960 224512 16260 224540
rect 6960 224288 7012 224512
rect 7956 224288 15660 224512
rect 16204 224288 16260 224512
rect 6960 224260 16260 224288
rect 616360 224512 625660 224540
rect 616360 224288 616416 224512
rect 616960 224288 624664 224512
rect 625608 224288 625660 224512
rect 616360 224260 625660 224288
rect 8160 223968 17220 223996
rect 8160 223744 8212 223968
rect 9156 223744 16620 223968
rect 17164 223744 17220 223968
rect 8160 223716 17220 223744
rect 615400 223968 624460 223996
rect 615400 223744 615456 223968
rect 616000 223744 623464 223968
rect 624408 223744 624460 223968
rect 615400 223716 624460 223744
rect 9360 223424 18170 223452
rect 9360 223200 9412 223424
rect 10356 223200 17580 223424
rect 18124 223200 18170 223424
rect 9360 223172 18170 223200
rect 614450 223424 623260 223452
rect 614450 223200 614496 223424
rect 615040 223200 622264 223424
rect 623208 223200 623260 223424
rect 614450 223172 623260 223200
rect 10560 222880 19160 222908
rect 10560 222656 10612 222880
rect 11556 222656 18540 222880
rect 19084 222656 19160 222880
rect 10560 222628 19160 222656
rect 613460 222880 622060 222908
rect 613460 222656 613536 222880
rect 614080 222656 621064 222880
rect 622008 222656 622060 222880
rect 613460 222628 622060 222656
rect 11760 222336 20120 222364
rect 11760 222112 11812 222336
rect 12756 222112 19500 222336
rect 20044 222112 20120 222336
rect 11760 222084 20120 222112
rect 612500 222336 620860 222364
rect 612500 222112 612576 222336
rect 613120 222112 619864 222336
rect 620808 222112 620860 222336
rect 612500 222084 620860 222112
rect 12960 221792 21060 221820
rect 12960 221568 13012 221792
rect 13956 221568 20460 221792
rect 21004 221568 21060 221792
rect 12960 221540 21060 221568
rect 611560 221792 619660 221820
rect 611560 221568 611616 221792
rect 612160 221568 618664 221792
rect 619608 221568 619660 221792
rect 611560 221540 619660 221568
rect 609647 212544 628047 212572
rect 609647 212320 609696 212544
rect 610240 212320 627064 212544
rect 628008 212320 628047 212544
rect 609647 212292 628047 212320
rect 610600 212000 626860 212028
rect 610600 211776 610656 212000
rect 611200 211776 625864 212000
rect 626808 211776 626860 212000
rect 610600 211748 626860 211776
rect 4573 211456 22973 211484
rect 4573 211232 4612 211456
rect 5556 211232 22380 211456
rect 22924 211232 22973 211456
rect 4573 211204 22973 211232
rect 616360 211456 625660 211484
rect 616360 211232 616416 211456
rect 616960 211232 624664 211456
rect 625608 211232 625660 211456
rect 616360 211204 625660 211232
rect 5760 210912 22020 210940
rect 5760 210688 5812 210912
rect 6756 210688 21420 210912
rect 21964 210688 22020 210912
rect 5760 210660 22020 210688
rect 615400 210912 624460 210940
rect 615400 210688 615456 210912
rect 616000 210688 623464 210912
rect 624408 210688 624460 210912
rect 615400 210660 624460 210688
rect 6960 210368 16260 210396
rect 6960 210144 7012 210368
rect 7956 210144 15660 210368
rect 16204 210144 16260 210368
rect 6960 210116 16260 210144
rect 614450 210368 623260 210396
rect 614450 210144 614496 210368
rect 615040 210144 622264 210368
rect 623208 210144 623260 210368
rect 614450 210116 623260 210144
rect 8160 209824 17220 209852
rect 8160 209600 8212 209824
rect 9156 209600 16620 209824
rect 17164 209600 17220 209824
rect 8160 209572 17220 209600
rect 613460 209824 622060 209852
rect 613460 209600 613536 209824
rect 614080 209600 621064 209824
rect 622008 209600 622060 209824
rect 613460 209572 622060 209600
rect 9360 209280 18170 209308
rect 9360 209056 9412 209280
rect 10356 209056 17580 209280
rect 18124 209056 18170 209280
rect 9360 209028 18170 209056
rect 612500 209280 620860 209308
rect 612500 209056 612576 209280
rect 613120 209056 619864 209280
rect 620808 209056 620860 209280
rect 612500 209028 620860 209056
rect 10560 208736 19160 208764
rect 10560 208512 10612 208736
rect 11556 208512 18540 208736
rect 19084 208512 19160 208736
rect 10560 208484 19160 208512
rect 611560 208736 619660 208764
rect 611560 208512 611616 208736
rect 612160 208512 618664 208736
rect 619608 208512 619660 208736
rect 611560 208484 619660 208512
rect 11760 208192 20120 208220
rect 11760 207968 11812 208192
rect 12756 207968 19500 208192
rect 20044 207968 20120 208192
rect 11760 207940 20120 207968
rect 12960 207648 21060 207676
rect 12960 207424 13012 207648
rect 13956 207424 20460 207648
rect 21004 207424 21060 207648
rect 12960 207396 21060 207424
rect -3216 40758 1182 40840
rect -3216 36134 -1777 40758
rect 1087 36134 1182 40758
rect -3216 36051 1182 36134
rect -3216 30718 1182 30800
rect -3216 26094 -1777 30718
rect 1087 26094 1182 30718
rect 208144 27328 212703 27373
rect 208144 27104 208191 27328
rect 209055 27104 212703 27328
rect 208144 27054 212703 27104
rect 226824 26900 227464 26936
rect 223584 26888 227464 26900
rect 223584 26664 226871 26888
rect 227415 26664 227464 26888
rect 223584 26653 227464 26664
rect 226824 26619 227464 26653
rect -3216 26011 1182 26094
rect 130944 7832 139976 7881
rect 130944 7608 130995 7832
rect 131859 7733 139976 7832
rect 131859 7608 139772 7733
rect 130944 7589 139772 7608
rect 139916 7589 139976 7733
rect 130944 7560 139976 7589
rect 132304 7169 138678 7214
rect 132304 7168 138472 7169
rect 132304 6944 132347 7168
rect 133211 7025 138472 7168
rect 138616 7025 138678 7169
rect 133211 6944 138678 7025
rect 132304 6894 138678 6944
rect 198943 -112 203749 -22
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -2938 203749 -1696
rect 208994 -112 213800 -22
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -2938 213800 -1696
<< via3 >>
rect 533467 952770 538091 954354
rect 543448 952770 548072 954354
rect 609696 910816 610240 911040
rect 627064 910816 628008 911040
rect 610656 910272 611200 910496
rect 625864 910272 626808 910496
rect 616416 909728 616960 909952
rect 624664 909728 625608 909952
rect 615456 909184 616000 909408
rect 623464 909184 624408 909408
rect 614496 908640 615040 908864
rect 622264 908640 623208 908864
rect 613536 908096 614080 908320
rect 621064 908096 622008 908320
rect 612576 907552 613120 907776
rect 619864 907552 620808 907776
rect 611616 907008 612160 907232
rect 618664 907008 619608 907232
rect 4612 905920 5556 906144
rect 22380 905920 22924 906144
rect 5812 905376 6756 905600
rect 21420 905376 21964 905600
rect 7012 904832 7956 905056
rect 15660 904832 16204 905056
rect 8212 904288 9156 904512
rect 16620 904288 17164 904512
rect 9412 903744 10356 903968
rect 17580 903744 18124 903968
rect 10612 903200 11556 903424
rect 18540 903200 19084 903424
rect 11812 902656 12756 902880
rect 19500 902656 20044 902880
rect 13012 902112 13956 902336
rect 20460 902112 21004 902336
rect 609696 896128 610240 896352
rect 627064 896128 628008 896352
rect 610656 895584 611200 895808
rect 625864 895584 626808 895808
rect 616416 895040 616960 895264
rect 624664 895040 625608 895264
rect 615456 894496 616000 894720
rect 623464 894496 624408 894720
rect 614496 893952 615040 894176
rect 622264 893952 623208 894176
rect 613536 893408 614080 893632
rect 621064 893408 622008 893632
rect 612576 892864 613120 893088
rect 619864 892864 620808 893088
rect 611616 892320 612160 892544
rect 618664 892320 619608 892544
rect 4612 891232 5556 891456
rect 22380 891232 22924 891456
rect 5812 890688 6756 890912
rect 21420 890688 21964 890912
rect 7012 890144 7956 890368
rect 15660 890144 16204 890368
rect 8212 889600 9156 889824
rect 16620 889600 17164 889824
rect 9412 889056 10356 889280
rect 17580 889056 18124 889280
rect 10612 888512 11556 888736
rect 18540 888512 19084 888736
rect 11812 887968 12756 888192
rect 19500 887968 20044 888192
rect 13012 887424 13956 887648
rect 20460 887424 21004 887648
rect -1777 880134 1087 884758
rect 609696 884704 610240 884928
rect 627064 884704 628008 884928
rect 610656 884160 611200 884384
rect 625864 884160 626808 884384
rect 616416 883616 616960 883840
rect 624664 883616 625608 883840
rect 615456 883072 616000 883296
rect 623464 883072 624408 883296
rect 614496 882528 615040 882752
rect 622264 882528 623208 882752
rect 613536 881984 614080 882208
rect 621064 881984 622008 882208
rect 612576 881440 613120 881664
rect 619864 881440 620808 881664
rect 611616 880896 612160 881120
rect 618664 880896 619608 881120
rect -1777 875184 1087 879648
rect 4612 878176 5556 878400
rect 22380 878176 22924 878400
rect 5812 877632 6756 877856
rect 21420 877632 21964 877856
rect 7012 877088 7956 877312
rect 15660 877088 16204 877312
rect 8212 876544 9156 876768
rect 16620 876544 17164 876768
rect 9412 876000 10356 876224
rect 17580 876000 18124 876224
rect 10612 875456 11556 875680
rect 18540 875456 19084 875680
rect 631301 875694 634165 880318
rect 11812 874912 12756 875136
rect 19500 874912 20044 875136
rect -1777 870094 1087 874718
rect 13012 874368 13956 874592
rect 20460 874368 21004 874592
rect 609696 871648 610240 871872
rect 627064 871648 628008 871872
rect 610656 871104 611200 871328
rect 625864 871104 626808 871328
rect 616416 870560 616960 870784
rect 624664 870560 625608 870784
rect 631301 870744 634165 875208
rect 615456 870016 616000 870240
rect 623464 870016 624408 870240
rect 614496 869472 615040 869696
rect 622264 869472 623208 869696
rect 613536 868928 614080 869152
rect 621064 868928 622008 869152
rect 612576 868384 613120 868608
rect 619864 868384 620808 868608
rect 611616 867840 612160 868064
rect 618664 867840 619608 868064
rect 631301 865643 634165 870267
rect 4612 865120 5556 865344
rect 22380 865120 22924 865344
rect 5812 864576 6756 864800
rect 21420 864576 21964 864800
rect 7012 864032 7956 864256
rect 15660 864032 16204 864256
rect 8212 863488 9156 863712
rect 16620 863488 17164 863712
rect 9412 862944 10356 863168
rect 17580 862944 18124 863168
rect 10612 862400 11556 862624
rect 18540 862400 19084 862624
rect 11812 861856 12756 862080
rect 19500 861856 20044 862080
rect 13012 861312 13956 861536
rect 20460 861312 21004 861536
rect 609696 858592 610240 858816
rect 627064 858592 628008 858816
rect 610656 858048 611200 858272
rect 625864 858048 626808 858272
rect 616416 857504 616960 857728
rect 624664 857504 625608 857728
rect 615456 856960 616000 857184
rect 623464 856960 624408 857184
rect 614496 856416 615040 856640
rect 622264 856416 623208 856640
rect 613536 855872 614080 856096
rect 621064 855872 622008 856096
rect 612576 855328 613120 855552
rect 619864 855328 620808 855552
rect 611616 854784 612160 855008
rect 618664 854784 619608 855008
rect 4612 852064 5556 852288
rect 22380 852064 22924 852288
rect 5812 851520 6756 851744
rect 21420 851520 21964 851744
rect 7012 850976 7956 851200
rect 15660 850976 16204 851200
rect 8212 850432 9156 850656
rect 16620 850432 17164 850656
rect 9412 849888 10356 850112
rect 17580 849888 18124 850112
rect 10612 849344 11556 849568
rect 18540 849344 19084 849568
rect 11812 848800 12756 849024
rect 19500 848800 20044 849024
rect 13012 848256 13956 848480
rect 20460 848256 21004 848480
rect 609696 845536 610240 845760
rect 627064 845536 628008 845760
rect 610656 844992 611200 845216
rect 625864 844992 626808 845216
rect 616416 844448 616960 844672
rect 624664 844448 625608 844672
rect 615456 843904 616000 844128
rect 623464 843904 624408 844128
rect 614496 843360 615040 843584
rect 622264 843360 623208 843584
rect 613536 842816 614080 843040
rect 621064 842816 622008 843040
rect 612576 842272 613120 842496
rect 619864 842272 620808 842496
rect 611616 841728 612160 841952
rect 618664 841728 619608 841952
rect 4612 839008 5556 839232
rect 22380 839008 22924 839232
rect 5812 838464 6756 838688
rect 21420 838464 21964 838688
rect 7012 837920 7956 838144
rect 15660 837920 16204 838144
rect 8212 837376 9156 837600
rect 16620 837376 17164 837600
rect 9412 836832 10356 837056
rect 17580 836832 18124 837056
rect 10612 836288 11556 836512
rect 18540 836288 19084 836512
rect 11812 835744 12756 835968
rect 19500 835744 20044 835968
rect 13012 835200 13956 835424
rect 20460 835200 21004 835424
rect 609696 832480 610240 832704
rect 627064 832480 628008 832704
rect 610656 831936 611200 832160
rect 625864 831936 626808 832160
rect 616416 831392 616960 831616
rect 624664 831392 625608 831616
rect 615456 830848 616000 831072
rect 623464 830848 624408 831072
rect 614496 830304 615040 830528
rect 622264 830304 623208 830528
rect 613536 829760 614080 829984
rect 621064 829760 622008 829984
rect 612576 829216 613120 829440
rect 619864 829216 620808 829440
rect 611616 828672 612160 828896
rect 618664 828672 619608 828896
rect 4612 825952 5556 826176
rect 22380 825952 22924 826176
rect 5812 825408 6756 825632
rect 21420 825408 21964 825632
rect 7012 824864 7956 825088
rect 15660 824864 16204 825088
rect 8212 824320 9156 824544
rect 16620 824320 17164 824544
rect 9412 823776 10356 824000
rect 17580 823776 18124 824000
rect 10612 823232 11556 823456
rect 18540 823232 19084 823456
rect 11812 822688 12756 822912
rect 19500 822688 20044 822912
rect 13012 822144 13956 822368
rect 20460 822144 21004 822368
rect 609696 819424 610240 819648
rect 627064 819424 628008 819648
rect 610656 818880 611200 819104
rect 625864 818880 626808 819104
rect 616416 818336 616960 818560
rect 624664 818336 625608 818560
rect 615456 817792 616000 818016
rect 623464 817792 624408 818016
rect 614496 817248 615040 817472
rect 622264 817248 623208 817472
rect 613536 816704 614080 816928
rect 621064 816704 622008 816928
rect 612576 816160 613120 816384
rect 619864 816160 620808 816384
rect 611616 815616 612160 815840
rect 618664 815616 619608 815840
rect 4612 812896 5556 813120
rect 22380 812896 22924 813120
rect 5812 812352 6756 812576
rect 21420 812352 21964 812576
rect 7012 811808 7956 812032
rect 15660 811808 16204 812032
rect 8212 811264 9156 811488
rect 16620 811264 17164 811488
rect 9412 810720 10356 810944
rect 17580 810720 18124 810944
rect 10612 810176 11556 810400
rect 18540 810176 19084 810400
rect 11812 809632 12756 809856
rect 19500 809632 20044 809856
rect 13012 809088 13956 809312
rect 20460 809088 21004 809312
rect 609696 806368 610240 806592
rect 627064 806368 628008 806592
rect 610656 805824 611200 806048
rect 625864 805824 626808 806048
rect 616416 805280 616960 805504
rect 624664 805280 625608 805504
rect 615456 804736 616000 804960
rect 623464 804736 624408 804960
rect 614496 804192 615040 804416
rect 622264 804192 623208 804416
rect 613536 803648 614080 803872
rect 621064 803648 622008 803872
rect 612576 803104 613120 803328
rect 619864 803104 620808 803328
rect 611616 802560 612160 802784
rect 618664 802560 619608 802784
rect -1777 795652 1087 800276
rect 4612 799840 5556 800064
rect 22380 799840 22924 800064
rect 5812 799296 6756 799520
rect 21420 799296 21964 799520
rect 7012 798752 7956 798976
rect 15660 798752 16204 798976
rect 8212 798208 9156 798432
rect 16620 798208 17164 798432
rect 9412 797664 10356 797888
rect 17580 797664 18124 797888
rect 10612 797120 11556 797344
rect 18540 797120 19084 797344
rect 11812 796576 12756 796800
rect 19500 796576 20044 796800
rect 13012 796032 13956 796256
rect 20460 796032 21004 796256
rect 609696 793312 610240 793536
rect 627064 793312 628008 793536
rect 610656 792768 611200 792992
rect 625864 792768 626808 792992
rect 616416 792224 616960 792448
rect 624664 792224 625608 792448
rect 615456 791680 616000 791904
rect 623464 791680 624408 791904
rect 614496 791136 615040 791360
rect 622264 791136 623208 791360
rect 613536 790592 614080 790816
rect 621064 790592 622008 790816
rect -1777 785673 1087 790297
rect 612576 790048 613120 790272
rect 619864 790048 620808 790272
rect 611616 789504 612160 789728
rect 618664 789504 619608 789728
rect 4612 786784 5556 787008
rect 22380 786784 22924 787008
rect 631301 786495 634165 791119
rect 5812 786240 6756 786464
rect 21420 786240 21964 786464
rect 7012 785696 7956 785920
rect 15660 785696 16204 785920
rect 8212 785152 9156 785376
rect 16620 785152 17164 785376
rect 9412 784608 10356 784832
rect 17580 784608 18124 784832
rect 10612 784064 11556 784288
rect 18540 784064 19084 784288
rect 11812 783520 12756 783744
rect 19500 783520 20044 783744
rect 13012 782976 13956 783200
rect 20460 782976 21004 783200
rect 609696 780256 610240 780480
rect 627064 780256 628008 780480
rect 610656 779712 611200 779936
rect 625864 779712 626808 779936
rect 616416 779168 616960 779392
rect 624664 779168 625608 779392
rect 615456 778624 616000 778848
rect 623464 778624 624408 778848
rect 614496 778080 615040 778304
rect 622264 778080 623208 778304
rect 613536 777536 614080 777760
rect 621064 777536 622008 777760
rect 612576 776992 613120 777216
rect 619864 776992 620808 777216
rect 611616 776448 612160 776672
rect 618664 776448 619608 776672
rect 631301 776512 634165 781136
rect 4612 773728 5556 773952
rect 22380 773728 22924 773952
rect 5812 773184 6756 773408
rect 21420 773184 21964 773408
rect 7012 772640 7956 772864
rect 15660 772640 16204 772864
rect 8212 772096 9156 772320
rect 16620 772096 17164 772320
rect 9412 771552 10356 771776
rect 17580 771552 18124 771776
rect 10612 771008 11556 771232
rect 18540 771008 19084 771232
rect 11812 770464 12756 770688
rect 19500 770464 20044 770688
rect 13012 769920 13956 770144
rect 20460 769920 21004 770144
rect 609696 767200 610240 767424
rect 627064 767200 628008 767424
rect 610656 766656 611200 766880
rect 625864 766656 626808 766880
rect 616416 766112 616960 766336
rect 624664 766112 625608 766336
rect 615456 765568 616000 765792
rect 623464 765568 624408 765792
rect 614496 765024 615040 765248
rect 622264 765024 623208 765248
rect 613536 764480 614080 764704
rect 621064 764480 622008 764704
rect 612576 763936 613120 764160
rect 619864 763936 620808 764160
rect 611616 763392 612160 763616
rect 618664 763392 619608 763616
rect 4612 760672 5556 760896
rect 22380 760672 22924 760896
rect 5812 760128 6756 760352
rect 21420 760128 21964 760352
rect 7012 759584 7956 759808
rect 15660 759584 16204 759808
rect 8212 759040 9156 759264
rect 16620 759040 17164 759264
rect 9412 758496 10356 758720
rect 17580 758496 18124 758720
rect 10612 757952 11556 758176
rect 18540 757952 19084 758176
rect 11812 757408 12756 757632
rect 19500 757408 20044 757632
rect 13012 756864 13956 757088
rect 20460 756864 21004 757088
rect 609696 754144 610240 754368
rect 627064 754144 628008 754368
rect 610656 753600 611200 753824
rect 625864 753600 626808 753824
rect 616416 753056 616960 753280
rect 624664 753056 625608 753280
rect 615456 752512 616000 752736
rect 623464 752512 624408 752736
rect 614496 751968 615040 752192
rect 622264 751968 623208 752192
rect 613536 751424 614080 751648
rect 621064 751424 622008 751648
rect 612576 750880 613120 751104
rect 619864 750880 620808 751104
rect 611616 750336 612160 750560
rect 618664 750336 619608 750560
rect 4612 747616 5556 747840
rect 22380 747616 22924 747840
rect 5812 747072 6756 747296
rect 21420 747072 21964 747296
rect 7012 746528 7956 746752
rect 15660 746528 16204 746752
rect 8212 745984 9156 746208
rect 16620 745984 17164 746208
rect 9412 745440 10356 745664
rect 17580 745440 18124 745664
rect 10612 744896 11556 745120
rect 18540 744896 19084 745120
rect 11812 744352 12756 744576
rect 19500 744352 20044 744576
rect 13012 743808 13956 744032
rect 20460 743808 21004 744032
rect 609696 741088 610240 741312
rect 627064 741088 628008 741312
rect 610656 740544 611200 740768
rect 625864 740544 626808 740768
rect 616416 740000 616960 740224
rect 624664 740000 625608 740224
rect 615456 739456 616000 739680
rect 623464 739456 624408 739680
rect 614496 738912 615040 739136
rect 622264 738912 623208 739136
rect 613536 738368 614080 738592
rect 621064 738368 622008 738592
rect 612576 737824 613120 738048
rect 619864 737824 620808 738048
rect 611616 737280 612160 737504
rect 618664 737280 619608 737504
rect 4612 736192 5556 736416
rect 22380 736192 22924 736416
rect 5812 735648 6756 735872
rect 21420 735648 21964 735872
rect 7012 735104 7956 735328
rect 15660 735104 16204 735328
rect 8212 734560 9156 734784
rect 16620 734560 17164 734784
rect 9412 734016 10356 734240
rect 17580 734016 18124 734240
rect 10612 733472 11556 733696
rect 18540 733472 19084 733696
rect 11812 732928 12756 733152
rect 19500 732928 20044 733152
rect 13012 732384 13956 732608
rect 20460 732384 21004 732608
rect 609696 728032 610240 728256
rect 627064 728032 628008 728256
rect 610656 727488 611200 727712
rect 625864 727488 626808 727712
rect 616416 726944 616960 727168
rect 624664 726944 625608 727168
rect 615456 726400 616000 726624
rect 623464 726400 624408 726624
rect 614496 725856 615040 726080
rect 622264 725856 623208 726080
rect 613536 725312 614080 725536
rect 621064 725312 622008 725536
rect 612576 724768 613120 724992
rect 619864 724768 620808 724992
rect 611616 724224 612160 724448
rect 618664 724224 619608 724448
rect 4612 721504 5556 721728
rect 22380 721504 22924 721728
rect 5812 720960 6756 721184
rect 21420 720960 21964 721184
rect 7012 720416 7956 720640
rect 15660 720416 16204 720640
rect 8212 719872 9156 720096
rect 16620 719872 17164 720096
rect 9412 719328 10356 719552
rect 17580 719328 18124 719552
rect 10612 718784 11556 719008
rect 18540 718784 19084 719008
rect 11812 718240 12756 718464
rect 19500 718240 20044 718464
rect 13012 717696 13956 717920
rect 20460 717696 21004 717920
rect 609696 713344 610240 713568
rect 627064 713344 628008 713568
rect 610656 712800 611200 713024
rect 625864 712800 626808 713024
rect 616416 712256 616960 712480
rect 624664 712256 625608 712480
rect 615456 711712 616000 711936
rect 623464 711712 624408 711936
rect 614496 711168 615040 711392
rect 622264 711168 623208 711392
rect 613536 710624 614080 710848
rect 621064 710624 622008 710848
rect 612576 710080 613120 710304
rect 619864 710080 620808 710304
rect 611616 709536 612160 709760
rect 618664 709536 619608 709760
rect 4612 708448 5556 708672
rect 22380 708448 22924 708672
rect 5812 707904 6756 708128
rect 21420 707904 21964 708128
rect 7012 707360 7956 707584
rect 15660 707360 16204 707584
rect 8212 706816 9156 707040
rect 16620 706816 17164 707040
rect 9412 706272 10356 706496
rect 17580 706272 18124 706496
rect 10612 705728 11556 705952
rect 18540 705728 19084 705952
rect 11812 705184 12756 705408
rect 19500 705184 20044 705408
rect 13012 704640 13956 704864
rect 20460 704640 21004 704864
rect 609696 701920 610240 702144
rect 627064 701920 628008 702144
rect 610656 701376 611200 701600
rect 625864 701376 626808 701600
rect 616416 700832 616960 701056
rect 624664 700832 625608 701056
rect 615456 700288 616000 700512
rect 623464 700288 624408 700512
rect 614496 699744 615040 699968
rect 622264 699744 623208 699968
rect 613536 699200 614080 699424
rect 621064 699200 622008 699424
rect 612576 698656 613120 698880
rect 619864 698656 620808 698880
rect 611616 698112 612160 698336
rect 618664 698112 619608 698336
rect 4612 692128 5556 692352
rect 22380 692128 22924 692352
rect 5812 691584 6756 691808
rect 21420 691584 21964 691808
rect 7012 691040 7956 691264
rect 15660 691040 16204 691264
rect 8212 690496 9156 690720
rect 16620 690496 17164 690720
rect 9412 689952 10356 690176
rect 17580 689952 18124 690176
rect 10612 689408 11556 689632
rect 18540 689408 19084 689632
rect 11812 688864 12756 689088
rect 19500 688864 20044 689088
rect 609696 688864 610240 689088
rect 627064 688864 628008 689088
rect 13012 688320 13956 688544
rect 20460 688320 21004 688544
rect 610656 688320 611200 688544
rect 625864 688320 626808 688544
rect 616416 687776 616960 688000
rect 624664 687776 625608 688000
rect 615456 687232 616000 687456
rect 623464 687232 624408 687456
rect 614496 686688 615040 686912
rect 622264 686688 623208 686912
rect 613536 686144 614080 686368
rect 621064 686144 622008 686368
rect 612576 685600 613120 685824
rect 619864 685600 620808 685824
rect 611616 685056 612160 685280
rect 618664 685056 619608 685280
rect 4612 682336 5556 682560
rect 22380 682336 22924 682560
rect 5812 681792 6756 682016
rect 21420 681792 21964 682016
rect 7012 681248 7956 681472
rect 15660 681248 16204 681472
rect 8212 680704 9156 680928
rect 16620 680704 17164 680928
rect 9412 680160 10356 680384
rect 17580 680160 18124 680384
rect 10612 679616 11556 679840
rect 18540 679616 19084 679840
rect 11812 679072 12756 679296
rect 19500 679072 20044 679296
rect 13012 678528 13956 678752
rect 20460 678528 21004 678752
rect 609696 675808 610240 676032
rect 627064 675808 628008 676032
rect 610656 675264 611200 675488
rect 625864 675264 626808 675488
rect 616416 674720 616960 674944
rect 624664 674720 625608 674944
rect 615456 674176 616000 674400
rect 623464 674176 624408 674400
rect 614496 673632 615040 673856
rect 622264 673632 623208 673856
rect 613536 673088 614080 673312
rect 621064 673088 622008 673312
rect 612576 672544 613120 672768
rect 619864 672544 620808 672768
rect 611616 672000 612160 672224
rect 618664 672000 619608 672224
rect 4612 669280 5556 669504
rect 22380 669280 22924 669504
rect 5812 668736 6756 668960
rect 21420 668736 21964 668960
rect 7012 668192 7956 668416
rect 15660 668192 16204 668416
rect 8212 667648 9156 667872
rect 16620 667648 17164 667872
rect 9412 667104 10356 667328
rect 17580 667104 18124 667328
rect 10612 666560 11556 666784
rect 18540 666560 19084 666784
rect 11812 666016 12756 666240
rect 19500 666016 20044 666240
rect 13012 665472 13956 665696
rect 20460 665472 21004 665696
rect 609696 662752 610240 662976
rect 627064 662752 628008 662976
rect 610656 662208 611200 662432
rect 625864 662208 626808 662432
rect 616416 661664 616960 661888
rect 624664 661664 625608 661888
rect 615456 661120 616000 661344
rect 623464 661120 624408 661344
rect 614496 660576 615040 660800
rect 622264 660576 623208 660800
rect 613536 660032 614080 660256
rect 621064 660032 622008 660256
rect 612576 659488 613120 659712
rect 619864 659488 620808 659712
rect 611616 658944 612160 659168
rect 618664 658944 619608 659168
rect 4612 656224 5556 656448
rect 22380 656224 22924 656448
rect 5812 655680 6756 655904
rect 21420 655680 21964 655904
rect 7012 655136 7956 655360
rect 15660 655136 16204 655360
rect 8212 654592 9156 654816
rect 16620 654592 17164 654816
rect 9412 654048 10356 654272
rect 17580 654048 18124 654272
rect 10612 653504 11556 653728
rect 18540 653504 19084 653728
rect 11812 652960 12756 653184
rect 19500 652960 20044 653184
rect 13012 652416 13956 652640
rect 20460 652416 21004 652640
rect 609696 649696 610240 649920
rect 627064 649696 628008 649920
rect 610656 649152 611200 649376
rect 625864 649152 626808 649376
rect 616416 648608 616960 648832
rect 624664 648608 625608 648832
rect 615456 648064 616000 648288
rect 623464 648064 624408 648288
rect 614496 647520 615040 647744
rect 622264 647520 623208 647744
rect 613536 646976 614080 647200
rect 621064 646976 622008 647200
rect 612576 646432 613120 646656
rect 619864 646432 620808 646656
rect 611616 645888 612160 646112
rect 618664 645888 619608 646112
rect 4612 641536 5556 641760
rect 22380 641536 22924 641760
rect 5812 640992 6756 641216
rect 21420 640992 21964 641216
rect 7012 640448 7956 640672
rect 15660 640448 16204 640672
rect 8212 639904 9156 640128
rect 16620 639904 17164 640128
rect 9412 639360 10356 639584
rect 17580 639360 18124 639584
rect 10612 638816 11556 639040
rect 18540 638816 19084 639040
rect 11812 638272 12756 638496
rect 19500 638272 20044 638496
rect 13012 637728 13956 637952
rect 20460 637728 21004 637952
rect 609696 636640 610240 636864
rect 627064 636640 628008 636864
rect 610656 636096 611200 636320
rect 625864 636096 626808 636320
rect 616416 635552 616960 635776
rect 624664 635552 625608 635776
rect 615456 635008 616000 635232
rect 623464 635008 624408 635232
rect 614496 634464 615040 634688
rect 622264 634464 623208 634688
rect 613536 633920 614080 634144
rect 621064 633920 622008 634144
rect 612576 633376 613120 633600
rect 619864 633376 620808 633600
rect 611616 632832 612160 633056
rect 618664 632832 619608 633056
rect 4612 630112 5556 630336
rect 22380 630112 22924 630336
rect 5812 629568 6756 629792
rect 21420 629568 21964 629792
rect 7012 629024 7956 629248
rect 15660 629024 16204 629248
rect 8212 628480 9156 628704
rect 16620 628480 17164 628704
rect 9412 627936 10356 628160
rect 17580 627936 18124 628160
rect 10612 627392 11556 627616
rect 18540 627392 19084 627616
rect 11812 626848 12756 627072
rect 19500 626848 20044 627072
rect 13012 626304 13956 626528
rect 20460 626304 21004 626528
rect 609696 623584 610240 623808
rect 627064 623584 628008 623808
rect 610656 623040 611200 623264
rect 625864 623040 626808 623264
rect 616416 622496 616960 622720
rect 624664 622496 625608 622720
rect 615456 621952 616000 622176
rect 623464 621952 624408 622176
rect 614496 621408 615040 621632
rect 622264 621408 623208 621632
rect 613536 620864 614080 621088
rect 621064 620864 622008 621088
rect 612576 620320 613120 620544
rect 619864 620320 620808 620544
rect 611616 619776 612160 620000
rect 618664 619776 619608 620000
rect 4612 617056 5556 617280
rect 22380 617056 22924 617280
rect 5812 616512 6756 616736
rect 21420 616512 21964 616736
rect 7012 615968 7956 616192
rect 15660 615968 16204 616192
rect 8212 615424 9156 615648
rect 16620 615424 17164 615648
rect 9412 614880 10356 615104
rect 17580 614880 18124 615104
rect 10612 614336 11556 614560
rect 18540 614336 19084 614560
rect 11812 613792 12756 614016
rect 19500 613792 20044 614016
rect 13012 613248 13956 613472
rect 20460 613248 21004 613472
rect 609696 610528 610240 610752
rect 627064 610528 628008 610752
rect 610656 609984 611200 610208
rect 625864 609984 626808 610208
rect 616416 609440 616960 609664
rect 624664 609440 625608 609664
rect 615456 608896 616000 609120
rect 623464 608896 624408 609120
rect 614496 608352 615040 608576
rect 622264 608352 623208 608576
rect 613536 607808 614080 608032
rect 621064 607808 622008 608032
rect 612576 607264 613120 607488
rect 619864 607264 620808 607488
rect 611616 606720 612160 606944
rect 618664 606720 619608 606944
rect 4612 606176 5556 606400
rect 22380 606176 22924 606400
rect 5812 605632 6756 605856
rect 21420 605632 21964 605856
rect 7012 605088 7956 605312
rect 15660 605088 16204 605312
rect 8212 604544 9156 604768
rect 16620 604544 17164 604768
rect 9412 604000 10356 604224
rect 17580 604000 18124 604224
rect 10612 603456 11556 603680
rect 18540 603456 19084 603680
rect 11812 602912 12756 603136
rect 19500 602912 20044 603136
rect 13012 602368 13956 602592
rect 20460 602368 21004 602592
rect 609696 597472 610240 597696
rect 627064 597472 628008 597696
rect 610656 596928 611200 597152
rect 625864 596928 626808 597152
rect 616416 596384 616960 596608
rect 624664 596384 625608 596608
rect 615456 595840 616000 596064
rect 623464 595840 624408 596064
rect 614496 595296 615040 595520
rect 622264 595296 623208 595520
rect 613536 594752 614080 594976
rect 621064 594752 622008 594976
rect 612576 594208 613120 594432
rect 619864 594208 620808 594432
rect 611616 593664 612160 593888
rect 618664 593664 619608 593888
rect 4612 590944 5556 591168
rect 22380 590944 22924 591168
rect 5812 590400 6756 590624
rect 21420 590400 21964 590624
rect 7012 589856 7956 590080
rect 15660 589856 16204 590080
rect 8212 589312 9156 589536
rect 16620 589312 17164 589536
rect 9412 588768 10356 588992
rect 17580 588768 18124 588992
rect 10612 588224 11556 588448
rect 18540 588224 19084 588448
rect 11812 587680 12756 587904
rect 19500 587680 20044 587904
rect 13012 587136 13956 587360
rect 20460 587136 21004 587360
rect 609696 584416 610240 584640
rect 627064 584416 628008 584640
rect 610656 583872 611200 584096
rect 625864 583872 626808 584096
rect 616416 583328 616960 583552
rect 624664 583328 625608 583552
rect 615456 582784 616000 583008
rect 623464 582784 624408 583008
rect 614496 582240 615040 582464
rect 622264 582240 623208 582464
rect 613536 581696 614080 581920
rect 621064 581696 622008 581920
rect 612576 581152 613120 581376
rect 619864 581152 620808 581376
rect 611616 580608 612160 580832
rect 618664 580608 619608 580832
rect 4612 577888 5556 578112
rect 22380 577888 22924 578112
rect 5812 577344 6756 577568
rect 21420 577344 21964 577568
rect 7012 576800 7956 577024
rect 15660 576800 16204 577024
rect 8212 576256 9156 576480
rect 16620 576256 17164 576480
rect 9412 575712 10356 575936
rect 17580 575712 18124 575936
rect 10612 575168 11556 575392
rect 18540 575168 19084 575392
rect 11812 574624 12756 574848
rect 19500 574624 20044 574848
rect 13012 574080 13956 574304
rect 20460 574080 21004 574304
rect 609696 571360 610240 571584
rect 627064 571360 628008 571584
rect 610656 570816 611200 571040
rect 625864 570816 626808 571040
rect 616416 570272 616960 570496
rect 624664 570272 625608 570496
rect 615456 569728 616000 569952
rect 623464 569728 624408 569952
rect 614496 569184 615040 569408
rect 622264 569184 623208 569408
rect 613536 568640 614080 568864
rect 621064 568640 622008 568864
rect 612576 568096 613120 568320
rect 619864 568096 620808 568320
rect 611616 567552 612160 567776
rect 618664 567552 619608 567776
rect 4612 567008 5556 567232
rect 22380 567008 22924 567232
rect 5812 566464 6756 566688
rect 21420 566464 21964 566688
rect 7012 565920 7956 566144
rect 15660 565920 16204 566144
rect 8212 565376 9156 565600
rect 16620 565376 17164 565600
rect 9412 564832 10356 565056
rect 17580 564832 18124 565056
rect 10612 564288 11556 564512
rect 18540 564288 19084 564512
rect 11812 563744 12756 563968
rect 19500 563744 20044 563968
rect 13012 563200 13956 563424
rect 20460 563200 21004 563424
rect 609696 558304 610240 558528
rect 627064 558304 628008 558528
rect 610656 557760 611200 557984
rect 625864 557760 626808 557984
rect 616416 557216 616960 557440
rect 624664 557216 625608 557440
rect 615456 556672 616000 556896
rect 623464 556672 624408 556896
rect 614496 556128 615040 556352
rect 622264 556128 623208 556352
rect 613536 555584 614080 555808
rect 621064 555584 622008 555808
rect 612576 555040 613120 555264
rect 619864 555040 620808 555264
rect 611616 554496 612160 554720
rect 618664 554496 619608 554720
rect 4612 551776 5556 552000
rect 22380 551776 22924 552000
rect 5812 551232 6756 551456
rect 21420 551232 21964 551456
rect 7012 550688 7956 550912
rect 15660 550688 16204 550912
rect 8212 550144 9156 550368
rect 16620 550144 17164 550368
rect 9412 549600 10356 549824
rect 17580 549600 18124 549824
rect 10612 549056 11556 549280
rect 18540 549056 19084 549280
rect 11812 548512 12756 548736
rect 19500 548512 20044 548736
rect 13012 547968 13956 548192
rect 20460 547968 21004 548192
rect 614496 543072 615040 543296
rect 622264 543072 623208 543296
rect 613536 542528 614080 542752
rect 621064 542528 622008 542752
rect 612576 541984 613120 542208
rect 619864 541984 620808 542208
rect 611616 541440 612160 541664
rect 618664 541440 619608 541664
rect 4612 538720 5556 538944
rect 22380 538720 22924 538944
rect 5812 538176 6756 538400
rect 21420 538176 21964 538400
rect 7012 537632 7956 537856
rect 15660 537632 16204 537856
rect 8212 537088 9156 537312
rect 16620 537088 17164 537312
rect 9412 536544 10356 536768
rect 17580 536544 18124 536768
rect 10612 536000 11556 536224
rect 18540 536000 19084 536224
rect 11812 535456 12756 535680
rect 19500 535456 20044 535680
rect 13012 534912 13956 535136
rect 20460 534912 21004 535136
rect 609696 530560 610240 530784
rect 627064 530560 628008 530784
rect 610656 530016 611200 530240
rect 625864 530016 626808 530240
rect 616416 529472 616960 529696
rect 624664 529472 625608 529696
rect 615456 528928 616000 529152
rect 623464 528928 624408 529152
rect 614496 528384 615040 528608
rect 622264 528384 623208 528608
rect 613536 527840 614080 528064
rect 621064 527840 622008 528064
rect 612576 527296 613120 527520
rect 619864 527296 620808 527520
rect 611616 526752 612160 526976
rect 618664 526752 619608 526976
rect 4612 525664 5556 525888
rect 22380 525664 22924 525888
rect 5812 525120 6756 525344
rect 21420 525120 21964 525344
rect 7012 524576 7956 524800
rect 15660 524576 16204 524800
rect 8212 524032 9156 524256
rect 16620 524032 17164 524256
rect 9412 523488 10356 523712
rect 17580 523488 18124 523712
rect 10612 522944 11556 523168
rect 18540 522944 19084 523168
rect 11812 522400 12756 522624
rect 19500 522400 20044 522624
rect 13012 521856 13956 522080
rect 20460 521856 21004 522080
rect 609696 517504 610240 517728
rect 627064 517504 628008 517728
rect 610656 516960 611200 517184
rect 625864 516960 626808 517184
rect 616416 516416 616960 516640
rect 624664 516416 625608 516640
rect 615456 515872 616000 516096
rect 623464 515872 624408 516096
rect 614496 515328 615040 515552
rect 622264 515328 623208 515552
rect 613536 514784 614080 515008
rect 621064 514784 622008 515008
rect 612576 514240 613120 514464
rect 619864 514240 620808 514464
rect 611616 513696 612160 513920
rect 618664 513696 619608 513920
rect 4612 512608 5556 512832
rect 22380 512608 22924 512832
rect 5812 512064 6756 512288
rect 21420 512064 21964 512288
rect 7012 511520 7956 511744
rect 15660 511520 16204 511744
rect 8212 510976 9156 511200
rect 16620 510976 17164 511200
rect 9412 510432 10356 510656
rect 17580 510432 18124 510656
rect 10612 509888 11556 510112
rect 18540 509888 19084 510112
rect 11812 509344 12756 509568
rect 19500 509344 20044 509568
rect 13012 508800 13956 509024
rect 20460 508800 21004 509024
rect 609696 504448 610240 504672
rect 627064 504448 628008 504672
rect 610656 503904 611200 504128
rect 625864 503904 626808 504128
rect 616416 503360 616960 503584
rect 624664 503360 625608 503584
rect 615456 502816 616000 503040
rect 623464 502816 624408 503040
rect 614496 502272 615040 502496
rect 622264 502272 623208 502496
rect 613536 501728 614080 501952
rect 621064 501728 622008 501952
rect 612576 501184 613120 501408
rect 619864 501184 620808 501408
rect 611616 500640 612160 500864
rect 618664 500640 619608 500864
rect 4612 499552 5556 499776
rect 22380 499552 22924 499776
rect 5812 499008 6756 499232
rect 21420 499008 21964 499232
rect 7012 498464 7956 498688
rect 15660 498464 16204 498688
rect 8212 497920 9156 498144
rect 16620 497920 17164 498144
rect 9412 497376 10356 497600
rect 17580 497376 18124 497600
rect 10612 496832 11556 497056
rect 18540 496832 19084 497056
rect 11812 496288 12756 496512
rect 19500 496288 20044 496512
rect 13012 495744 13956 495968
rect 20460 495744 21004 495968
rect 609696 491392 610240 491616
rect 627064 491392 628008 491616
rect 610656 490848 611200 491072
rect 625864 490848 626808 491072
rect 616416 490304 616960 490528
rect 624664 490304 625608 490528
rect 615456 489760 616000 489984
rect 623464 489760 624408 489984
rect 614496 489216 615040 489440
rect 622264 489216 623208 489440
rect 613536 488672 614080 488896
rect 621064 488672 622008 488896
rect 612576 488128 613120 488352
rect 619864 488128 620808 488352
rect 611616 487584 612160 487808
rect 618664 487584 619608 487808
rect 4612 486496 5556 486720
rect 22380 486496 22924 486720
rect 5812 485952 6756 486176
rect 21420 485952 21964 486176
rect 7012 485408 7956 485632
rect 15660 485408 16204 485632
rect 8212 484864 9156 485088
rect 16620 484864 17164 485088
rect 9412 484320 10356 484544
rect 17580 484320 18124 484544
rect 10612 483776 11556 484000
rect 18540 483776 19084 484000
rect 11812 483232 12756 483456
rect 19500 483232 20044 483456
rect 13012 482688 13956 482912
rect 20460 482688 21004 482912
rect 609696 476704 610240 476928
rect 627064 476704 628008 476928
rect 610656 476160 611200 476384
rect 625864 476160 626808 476384
rect 616416 475616 616960 475840
rect 624664 475616 625608 475840
rect 615456 475072 616000 475296
rect 623464 475072 624408 475296
rect 614496 474528 615040 474752
rect 622264 474528 623208 474752
rect 613536 473984 614080 474208
rect 621064 473984 622008 474208
rect 612576 473440 613120 473664
rect 619864 473440 620808 473664
rect 611616 472896 612160 473120
rect 618664 472896 619608 473120
rect 631301 471895 634165 476519
rect 4612 471264 5556 471488
rect 22380 471264 22924 471488
rect 5812 470720 6756 470944
rect 21420 470720 21964 470944
rect 7012 470176 7956 470400
rect 15660 470176 16204 470400
rect 8212 469632 9156 469856
rect 16620 469632 17164 469856
rect 9412 469088 10356 469312
rect 17580 469088 18124 469312
rect 10612 468544 11556 468768
rect 18540 468544 19084 468768
rect 11812 468000 12756 468224
rect 19500 468000 20044 468224
rect 13012 467456 13956 467680
rect 20460 467456 21004 467680
rect 609696 463648 610240 463872
rect 627064 463648 628008 463872
rect 610656 463104 611200 463328
rect 625864 463104 626808 463328
rect 616416 462560 616960 462784
rect 624664 462560 625608 462784
rect 615456 462016 616000 462240
rect 623464 462016 624408 462240
rect 631301 461912 634165 466536
rect 614496 461472 615040 461696
rect 622264 461472 623208 461696
rect 613536 460928 614080 461152
rect 621064 460928 622008 461152
rect 4612 460384 5556 460608
rect 22380 460384 22924 460608
rect 612576 460384 613120 460608
rect 619864 460384 620808 460608
rect 5812 459840 6756 460064
rect 21420 459840 21964 460064
rect 611616 459840 612160 460064
rect 618664 459840 619608 460064
rect 7012 459296 7956 459520
rect 15660 459296 16204 459520
rect 8212 458752 9156 458976
rect 16620 458752 17164 458976
rect 9412 458208 10356 458432
rect 17580 458208 18124 458432
rect 10612 457664 11556 457888
rect 18540 457664 19084 457888
rect 11812 457120 12756 457344
rect 19500 457120 20044 457344
rect 13012 456576 13956 456800
rect 20460 456576 21004 456800
rect -1777 451052 1087 455676
rect 609696 450592 610240 450816
rect 627064 450592 628008 450816
rect 610656 450048 611200 450272
rect 625864 450048 626808 450272
rect 616416 449504 616960 449728
rect 624664 449504 625608 449728
rect 615456 448960 616000 449184
rect 623464 448960 624408 449184
rect 614496 448416 615040 448640
rect 622264 448416 623208 448640
rect 613536 447872 614080 448096
rect 621064 447872 622008 448096
rect 4612 447328 5556 447552
rect 22380 447328 22924 447552
rect 612576 447328 613120 447552
rect 619864 447328 620808 447552
rect 5812 446784 6756 447008
rect 21420 446784 21964 447008
rect 611616 446784 612160 447008
rect 618664 446784 619608 447008
rect 7012 446240 7956 446464
rect 15660 446240 16204 446464
rect -1777 441073 1087 445697
rect 8212 445696 9156 445920
rect 16620 445696 17164 445920
rect 9412 445152 10356 445376
rect 17580 445152 18124 445376
rect 10612 444608 11556 444832
rect 18540 444608 19084 444832
rect 11812 444064 12756 444288
rect 19500 444064 20044 444288
rect 13012 443520 13956 443744
rect 20460 443520 21004 443744
rect 609696 437536 610240 437760
rect 627064 437536 628008 437760
rect 610656 436992 611200 437216
rect 625864 436992 626808 437216
rect 616416 436448 616960 436672
rect 624664 436448 625608 436672
rect 615456 435904 616000 436128
rect 623464 435904 624408 436128
rect 614496 435360 615040 435584
rect 622264 435360 623208 435584
rect 613536 434816 614080 435040
rect 621064 434816 622008 435040
rect 4612 434272 5556 434496
rect 22380 434272 22924 434496
rect 612576 434272 613120 434496
rect 619864 434272 620808 434496
rect 5812 433728 6756 433952
rect 21420 433728 21964 433952
rect 611616 433728 612160 433952
rect 618664 433728 619608 433952
rect 7012 433184 7956 433408
rect 15660 433184 16204 433408
rect 8212 432640 9156 432864
rect 16620 432640 17164 432864
rect 9412 432096 10356 432320
rect 17580 432096 18124 432320
rect 10612 431552 11556 431776
rect 18540 431552 19084 431776
rect 11812 431008 12756 431232
rect 19500 431008 20044 431232
rect 13012 430464 13956 430688
rect 20460 430464 21004 430688
rect 631301 427894 634165 432518
rect 609696 424480 610240 424704
rect 627064 424480 628008 424704
rect 610656 423936 611200 424160
rect 625864 423936 626808 424160
rect 616416 423392 616960 423616
rect 624664 423392 625608 423616
rect 615456 422848 616000 423072
rect 623464 422848 624408 423072
rect 631301 422944 634165 427408
rect 614496 422304 615040 422528
rect 622264 422304 623208 422528
rect 613536 421760 614080 421984
rect 621064 421760 622008 421984
rect 4612 421216 5556 421440
rect 22380 421216 22924 421440
rect 612576 421216 613120 421440
rect 619864 421216 620808 421440
rect 5812 420672 6756 420896
rect 21420 420672 21964 420896
rect 611616 420672 612160 420896
rect 618664 420672 619608 420896
rect 7012 420128 7956 420352
rect 15660 420128 16204 420352
rect 8212 419584 9156 419808
rect 16620 419584 17164 419808
rect 9412 419040 10356 419264
rect 17580 419040 18124 419264
rect 10612 418496 11556 418720
rect 18540 418496 19084 418720
rect 11812 417952 12756 418176
rect 19500 417952 20044 418176
rect 631301 417843 634165 422467
rect 13012 417408 13956 417632
rect 20460 417408 21004 417632
rect -1777 408934 1087 413558
rect 609696 411424 610240 411648
rect 627064 411424 628008 411648
rect 610656 410880 611200 411104
rect 625864 410880 626808 411104
rect 616416 410336 616960 410560
rect 624664 410336 625608 410560
rect 615456 409792 616000 410016
rect 623464 409792 624408 410016
rect 614496 409248 615040 409472
rect 622264 409248 623208 409472
rect 613536 408704 614080 408928
rect 621064 408704 622008 408928
rect -1777 403984 1087 408448
rect 4612 408160 5556 408384
rect 22380 408160 22924 408384
rect 612576 408160 613120 408384
rect 619864 408160 620808 408384
rect 5812 407616 6756 407840
rect 21420 407616 21964 407840
rect 611616 407616 612160 407840
rect 618664 407616 619608 407840
rect 7012 407072 7956 407296
rect 15660 407072 16204 407296
rect 8212 406528 9156 406752
rect 16620 406528 17164 406752
rect 9412 405984 10356 406208
rect 17580 405984 18124 406208
rect 10612 405440 11556 405664
rect 18540 405440 19084 405664
rect 11812 404896 12756 405120
rect 19500 404896 20044 405120
rect 13012 404352 13956 404576
rect 20460 404352 21004 404576
rect -1777 398894 1087 403518
rect 609696 398368 610240 398592
rect 627064 398368 628008 398592
rect 610656 397824 611200 398048
rect 625864 397824 626808 398048
rect 616416 397280 616960 397504
rect 624664 397280 625608 397504
rect 615456 396736 616000 396960
rect 623464 396736 624408 396960
rect 614496 396192 615040 396416
rect 622264 396192 623208 396416
rect 613536 395648 614080 395872
rect 621064 395648 622008 395872
rect 4612 395104 5556 395328
rect 22380 395104 22924 395328
rect 612576 395104 613120 395328
rect 619864 395104 620808 395328
rect 5812 394560 6756 394784
rect 21420 394560 21964 394784
rect 611616 394560 612160 394784
rect 618664 394560 619608 394784
rect 7012 394016 7956 394240
rect 15660 394016 16204 394240
rect 8212 393472 9156 393696
rect 16620 393472 17164 393696
rect 9412 392928 10356 393152
rect 17580 392928 18124 393152
rect 10612 392384 11556 392608
rect 18540 392384 19084 392608
rect 11812 391840 12756 392064
rect 19500 391840 20044 392064
rect 13012 391296 13956 391520
rect 20460 391296 21004 391520
rect 609696 385312 610240 385536
rect 627064 385312 628008 385536
rect 610656 384768 611200 384992
rect 625864 384768 626808 384992
rect 616416 384224 616960 384448
rect 624664 384224 625608 384448
rect 615456 383680 616000 383904
rect 623464 383680 624408 383904
rect 631301 383703 634165 388327
rect 614496 383136 615040 383360
rect 622264 383136 623208 383360
rect 613536 382592 614080 382816
rect 621064 382592 622008 382816
rect 4612 382048 5556 382272
rect 22380 382048 22924 382272
rect 612576 382048 613120 382272
rect 619864 382048 620808 382272
rect 5812 381504 6756 381728
rect 21420 381504 21964 381728
rect 611616 381504 612160 381728
rect 618664 381504 619608 381728
rect 7012 380960 7956 381184
rect 15660 380960 16204 381184
rect 8212 380416 9156 380640
rect 16620 380416 17164 380640
rect 9412 379872 10356 380096
rect 17580 379872 18124 380096
rect 10612 379328 11556 379552
rect 18540 379328 19084 379552
rect 11812 378784 12756 379008
rect 19500 378784 20044 379008
rect 13012 378240 13956 378464
rect 20460 378240 21004 378464
rect 631301 373720 634165 378344
rect 4612 368992 5556 369216
rect 22380 368992 22924 369216
rect 609696 368992 610240 369216
rect 627064 368992 628008 369216
rect 5812 368448 6756 368672
rect 21420 368448 21964 368672
rect 610656 368448 611200 368672
rect 625864 368448 626808 368672
rect 7012 367904 7956 368128
rect 15660 367904 16204 368128
rect 616416 367904 616960 368128
rect 624664 367904 625608 368128
rect 8212 367360 9156 367584
rect 16620 367360 17164 367584
rect 615456 367360 616000 367584
rect 623464 367360 624408 367584
rect 9412 366816 10356 367040
rect 17580 366816 18124 367040
rect 614496 366816 615040 367040
rect 622264 366816 623208 367040
rect 10612 366272 11556 366496
rect 18540 366272 19084 366496
rect 613536 366272 614080 366496
rect 621064 366272 622008 366496
rect 11812 365728 12756 365952
rect 19500 365728 20044 365952
rect 612576 365728 613120 365952
rect 619864 365728 620808 365952
rect 13012 365184 13956 365408
rect 20460 365184 21004 365408
rect 611616 365184 612160 365408
rect 618664 365184 619608 365408
rect 4612 355936 5556 356160
rect 22380 355936 22924 356160
rect 609696 355936 610240 356160
rect 627064 355936 628008 356160
rect 5812 355392 6756 355616
rect 21420 355392 21964 355616
rect 610656 355392 611200 355616
rect 625864 355392 626808 355616
rect 7012 354848 7956 355072
rect 15660 354848 16204 355072
rect 616416 354848 616960 355072
rect 624664 354848 625608 355072
rect 8212 354304 9156 354528
rect 16620 354304 17164 354528
rect 615456 354304 616000 354528
rect 623464 354304 624408 354528
rect 9412 353760 10356 353984
rect 17580 353760 18124 353984
rect 614496 353760 615040 353984
rect 622264 353760 623208 353984
rect 10612 353216 11556 353440
rect 18540 353216 19084 353440
rect 613536 353216 614080 353440
rect 621064 353216 622008 353440
rect 11812 352672 12756 352896
rect 19500 352672 20044 352896
rect 612576 352672 613120 352896
rect 619864 352672 620808 352896
rect 13012 352128 13956 352352
rect 20460 352128 21004 352352
rect 611616 352128 612160 352352
rect 618664 352128 619608 352352
rect 609696 342880 610240 343104
rect 627064 342880 628008 343104
rect 610656 342336 611200 342560
rect 625864 342336 626808 342560
rect 616416 341792 616960 342016
rect 624664 341792 625608 342016
rect 615456 341248 616000 341472
rect 623464 341248 624408 341472
rect 4612 340704 5556 340928
rect 22380 340704 22924 340928
rect 614496 340704 615040 340928
rect 622264 340704 623208 340928
rect 5812 340160 6756 340384
rect 21420 340160 21964 340384
rect 613536 340160 614080 340384
rect 621064 340160 622008 340384
rect 7012 339616 7956 339840
rect 15660 339616 16204 339840
rect 612576 339616 613120 339840
rect 619864 339616 620808 339840
rect 8212 339072 9156 339296
rect 16620 339072 17164 339296
rect 611616 339072 612160 339296
rect 618664 339072 619608 339296
rect 9412 338528 10356 338752
rect 17580 338528 18124 338752
rect 10612 337984 11556 338208
rect 18540 337984 19084 338208
rect 11812 337440 12756 337664
rect 19500 337440 20044 337664
rect 13012 336896 13956 337120
rect 20460 336896 21004 337120
rect 4612 329824 5556 330048
rect 22380 329824 22924 330048
rect 609696 329824 610240 330048
rect 627064 329824 628008 330048
rect 5812 329280 6756 329504
rect 21420 329280 21964 329504
rect 610656 329280 611200 329504
rect 625864 329280 626808 329504
rect 7012 328736 7956 328960
rect 15660 328736 16204 328960
rect 616416 328736 616960 328960
rect 624664 328736 625608 328960
rect 8212 328192 9156 328416
rect 16620 328192 17164 328416
rect 615456 328192 616000 328416
rect 623464 328192 624408 328416
rect 9412 327648 10356 327872
rect 17580 327648 18124 327872
rect 614496 327648 615040 327872
rect 622264 327648 623208 327872
rect 10612 327104 11556 327328
rect 18540 327104 19084 327328
rect 613536 327104 614080 327328
rect 621064 327104 622008 327328
rect 11812 326560 12756 326784
rect 19500 326560 20044 326784
rect 612576 326560 613120 326784
rect 619864 326560 620808 326784
rect 13012 326016 13956 326240
rect 20460 326016 21004 326240
rect 611616 326016 612160 326240
rect 618664 326016 619608 326240
rect 609696 318400 610240 318624
rect 627064 318400 628008 318624
rect 610656 317856 611200 318080
rect 625864 317856 626808 318080
rect 616416 317312 616960 317536
rect 624664 317312 625608 317536
rect 4612 316768 5556 316992
rect 22380 316768 22924 316992
rect 615456 316768 616000 316992
rect 623464 316768 624408 316992
rect 5812 316224 6756 316448
rect 21420 316224 21964 316448
rect 614496 316224 615040 316448
rect 622264 316224 623208 316448
rect 7012 315680 7956 315904
rect 15660 315680 16204 315904
rect 613536 315680 614080 315904
rect 621064 315680 622008 315904
rect 8212 315136 9156 315360
rect 16620 315136 17164 315360
rect 612576 315136 613120 315360
rect 619864 315136 620808 315360
rect 9412 314592 10356 314816
rect 17580 314592 18124 314816
rect 611616 314592 612160 314816
rect 618664 314592 619608 314816
rect 10612 314048 11556 314272
rect 18540 314048 19084 314272
rect 11812 313504 12756 313728
rect 19500 313504 20044 313728
rect 13012 312960 13956 313184
rect 20460 312960 21004 313184
rect 4612 305888 5556 306112
rect 22380 305888 22924 306112
rect 5812 305344 6756 305568
rect 21420 305344 21964 305568
rect 7012 304800 7956 305024
rect 15660 304800 16204 305024
rect 8212 304256 9156 304480
rect 16620 304256 17164 304480
rect 9412 303712 10356 303936
rect 17580 303712 18124 303936
rect 609696 303712 610240 303936
rect 627064 303712 628008 303936
rect 10612 303168 11556 303392
rect 18540 303168 19084 303392
rect 610656 303168 611200 303392
rect 625864 303168 626808 303392
rect 11812 302624 12756 302848
rect 19500 302624 20044 302848
rect 616416 302624 616960 302848
rect 624664 302624 625608 302848
rect 13012 302080 13956 302304
rect 20460 302080 21004 302304
rect 615456 302080 616000 302304
rect 623464 302080 624408 302304
rect 614496 301536 615040 301760
rect 622264 301536 623208 301760
rect 613536 300992 614080 301216
rect 621064 300992 622008 301216
rect 612576 300448 613120 300672
rect 619864 300448 620808 300672
rect 611616 299904 612160 300128
rect 618664 299904 619608 300128
rect 4612 290656 5556 290880
rect 22380 290656 22924 290880
rect 609696 290656 610240 290880
rect 627064 290656 628008 290880
rect 5812 290112 6756 290336
rect 21420 290112 21964 290336
rect 610656 290112 611200 290336
rect 625864 290112 626808 290336
rect 7012 289568 7956 289792
rect 15660 289568 16204 289792
rect 616416 289568 616960 289792
rect 624664 289568 625608 289792
rect 8212 289024 9156 289248
rect 16620 289024 17164 289248
rect 615456 289024 616000 289248
rect 623464 289024 624408 289248
rect 9412 288480 10356 288704
rect 17580 288480 18124 288704
rect 614496 288480 615040 288704
rect 622264 288480 623208 288704
rect 10612 287936 11556 288160
rect 18540 287936 19084 288160
rect 613536 287936 614080 288160
rect 621064 287936 622008 288160
rect 11812 287392 12756 287616
rect 19500 287392 20044 287616
rect 612576 287392 613120 287616
rect 619864 287392 620808 287616
rect 13012 286848 13956 287072
rect 20460 286848 21004 287072
rect 611616 286848 612160 287072
rect 618664 286848 619608 287072
rect 4612 277600 5556 277824
rect 22380 277600 22924 277824
rect 609696 277600 610240 277824
rect 627064 277600 628008 277824
rect 5812 277056 6756 277280
rect 21420 277056 21964 277280
rect 610656 277056 611200 277280
rect 625864 277056 626808 277280
rect 7012 276512 7956 276736
rect 15660 276512 16204 276736
rect 616416 276512 616960 276736
rect 624664 276512 625608 276736
rect 8212 275968 9156 276192
rect 16620 275968 17164 276192
rect 615456 275968 616000 276192
rect 623464 275968 624408 276192
rect 9412 275424 10356 275648
rect 17580 275424 18124 275648
rect 614496 275424 615040 275648
rect 622264 275424 623208 275648
rect 10612 274880 11556 275104
rect 18540 274880 19084 275104
rect 613536 274880 614080 275104
rect 621064 274880 622008 275104
rect 11812 274336 12756 274560
rect 19500 274336 20044 274560
rect 612576 274336 613120 274560
rect 619864 274336 620808 274560
rect 13012 273792 13956 274016
rect 20460 273792 21004 274016
rect 611616 273792 612160 274016
rect 618664 273792 619608 274016
rect 4612 266720 5556 266944
rect 22380 266720 22924 266944
rect 5812 266176 6756 266400
rect 21420 266176 21964 266400
rect 7012 265632 7956 265856
rect 15660 265632 16204 265856
rect 8212 265088 9156 265312
rect 16620 265088 17164 265312
rect 9412 264544 10356 264768
rect 17580 264544 18124 264768
rect 10612 264000 11556 264224
rect 18540 264000 19084 264224
rect 11812 263456 12756 263680
rect 19500 263456 20044 263680
rect 13012 262912 13956 263136
rect 20460 262912 21004 263136
rect 609696 262912 610240 263136
rect 627064 262912 628008 263136
rect 610656 262368 611200 262592
rect 625864 262368 626808 262592
rect 616416 261824 616960 262048
rect 624664 261824 625608 262048
rect 615456 261280 616000 261504
rect 623464 261280 624408 261504
rect 614496 260736 615040 260960
rect 622264 260736 623208 260960
rect 613536 260192 614080 260416
rect 621064 260192 622008 260416
rect 612576 259648 613120 259872
rect 619864 259648 620808 259872
rect 611616 259104 612160 259328
rect 618664 259104 619608 259328
rect 4612 251488 5556 251712
rect 22380 251488 22924 251712
rect 609696 251488 610240 251712
rect 627064 251488 628008 251712
rect 5812 250944 6756 251168
rect 21420 250944 21964 251168
rect 610656 250944 611200 251168
rect 625864 250944 626808 251168
rect 7012 250400 7956 250624
rect 15660 250400 16204 250624
rect 616416 250400 616960 250624
rect 624664 250400 625608 250624
rect 8212 249856 9156 250080
rect 16620 249856 17164 250080
rect 615456 249856 616000 250080
rect 623464 249856 624408 250080
rect 9412 249312 10356 249536
rect 17580 249312 18124 249536
rect 614496 249312 615040 249536
rect 622264 249312 623208 249536
rect 10612 248768 11556 248992
rect 18540 248768 19084 248992
rect 613536 248768 614080 248992
rect 621064 248768 622008 248992
rect 11812 248224 12756 248448
rect 19500 248224 20044 248448
rect 612576 248224 613120 248448
rect 619864 248224 620808 248448
rect 13012 247680 13956 247904
rect 20460 247680 21004 247904
rect 611616 247680 612160 247904
rect 618664 247680 619608 247904
rect 4612 238432 5556 238656
rect 22380 238432 22924 238656
rect 609696 238432 610240 238656
rect 627064 238432 628008 238656
rect 5812 237888 6756 238112
rect 21420 237888 21964 238112
rect 610656 237888 611200 238112
rect 625864 237888 626808 238112
rect 7012 237344 7956 237568
rect 15660 237344 16204 237568
rect 616416 237344 616960 237568
rect 624664 237344 625608 237568
rect 8212 236800 9156 237024
rect 16620 236800 17164 237024
rect 615456 236800 616000 237024
rect 623464 236800 624408 237024
rect 9412 236256 10356 236480
rect 17580 236256 18124 236480
rect 614496 236256 615040 236480
rect 622264 236256 623208 236480
rect 10612 235712 11556 235936
rect 18540 235712 19084 235936
rect 613536 235712 614080 235936
rect 621064 235712 622008 235936
rect 11812 235168 12756 235392
rect 19500 235168 20044 235392
rect 612576 235168 613120 235392
rect 619864 235168 620808 235392
rect 13012 234624 13956 234848
rect 20460 234624 21004 234848
rect 611616 234624 612160 234848
rect 618664 234624 619608 234848
rect 4612 225376 5556 225600
rect 22380 225376 22924 225600
rect 609696 225376 610240 225600
rect 627064 225376 628008 225600
rect 5812 224832 6756 225056
rect 21420 224832 21964 225056
rect 610656 224832 611200 225056
rect 625864 224832 626808 225056
rect 7012 224288 7956 224512
rect 15660 224288 16204 224512
rect 616416 224288 616960 224512
rect 624664 224288 625608 224512
rect 8212 223744 9156 223968
rect 16620 223744 17164 223968
rect 615456 223744 616000 223968
rect 623464 223744 624408 223968
rect 9412 223200 10356 223424
rect 17580 223200 18124 223424
rect 614496 223200 615040 223424
rect 622264 223200 623208 223424
rect 10612 222656 11556 222880
rect 18540 222656 19084 222880
rect 613536 222656 614080 222880
rect 621064 222656 622008 222880
rect 11812 222112 12756 222336
rect 19500 222112 20044 222336
rect 612576 222112 613120 222336
rect 619864 222112 620808 222336
rect 13012 221568 13956 221792
rect 20460 221568 21004 221792
rect 611616 221568 612160 221792
rect 618664 221568 619608 221792
rect 609696 212320 610240 212544
rect 627064 212320 628008 212544
rect 610656 211776 611200 212000
rect 625864 211776 626808 212000
rect 4612 211232 5556 211456
rect 22380 211232 22924 211456
rect 616416 211232 616960 211456
rect 624664 211232 625608 211456
rect 5812 210688 6756 210912
rect 21420 210688 21964 210912
rect 615456 210688 616000 210912
rect 623464 210688 624408 210912
rect 7012 210144 7956 210368
rect 15660 210144 16204 210368
rect 614496 210144 615040 210368
rect 622264 210144 623208 210368
rect 8212 209600 9156 209824
rect 16620 209600 17164 209824
rect 613536 209600 614080 209824
rect 621064 209600 622008 209824
rect 9412 209056 10356 209280
rect 17580 209056 18124 209280
rect 612576 209056 613120 209280
rect 619864 209056 620808 209280
rect 10612 208512 11556 208736
rect 18540 208512 19084 208736
rect 611616 208512 612160 208736
rect 618664 208512 619608 208736
rect 11812 207968 12756 208192
rect 19500 207968 20044 208192
rect 13012 207424 13956 207648
rect 20460 207424 21004 207648
rect -1777 36134 1087 40758
rect -1777 26094 1087 30718
rect 208191 27104 209055 27328
rect 226871 26664 227415 26888
rect 130995 7608 131859 7832
rect 139772 7589 139916 7733
rect 132347 6944 133211 7168
rect 138472 7025 138616 7169
rect 199023 -1696 203647 -112
rect 209074 -1696 213698 -112
<< metal4 >>
rect 533387 954354 538193 954482
rect 533387 952770 533467 954354
rect 538091 952770 538193 954354
rect 533387 931860 538193 952770
rect 533387 929704 533550 931860
rect 537946 929704 538193 931860
rect 533387 929492 538193 929704
rect 543368 954354 548174 954482
rect 543368 952770 543448 954354
rect 548072 952770 548174 954354
rect 543368 931860 548174 952770
rect 543368 929704 543531 931860
rect 547927 929704 548174 931860
rect 543368 929492 548174 929704
rect -1858 884758 1182 884840
rect -1858 880134 -1777 884758
rect 1087 880134 1182 884758
rect 631206 880318 634246 880400
rect -1858 880051 1182 880134
rect -1858 879648 1182 879730
rect -1858 875184 -1777 879648
rect 1087 875184 1182 879648
rect 631206 875694 631301 880318
rect 634165 875694 634246 880318
rect 631206 875611 634246 875694
rect -1858 875120 1182 875184
rect 631206 875208 634246 875290
rect -1858 874718 1182 874800
rect -1858 870094 -1777 874718
rect 1087 870094 1182 874718
rect 631206 870744 631301 875208
rect 634165 870744 634246 875208
rect 631206 870669 634246 870744
rect 631206 870267 634246 870349
rect -1858 870011 1182 870094
rect 631206 865643 631301 870267
rect 634165 865643 634246 870267
rect 631206 865560 634246 865643
rect -1858 800276 1182 800358
rect -1858 795652 -1777 800276
rect 1087 795652 1182 800276
rect -1858 795569 1182 795652
rect 631206 791119 634246 791201
rect -1858 790297 1182 790318
rect -1858 785673 -1777 790297
rect 1087 785673 1182 790297
rect 631206 786495 631301 791119
rect 634165 786495 634246 791119
rect 631206 786412 634246 786495
rect -1858 785589 1182 785673
rect 631206 781136 634246 781218
rect 631206 776512 631301 781136
rect 634165 776512 634246 781136
rect 631206 776429 634246 776512
rect 631206 476519 634246 476601
rect 631206 471895 631301 476519
rect 634165 471895 634246 476519
rect 631206 471812 634246 471895
rect 631206 466536 634246 466618
rect 631206 461912 631301 466536
rect 634165 461912 634246 466536
rect 631206 461829 634246 461912
rect -1858 455676 1182 455758
rect -1858 451052 -1777 455676
rect 1087 451052 1182 455676
rect -1858 450969 1182 451052
rect -1858 445697 1182 445718
rect -1858 441073 -1777 445697
rect 1087 441073 1182 445697
rect -1858 440989 1182 441073
rect 631206 432518 634246 432600
rect 631206 427894 631301 432518
rect 634165 427894 634246 432518
rect 631206 427811 634246 427894
rect 631206 427408 634246 427490
rect 631206 422944 631301 427408
rect 634165 422944 634246 427408
rect 631206 422869 634246 422944
rect 631206 422467 634246 422549
rect 631206 417843 631301 422467
rect 634165 417843 634246 422467
rect 631206 417760 634246 417843
rect -1858 413558 1182 413640
rect -1858 408934 -1777 413558
rect 1087 408934 1182 413558
rect -1858 408851 1182 408934
rect -1858 408448 1182 408530
rect -1858 403984 -1777 408448
rect 1087 403984 1182 408448
rect -1858 403920 1182 403984
rect -1858 403518 1182 403600
rect -1858 398894 -1777 403518
rect 1087 398894 1182 403518
rect -1858 398811 1182 398894
rect 631206 388327 634246 388409
rect 631206 383703 631301 388327
rect 634165 383703 634246 388327
rect 631206 383620 634246 383703
rect 631206 378344 634246 378426
rect 631206 373720 631301 378344
rect 634165 373720 634246 378344
rect 631206 373637 634246 373720
rect -1858 40758 1182 40840
rect -1858 36134 -1777 40758
rect 1087 36134 1182 40758
rect -1858 36051 1182 36134
rect -1858 30718 1182 30800
rect -1858 26094 -1777 30718
rect 1087 26094 1182 30718
rect 209504 27682 212862 28083
rect 223604 27047 226064 27376
rect -1858 26011 1182 26094
rect 137400 6414 137791 6496
rect 137400 6178 137476 6414
rect 137712 6178 137791 6414
rect 137400 6094 137791 6178
rect 137400 5858 137476 6094
rect 137712 5858 137791 6094
rect 137400 5774 137791 5858
rect 137400 5538 137476 5774
rect 137712 5538 137791 5774
rect 137400 5454 137791 5538
rect 137400 5218 137476 5454
rect 137712 5218 137791 5454
rect 137400 5134 137791 5218
rect 137400 4898 137476 5134
rect 137712 4898 137791 5134
rect 137400 4814 137791 4898
rect 137400 4578 137476 4814
rect 137712 4578 137791 4814
rect 137400 4497 137791 4578
rect 138800 4094 139282 6496
rect 138800 3858 138932 4094
rect 139168 3858 139282 4094
rect 138800 3774 139282 3858
rect 138800 3538 138932 3774
rect 139168 3538 139282 3774
rect 138800 3454 139282 3538
rect 138800 3218 138932 3454
rect 139168 3218 139282 3454
rect 138800 3134 139282 3218
rect 138800 2898 138932 3134
rect 139168 2898 139282 3134
rect 138800 2814 139282 2898
rect 138800 2578 138932 2814
rect 139168 2578 139282 2814
rect 138800 2494 139282 2578
rect 138800 2258 138932 2494
rect 139168 2258 139282 2494
rect 138800 2176 139282 2258
rect 198943 6414 203749 6496
rect 198943 4578 199106 6414
rect 203502 4578 203749 6414
rect 198943 -112 203749 4578
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -1824 203749 -1696
rect 208994 6414 213800 6496
rect 208994 4578 209157 6414
rect 213553 4578 213800 6414
rect 208994 -112 213800 4578
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -1824 213800 -1696
<< via4 >>
rect 533550 929704 537946 931860
rect 543531 929704 547927 931860
rect -1736 880322 1060 884718
rect 13046 880322 13922 884718
rect -1736 875212 1060 879608
rect 11846 875212 12722 879608
rect 627098 875882 627974 880278
rect 631328 875882 634124 880278
rect -1736 870282 1060 874678
rect 13046 874592 13922 874678
rect 13046 874368 13922 874592
rect 13046 870282 13922 874368
rect 625898 871328 626774 875168
rect 625898 871104 626774 871328
rect 625898 870772 626774 871104
rect 631328 870772 634124 875168
rect 627098 865831 627974 870227
rect 631328 865831 634124 870227
rect -1736 795840 1060 800236
rect 7046 798976 7922 800236
rect 7046 798752 7922 798976
rect 7046 795840 7922 798752
rect 621098 790816 621974 791079
rect 621098 790592 621974 790816
rect -1736 785861 1060 790257
rect 7046 785920 7922 790257
rect 621098 786683 621974 790592
rect 631328 786683 634124 791079
rect 7046 785861 7922 785920
rect 621098 777760 621974 781096
rect 621098 777536 621974 777760
rect 621098 776700 621974 777536
rect 631328 776700 634124 781096
rect 621098 474208 621974 476479
rect 621098 473984 621974 474208
rect 621098 472083 621974 473984
rect 631328 472083 634124 476479
rect 621098 462100 621974 466496
rect 631328 462100 634124 466496
rect -1736 451240 1060 455636
rect 8246 451240 9122 455636
rect -1736 441261 1060 445657
rect 8246 441261 9122 445657
rect 625898 428082 626774 432478
rect 631328 428082 634124 432478
rect 627098 424704 627974 427368
rect 627098 424480 627974 424704
rect 627098 422972 627974 424480
rect 631328 422972 634124 427368
rect 625898 418031 626774 422427
rect 631328 418031 634124 422427
rect -1736 409122 1060 413518
rect 11846 409122 12722 413518
rect -1736 404012 1060 408408
rect 13046 404576 13922 408408
rect 13046 404352 13922 404576
rect 13046 404012 13922 404352
rect -1736 399082 1060 403478
rect 11846 399082 12722 403478
rect 622298 383891 623174 388287
rect 631328 383891 634124 388287
rect 622298 373908 623174 378304
rect 631328 373908 634124 378304
rect -1736 36322 1060 40718
rect 2246 36322 3122 40718
rect -1736 26282 1060 30678
rect 2246 26282 3122 30678
rect 137476 6178 137712 6414
rect 137476 5858 137712 6094
rect 137476 5538 137712 5774
rect 137476 5218 137712 5454
rect 137476 4898 137712 5134
rect 137476 4578 137712 4814
rect 138932 3858 139168 4094
rect 138932 3538 139168 3774
rect 138932 3218 139168 3454
rect 138932 2898 139168 3134
rect 138932 2578 139168 2814
rect 138932 2258 139168 2494
rect 199106 4578 203502 6414
rect 209157 4578 213553 6414
<< metal5 >>
rect -1858 884718 13984 884840
rect -1858 880322 -1736 884718
rect 1060 880322 13046 884718
rect 13922 880322 13984 884718
rect -1858 880050 13984 880322
rect 627036 880278 634246 880400
rect -1858 879608 12784 879730
rect -1858 875212 -1736 879608
rect 1060 875212 11846 879608
rect 12722 875212 12784 879608
rect 627036 875882 627098 880278
rect 627974 875882 631328 880278
rect 634124 875882 634246 880278
rect 627036 875610 634246 875882
rect -1858 875120 12784 875212
rect 625836 875168 634246 875290
rect -1858 874678 13984 874800
rect -1858 870282 -1736 874678
rect 1060 870282 13046 874678
rect 13922 870282 13984 874678
rect 625836 870772 625898 875168
rect 626774 870772 631328 875168
rect 634124 870772 634246 875168
rect 625836 870669 634246 870772
rect -1858 870010 13984 870282
rect 627036 870227 634246 870349
rect 627036 865831 627098 870227
rect 627974 865831 631328 870227
rect 634124 865831 634246 870227
rect 627036 865559 634246 865831
rect -1858 800236 7984 800358
rect -1858 795840 -1736 800236
rect 1060 795840 7046 800236
rect 7922 795840 7984 800236
rect -1858 795568 7984 795840
rect 621036 791079 634246 791201
rect -1858 790257 7984 790379
rect -1858 785861 -1736 790257
rect 1060 785861 7046 790257
rect 7922 785861 7984 790257
rect 621036 786683 621098 791079
rect 621974 786683 631328 791079
rect 634124 786683 634246 791079
rect 621036 786411 634246 786683
rect -1858 785589 7984 785861
rect 621036 781096 634246 781218
rect 621036 776700 621098 781096
rect 621974 776700 631328 781096
rect 634124 776700 634246 781096
rect 621036 776428 634246 776700
rect 621036 476479 634246 476601
rect 621036 472083 621098 476479
rect 621974 472083 631328 476479
rect 634124 472083 634246 476479
rect 621036 471811 634246 472083
rect 621036 466496 634246 466618
rect 621036 462100 621098 466496
rect 621974 462100 631328 466496
rect 634124 462100 634246 466496
rect 621036 461828 634246 462100
rect -1858 455636 9184 455758
rect -1858 451240 -1736 455636
rect 1060 451240 8246 455636
rect 9122 451240 9184 455636
rect -1858 450968 9184 451240
rect -1858 445657 9184 445779
rect -1858 441261 -1736 445657
rect 1060 441261 8246 445657
rect 9122 441261 9184 445657
rect -1858 440989 9184 441261
rect 625836 432478 634246 432600
rect 625836 428082 625898 432478
rect 626774 428082 631328 432478
rect 634124 428082 634246 432478
rect 625836 427810 634246 428082
rect 627036 427368 634246 427490
rect 627036 422972 627098 427368
rect 627974 422972 631328 427368
rect 634124 422972 634246 427368
rect 627036 422869 634246 422972
rect 625836 422427 634246 422549
rect 625836 418031 625898 422427
rect 626774 418031 631328 422427
rect 634124 418031 634246 422427
rect 625836 417759 634246 418031
rect -1858 413518 12784 413640
rect -1858 409122 -1736 413518
rect 1060 409122 11846 413518
rect 12722 409122 12784 413518
rect -1858 408850 12784 409122
rect -1858 408408 13984 408530
rect -1858 404012 -1736 408408
rect 1060 404012 13046 408408
rect 13922 404012 13984 408408
rect -1858 403920 13984 404012
rect -1858 403478 12784 403600
rect -1858 399082 -1736 403478
rect 1060 399082 11846 403478
rect 12722 399082 12784 403478
rect -1858 398810 12784 399082
rect 622236 388287 634246 388409
rect 622236 383891 622298 388287
rect 623174 383891 631328 388287
rect 634124 383891 634246 388287
rect 622236 383619 634246 383891
rect 622236 378304 634246 378426
rect 622236 373908 622298 378304
rect 623174 373908 631328 378304
rect 634124 373908 634246 378304
rect 622236 373636 634246 373908
rect -1858 40718 3184 40840
rect -1858 36322 -1736 40718
rect 1060 36322 2246 40718
rect 3122 36322 3184 40718
rect -1858 36050 3184 36322
rect -1858 30678 3184 30800
rect -1858 26282 -1736 30678
rect 1060 26282 2246 30678
rect 3122 26282 3184 30678
rect -1858 26010 3184 26282
<< properties >>
string FIXED_BBOX 0 0 633000 953400
<< end >>
