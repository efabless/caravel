magic
tech sky130A
magscale 1 2
timestamp 1512359325
<< checkpaint >>
rect 38504 414288 679066 999106
<< metal3 >>
tri 81502 983518 82144 984160 se
rect 82144 984060 87144 997762
rect 82144 983518 86602 984060
tri 86602 983518 87144 984060 nw
rect 133544 983518 138544 997772
rect 81502 982718 86502 983518
tri 86502 983418 86602 983518 nw
rect 133502 983382 138544 983518
rect 184944 983518 189944 997736
rect 221000 995592 235279 997736
rect 221000 993848 221427 995592
rect 234851 993848 235279 995592
rect 221000 993420 235279 993848
tri 221000 984160 230260 993420 ne
rect 230260 984160 235279 993420
tri 230260 984060 230360 984160 ne
rect 230360 984060 235279 984160
tri 230360 983518 230902 984060 ne
rect 230902 983518 235279 984060
rect 235579 984141 237779 997736
rect 237978 984242 240178 997736
tri 237978 984141 238079 984242 ne
rect 238079 984141 240178 984242
tri 235579 983518 236202 984141 ne
rect 236202 983518 237779 984141
tri 238079 983868 238352 984141 ne
rect 238352 983868 240178 984141
rect 240478 995592 254800 997736
rect 240478 993848 240905 995592
rect 254329 993848 254800 995592
rect 240478 992116 254800 993848
rect 273600 995592 287879 997754
rect 273600 993848 274027 995592
rect 287451 993848 287879 995592
rect 273600 992520 287879 993848
tri 273600 992116 274004 992520 ne
rect 274004 992116 287879 992520
rect 240478 984242 246926 992116
tri 246926 984242 254800 992116 nw
tri 274004 984242 281878 992116 ne
rect 281878 984242 287879 992116
tri 240478 983868 240852 984242 ne
rect 240852 983868 246552 984242
tri 246552 983868 246926 984242 nw
tri 281878 983868 282252 984242 ne
rect 282252 983868 287879 984242
tri 237779 983518 238129 983868 sw
tri 238352 983518 238702 983868 ne
rect 238702 983518 240178 983868
tri 240178 983518 240528 983868 sw
tri 240852 983518 241202 983868 ne
rect 184944 983452 190502 983518
rect 133502 982718 138502 983382
rect 185502 982718 190502 983452
rect 230902 982718 235902 983518
rect 236202 982718 238402 983518
rect 238702 982718 240902 983518
rect 241202 982718 246202 983868
tri 246202 983518 246552 983868 nw
tri 282252 983518 282602 983868 ne
rect 282602 983795 287879 983868
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 288179 983795 290379 997754
rect 288179 983718 290302 983795
tri 290302 983718 290379 983795 nw
tri 287979 983518 288179 983718 se
rect 288179 983518 290102 983718
tri 290102 983518 290302 983718 nw
rect 290578 983694 292778 997754
tri 290402 983518 290578 983694 se
rect 290578 983518 292602 983694
tri 292602 983518 292778 983694 nw
rect 293078 995592 307400 997754
rect 293078 993848 293505 995592
rect 306929 993848 307400 995592
rect 293078 993016 307400 993848
rect 293078 992520 306904 993016
tri 306904 992520 307400 993016 nw
rect 375400 995592 389679 997722
rect 375400 993848 375827 995592
rect 389251 993848 389679 995592
rect 293078 983795 298179 992520
tri 298179 983795 306904 992520 nw
rect 375400 992420 389679 993848
tri 375400 983795 384025 992420 ne
rect 384025 983895 389679 992420
rect 384025 983795 389302 983895
rect 293078 983718 298102 983795
tri 298102 983718 298179 983795 nw
tri 384025 983718 384102 983795 ne
rect 384102 983718 389302 983795
rect 293078 983694 298078 983718
tri 298078 983694 298102 983718 nw
tri 384102 983694 384126 983718 ne
rect 384126 983694 389302 983718
rect 293078 983518 297902 983694
tri 297902 983518 298078 983694 nw
tri 384126 983518 384302 983694 ne
rect 287902 982718 290102 983518
rect 290402 982718 292602 983518
rect 292902 982718 297902 983518
rect 384302 982718 389302 983694
tri 389302 983518 389679 983895 nw
rect 389979 983895 392179 997722
rect 389979 983798 392082 983895
tri 392082 983798 392179 983895 nw
tri 389699 983518 389979 983798 se
rect 389979 983794 392078 983798
tri 392078 983794 392082 983798 nw
rect 392378 983794 394578 997722
rect 389979 983518 391802 983794
tri 391802 983518 392078 983794 nw
tri 392102 983518 392378 983794 se
rect 392378 983518 394302 983794
tri 394302 983518 394578 983794 nw
rect 394878 995592 409200 997722
rect 394878 993848 395305 995592
rect 408729 993848 409200 995592
rect 394878 993116 409200 993848
rect 394878 993016 409100 993116
tri 409100 993016 409200 993116 nw
rect 394878 992520 408604 993016
tri 408604 992520 409100 993016 nw
rect 394878 992420 408504 992520
tri 408504 992420 408604 992520 nw
rect 394878 983895 399979 992420
tri 399979 983895 408504 992420 nw
rect 394878 983798 399882 983895
tri 399882 983798 399979 983895 nw
rect 394878 983794 399878 983798
tri 399878 983794 399882 983798 nw
rect 394878 983518 399602 983794
tri 399602 983518 399878 983794 nw
rect 478744 983518 483744 997704
rect 530144 984064 535144 997792
tri 535144 984064 535156 984076 sw
tri 530144 983895 530313 984064 ne
rect 530313 983895 535156 984064
tri 530313 983798 530410 983895 ne
rect 530410 983798 535156 983895
tri 530410 983794 530414 983798 ne
rect 530414 983794 535156 983798
tri 530414 983518 530690 983794 ne
rect 530690 983518 535156 983794
tri 535156 983518 535702 984064 sw
rect 575700 983678 580479 997692
rect 585678 983741 590458 997692
tri 590458 983741 590479 983762 sw
tri 580479 983678 580542 983741 sw
rect 585678 983700 590479 983741
tri 590479 983700 590520 983741 sw
tri 585678 983678 585700 983700 ne
rect 585700 983678 590520 983700
tri 575700 983518 575860 983678 ne
rect 575860 983518 580542 983678
tri 580542 983518 580702 983678 sw
tri 585700 983518 585860 983678 ne
rect 585860 983518 590520 983678
tri 590520 983518 590702 983700 sw
rect 631944 983518 636944 997846
rect 389602 982718 391802 983518
rect 392102 982718 394302 983518
rect 394602 982718 399602 983518
rect 478702 983384 483744 983518
tri 530690 983506 530702 983518 ne
rect 478702 982718 483702 983384
rect 530702 982718 535702 983518
tri 575860 983506 575872 983518 ne
rect 575872 983506 580702 983518
tri 575872 983476 575902 983506 ne
rect 575902 982718 580702 983506
tri 585860 983476 585902 983518 ne
rect 585902 982718 590702 983518
rect 631902 983374 636944 983518
rect 631902 982718 636902 983374
rect 39764 963960 63464 965144
tri 63464 963960 64648 965144 sw
rect 39764 960144 65308 963960
tri 63325 958961 64508 960144 ne
rect 64508 958960 65308 960144
rect 649308 961656 650108 961702
rect 649308 956702 677806 961656
rect 650016 956656 677806 956702
rect 64508 926940 65308 927360
rect 41056 922560 65308 926940
rect 41056 922151 64552 922560
rect 649308 922502 650108 923302
tri 650108 922502 650908 923302 sw
rect 649308 918502 676480 922502
tri 649926 917700 650728 918502 ne
rect 650728 917700 676480 918502
rect 64508 916900 65308 917361
rect 41056 912560 65308 916900
rect 41056 912100 64560 912560
rect 649308 912449 650108 913302
tri 650108 912449 650961 913302 sw
rect 649308 908502 676480 912449
tri 649934 907660 650776 908502 ne
rect 650776 907660 676480 908502
tri 64006 842458 64508 842960 se
rect 64508 842458 65308 842960
rect 39900 838160 65308 842458
rect 39900 837678 64152 838160
tri 64152 837678 64634 838160 nw
rect 649308 833301 650108 834080
tri 64027 832479 64508 832960 se
rect 64508 832479 65308 832960
rect 39900 828160 65308 832479
rect 649308 829280 677632 833301
rect 649858 828521 677632 829280
rect 49892 828159 64634 828160
rect 39900 827699 64174 828159
tri 64174 827699 64634 828159 nw
rect 649308 823322 650108 824080
rect 649308 819280 677632 823322
rect 649858 818542 677632 819280
rect 649308 518701 650108 518748
rect 649308 513948 677632 518701
rect 650058 513921 667116 513948
rect 649308 508722 650108 508748
rect 649308 503948 677632 508722
rect 650066 503942 667124 503948
tri 63960 497858 64508 498406 se
rect 64508 497858 65308 498406
rect 39900 493606 65308 497858
rect 39900 493078 64012 493606
tri 64012 493078 64540 493606 nw
tri 63982 487879 64508 488405 se
rect 64508 487879 65308 488406
rect 39900 483606 65308 487879
rect 39900 483099 64041 483606
tri 64041 483099 64548 483606 nw
rect 649308 474700 650108 474948
rect 649308 470148 676178 474700
rect 650042 469900 676178 470148
rect 649308 464649 650108 464948
rect 649308 460148 676178 464649
rect 650042 459860 676178 460148
tri 63842 455740 64508 456406 se
rect 64508 455740 65308 456406
rect 41400 451606 65308 455740
rect 41400 450951 63927 451606
tri 63927 450951 64582 451606 nw
tri 63802 445700 64508 446406 se
rect 64508 445700 65308 446406
rect 41400 441606 65308 445700
rect 41400 440900 63858 441606
tri 63858 440900 64564 441606 nw
rect 650068 430348 677676 430501
rect 649308 425721 677676 430348
rect 649308 425562 677024 425721
rect 649308 425548 650108 425562
rect 650058 420348 677676 420522
rect 649308 415742 677676 420348
rect 649308 415548 650108 415742
<< via3 >>
rect 221427 993848 234851 995592
rect 240905 993848 254329 995592
rect 274027 993848 287451 995592
rect 293505 993848 306929 995592
rect 375827 993848 389251 995592
rect 395305 993848 408729 995592
<< metal4 >>
rect 221000 995592 235279 996020
rect 221000 993848 221427 995592
rect 234851 993848 235279 995592
rect 221000 993420 235279 993848
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995592 254757 996020
rect 240478 993848 240905 995592
rect 254329 993848 254757 995592
rect 240478 993820 254757 993848
rect 273600 995592 287879 996020
rect 273600 993848 274027 995592
rect 287451 993848 287879 995592
rect 240478 992116 254800 993820
rect 273600 992520 287879 993848
tri 273600 992116 274004 992520 ne
rect 274004 992116 287879 992520
rect 240478 984242 246926 992116
tri 246926 984242 254800 992116 nw
tri 274004 984242 281878 992116 ne
rect 281878 984242 287879 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 246926 984242 nw
tri 281878 983518 282602 984242 ne
rect 282602 983795 287879 984242
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995592 307357 996020
rect 293078 993848 293505 995592
rect 306929 993848 307357 995592
rect 293078 993820 307357 993848
rect 375400 995592 389679 996020
rect 375400 993848 375827 995592
rect 389251 993848 389679 995592
rect 293078 993016 307400 993820
rect 293078 992520 306904 993016
tri 306904 992520 307400 993016 nw
rect 293078 983795 298179 992520
tri 298179 983795 306904 992520 nw
rect 375400 992420 389679 993848
tri 375400 983795 384025 992420 ne
rect 384025 983895 389679 992420
rect 384025 983795 389302 983895
rect 293078 983518 297902 983795
tri 297902 983518 298179 983795 nw
tri 384025 983518 384302 983795 ne
rect 292902 982718 297902 983518
rect 384302 982718 389302 983795
tri 389302 983518 389679 983895 nw
rect 394878 995592 409157 996020
rect 394878 993848 395305 995592
rect 408729 993848 409157 995592
rect 394878 993820 409157 993848
rect 394878 993116 409200 993820
rect 394878 993016 409100 993116
tri 409100 993016 409200 993116 nw
rect 394878 992520 408604 993016
tri 408604 992520 409100 993016 nw
rect 394878 992420 408504 992520
tri 408504 992420 408604 992520 nw
rect 394878 983895 399979 992420
tri 399979 983895 408504 992420 nw
rect 394878 983518 399602 983895
tri 399602 983518 399979 983895 nw
rect 394602 982718 399602 983518
<< via4 >>
rect 221461 993962 234817 995478
rect 240939 993962 254295 995478
rect 274061 993962 287417 995478
rect 293539 993962 306895 995478
rect 375861 993962 389217 995478
rect 395339 993962 408695 995478
<< metal5 >>
rect 221000 995478 235279 996020
rect 221000 993962 221461 995478
rect 234817 993962 235279 995478
rect 221000 993420 235279 993962
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995478 254757 996020
rect 240478 993962 240939 995478
rect 254295 993962 254757 995478
rect 240478 993820 254757 993962
rect 273600 995478 287879 996020
rect 273600 993962 274061 995478
rect 287417 993962 287879 995478
rect 240478 992116 254800 993820
rect 273600 992520 287879 993962
tri 273600 992116 274004 992520 ne
rect 274004 992116 287879 992520
rect 240478 984242 246926 992116
tri 246926 984242 254800 992116 nw
tri 274004 984242 281878 992116 ne
rect 281878 984242 287879 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 246926 984242 nw
tri 281878 983518 282602 984242 ne
rect 282602 983795 287879 984242
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995478 307357 996020
rect 293078 993962 293539 995478
rect 306895 993962 307357 995478
rect 293078 993820 307357 993962
rect 375400 995478 389679 996020
rect 375400 993962 375861 995478
rect 389217 993962 389679 995478
rect 293078 993016 307400 993820
rect 293078 992520 306904 993016
tri 306904 992520 307400 993016 nw
rect 293078 983795 298179 992520
tri 298179 983795 306904 992520 nw
rect 375400 992420 389679 993962
tri 375400 983795 384025 992420 ne
rect 384025 983895 389679 992420
rect 384025 983795 389302 983895
rect 293078 983518 297902 983795
tri 297902 983518 298179 983795 nw
tri 384025 983518 384302 983795 ne
rect 292902 982718 297902 983518
rect 384302 982718 389302 983795
tri 389302 983518 389679 983895 nw
rect 394878 995478 409157 996020
rect 394878 993962 395339 995478
rect 408695 993962 409157 995478
rect 394878 993820 409157 993962
rect 394878 993116 409200 993820
rect 394878 993016 409100 993116
tri 409100 993016 409200 993116 nw
rect 394878 992520 408604 993016
tri 408604 992520 409100 993016 nw
rect 394878 992420 408504 992520
tri 408504 992420 408604 992520 nw
rect 394878 983895 399979 992420
tri 399979 983895 408504 992420 nw
rect 394878 983518 399602 983895
tri 399602 983518 399979 983895 nw
rect 394602 982718 399602 983518
<< properties >>
string FIXED_BBOX 19763 897847 697807 1017847
<< end >>
